module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
output n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 ;
wire n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
 n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
 n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
 n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
 n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
 n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
 n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
 n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
 n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
 n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
 n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
 n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , 
 n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
 n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , 
 n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , 
 n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , 
 n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , 
 n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , 
 n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , 
 n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , 
 n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , 
 n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , 
 n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , 
 n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , 
 n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , 
 n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , 
 n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , 
 n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , 
 n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , 
 n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
 n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , 
 n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
 n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , 
 n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , 
 n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , 
 n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
 n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
 n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
 n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , 
 n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , 
 n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , 
 n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
 n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , 
 n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , 
 n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , 
 n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
 n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
 n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
 n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , 
 n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , 
 n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
 n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , 
 n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , 
 n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , 
 n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
 n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
 n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , 
 n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
 n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
 n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , 
 n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , 
 n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , 
 n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , 
 n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , 
 n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , 
 n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , 
 n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
 n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , 
 n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , 
 n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , 
 n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , 
 n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , 
 n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , 
 n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , 
 n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , 
 n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , 
 n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , 
 n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
 n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , 
 n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , 
 n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , 
 n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
 n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
 n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , 
 n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , 
 n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , 
 n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , 
 n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , 
 n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , 
 n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , 
 n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , 
 n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , 
 n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , 
 n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , 
 n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
 n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
 n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
 n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
 n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
 n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
 n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , 
 n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , 
 n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , 
 n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
 n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
 n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
 n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
 n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
 n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
 n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
 n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
 n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
 n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
 n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
 n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
 n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
 n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , 
 n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , 
 n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , 
 n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , 
 n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , 
 n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
 n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , 
 n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , 
 n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , 
 n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , 
 n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
 n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
 n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
 n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , 
 n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , 
 n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , 
 n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , 
 n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
 n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , 
 n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , 
 n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , 
 n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , 
 n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , 
 n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , 
 n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , 
 n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , 
 n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , 
 n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , 
 n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , 
 n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
 n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , 
 n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , 
 n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , 
 n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , 
 n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , 
 n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , 
 n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , 
 n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , 
 n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , 
 n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , 
 n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , 
 n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , 
 n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , 
 n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , 
 n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
 n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , 
 n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
 n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , 
 n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , 
 n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , 
 n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , 
 n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
 n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , 
 n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , 
 n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , 
 n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , 
 n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , 
 n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , 
 n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
 n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
 n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , 
 n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , 
 n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , 
 n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , 
 n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , 
 n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
 n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , 
 n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , 
 n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , 
 n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , 
 n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , 
 n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , 
 n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , 
 n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , 
 n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , 
 n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
 n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
 n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , 
 n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , 
 n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , 
 n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , 
 n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , 
 n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , 
 n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , 
 n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , 
 n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
 n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
 n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , 
 n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , 
 n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
 n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
 n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
 n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
 n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , 
 n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , 
 n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , 
 n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , 
 n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , 
 n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , 
 n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , 
 n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , 
 n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , 
 n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , 
 n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , 
 n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , 
 n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , 
 n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , 
 n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , 
 n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , 
 n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , 
 n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , 
 n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , 
 n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , 
 n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , 
 n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , 
 n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , 
 n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , 
 n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , 
 n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , 
 n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , 
 n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , 
 n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , 
 n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , 
 n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , 
 n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , 
 n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , 
 n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , 
 n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , 
 n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , 
 n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , 
 n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , 
 n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , 
 n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , 
 n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , 
 n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , 
 n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , 
 n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , 
 n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
 n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
 n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , 
 n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , 
 n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , 
 n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , 
 n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , 
 n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , 
 n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , 
 n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , 
 n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , 
 n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , 
 n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , 
 n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , 
 n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , 
 n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , 
 n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , 
 n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , 
 n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , 
 n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , 
 n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , 
 n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , 
 n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , 
 n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , 
 n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , 
 n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , 
 n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , 
 n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , 
 n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , 
 n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
 n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , 
 n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
 n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
 n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
 n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
 n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , 
 n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
 n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , 
 n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
 n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , 
 n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , 
 n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , 
 n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , 
 n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , 
 n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , 
 n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , 
 n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , 
 n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , 
 n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , 
 n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , 
 n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , 
 n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , 
 n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , 
 n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , 
 n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
 n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
 n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
 n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , 
 n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , 
 n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , 
 n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , 
 n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , 
 n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , 
 n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , 
 n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
 n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , 
 n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
 n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
 n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
 n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
 n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
 n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
 n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
 n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , 
 n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , 
 n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
 n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , 
 n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
 n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
 n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
 n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
 n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
 n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , 
 n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , 
 n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , 
 n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , 
 n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , 
 n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
 n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , 
 n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , 
 n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , 
 n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , 
 n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , 
 n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , 
 n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , 
 n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , 
 n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , 
 n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
 n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , 
 n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , 
 n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , 
 n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , 
 n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , 
 n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , 
 n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , 
 n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , 
 n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , 
 n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , 
 n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , 
 n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , 
 n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , 
 n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , 
 n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , 
 n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , 
 n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , 
 n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , 
 n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , 
 n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , 
 n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , 
 n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , 
 n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , 
 n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , 
 n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , 
 n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , 
 n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , 
 n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , 
 n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , 
 n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , 
 n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , 
 n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , 
 n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , 
 n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , 
 n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , 
 n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , 
 n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , 
 n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , 
 n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , 
 n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , 
 n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , 
 n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , 
 n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , 
 n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , 
 n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , 
 n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , 
 n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , 
 n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , 
 n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , 
 n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , 
 n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , 
 n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , 
 n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , 
 n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , 
 n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , 
 n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , 
 n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , 
 n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , 
 n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , 
 n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , 
 n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , 
 n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , 
 n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , 
 n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , 
 n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , 
 n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , 
 n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
 n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , 
 n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , 
 n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , 
 n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , 
 n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , 
 n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , 
 n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
 n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , 
 n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , 
 n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
 n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
 n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , 
 n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , 
 n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , 
 n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , 
 n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , 
 n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , 
 n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , 
 n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , 
 n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , 
 n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , 
 n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , 
 n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
 n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , 
 n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , 
 n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , 
 n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , 
 n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , 
 n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , 
 n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , 
 n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , 
 n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , 
 n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , 
 n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , 
 n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , 
 n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , 
 n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , 
 n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , 
 n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , 
 n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , 
 n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , 
 n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , 
 n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , 
 n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , 
 n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , 
 n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , 
 n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , 
 n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , 
 n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , 
 n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , 
 n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , 
 n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , 
 n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , 
 n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , 
 n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , 
 n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , 
 n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , 
 n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , 
 n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , 
 n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , 
 n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , 
 n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , 
 n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , 
 n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , 
 n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , 
 n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , 
 n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , 
 n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , 
 n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , 
 n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , 
 n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , 
 n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , 
 n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , 
 n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , 
 n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , 
 n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , 
 n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , 
 n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , 
 n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , 
 n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , 
 n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , 
 n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , 
 n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , 
 n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , 
 n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , 
 n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , 
 n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , 
 n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , 
 n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , 
 n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , 
 n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , 
 n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , 
 n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , 
 n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
 n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
 n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , 
 n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , 
 n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , 
 n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , 
 n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , 
 n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , 
 n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , 
 n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , 
 n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , 
 n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , 
 n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , 
 n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , 
 n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , 
 n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , 
 n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , 
 n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , 
 n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , 
 n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , 
 n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , 
 n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , 
 n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , 
 n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , 
 n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , 
 n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , 
 n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , 
 n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , 
 n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , 
 n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , 
 n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , 
 n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , 
 n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , 
 n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , 
 n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , 
 n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , 
 n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , 
 n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , 
 n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , 
 n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , 
 n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , 
 n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , 
 n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , 
 n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , 
 n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , 
 n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , 
 n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , 
 n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , 
 n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , 
 n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , 
 n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , 
 n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , 
 n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , 
 n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , 
 n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , 
 n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , 
 n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , 
 n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , 
 n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , 
 n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , 
 n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , 
 n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , 
 n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , 
 n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , 
 n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , 
 n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , 
 n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , 
 n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , 
 n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , 
 n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
 n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , 
 n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , 
 n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , 
 n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , 
 n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , 
 n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , 
 n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , 
 n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , 
 n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
 n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
 n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
 n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
 n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
 n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , 
 n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , 
 n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , 
 n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , 
 n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , 
 n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , 
 n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , 
 n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , 
 n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , 
 n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , 
 n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , 
 n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , 
 n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , 
 n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , 
 n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , 
 n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , 
 n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
 n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
 n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , 
 n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , 
 n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , 
 n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , 
 n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , 
 n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , 
 n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , 
 n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , 
 n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , 
 n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , 
 n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , 
 n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , 
 n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , 
 n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , 
 n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , 
 n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , 
 n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , 
 n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , 
 n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , 
 n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , 
 n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , 
 n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , 
 n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , 
 n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , 
 n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , 
 n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , 
 n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , 
 n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , 
 n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , 
 n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , 
 n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , 
 n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , 
 n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , 
 n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , 
 n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , 
 n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , 
 n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
 n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
 n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
 n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , 
 n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , 
 n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , 
 n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , 
 n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , 
 n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , 
 n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , 
 n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , 
 n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , 
 n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , 
 n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , 
 n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , 
 n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , 
 n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
 n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , 
 n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , 
 n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , 
 n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , 
 n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , 
 n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , 
 n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , 
 n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
 n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
 n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
 n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
 n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , 
 n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , 
 n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
 n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
 n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
 n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
 n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
 n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
 n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
 n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
 n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
 n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
 n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , 
 n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , 
 n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , 
 n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , 
 n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , 
 n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , 
 n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , 
 n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , 
 n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , 
 n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , 
 n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , 
 n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , 
 n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , 
 n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , 
 n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , 
 n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , 
 n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , 
 n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , 
 n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , 
 n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , 
 n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , 
 n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , 
 n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , 
 n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , 
 n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , 
 n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , 
 n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , 
 n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , 
 n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , 
 n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , 
 n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , 
 n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , 
 n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , 
 n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , 
 n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , 
 n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , 
 n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , 
 n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , 
 n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , 
 n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , 
 n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , 
 n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , 
 n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , 
 n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , 
 n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , 
 n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , 
 n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , 
 n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , 
 n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , 
 n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , 
 n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
 n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , 
 n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , 
 n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , 
 n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , 
 n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , 
 n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , 
 n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , 
 n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , 
 n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , 
 n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , 
 n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , 
 n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , 
 n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , 
 n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , 
 n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , 
 n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , 
 n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , 
 n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , 
 n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , 
 n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , 
 n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , 
 n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , 
 n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , 
 n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , 
 n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , 
 n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , 
 n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , 
 n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , 
 n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , 
 n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , 
 n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , 
 n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , 
 n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , 
 n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , 
 n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , 
 n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , 
 n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , 
 n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , 
 n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , 
 n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , 
 n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , 
 n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , 
 n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , 
 n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , 
 n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , 
 n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , 
 n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , 
 n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , 
 n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , 
 n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , 
 n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , 
 n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , 
 n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , 
 n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , 
 n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , 
 n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , 
 n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , 
 n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , 
 n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , 
 n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , 
 n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , 
 n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , 
 n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , 
 n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , 
 n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , 
 n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , 
 n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , 
 n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , 
 n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , 
 n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , 
 n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , 
 n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , 
 n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , 
 n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , 
 n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , 
 n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , 
 n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , 
 n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , 
 n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , 
 n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , 
 n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , 
 n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , 
 n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , 
 n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , 
 n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , 
 n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , 
 n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , 
 n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , 
 n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , 
 n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , 
 n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , 
 n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , 
 n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , 
 n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , 
 n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , 
 n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , 
 n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , 
 n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , 
 n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , 
 n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , 
 n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , 
 n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , 
 n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , 
 n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , 
 n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , 
 n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , 
 n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , 
 n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , 
 n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , 
 n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , 
 n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , 
 n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , 
 n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , 
 n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , 
 n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , 
 n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , 
 n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , 
 n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , 
 n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , 
 n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , 
 n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , 
 n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , 
 n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , 
 n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , 
 n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , 
 n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , 
 n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , 
 n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , 
 n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , 
 n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , 
 n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , 
 n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , 
 n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , 
 n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , 
 n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , 
 n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , 
 n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , 
 n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , 
 n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , 
 n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , 
 n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , 
 n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , 
 n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , 
 n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , 
 n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , 
 n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
 n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , 
 n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , 
 n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , 
 n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
 n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , 
 n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
 n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
 n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , 
 n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , 
 n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , 
 n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , 
 n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , 
 n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , 
 n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , 
 n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , 
 n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , 
 n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , 
 n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , 
 n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , 
 n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , 
 n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , 
 n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , 
 n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , 
 n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , 
 n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , 
 n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , 
 n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , 
 n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , 
 n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , 
 n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , 
 n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , 
 n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , 
 n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , 
 n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , 
 n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , 
 n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , 
 n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , 
 n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , 
 n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , 
 n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , 
 n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , 
 n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , 
 n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , 
 n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , 
 n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , 
 n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , 
 n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , 
 n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , 
 n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , 
 n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , 
 n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , 
 n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , 
 n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , 
 n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , 
 n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , 
 n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , 
 n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , 
 n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , 
 n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , 
 n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , 
 n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , 
 n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , 
 n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , 
 n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , 
 n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , 
 n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , 
 n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , 
 n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , 
 n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , 
 n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , 
 n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , 
 n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , 
 n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , 
 n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , 
 n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , 
 n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , 
 n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , 
 n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , 
 n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , 
 n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , 
 n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , 
 n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , 
 n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , 
 n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , 
 n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , 
 n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , 
 n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , 
 n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , 
 n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , 
 n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , 
 n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , 
 n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , 
 n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , 
 n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , 
 n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , 
 n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , 
 n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , 
 n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , 
 n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , 
 n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , 
 n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , 
 n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , 
 n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , 
 n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , 
 n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , 
 n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , 
 n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , 
 n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , 
 n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , 
 n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , 
 n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , 
 n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , 
 n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , 
 n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , 
 n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , 
 n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , 
 n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , 
 n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , 
 n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , 
 n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , 
 n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , 
 n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , 
 n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , 
 n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , 
 n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , 
 n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , 
 n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , 
 n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , 
 n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , 
 n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , 
 n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , 
 n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , 
 n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , 
 n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , 
 n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , 
 n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , 
 n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , 
 n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , 
 n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , 
 n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , 
 n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , 
 n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , 
 n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , 
 n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , 
 n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , 
 n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , 
 n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , 
 n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , 
 n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , 
 n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , 
 n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , 
 n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , 
 n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , 
 n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , 
 n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , 
 n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , 
 n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , 
 n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , 
 n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , 
 n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , 
 n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , 
 n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , 
 n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , 
 n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , 
 n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , 
 n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , 
 n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , 
 n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , 
 n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , 
 n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , 
 n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , 
 n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , 
 n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , 
 n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , 
 n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , 
 n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , 
 n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , 
 n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , 
 n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , 
 n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , 
 n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , 
 n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , 
 n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , 
 n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , 
 n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , 
 n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , 
 n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , 
 n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , 
 n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , 
 n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , 
 n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , 
 n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , 
 n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , 
 n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , 
 n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , 
 n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , 
 n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , 
 n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , 
 n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , 
 n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , 
 n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , 
 n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , 
 n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , 
 n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , 
 n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , 
 n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , 
 n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , 
 n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , 
 n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , 
 n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , 
 n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , 
 n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , 
 n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , 
 n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , 
 n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , 
 n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , 
 n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , 
 n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , 
 n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , 
 n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , 
 n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , 
 n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , 
 n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , 
 n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , 
 n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , 
 n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , 
 n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , 
 n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , 
 n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , 
 n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , 
 n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , 
 n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , 
 n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , 
 n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , 
 n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , 
 n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , 
 n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , 
 n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , 
 n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , 
 n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , 
 n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , 
 n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , 
 n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , 
 n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , 
 n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , 
 n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , 
 n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , 
 n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , 
 n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , 
 n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , 
 n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , 
 n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , 
 n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , 
 n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , 
 n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , 
 n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , 
 n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , 
 n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , 
 n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , 
 n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , 
 n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , 
 n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , 
 n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , 
 n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , 
 n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , 
 n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , 
 n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , 
 n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , 
 n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , 
 n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , 
 n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , 
 n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , 
 n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , 
 n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , 
 n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , 
 n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , 
 n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , 
 n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , 
 n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , 
 n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , 
 n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , 
 n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , 
 n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , 
 n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , 
 n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , 
 n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , 
 n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , 
 n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , 
 n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , 
 n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , 
 n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , 
 n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , 
 n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , 
 n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , 
 n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , 
 n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , 
 n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , 
 n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , 
 n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , 
 n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , 
 n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , 
 n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , 
 n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , 
 n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , 
 n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , 
 n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , 
 n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , 
 n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , 
 n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , 
 n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , 
 n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , 
 n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , 
 n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , 
 n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , 
 n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , 
 n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , 
 n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , 
 n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , 
 n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , 
 n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , 
 n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , 
 n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , 
 n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , 
 n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , 
 n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , 
 n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , 
 n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , 
 n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , 
 n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , 
 n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , 
 n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , 
 n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , 
 n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , 
 n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , 
 n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , 
 n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , 
 n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , 
 n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , 
 n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , 
 n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , 
 n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , 
 n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , 
 n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , 
 n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , 
 n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , 
 n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , 
 n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , 
 n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , 
 n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , 
 n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , 
 n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , 
 n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , 
 n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , 
 n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , 
 n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , 
 n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
 n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , 
 n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , 
 n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , 
 n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , 
 n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , 
 n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , 
 n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , 
 n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , 
 n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , 
 n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , 
 n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , 
 n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , 
 n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , 
 n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , 
 n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , 
 n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , 
 n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , 
 n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , 
 n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , 
 n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , 
 n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , 
 n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , 
 n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , 
 n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , 
 n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , 
 n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , 
 n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , 
 n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , 
 n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , 
 n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , 
 n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , 
 n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , 
 n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , 
 n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , 
 n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , 
 n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , 
 n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , 
 n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , 
 n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , 
 n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , 
 n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , 
 n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , 
 n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , 
 n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , 
 n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , 
 n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , 
 n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , 
 n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , 
 n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , 
 n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , 
 n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , 
 n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , 
 n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , 
 n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , 
 n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , 
 n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , 
 n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , 
 n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , 
 n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , 
 n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , 
 n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , 
 n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , 
 n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , 
 n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , 
 n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , 
 n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , 
 n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , 
 n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , 
 n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , 
 n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , 
 n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , 
 n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , 
 n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , 
 n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , 
 n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , 
 n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , 
 n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , 
 n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , 
 n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , 
 n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , 
 n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , 
 n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , 
 n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , 
 n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , 
 n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , 
 n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , 
 n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , 
 n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , 
 n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , 
 n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , 
 n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , 
 n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , 
 n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , 
 n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , 
 n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , 
 n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , 
 n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , 
 n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , 
 n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , 
 n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , 
 n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , 
 n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , 
 n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , 
 n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , 
 n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , 
 n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , 
 n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , 
 n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , 
 n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , 
 n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , 
 n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , 
 n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , 
 n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , 
 n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , 
 n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , 
 n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , 
 n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , 
 n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , 
 n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , 
 n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , 
 n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , 
 n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , 
 n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , 
 n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , 
 n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , 
 n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , 
 n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , 
 n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , 
 n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , 
 n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , 
 n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , 
 n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , 
 n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , 
 n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , 
 n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , 
 n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , 
 n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , 
 n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , 
 n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , 
 n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , 
 n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , 
 n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , 
 n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , 
 n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , 
 n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , 
 n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , 
 n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , 
 n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , 
 n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , 
 n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , 
 n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , 
 n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , 
 n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , 
 n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , 
 n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , 
 n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , 
 n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , 
 n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , 
 n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , 
 n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , 
 n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , 
 n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , 
 n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , 
 n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , 
 n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , 
 n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , 
 n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , 
 n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , 
 n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , 
 n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , 
 n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , 
 n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , 
 n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , 
 n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , 
 n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , 
 n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , 
 n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , 
 n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , 
 n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , 
 n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , 
 n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , 
 n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , 
 n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , 
 n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , 
 n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , 
 n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , 
 n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , 
 n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , 
 n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , 
 n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , 
 n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , 
 n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , 
 n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , 
 n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , 
 n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , 
 n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , 
 n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , 
 n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , 
 n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , 
 n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , 
 n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , 
 n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , 
 n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , 
 n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , 
 n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , 
 n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , 
 n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , 
 n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , 
 n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , 
 n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , 
 n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , 
 n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , 
 n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , 
 n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , 
 n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , 
 n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , 
 n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , 
 n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , 
 n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , 
 n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , 
 n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , 
 n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , 
 n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , 
 n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , 
 n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , 
 n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , 
 n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , 
 n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , 
 n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , 
 n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , 
 n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , 
 n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , 
 n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , 
 n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , 
 n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , 
 n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , 
 n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , 
 n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , 
 n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , 
 n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , 
 n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , 
 n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , 
 n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , 
 n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , 
 n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , 
 n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , 
 n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , 
 n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , 
 n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , 
 n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , 
 n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , 
 n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , 
 n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , 
 n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , 
 n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , 
 n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , 
 n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , 
 n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , 
 n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , 
 n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , 
 n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , 
 n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , 
 n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , 
 n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , 
 n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , 
 n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , 
 n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , 
 n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , 
 n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , 
 n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , 
 n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , 
 n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , 
 n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , 
 n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , 
 n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , 
 n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , 
 n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , 
 n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , 
 n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , 
 n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , 
 n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , 
 n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , 
 n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , 
 n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , 
 n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , 
 n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , 
 n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , 
 n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , 
 n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , 
 n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , 
 n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , 
 n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , 
 n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , 
 n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , 
 n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , 
 n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , 
 n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , 
 n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , 
 n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , 
 n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , 
 n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , 
 n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , 
 n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , 
 n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , 
 n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , 
 n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , 
 n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , 
 n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , 
 n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , 
 n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , 
 n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , 
 n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , 
 n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , 
 n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , 
 n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , 
 n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , 
 n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , 
 n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , 
 n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , 
 n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , 
 n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , 
 n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , 
 n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , 
 n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , 
 n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , 
 n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , 
 n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , 
 n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , 
 n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , 
 n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , 
 n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , 
 n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , 
 n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , 
 n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , 
 n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , 
 n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , 
 n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , 
 n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , 
 n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , 
 n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , 
 n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , 
 n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , 
 n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , 
 n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , 
 n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , 
 n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , 
 n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , 
 n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , 
 n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , 
 n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , 
 n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , 
 n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , 
 n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , 
 n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , 
 n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , 
 n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , 
 n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , 
 n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , 
 n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , 
 n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , 
 n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , 
 n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , 
 n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , 
 n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , 
 n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , 
 n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , 
 n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , 
 n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , 
 n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , 
 n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , 
 n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , 
 n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , 
 n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , 
 n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , 
 n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , 
 n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , 
 n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , 
 n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , 
 n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , 
 n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , 
 n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , 
 n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , 
 n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , 
 n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , 
 n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , 
 n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , 
 n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , 
 n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , 
 n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , 
 n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , 
 n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , 
 n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , 
 n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , 
 n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , 
 n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , 
 n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , 
 n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , 
 n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , 
 n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , 
 n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , 
 n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , 
 n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , 
 n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , 
 n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , 
 n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , 
 n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , 
 n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , 
 n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , 
 n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , 
 n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , 
 n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , 
 n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , 
 n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , 
 n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , 
 n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , 
 n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , 
 n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , 
 n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , 
 n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , 
 n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , 
 n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , 
 n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , 
 n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , 
 n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , 
 n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , 
 n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , 
 n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , 
 n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , 
 n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , 
 n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , 
 n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , 
 n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , 
 n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , 
 n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , 
 n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , 
 n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , 
 n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , 
 n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , 
 n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , 
 n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , 
 n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , 
 n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , 
 n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , 
 n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , 
 n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , 
 n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , 
 n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , 
 n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , 
 n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , 
 n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , 
 n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , 
 n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , 
 n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , 
 n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , 
 n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , 
 n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , 
 n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , 
 n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , 
 n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , 
 n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , 
 n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , 
 n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , 
 n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , 
 n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , 
 n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , 
 n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , 
 n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , 
 n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , 
 n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , 
 n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , 
 n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , 
 n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , 
 n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , 
 n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , 
 n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , 
 n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , 
 n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , 
 n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , 
 n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , 
 n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , 
 n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , 
 n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , 
 n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , 
 n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , 
 n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , 
 n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , 
 n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , 
 n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , 
 n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , 
 n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , 
 n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , 
 n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , 
 n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , 
 n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , 
 n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , 
 n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , 
 n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , 
 n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , 
 n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , 
 n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , 
 n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , 
 n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , 
 n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , 
 n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , 
 n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , 
 n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , 
 n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , 
 n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , 
 n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , 
 n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , 
 n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , 
 n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , 
 n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , 
 n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , 
 n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , 
 n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , 
 n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , 
 n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , 
 n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , 
 n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , 
 n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , 
 n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , 
 n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , 
 n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , 
 n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , 
 n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , 
 n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , 
 n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , 
 n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , 
 n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , 
 n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , 
 n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , 
 n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , 
 n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , 
 n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , 
 n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , 
 n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , 
 n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , 
 n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , 
 n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , 
 n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , 
 n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , 
 n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , 
 n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , 
 n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , 
 n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , 
 n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , 
 n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , 
 n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , 
 n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , 
 n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , 
 n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , 
 n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , 
 n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , 
 n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , 
 n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , 
 n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , 
 n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , 
 n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , 
 n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , 
 n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , 
 n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , 
 n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , 
 n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , 
 n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , 
 n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , 
 n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , 
 n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , 
 n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , 
 n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , 
 n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , 
 n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , 
 n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , 
 n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , 
 n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , 
 n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , 
 n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , 
 n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , 
 n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , 
 n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , 
 n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , 
 n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , 
 n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , 
 n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , 
 n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , 
 n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , 
 n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , 
 n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , 
 n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , 
 n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , 
 n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , 
 n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , 
 n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , 
 n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , 
 n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , 
 n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , 
 n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , 
 n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , 
 n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , 
 n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , 
 n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , 
 n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , 
 n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , 
 n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , 
 n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , 
 n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , 
 n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , 
 n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , 
 n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , 
 n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , 
 n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , 
 n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , 
 n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , 
 n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , 
 n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , 
 n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , 
 n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , 
 n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , 
 n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , 
 n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , 
 n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , 
 n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , 
 n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , 
 n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , 
 n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , 
 n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , 
 n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , 
 n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , 
 n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , 
 n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , 
 n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , 
 n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , 
 n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , 
 n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , 
 n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , 
 n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , 
 n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , 
 n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , 
 n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , 
 n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , 
 n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , 
 n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , 
 n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , 
 n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , 
 n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , 
 n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , 
 n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , 
 n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , 
 n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , 
 n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , 
 n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , 
 n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , 
 n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , 
 n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , 
 n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , 
 n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , 
 n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , 
 n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , 
 n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , 
 n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , 
 n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , 
 n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , 
 n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , 
 n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , 
 n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , 
 n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , 
 n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , 
 n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , 
 n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , 
 n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , 
 n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , 
 n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , 
 n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , 
 n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , 
 n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , 
 n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , 
 n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , 
 n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , 
 n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , 
 n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , 
 n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , 
 n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , 
 n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , 
 n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , 
 n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , 
 n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , 
 n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , 
 n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , 
 n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , 
 n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , 
 n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , 
 n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , 
 n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , 
 n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , 
 n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , 
 n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , 
 n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , 
 n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , 
 n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , 
 n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , 
 n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , 
 n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , 
 n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , 
 n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , 
 n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , 
 n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , 
 n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , 
 n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , 
 n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , 
 n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , 
 n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , 
 n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , 
 n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , 
 n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , 
 n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , 
 n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , 
 n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , 
 n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , 
 n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , 
 n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , 
 n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , 
 n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , 
 n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , 
 n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , 
 n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , 
 n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , 
 n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , 
 n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , 
 n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , 
 n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , 
 n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , 
 n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , 
 n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , 
 n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , 
 n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , 
 n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , 
 n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , 
 n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , 
 n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , 
 n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , 
 n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , 
 n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , 
 n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , 
 n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , 
 n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , 
 n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , 
 n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , 
 n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , 
 n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , 
 n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , 
 n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , 
 n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , 
 n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , 
 n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , 
 n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , 
 n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , 
 n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , 
 n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , 
 n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , 
 n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , 
 n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , 
 n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , 
 n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , 
 n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , 
 n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , 
 n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , 
 n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , 
 n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , 
 n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , 
 n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , 
 n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , 
 n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , 
 n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , 
 n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , 
 n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , 
 n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , 
 n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , 
 n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , 
 n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , 
 n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , 
 n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , 
 n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , 
 n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , 
 n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , 
 n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , 
 n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , 
 n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , 
 n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , 
 n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , 
 n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , 
 n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , 
 n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , 
 n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , 
 n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , 
 n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , 
 n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , 
 n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , 
 n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , 
 n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , 
 n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , 
 n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , 
 n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , 
 n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , 
 n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , 
 n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , 
 n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , 
 n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , 
 n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , 
 n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , 
 n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , 
 n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , 
 n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , 
 n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , 
 n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , 
 n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , 
 n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , 
 n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , 
 n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , 
 n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , 
 n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , 
 n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , 
 n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , 
 n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , 
 n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , 
 n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , 
 n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , 
 n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , 
 n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , 
 n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , 
 n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , 
 n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , 
 n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , 
 n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , 
 n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , 
 n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , 
 n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , 
 n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , 
 n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , 
 n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , 
 n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , 
 n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , 
 n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , 
 n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , 
 n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , 
 n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , 
 n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , 
 n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , 
 n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , 
 n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , 
 n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , 
 n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , 
 n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , 
 n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , 
 n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , 
 n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , 
 n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , 
 n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , 
 n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , 
 n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , 
 n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , 
 n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , 
 n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , 
 n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , 
 n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , 
 n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , 
 n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , 
 n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , 
 n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , 
 n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , 
 n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , 
 n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , 
 n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , 
 n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , 
 n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , 
 n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , 
 n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , 
 n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , 
 n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , 
 n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , 
 n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , 
 n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , 
 n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , 
 n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , 
 n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , 
 n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , 
 n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , 
 n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , 
 n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , 
 n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , 
 n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , 
 n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , 
 n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , 
 n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , 
 n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , 
 n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , 
 n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , 
 n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , 
 n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , 
 n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , 
 n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , 
 n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , 
 n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , 
 n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , 
 n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , 
 n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , 
 n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , 
 n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , 
 n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , 
 n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , 
 n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , 
 n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , 
 n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , 
 n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , 
 n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , 
 n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , 
 n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , 
 n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , 
 n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , 
 n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , 
 n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , 
 n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , 
 n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , 
 n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , 
 n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , 
 n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , 
 n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , 
 n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , 
 n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , 
 n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , 
 n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , 
 n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , 
 n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , 
 n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , 
 n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , 
 n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , 
 n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , 
 n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , 
 n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , 
 n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , 
 n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , 
 n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , 
 n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , 
 n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , 
 n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , 
 n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , 
 n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , 
 n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , 
 n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , 
 n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , 
 n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , 
 n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , 
 n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , 
 n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , 
 n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , 
 n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , 
 n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , 
 n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , 
 n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , 
 n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , 
 n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , 
 n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , 
 n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , 
 n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , 
 n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , 
 n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , 
 n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , 
 n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , 
 n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , 
 n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , 
 n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , 
 n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , 
 n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , 
 n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , 
 n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , 
 n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , 
 n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , 
 n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , 
 n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , 
 n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , 
 n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , 
 n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , 
 n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , 
 n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , 
 n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , 
 n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , 
 n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , 
 n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , 
 n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , 
 n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , 
 n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , 
 n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , 
 n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , 
 n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , 
 n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , 
 n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , 
 n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , 
 n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , 
 n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , 
 n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , 
 n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , 
 n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , 
 n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , 
 n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , 
 n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , 
 n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , 
 n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , 
 n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , 
 n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , 
 n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , 
 n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , 
 n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , 
 n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , 
 n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , 
 n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , 
 n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , 
 n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , 
 n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , 
 n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , 
 n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , 
 n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , 
 n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , 
 n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , 
 n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , 
 n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , 
 n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , 
 n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , 
 n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , 
 n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , 
 n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , 
 n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , 
 n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , 
 n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , 
 n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , 
 n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , 
 n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , 
 n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , 
 n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , 
 n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , 
 n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , 
 n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , 
 n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , 
 n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , 
 n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , 
 n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , 
 n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , 
 n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , 
 n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , 
 n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , 
 n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , 
 n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , 
 n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , 
 n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , 
 n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , 
 n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , 
 n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , 
 n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , 
 n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , 
 n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , 
 n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , 
 n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , 
 n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , 
 n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , 
 n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , 
 n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , 
 n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , 
 n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , 
 n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , 
 n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , 
 n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , 
 n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , 
 n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , 
 n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , 
 n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , 
 n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , 
 n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , 
 n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , 
 n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , 
 n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , 
 n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , 
 n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , 
 n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , 
 n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , 
 n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , 
 n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , 
 n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , 
 n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , 
 n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , 
 n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , 
 n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , 
 n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , 
 n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , 
 n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , 
 n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , 
 n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , 
 n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , 
 n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , 
 n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , 
 n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , 
 n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , 
 n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , 
 n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , 
 n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , 
 n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , 
 n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , 
 n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , 
 n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , 
 n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , 
 n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , 
 n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , 
 n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , 
 n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , 
 n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , 
 n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , 
 n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , 
 n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , 
 n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , 
 n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , 
 n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , 
 n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , 
 n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , 
 n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , 
 n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , 
 n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , 
 n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , 
 n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , 
 n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , 
 n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , 
 n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , 
 n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , 
 n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , 
 n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , 
 n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , 
 n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , 
 n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , 
 n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , 
 n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , 
 n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , 
 n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , 
 n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , 
 n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , 
 n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , 
 n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , 
 n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , 
 n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , 
 n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , 
 n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , 
 n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , 
 n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , 
 n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , 
 n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , 
 n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , 
 n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , 
 n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , 
 n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , 
 n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , 
 n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , 
 n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , 
 n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , 
 n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , 
 n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , 
 n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , 
 n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , 
 n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , 
 n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , 
 n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , 
 n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , 
 n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , 
 n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , 
 n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , 
 n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , 
 n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , 
 n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , 
 n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , 
 n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , 
 n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , 
 n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , 
 n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , 
 n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , 
 n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , 
 n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , 
 n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , 
 n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , 
 n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , 
 n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , 
 n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , 
 n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , 
 n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , 
 n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , 
 n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , 
 n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , 
 n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , 
 n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , 
 n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , 
 n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , 
 n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , 
 n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , 
 n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , 
 n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , 
 n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , 
 n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , 
 n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , 
 n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , 
 n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , 
 n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , 
 n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , 
 n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , 
 n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , 
 n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , 
 n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , 
 n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , 
 n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , 
 n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , 
 n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , 
 n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , 
 n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , 
 n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , 
 n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , 
 n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , 
 n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , 
 n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , 
 n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , 
 n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , 
 n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , 
 n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , 
 n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , 
 n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , 
 n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , 
 n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , 
 n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , 
 n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , 
 n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , 
 n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , 
 n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , 
 n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , 
 n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , 
 n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , 
 n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , 
 n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , 
 n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , 
 n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , 
 n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , 
 n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , 
 n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , 
 n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , 
 n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , 
 n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , 
 n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , 
 n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , 
 n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , 
 n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , 
 n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , 
 n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
 n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
 n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
 n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
 n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
 n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
 n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
 n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
 n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , 
 n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , 
 n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , 
 n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , 
 n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , 
 n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , 
 n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , 
 n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , 
 n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , 
 n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , 
 n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , 
 n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
 n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , 
 n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , 
 n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , 
 n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , 
 n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , 
 n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , 
 n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , 
 n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , 
 n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , 
 n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , 
 n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , 
 n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , 
 n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , 
 n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , 
 n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , 
 n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , 
 n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , 
 n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , 
 n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , 
 n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , 
 n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , 
 n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , 
 n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , 
 n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , 
 n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , 
 n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , 
 n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , 
 n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , 
 n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , 
 n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , 
 n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , 
 n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , 
 n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , 
 n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , 
 n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , 
 n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , 
 n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , 
 n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , 
 n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , 
 n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , 
 n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , 
 n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , 
 n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , 
 n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , 
 n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , 
 n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , 
 n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , 
 n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , 
 n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , 
 n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , 
 n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , 
 n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , 
 n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , 
 n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , 
 n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , 
 n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , 
 n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , 
 n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , 
 n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , 
 n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , 
 n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , 
 n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , 
 n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , 
 n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , 
 n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , 
 n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , 
 n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , 
 n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , 
 n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , 
 n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , 
 n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , 
 n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , 
 n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , 
 n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , 
 n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , 
 n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , 
 n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , 
 n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , 
 n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , 
 n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , 
 n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , 
 n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , 
 n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , 
 n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , 
 n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , 
 n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , 
 n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , 
 n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , 
 n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , 
 n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , 
 n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , 
 n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , 
 n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , 
 n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , 
 n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , 
 n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , 
 n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , 
 n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , 
 n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , 
 n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , 
 n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , 
 n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , 
 n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , 
 n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , 
 n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , 
 n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , 
 n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , 
 n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , 
 n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , 
 n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , 
 n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , 
 n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , 
 n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , 
 n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , 
 n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , 
 n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , 
 n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , 
 n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , 
 n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , 
 n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , 
 n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , 
 n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , 
 n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , 
 n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , 
 n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , 
 n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , 
 n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , 
 n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , 
 n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , 
 n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , 
 n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , 
 n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , 
 n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , 
 n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , 
 n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , 
 n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , 
 n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , 
 n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , 
 n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , 
 n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , 
 n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , 
 n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , 
 n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , 
 n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , 
 n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , 
 n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , 
 n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , 
 n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , 
 n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , 
 n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , 
 n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , 
 n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , 
 n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , 
 n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , 
 n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , 
 n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , 
 n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , 
 n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , 
 n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , 
 n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , 
 n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , 
 n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , 
 n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , 
 n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , 
 n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , 
 n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , 
 n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , 
 n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , 
 n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , 
 n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , 
 n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , 
 n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , 
 n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , 
 n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , 
 n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , 
 n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , 
 n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , 
 n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , 
 n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , 
 n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , 
 n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , 
 n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , 
 n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , 
 n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , 
 n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , 
 n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , 
 n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , 
 n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , 
 n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , 
 n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , 
 n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , 
 n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , 
 n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , 
 n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , 
 n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , 
 n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , 
 n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , 
 n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , 
 n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , 
 n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , 
 n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , 
 n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , 
 n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , 
 n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , 
 n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , 
 n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , 
 n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , 
 n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , 
 n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , 
 n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , 
 n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , 
 n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , 
 n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , 
 n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , 
 n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , 
 n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , 
 n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , 
 n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , 
 n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , 
 n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , 
 n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , 
 n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , 
 n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , 
 n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , 
 n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , 
 n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , 
 n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , 
 n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , 
 n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , 
 n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , 
 n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , 
 n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , 
 n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , 
 n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , 
 n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , 
 n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , 
 n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , 
 n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , 
 n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , 
 n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , 
 n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , 
 n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , 
 n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , 
 n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , 
 n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , 
 n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , 
 n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , 
 n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , 
 n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , 
 n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , 
 n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , 
 n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , 
 n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , 
 n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , 
 n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , 
 n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , 
 n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , 
 n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , 
 n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , 
 n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , 
 n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , 
 n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , 
 n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , 
 n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , 
 n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , 
 n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , 
 n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , 
 n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , 
 n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , 
 n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , 
 n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , 
 n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , 
 n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , 
 n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , 
 n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , 
 n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , 
 n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , 
 n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , 
 n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , 
 n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , 
 n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , 
 n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , 
 n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , 
 n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , 
 n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , 
 n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , 
 n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , 
 n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , 
 n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , 
 n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , 
 n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , 
 n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , 
 n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , 
 n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , 
 n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , 
 n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , 
 n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , 
 n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , 
 n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , 
 n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , 
 n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , 
 n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
 n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , 
 n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , 
 n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , 
 n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , 
 n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , 
 n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , 
 n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , 
 n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , 
 n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , 
 n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , 
 n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , 
 n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , 
 n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , 
 n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , 
 n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , 
 n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , 
 n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , 
 n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , 
 n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , 
 n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , 
 n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , 
 n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , 
 n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , 
 n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , 
 n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , 
 n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , 
 n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , 
 n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , 
 n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , 
 n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , 
 n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , 
 n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , 
 n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , 
 n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , 
 n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , 
 n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , 
 n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , 
 n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , 
 n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , 
 n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , 
 n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , 
 n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , 
 n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , 
 n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , 
 n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , 
 n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , 
 n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , 
 n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , 
 n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , 
 n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , 
 n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , 
 n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , 
 n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , 
 n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , 
 n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , 
 n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , 
 n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , 
 n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , 
 n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , 
 n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , 
 n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , 
 n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , 
 n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , 
 n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , 
 n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , 
 n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , 
 n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , 
 n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , 
 n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , 
 n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , 
 n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , 
 n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , 
 n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , 
 n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , 
 n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , 
 n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , 
 n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , 
 n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , 
 n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , 
 n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , 
 n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , 
 n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , 
 n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , 
 n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , 
 n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , 
 n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , 
 n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , 
 n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , 
 n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , 
 n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , 
 n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , 
 n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , 
 n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , 
 n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , 
 n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , 
 n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , 
 n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , 
 n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , 
 n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , 
 n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , 
 n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , 
 n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , 
 n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , 
 n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , 
 n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , 
 n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , 
 n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , 
 n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , 
 n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , 
 n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , 
 n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , 
 n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , 
 n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , 
 n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , 
 n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , 
 n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , 
 n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , 
 n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , 
 n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , 
 n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , 
 n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , 
 n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , 
 n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , 
 n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , 
 n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , 
 n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , 
 n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , 
 n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , 
 n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , 
 n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , 
 n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , 
 n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , 
 n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , 
 n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , 
 n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , 
 n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , 
 n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , 
 n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , 
 n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , 
 n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , 
 n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , 
 n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , 
 n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , 
 n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , 
 n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , 
 n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , 
 n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , 
 n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , 
 n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , 
 n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , 
 n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , 
 n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , 
 n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , 
 n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , 
 n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , 
 n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , 
 n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , 
 n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , 
 n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , 
 n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , 
 n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , 
 n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , 
 n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , 
 n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , 
 n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , 
 n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , 
 n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , 
 n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , 
 n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , 
 n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , 
 n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , 
 n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , 
 n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , 
 n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , 
 n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , 
 n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , 
 n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , 
 n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , 
 n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , 
 n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , 
 n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , 
 n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , 
 n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , 
 n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , 
 n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , 
 n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , 
 n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , 
 n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , 
 n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , 
 n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , 
 n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , 
 n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , 
 n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , 
 n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , 
 n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , 
 n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , 
 n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , 
 n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , 
 n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , 
 n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , 
 n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , 
 n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , 
 n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , 
 n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , 
 n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , 
 n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , 
 n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , 
 n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , 
 n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , 
 n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , 
 n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , 
 n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , 
 n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , 
 n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , 
 n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , 
 n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , 
 n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , 
 n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , 
 n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , 
 n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , 
 n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , 
 n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , 
 n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , 
 n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , 
 n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , 
 n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , 
 n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , 
 n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , 
 n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , 
 n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , 
 n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , 
 n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , 
 n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , 
 n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , 
 n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , 
 n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , 
 n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , 
 n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , 
 n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , 
 n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , 
 n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , 
 n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , 
 n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , 
 n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , 
 n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , 
 n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , 
 n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , 
 n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , 
 n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , 
 n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , 
 n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , 
 n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , 
 n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , 
 n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , 
 n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , 
 n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , 
 n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , 
 n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , 
 n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , 
 n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , 
 n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , 
 n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , 
 n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , 
 n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , 
 n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , 
 n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , 
 n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , 
 n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , 
 n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , 
 n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , 
 n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , 
 n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , 
 n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , 
 n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , 
 n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , 
 n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , 
 n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , 
 n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , 
 n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , 
 n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , 
 n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , 
 n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , 
 n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , 
 n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , 
 n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , 
 n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , 
 n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , 
 n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , 
 n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , 
 n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , 
 n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , 
 n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , 
 n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , 
 n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , 
 n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , 
 n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , 
 n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , 
 n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , 
 n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , 
 n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , 
 n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , 
 n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , 
 n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , 
 n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , 
 n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , 
 n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , 
 n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , 
 n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , 
 n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , 
 n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , 
 n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , 
 n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , 
 n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , 
 n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , 
 n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , 
 n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , 
 n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , 
 n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , 
 n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , 
 n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , 
 n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , 
 n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , 
 n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , 
 n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , 
 n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , 
 n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , 
 n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , 
 n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , 
 n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , 
 n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , 
 n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , 
 n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , 
 n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , 
 n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , 
 n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , 
 n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , 
 n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , 
 n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , 
 n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , 
 n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , 
 n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , 
 n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , 
 n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , 
 n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , 
 n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , 
 n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , 
 n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , 
 n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , 
 n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , 
 n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , 
 n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , 
 n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , 
 n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , 
 n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , 
 n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , 
 n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , 
 n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , 
 n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , 
 n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , 
 n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , 
 n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , 
 n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , 
 n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , 
 n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , 
 n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , 
 n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , 
 n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , 
 n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , 
 n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , 
 n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , 
 n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , 
 n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , 
 n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , 
 n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , 
 n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , 
 n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , 
 n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , 
 n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , 
 n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , 
 n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , 
 n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , 
 n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , 
 n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , 
 n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , 
 n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , 
 n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , 
 n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , 
 n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , 
 n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , 
 n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , 
 n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , 
 n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , 
 n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , 
 n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , 
 n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , 
 n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , 
 n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , 
 n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , 
 n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , 
 n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , 
 n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , 
 n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , 
 n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , 
 n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , 
 n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , 
 n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , 
 n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , 
 n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , 
 n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , 
 n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , 
 n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , 
 n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , 
 n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , 
 n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , 
 n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , 
 n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , 
 n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , 
 n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , 
 n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , 
 n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , 
 n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , 
 n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , 
 n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , 
 n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , 
 n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , 
 n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , 
 n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , 
 n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , 
 n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , 
 n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , 
 n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , 
 n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , 
 n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , 
 n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , 
 n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , 
 n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , 
 n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , 
 n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , 
 n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , 
 n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , 
 n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , 
 n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , 
 n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , 
 n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , 
 n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , 
 n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , 
 n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , 
 n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , 
 n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , 
 n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , 
 n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , 
 n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , 
 n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , 
 n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , 
 n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , 
 n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , 
 n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , 
 n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , 
 n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , 
 n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , 
 n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , 
 n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , 
 n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , 
 n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , 
 n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , 
 n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , 
 n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , 
 n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , 
 n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , 
 n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , 
 n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , 
 n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , 
 n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , 
 n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , 
 n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , 
 n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , 
 n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , 
 n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , 
 n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , 
 n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , 
 n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , 
 n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , 
 n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , 
 n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , 
 n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , 
 n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , 
 n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , 
 n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , 
 n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , 
 n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , 
 n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , 
 n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , 
 n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , 
 n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , 
 n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , 
 n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , 
 n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , 
 n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , 
 n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , 
 n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , 
 n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , 
 n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , 
 n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , 
 n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , 
 n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , 
 n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , 
 n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , 
 n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , 
 n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , 
 n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , 
 n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , 
 n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , 
 n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , 
 n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , 
 n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , 
 n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , 
 n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , 
 n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , 
 n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , 
 n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , 
 n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , 
 n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , 
 n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , 
 n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , 
 n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , 
 n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , 
 n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , 
 n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , 
 n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , 
 n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , 
 n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , 
 n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , 
 n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , 
 n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , 
 n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , 
 n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , 
 n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , 
 n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , 
 n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , 
 n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , 
 n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , 
 n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , 
 n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , 
 n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , 
 n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , 
 n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , 
 n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , 
 n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , 
 n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , 
 n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , 
 n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , 
 n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , 
 n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , 
 n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , 
 n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , 
 n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , 
 n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , 
 n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , 
 n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , 
 n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , 
 n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , 
 n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , 
 n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , 
 n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , 
 n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , 
 n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , 
 n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , 
 n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , 
 n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , 
 n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , 
 n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , 
 n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , 
 n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , 
 n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , 
 n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , 
 n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , 
 n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , 
 n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , 
 n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , 
 n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , 
 n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , 
 n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , 
 n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , 
 n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , 
 n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , 
 n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , 
 n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , 
 n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , 
 n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , 
 n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , 
 n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , 
 n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , 
 n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , 
 n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , 
 n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , 
 n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , 
 n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , 
 n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , 
 n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , 
 n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , 
 n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , 
 n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , 
 n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , 
 n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , 
 n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , 
 n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , 
 n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , 
 n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , 
 n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , 
 n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , 
 n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , 
 n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , 
 n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , 
 n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , 
 n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , 
 n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , 
 n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , 
 n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , 
 n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , 
 n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , 
 n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , 
 n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , 
 n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , 
 n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , 
 n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , 
 n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , 
 n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , 
 n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , 
 n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , 
 n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , 
 n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , 
 n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , 
 n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , 
 n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , 
 n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , 
 n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , 
 n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , 
 n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , 
 n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , 
 n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , 
 n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , 
 n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , 
 n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , 
 n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , 
 n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , 
 n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , 
 n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , 
 n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , 
 n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , 
 n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , 
 n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , 
 n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , 
 n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , 
 n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , 
 n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , 
 n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , 
 n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , 
 n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , 
 n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , 
 n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , 
 n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , 
 n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , 
 n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , 
 n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , 
 n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , 
 n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , 
 n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , 
 n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , 
 n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , 
 n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , 
 n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , 
 n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , 
 n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , 
 n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , 
 n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , 
 n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , 
 n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , 
 n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , 
 n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , 
 n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , 
 n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , 
 n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , 
 n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , 
 n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , 
 n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , 
 n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , 
 n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , 
 n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , 
 n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , 
 n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , 
 n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , 
 n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , 
 n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , 
 n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , 
 n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , 
 n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , 
 n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , 
 n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , 
 n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , 
 n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , 
 n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , 
 n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , 
 n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , 
 n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , 
 n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , 
 n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , 
 n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , 
 n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , 
 n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , 
 n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , 
 n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , 
 n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , 
 n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , 
 n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , 
 n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , 
 n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , 
 n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , 
 n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , 
 n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , 
 n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , 
 n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , 
 n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , 
 n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , 
 n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , 
 n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , 
 n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , 
 n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , 
 n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , 
 n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , 
 n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , 
 n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , 
 n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , 
 n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , 
 n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , 
 n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , 
 n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , 
 n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , 
 n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , 
 n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , 
 n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , 
 n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , 
 n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , 
 n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , 
 n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , 
 n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , 
 n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , 
 n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , 
 n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , 
 n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , 
 n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , 
 n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , 
 n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , 
 n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , 
 n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , 
 n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , 
 n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , 
 n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , 
 n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , 
 n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , 
 n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , 
 n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , 
 n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , 
 n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , 
 n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , 
 n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , 
 n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , 
 n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , 
 n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , 
 n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , 
 n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , 
 n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , 
 n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , 
 n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , 
 n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , 
 n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , 
 n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , 
 n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , 
 n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , 
 n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , 
 n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , 
 n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , 
 n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , 
 n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , 
 n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , 
 n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , 
 n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , 
 n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , 
 n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , 
 n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , 
 n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , 
 n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , 
 n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , 
 n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , 
 n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , 
 n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , 
 n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , 
 n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , 
 n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , 
 n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , 
 n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , 
 n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , 
 n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , 
 n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , 
 n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , 
 n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , 
 n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , 
 n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , 
 n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , 
 n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , 
 n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , 
 n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , 
 n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , 
 n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , 
 n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , 
 n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , 
 n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , 
 n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , 
 n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , 
 n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , 
 n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , 
 n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , 
 n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , 
 n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , 
 n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , 
 n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , 
 n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , 
 n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , 
 n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , 
 n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , 
 n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , 
 n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , 
 n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , 
 n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , 
 n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , 
 n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , 
 n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , 
 n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , 
 n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , 
 n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , 
 n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , 
 n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , 
 n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , 
 n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , 
 n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , 
 n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , 
 n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , 
 n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , 
 n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , 
 n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , 
 n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , 
 n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , 
 n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , 
 n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , 
 n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , 
 n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , 
 n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , 
 n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , 
 n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , 
 n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , 
 n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , 
 n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , 
 n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , 
 n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , 
 n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , 
 n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , 
 n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , 
 n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , 
 n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , 
 n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , 
 n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , 
 n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , 
 n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , 
 n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , 
 n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , 
 n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , 
 n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , 
 n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , 
 n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , 
 n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , 
 n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , 
 n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , 
 n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , 
 n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , 
 n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , 
 n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , 
 n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , 
 n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , 
 n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , 
 n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , 
 n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , 
 n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , 
 n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , 
 n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , 
 n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , 
 n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , 
 n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , 
 n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , 
 n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , 
 n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , 
 n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , 
 n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , 
 n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , 
 n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , 
 n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , 
 n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , 
 n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , 
 n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , 
 n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , 
 n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , 
 n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , 
 n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , 
 n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , 
 n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , 
 n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , 
 n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , 
 n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , 
 n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , 
 n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , 
 n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , 
 n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , 
 n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , 
 n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , 
 n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , 
 n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , 
 n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , 
 n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , 
 n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , 
 n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , 
 n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , 
 n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , 
 n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , 
 n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , 
 n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , 
 n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , 
 n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , 
 n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , 
 n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , 
 n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , 
 n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , 
 n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , 
 n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , 
 n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , 
 n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , 
 n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , 
 n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , 
 n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , 
 n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , 
 n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , 
 n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , 
 n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , 
 n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , 
 n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , 
 n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , 
 n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , 
 n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , 
 n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , 
 n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , 
 n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , 
 n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , 
 n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , 
 n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , 
 n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , 
 n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , 
 n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , 
 n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , 
 n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , 
 n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , 
 n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , 
 n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , 
 n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , 
 n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , 
 n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , 
 n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , 
 n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , 
 n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , 
 n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , 
 n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , 
 n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , 
 n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , 
 n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , 
 n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , 
 n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , 
 n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , 
 n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , 
 n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , 
 n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , 
 n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , 
 n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , 
 n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , 
 n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , 
 n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , 
 n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , 
 n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , 
 n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , 
 n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , 
 n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , 
 n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , 
 n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , 
 n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , 
 n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , 
 n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , 
 n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , 
 n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , 
 n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , 
 n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , 
 n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , 
 n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , 
 n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , 
 n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , 
 n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , 
 n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , 
 n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , 
 n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , 
 n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , 
 n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , 
 n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , 
 n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , 
 n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , 
 n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , 
 n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , 
 n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , 
 n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , 
 n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , 
 n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , 
 n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , 
 n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , 
 n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , 
 n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , 
 n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , 
 n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , 
 n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , 
 n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , 
 n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , 
 n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , 
 n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , 
 n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , 
 n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , 
 n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , 
 n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , 
 n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , 
 n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , 
 n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , 
 n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , 
 n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , 
 n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , 
 n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , 
 n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , 
 n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , 
 n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , 
 n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , 
 n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , 
 n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , 
 n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , 
 n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , 
 n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , 
 n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , 
 n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , 
 n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , 
 n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , 
 n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , 
 n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , 
 n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , 
 n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , 
 n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , 
 n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , 
 n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , 
 n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , 
 n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , 
 n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , 
 n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , 
 n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , 
 n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , 
 n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , 
 n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , 
 n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , 
 n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , 
 n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , 
 n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , 
 n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , 
 n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , 
 n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , 
 n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , 
 n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , 
 n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , 
 n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , 
 n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , 
 n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , 
 n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , 
 n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , 
 n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , 
 n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , 
 n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , 
 n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , 
 n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , 
 n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , 
 n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , 
 n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , 
 n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , 
 n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , 
 n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , 
 n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , 
 n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , 
 n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , 
 n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , 
 n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , 
 n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , 
 n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , 
 n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , 
 n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , 
 n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , 
 n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , 
 n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , 
 n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , 
 n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , 
 n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , 
 n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , 
 n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , 
 n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , 
 n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , 
 n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , 
 n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , 
 n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , 
 n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , 
 n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , 
 n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , 
 n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , 
 n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , 
 n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , 
 n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , 
 n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , 
 n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , 
 n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , 
 n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , 
 n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , 
 n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , 
 n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , 
 n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , 
 n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , 
 n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , 
 n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , 
 n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , 
 n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , 
 n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , 
 n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , 
 n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , 
 n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , 
 n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , 
 n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , 
 n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , 
 n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , 
 n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , 
 n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , 
 n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , 
 n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , 
 n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , 
 n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , 
 n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , 
 n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , 
 n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , 
 n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , 
 n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , 
 n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , 
 n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , 
 n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , 
 n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , 
 n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , 
 n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , 
 n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , 
 n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , 
 n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , 
 n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , 
 n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , 
 n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , 
 n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , 
 n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , 
 n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , 
 n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , 
 n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , 
 n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , 
 n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , 
 n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , 
 n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , 
 n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , 
 n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , 
 n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , 
 n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , 
 n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , 
 n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , 
 n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , 
 n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , 
 n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , 
 n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , 
 n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , 
 n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , 
 n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , 
 n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , 
 n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , 
 n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , 
 n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , 
 n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , 
 n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , 
 n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , 
 n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , 
 n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , 
 n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , 
 n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , 
 n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , 
 n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , 
 n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , 
 n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , 
 n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , 
 n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , 
 n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , 
 n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , 
 n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , 
 n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , 
 n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , 
 n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , 
 n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , 
 n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , 
 n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , 
 n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , 
 n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , 
 n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , 
 n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , 
 n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , 
 n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , 
 n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , 
 n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , 
 n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , 
 n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , 
 n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , 
 n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , 
 n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , 
 n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , 
 n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , 
 n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , 
 n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , 
 n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , 
 n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , 
 n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , 
 n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , 
 n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , 
 n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , 
 n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , 
 n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , 
 n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , 
 n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , 
 n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , 
 n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , 
 n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , 
 n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , 
 n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , 
 n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , 
 n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , 
 n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , 
 n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , 
 n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , 
 n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , 
 n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , 
 n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , 
 n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , 
 n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , 
 n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , 
 n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , 
 n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , 
 n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , 
 n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , 
 n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , 
 n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , 
 n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , 
 n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , 
 n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , 
 n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , 
 n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , 
 n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , 
 n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , 
 n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , 
 n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , 
 n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , 
 n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , 
 n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , 
 n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , 
 n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , 
 n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , 
 n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , 
 n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , 
 n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , 
 n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , 
 n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , 
 n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , 
 n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , 
 n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , 
 n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , 
 n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , 
 n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , 
 n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , 
 n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , 
 n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , 
 n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , 
 n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , 
 n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , 
 n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , 
 n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , 
 n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , 
 n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , 
 n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , 
 n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , 
 n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , 
 n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , 
 n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , 
 n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , 
 n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , 
 n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , 
 n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , 
 n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , 
 n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , 
 n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , 
 n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , 
 n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , 
 n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , 
 n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , 
 n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , 
 n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , 
 n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , 
 n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , 
 n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , 
 n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , 
 n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , 
 n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , 
 n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , 
 n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , 
 n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , 
 n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , 
 n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , 
 n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , 
 n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , 
 n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , 
 n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , 
 n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , 
 n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , 
 n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , 
 n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , 
 n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , 
 n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , 
 n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , 
 n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , 
 n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , 
 n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , 
 n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , 
 n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , 
 n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , 
 n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , 
 n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , 
 n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , 
 n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , 
 n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , 
 n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , 
 n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , 
 n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , 
 n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , 
 n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , 
 n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , 
 n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , 
 n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , 
 n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , 
 n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , 
 n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , 
 n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , 
 n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , 
 n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , 
 n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , 
 n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , 
 n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , 
 n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , 
 n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , 
 n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , 
 n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , 
 n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , 
 n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , 
 n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , 
 n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , 
 n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , 
 n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , 
 n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , 
 n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , 
 n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , 
 n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , 
 n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , 
 n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , 
 n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , 
 n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , 
 n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , 
 n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , 
 n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , 
 n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , 
 n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , 
 n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , 
 n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , 
 n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , 
 n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , 
 n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , 
 n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , 
 n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , 
 n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , 
 n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , 
 n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , 
 n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , 
 n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , 
 n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , 
 n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , 
 n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , 
 n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , 
 n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , 
 n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , 
 n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , 
 n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , 
 n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , 
 n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , 
 n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , 
 n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , 
 n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , 
 n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , 
 n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , 
 n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , 
 n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , 
 n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , 
 n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , 
 n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , 
 n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , 
 n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , 
 n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , 
 n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , 
 n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , 
 n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , 
 n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , 
 n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , 
 n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , 
 n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , 
 n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , 
 n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , 
 n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , 
 n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , 
 n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , 
 n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , 
 n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , 
 n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , 
 n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , 
 n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , 
 n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , 
 n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , 
 n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , 
 n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , 
 n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , 
 n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , 
 n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , 
 n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , 
 n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , 
 n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , 
 n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , 
 n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , 
 n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , 
 n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , 
 n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , 
 n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , 
 n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , 
 n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , 
 n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , 
 n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , 
 n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , 
 n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , 
 n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , 
 n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , 
 n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , 
 n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , 
 n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , 
 n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , 
 n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , 
 n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , 
 n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , 
 n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , 
 n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , 
 n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , 
 n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , 
 n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , 
 n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , 
 n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , 
 n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , 
 n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , 
 n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , 
 n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , 
 n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , 
 n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , 
 n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , 
 n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , 
 n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , 
 n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , 
 n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , 
 n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , 
 n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , 
 n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , 
 n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , 
 n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , 
 n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , 
 n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , 
 n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , 
 n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , 
 n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , 
 n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , 
 n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , 
 n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , 
 n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , 
 n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , 
 n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , 
 n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , 
 n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , 
 n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , 
 n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , 
 n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , 
 n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , 
 n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , 
 n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , 
 n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , 
 n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , 
 n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , 
 n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , 
 n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , 
 n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , 
 n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , 
 n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , 
 n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , 
 n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , 
 n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , 
 n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , 
 n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , 
 n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , 
 n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , 
 n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , 
 n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , 
 n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , 
 n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , 
 n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , 
 n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , 
 n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , 
 n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , 
 n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , 
 n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , 
 n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , 
 n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , 
 n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , 
 n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , 
 n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , 
 n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , 
 n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , 
 n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , 
 n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , 
 n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , 
 n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , 
 n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , 
 n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , 
 n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , 
 n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , 
 n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , 
 n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , 
 n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , 
 n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , 
 n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , 
 n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , 
 n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , 
 n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , 
 n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , 
 n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , 
 n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , 
 n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , 
 n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , 
 n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , 
 n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , 
 n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , 
 n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , 
 n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , 
 n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , 
 n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , 
 n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , 
 n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , 
 n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , 
 n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , 
 n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , 
 n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , 
 n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , 
 n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , 
 n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , 
 n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , 
 n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , 
 n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , 
 n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , 
 n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , 
 n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , 
 n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , 
 n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , 
 n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , 
 n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , 
 n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , 
 n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , 
 n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , 
 n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , 
 n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , 
 n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , 
 n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , 
 n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , 
 n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , 
 n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , 
 n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , 
 n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , 
 n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , 
 n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , 
 n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , 
 n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , 
 n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , 
 n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , 
 n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , 
 n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , 
 n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , 
 n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , 
 n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , 
 n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , 
 n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , 
 n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , 
 n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , 
 n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , 
 n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , 
 n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , 
 n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , 
 n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , 
 n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , 
 n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , 
 n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , 
 n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , 
 n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , 
 n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , 
 n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , 
 n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , 
 n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , 
 n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , 
 n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , 
 n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , 
 n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , 
 n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , 
 n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , 
 n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , 
 n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , 
 n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , 
 n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , 
 n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , 
 n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , 
 n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , 
 n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , 
 n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , 
 n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , 
 n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , 
 n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , 
 n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , 
 n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , 
 n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , 
 n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , 
 n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , 
 n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , 
 n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , 
 n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , 
 n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , 
 n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , 
 n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , 
 n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , 
 n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , 
 n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , 
 n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , 
 n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , 
 n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , 
 n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , 
 n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , 
 n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , 
 n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , 
 n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , 
 n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , 
 n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , 
 n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , 
 n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , 
 n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , 
 n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , 
 n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , 
 n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , 
 n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , 
 n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , 
 n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , 
 n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , 
 n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , 
 n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , 
 n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , 
 n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , 
 n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , 
 n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , 
 n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , 
 n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , 
 n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , 
 n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , 
 n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , 
 n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , 
 n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , 
 n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , 
 n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , 
 n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , 
 n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , 
 n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , 
 n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , 
 n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , 
 n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , 
 n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , 
 n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , 
 n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , 
 n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , 
 n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , 
 n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , 
 n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , 
 n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , 
 n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , 
 n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , 
 n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , 
 n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , 
 n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , 
 n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , 
 n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , 
 n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , 
 n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , 
 n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , 
 n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , 
 n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , 
 n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , 
 n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , 
 n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , 
 n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , 
 n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , 
 n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , 
 n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , 
 n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , 
 n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , 
 n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , 
 n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , 
 n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , 
 n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , 
 n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , 
 n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , 
 n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , 
 n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , 
 n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , 
 n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , 
 n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , 
 n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , 
 n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , 
 n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , 
 n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , 
 n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , 
 n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , 
 n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , 
 n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , 
 n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , 
 n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , 
 n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , 
 n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , 
 n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , 
 n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , 
 n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , 
 n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , 
 n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , 
 n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , 
 n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , 
 n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , 
 n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , 
 n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , 
 n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , 
 n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , 
 n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , 
 n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , 
 n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , 
 n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , 
 n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , 
 n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , 
 n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , 
 n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , 
 n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , 
 n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , 
 n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , 
 n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , 
 n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , 
 n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , 
 n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , 
 n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , 
 n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , 
 n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , 
 n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , 
 n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , 
 n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , 
 n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , 
 n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , 
 n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , 
 n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , 
 n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , 
 n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , 
 n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , 
 n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , 
 n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , 
 n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , 
 n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , 
 n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , 
 n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , 
 n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , 
 n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , 
 n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , 
 n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , 
 n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , 
 n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , 
 n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , 
 n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , 
 n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , 
 n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , 
 n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , 
 n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , 
 n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , 
 n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , 
 n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , 
 n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , 
 n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , 
 n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , 
 n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , 
 n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , 
 n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , 
 n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , 
 n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , 
 n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , 
 n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , 
 n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , 
 n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , 
 n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , 
 n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , 
 n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , 
 n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , 
 n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , 
 n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , 
 n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , 
 n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , 
 n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , 
 n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , 
 n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , 
 n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , 
 n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , 
 n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , 
 n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , 
 n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , 
 n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , 
 n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , 
 n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , 
 n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , 
 n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , 
 n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , 
 n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , 
 n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , 
 n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , 
 n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , 
 n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , 
 n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , 
 n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , 
 n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , 
 n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , 
 n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , 
 n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , 
 n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , 
 n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , 
 n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , 
 n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , 
 n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , 
 n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , 
 n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , 
 n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , 
 n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , 
 n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , 
 n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , 
 n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , 
 n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , 
 n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , 
 n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , 
 n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , 
 n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , 
 n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , 
 n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , 
 n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , 
 n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , 
 n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , 
 n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , 
 n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , 
 n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , 
 n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , 
 n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , 
 n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , 
 n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , 
 n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , 
 n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , 
 n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , 
 n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , 
 n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , 
 n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , 
 n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , 
 n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , 
 n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , 
 n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , 
 n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , 
 n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , 
 n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , 
 n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , 
 n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , 
 n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , 
 n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , 
 n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , 
 n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , 
 n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , 
 n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , 
 n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , 
 n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , 
 n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , 
 n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , 
 n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , 
 n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , 
 n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , 
 n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , 
 n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , 
 n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , 
 n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , 
 n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , 
 n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , 
 n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , 
 n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , 
 n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , 
 n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , 
 n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , 
 n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , 
 n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , 
 n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , 
 n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , 
 n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , 
 n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , 
 n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , 
 n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , 
 n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , 
 n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , 
 n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , 
 n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , 
 n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , 
 n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , 
 n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , 
 n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , 
 n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , 
 n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , 
 n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , 
 n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , 
 n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , 
 n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , 
 n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , 
 n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , 
 n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , 
 n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , 
 n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , 
 n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , 
 n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , 
 n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , 
 n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , 
 n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , 
 n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , 
 n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , 
 n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , 
 n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , 
 n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , 
 n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , 
 n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , 
 n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , 
 n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , 
 n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , 
 n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , 
 n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , 
 n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , 
 n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , 
 n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , 
 n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , 
 n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , 
 n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , 
 n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , 
 n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , 
 n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , 
 n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , 
 n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , 
 n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , 
 n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , 
 n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , 
 n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , 
 n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , 
 n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , 
 n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , 
 n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , 
 n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , 
 n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , 
 n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , 
 n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , 
 n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , 
 n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , 
 n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , 
 n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , 
 n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , 
 n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , 
 n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , 
 n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , 
 n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , 
 n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , 
 n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , 
 n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , 
 n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , 
 n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , 
 n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , 
 n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , 
 n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , 
 n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , 
 n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , 
 n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , 
 n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , 
 n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , 
 n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , 
 n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , 
 n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , 
 n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , 
 n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , 
 n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , 
 n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , 
 n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , 
 n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , 
 n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , 
 n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , 
 n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , 
 n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , 
 n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , 
 n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , 
 n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , 
 n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , 
 n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , 
 n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , 
 n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , 
 n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , 
 n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , 
 n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , 
 n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , 
 n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , 
 n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , 
 n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , 
 n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , 
 n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , 
 n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , 
 n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , 
 n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , 
 n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , 
 n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , 
 n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , 
 n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , 
 n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , 
 n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , 
 n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , 
 n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , 
 n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , 
 n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , 
 n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , 
 n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , 
 n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , 
 n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , 
 n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , 
 n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , 
 n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , 
 n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , 
 n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , 
 n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , 
 n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , 
 n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , 
 n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , 
 n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , 
 n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , 
 n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , 
 n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , 
 n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , 
 n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , 
 n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , 
 n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , 
 n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , 
 n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , 
 n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , 
 n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , 
 n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , 
 n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , 
 n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , 
 n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , 
 n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , 
 n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , 
 n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , 
 n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , 
 n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , 
 n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , 
 n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , 
 n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , 
 n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , 
 n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , 
 n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , 
 n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , 
 n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , 
 n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , 
 n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , 
 n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , 
 n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , 
 n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , 
 n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , 
 n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , 
 n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , 
 n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , 
 n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , 
 n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , 
 n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , 
 n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , 
 n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , 
 n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , 
 n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , 
 n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , 
 n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , 
 n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , 
 n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , 
 n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , 
 n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , 
 n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , 
 n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , 
 n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , 
 n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , 
 n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , 
 n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , 
 n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , 
 n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , 
 n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , 
 n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , 
 n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , 
 n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , 
 n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , 
 n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , 
 n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , 
 n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , 
 n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , 
 n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , 
 n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , 
 n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , 
 n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , 
 n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , 
 n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , 
 n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , 
 n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , 
 n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , 
 n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , 
 n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , 
 n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , 
 n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , 
 n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , 
 n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , 
 n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , 
 n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , 
 n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , 
 n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , 
 n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , 
 n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , 
 n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , 
 n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , 
 n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , 
 n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , 
 n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , 
 n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , 
 n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , 
 n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , 
 n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , 
 n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , 
 n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , 
 n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , 
 n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , 
 n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , 
 n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , 
 n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , 
 n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , 
 n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , 
 n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , 
 n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , 
 n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , 
 n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , 
 n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , 
 n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , 
 n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , 
 n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , 
 n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , 
 n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , 
 n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , 
 n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , 
 n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , 
 n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , 
 n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , 
 n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , 
 n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , 
 n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , 
 n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , 
 n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , 
 n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , 
 n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , 
 n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , 
 n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , 
 n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , 
 n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , 
 n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , 
 n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , 
 n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , 
 n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , 
 n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , 
 n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , 
 n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , 
 n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , 
 n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , 
 n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , 
 n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , 
 n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , 
 n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , 
 n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , 
 n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , 
 n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , 
 n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , 
 n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , 
 n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , 
 n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , 
 n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , 
 n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , 
 n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , 
 n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , 
 n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , 
 n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , 
 n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , 
 n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , 
 n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , 
 n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , 
 n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , 
 n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , 
 n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , 
 n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , 
 n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , 
 n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , 
 n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , 
 n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , 
 n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , 
 n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , 
 n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , 
 n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , 
 n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , 
 n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , 
 n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , 
 n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , 
 n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , 
 n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , 
 n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , 
 n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , 
 n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , 
 n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , 
 n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , 
 n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , 
 n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , 
 n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , 
 n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , 
 n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , 
 n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , 
 n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , 
 n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , 
 n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , 
 n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , 
 n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , 
 n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , 
 n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , 
 n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , 
 n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , 
 n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , 
 n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , 
 n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , 
 n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , 
 n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , 
 n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , 
 n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , 
 n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , 
 n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , 
 n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , 
 n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , 
 n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , 
 n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , 
 n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , 
 n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , 
 n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , 
 n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , 
 n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , 
 n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , 
 n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , 
 n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , 
 n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , 
 n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , 
 n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , 
 n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , 
 n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , 
 n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , 
 n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , 
 n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , 
 n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , 
 n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , 
 n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , 
 n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , 
 n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , 
 n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , 
 n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , 
 n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , 
 n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , 
 n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , 
 n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , 
 n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , 
 n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , 
 n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , 
 n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , 
 n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , 
 n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , 
 n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , 
 n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , 
 n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , 
 n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , 
 n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , 
 n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , 
 n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , 
 n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , 
 n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , 
 n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , 
 n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , 
 n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , 
 n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , 
 n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , 
 n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , 
 n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , 
 n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , 
 n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , 
 n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , 
 n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , 
 n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , 
 n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , 
 n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , 
 n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , 
 n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , 
 n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , 
 n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , 
 n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , 
 n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , 
 n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , 
 n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , 
 n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , 
 n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , 
 n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , 
 n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , 
 n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , 
 n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , 
 n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , 
 n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , 
 n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , 
 n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , 
 n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , 
 n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , 
 n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , 
 n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , 
 n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , 
 n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , 
 n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , 
 n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , 
 n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , 
 n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , 
 n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , 
 n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , 
 n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , 
 n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , 
 n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , 
 n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , 
 n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , 
 n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , 
 n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , 
 n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , 
 n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , 
 n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , 
 n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , 
 n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , 
 n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , 
 n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , 
 n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , 
 n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , 
 n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , 
 n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , 
 n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , 
 n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , 
 n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , 
 n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , 
 n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , 
 n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , 
 n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , 
 n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , 
 n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , 
 n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , 
 n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , 
 n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , 
 n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , 
 n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , 
 n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , 
 n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , 
 n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , 
 n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , 
 n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , 
 n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , 
 n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , 
 n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , 
 n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , 
 n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , 
 n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , 
 n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , 
 n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , 
 n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , 
 n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , 
 n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , 
 n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , 
 n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , 
 n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , 
 n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , 
 n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , 
 n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , 
 n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , 
 n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , 
 n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , 
 n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , 
 n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , 
 n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , 
 n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , 
 n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , 
 n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , 
 n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , 
 n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , 
 n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , 
 n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , 
 n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , 
 n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , 
 n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , 
 n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , 
 n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , 
 n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , 
 n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , 
 n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , 
 n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , 
 n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , 
 n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , 
 n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , 
 n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , 
 n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , 
 n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , 
 n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , 
 n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , 
 n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , 
 n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , 
 n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , 
 n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , 
 n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , 
 n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , 
 n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , 
 n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , 
 n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , 
 n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , 
 n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , 
 n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , 
 n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , 
 n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , 
 n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , 
 n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , 
 n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , 
 n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , 
 n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , 
 n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , 
 n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , 
 n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , 
 n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , 
 n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , 
 n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , 
 n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , 
 n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , 
 n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , 
 n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , 
 n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , 
 n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , 
 n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , 
 n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , 
 n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , 
 n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , 
 n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , 
 n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , 
 n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , 
 n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , 
 n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , 
 n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , 
 n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , 
 n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , 
 n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , 
 n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , 
 n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , 
 n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , 
 n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , 
 n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , 
 n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , 
 n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , 
 n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , 
 n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , 
 n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , 
 n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , 
 n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , 
 n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , 
 n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , 
 n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , 
 n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , 
 n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , 
 n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , 
 n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , 
 n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , 
 n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , 
 n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , 
 n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , 
 n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , 
 n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , 
 n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , 
 n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , 
 n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , 
 n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , 
 n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , 
 n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , 
 n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , 
 n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , 
 n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , 
 n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , 
 n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , 
 n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , 
 n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , 
 n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , 
 n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , 
 n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , 
 n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , 
 n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , 
 n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , 
 n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , 
 n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , 
 n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , 
 n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , 
 n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , 
 n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , 
 n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , 
 n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , 
 n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , 
 n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , 
 n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , 
 n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , 
 n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , 
 n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , 
 n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , 
 n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , 
 n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , 
 n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , 
 n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , 
 n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , 
 n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , 
 n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , 
 n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , 
 n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , 
 n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , 
 n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , 
 n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , 
 n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , 
 n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , 
 n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , 
 n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , 
 n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , 
 n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , 
 n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , 
 n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , 
 n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , 
 n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , 
 n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , 
 n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , 
 n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , 
 n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , 
 n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , 
 n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , 
 n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , 
 n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , 
 n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , 
 n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , 
 n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , 
 n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , 
 n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , 
 n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , 
 n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , 
 n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , 
 n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , 
 n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , 
 n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , 
 n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , 
 n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , 
 n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , 
 n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , 
 n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , 
 n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , 
 n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , 
 n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , 
 n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , 
 n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , 
 n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , 
 n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , 
 n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , 
 n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , 
 n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , 
 n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , 
 n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , 
 n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , 
 n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , 
 n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , 
 n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , 
 n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , 
 n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , 
 n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , 
 n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , 
 n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , 
 n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , 
 n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , 
 n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , 
 n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , 
 n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , 
 n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , 
 n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , 
 n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , 
 n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , 
 n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , 
 n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , 
 n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , 
 n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , 
 n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , 
 n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , 
 n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , 
 n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , 
 n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , 
 n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , 
 n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , 
 n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , 
 n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , 
 n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , 
 n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , 
 n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , 
 n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , 
 n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , 
 n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , 
 n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , 
 n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , 
 n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , 
 n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , 
 n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , 
 n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , 
 n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , 
 n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , 
 n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , 
 n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , 
 n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , 
 n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , 
 n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , 
 n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , 
 n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , 
 n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , 
 n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , 
 n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , 
 n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , 
 n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , 
 n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , 
 n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , 
 n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , 
 n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , 
 n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , 
 n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , 
 n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , 
 n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , 
 n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , 
 n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , 
 n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , 
 n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , 
 n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , 
 n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , 
 n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , 
 n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , 
 n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , 
 n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , 
 n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , 
 n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , 
 n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , 
 n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , 
 n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , 
 n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , 
 n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , 
 n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , 
 n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , 
 n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , 
 n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , 
 n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , 
 n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , 
 n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , 
 n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , 
 n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , 
 n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , 
 n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , 
 n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , 
 n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , 
 n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , 
 n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , 
 n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , 
 n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , 
 n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , 
 n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , 
 n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , 
 n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , 
 n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , 
 n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , 
 n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , 
 n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , 
 n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , 
 n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , 
 n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , 
 n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , 
 n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , 
 n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , 
 n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , 
 n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , 
 n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , 
 n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , 
 n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , 
 n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , 
 n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , 
 n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , 
 n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , 
 n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , 
 n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , 
 n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , 
 n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , 
 n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , 
 n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , 
 n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , 
 n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , 
 n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , 
 n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , 
 n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , 
 n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , 
 n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , 
 n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , 
 n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , 
 n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , 
 n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , 
 n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , 
 n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , 
 n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , 
 n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , 
 n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , 
 n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , 
 n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , 
 n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , 
 n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , 
 n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , 
 n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , 
 n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , 
 n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , 
 n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , 
 n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , 
 n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , 
 n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , 
 n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , 
 n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , 
 n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , 
 n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , 
 n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , 
 n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , 
 n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , 
 n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , 
 n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , 
 n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , 
 n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , 
 n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , 
 n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , 
 n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , 
 n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , 
 n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , 
 n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , 
 n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , 
 n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , 
 n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , 
 n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , 
 n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , 
 n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , 
 n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , 
 n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , 
 n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , 
 n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , 
 n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , 
 n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , 
 n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , 
 n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , 
 n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , 
 n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , 
 n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , 
 n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , 
 n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , 
 n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , 
 n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , 
 n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , 
 n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , 
 n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , 
 n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , 
 n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , 
 n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , 
 n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , 
 n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , 
 n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , 
 n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , 
 n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , 
 n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , 
 n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , 
 n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , 
 n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , 
 n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , 
 n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , 
 n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , 
 n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , 
 n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , 
 n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , 
 n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , 
 n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , 
 n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , 
 n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , 
 n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , 
 n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , 
 n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , 
 n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , 
 n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , 
 n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , 
 n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , 
 n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , 
 n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , 
 n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , 
 n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , 
 n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , 
 n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , 
 n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , 
 n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , 
 n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , 
 n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , 
 n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , 
 n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , 
 n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , 
 n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , 
 n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , 
 n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , 
 n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , 
 n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , 
 n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , 
 n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , 
 n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , 
 n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , 
 n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , 
 n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , 
 n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , 
 n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , 
 n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , 
 n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , 
 n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , 
 n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , 
 n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , 
 n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , 
 n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , 
 n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , 
 n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , 
 n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , 
 n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , 
 n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , 
 n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , 
 n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , 
 n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , 
 n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , 
 n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , 
 n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , 
 n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , 
 n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , 
 n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , 
 n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , 
 n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , 
 n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , 
 n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , 
 n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , 
 n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , 
 n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , 
 n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , 
 n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , 
 n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , 
 n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , 
 n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , 
 n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , 
 n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , 
 n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , 
 n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , 
 n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , 
 n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , 
 n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , 
 n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , 
 n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , 
 n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , 
 n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , 
 n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , 
 n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , 
 n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , 
 n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , 
 n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , 
 n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , 
 n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , 
 n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , 
 n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , 
 n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , 
 n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , 
 n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , 
 n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , 
 n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , 
 n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , 
 n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , 
 n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , 
 n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , 
 n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , 
 n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , 
 n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , 
 n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , 
 n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , 
 n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , 
 n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , 
 n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , 
 n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , 
 n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , 
 n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , 
 n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , 
 n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , 
 n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , 
 n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , 
 n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , 
 n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , 
 n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , 
 n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , 
 n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , 
 n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , 
 n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , 
 n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , 
 n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , 
 n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , 
 n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , 
 n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , 
 n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , 
 n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , 
 n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , 
 n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , 
 n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , 
 n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , 
 n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , 
 n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , 
 n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , 
 n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , 
 n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , 
 n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , 
 n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , 
 n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , 
 n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , 
 n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , 
 n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , 
 n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , 
 n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , 
 n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , 
 n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , 
 n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , 
 n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , 
 n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , 
 n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , 
 n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , 
 n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , 
 n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , 
 n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , 
 n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , 
 n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , 
 n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , 
 n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , 
 n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , 
 n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , 
 n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , 
 n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , 
 n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , 
 n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , 
 n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , 
 n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , 
 n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , 
 n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , 
 n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , 
 n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , 
 n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , 
 n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , 
 n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , 
 n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , 
 n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , 
 n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , 
 n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , 
 n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , 
 n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , 
 n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , 
 n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , 
 n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , 
 n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , 
 n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , 
 n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , 
 n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , 
 n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , 
 n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , 
 n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , 
 n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , 
 n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , 
 n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , 
 n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , 
 n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , 
 n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , 
 n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , 
 n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , 
 n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , 
 n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , 
 n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , 
 n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , 
 n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , 
 n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , 
 n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , 
 n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , 
 n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , 
 n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , 
 n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , 
 n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , 
 n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , 
 n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , 
 n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , 
 n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , 
 n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , 
 n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , 
 n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , 
 n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , 
 n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , 
 n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , 
 n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , 
 n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , 
 n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , 
 n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , 
 n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , 
 n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , 
 n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , 
 n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , 
 n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , 
 n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , 
 n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , 
 n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , 
 n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , 
 n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , 
 n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , 
 n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , 
 n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , 
 n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , 
 n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , 
 n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , 
 n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , 
 n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , 
 n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , 
 n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , 
 n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , 
 n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , 
 n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , 
 n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , 
 n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , 
 n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , 
 n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , 
 n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , 
 n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , 
 n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , 
 n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , 
 n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , 
 n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , 
 n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , 
 n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , 
 n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , 
 n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , 
 n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , 
 n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , 
 n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , 
 n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , 
 n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , 
 n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , 
 n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , 
 n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , 
 n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , 
 n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , 
 n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , 
 n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , 
 n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , 
 n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , 
 n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , 
 n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , 
 n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , 
 n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , 
 n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , 
 n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , 
 n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , 
 n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , 
 n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , 
 n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , 
 n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , 
 n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , 
 n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , 
 n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , 
 n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , 
 n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , 
 n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , 
 n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , 
 n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , 
 n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , 
 n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , 
 n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , 
 n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , 
 n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , 
 n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , 
 n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , 
 n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , 
 n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , 
 n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , 
 n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , 
 n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , 
 n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , 
 n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , 
 n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , 
 n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , 
 n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , 
 n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , 
 n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , 
 n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , 
 n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , 
 n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , 
 n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , 
 n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , 
 n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , 
 n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , 
 n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , 
 n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , 
 n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , 
 n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , 
 n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , 
 n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , 
 n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , 
 n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , 
 n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , 
 n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , 
 n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , 
 n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , 
 n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , 
 n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , 
 n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , 
 n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , 
 n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , 
 n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , 
 n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , 
 n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , 
 n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , 
 n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , 
 n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , 
 n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , 
 n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , 
 n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , 
 n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , 
 n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , 
 n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , 
 n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , 
 n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , 
 n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , 
 n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , 
 n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , 
 n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , 
 n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , 
 n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , 
 n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , 
 n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , 
 n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , 
 n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , 
 n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , 
 n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , 
 n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , 
 n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , 
 n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , 
 n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , 
 n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , 
 n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , 
 n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , 
 n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , 
 n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , 
 n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , 
 n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , 
 n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , 
 n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , 
 n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , 
 n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , 
 n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , 
 n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , 
 n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , 
 n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , 
 n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , 
 n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , 
 n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , 
 n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , 
 n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , 
 n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , 
 n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , 
 n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , 
 n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , 
 n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , 
 n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , 
 n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , 
 n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , 
 n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , 
 n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , 
 n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , 
 n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , 
 n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , 
 n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , 
 n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , 
 n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , 
 n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , 
 n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , 
 n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , 
 n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , 
 n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , 
 n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , 
 n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , 
 n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , 
 n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , 
 n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , 
 n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , 
 n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , 
 n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , 
 n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , 
 n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , 
 n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , 
 n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , 
 n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , 
 n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , 
 n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , 
 n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , 
 n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , 
 n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , 
 n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , 
 n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , 
 n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , 
 n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , 
 n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , 
 n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , 
 n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , 
 n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , 
 n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , 
 n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , 
 n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , 
 n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , 
 n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , 
 n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , 
 n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , 
 n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , 
 n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , 
 n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , 
 n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , 
 n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , 
 n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , 
 n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , 
 n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , 
 n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , 
 n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , 
 n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , 
 n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , 
 n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , 
 n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , 
 n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , 
 n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , 
 n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , 
 n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , 
 n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , 
 n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , 
 n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , 
 n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , 
 n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , 
 n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , 
 n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , 
 n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , 
 n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , 
 n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , 
 n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , 
 n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , 
 n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , 
 n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , 
 n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , 
 n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , 
 n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , 
 n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , 
 n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , 
 n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , 
 n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , 
 n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , 
 n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , 
 n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , 
 n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , 
 n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , 
 n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , 
 n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , 
 n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , 
 n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , 
 n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , 
 n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , 
 n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , 
 n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , 
 n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , 
 n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , 
 n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , 
 n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , 
 n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , 
 n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , 
 n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , 
 n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , 
 n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , 
 n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , 
 n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , 
 n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , 
 n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , 
 n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , 
 n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , 
 n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , 
 n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , 
 n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , 
 n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , 
 n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , 
 n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , 
 n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , 
 n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , 
 n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , 
 n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , 
 n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , 
 n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , 
 n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , 
 n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , 
 n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , 
 n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , 
 n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , 
 n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , 
 n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , 
 n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , 
 n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , 
 n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , 
 n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , 
 n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , 
 n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , 
 n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , 
 n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , 
 n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , 
 n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , 
 n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , 
 n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , 
 n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , 
 n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , 
 n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , 
 n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , 
 n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , 
 n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , 
 n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , 
 n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , 
 n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , 
 n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , 
 n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , 
 n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , 
 n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , 
 n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , 
 n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , 
 n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , 
 n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , 
 n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , 
 n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , 
 n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , 
 n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , 
 n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , 
 n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , 
 n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , 
 n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , 
 n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , 
 n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , 
 n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , 
 n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , 
 n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , 
 n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , 
 n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , 
 n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , 
 n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , 
 n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , 
 n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , 
 n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , 
 n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , 
 n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , 
 n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , 
 n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , 
 n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , 
 n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , 
 n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , 
 n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , 
 n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , 
 n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , 
 n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , 
 n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , 
 n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , 
 n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , 
 n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , 
 n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , 
 n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , 
 n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , 
 n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , 
 n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , 
 n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , 
 n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , 
 n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , 
 n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , 
 n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , 
 n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , 
 n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , 
 n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , 
 n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , 
 n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , 
 n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , 
 n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , 
 n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , 
 n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , 
 n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , 
 n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , 
 n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , 
 n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , 
 n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , 
 n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , 
 n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , 
 n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , 
 n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , 
 n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , 
 n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , 
 n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , 
 n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , 
 n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , 
 n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , 
 n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , 
 n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , 
 n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , 
 n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , 
 n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , 
 n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , 
 n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , 
 n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , 
 n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , 
 n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , 
 n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , 
 n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , 
 n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , 
 n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , 
 n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , 
 n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , 
 n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , 
 n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , 
 n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , 
 n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , 
 n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , 
 n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , 
 n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , 
 n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , 
 n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , 
 n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , 
 n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , 
 n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , 
 n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , 
 n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , 
 n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , 
 n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , 
 n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , 
 n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , 
 n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , 
 n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , 
 n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , 
 n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , 
 n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , 
 n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , 
 n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , 
 n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , 
 n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , 
 n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , 
 n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , 
 n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , 
 n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , 
 n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , 
 n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , 
 n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , 
 n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , 
 n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , 
 n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , 
 n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , 
 n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , 
 n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , 
 n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , 
 n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , 
 n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , 
 n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , 
 n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , 
 n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , 
 n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , 
 n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , 
 n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , 
 n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , 
 n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , 
 n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , 
 n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , 
 n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , 
 n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , 
 n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , 
 n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , 
 n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , 
 n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , 
 n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , 
 n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , 
 n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , 
 n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , 
 n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , 
 n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , 
 n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , 
 n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , 
 n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , 
 n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , 
 n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , 
 n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , 
 n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , 
 n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , 
 n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , 
 n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , 
 n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , 
 n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , 
 n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , 
 n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , 
 n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , 
 n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , 
 n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , 
 n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , 
 n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , 
 n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , 
 n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , 
 n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , 
 n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , 
 n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , 
 n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , 
 n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , 
 n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , 
 n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , 
 n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , 
 n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , 
 n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , 
 n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , 
 n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , 
 n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , 
 n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , 
 n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , 
 n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , 
 n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , 
 n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , 
 n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , 
 n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , 
 n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , 
 n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , 
 n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , 
 n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , 
 n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , 
 n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , 
 n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , 
 n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , n64901 , n64902 , n64903 , n64904 , 
 n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , n64911 , n64912 , n64913 , n64914 , 
 n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , n64921 , n64922 , n64923 , n64924 , 
 n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , n64931 , n64932 , n64933 , n64934 , 
 n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , n64941 , n64942 , n64943 , n64944 , 
 n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , n64951 , n64952 , n64953 , n64954 , 
 n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , n64961 , n64962 , n64963 , n64964 , 
 n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , n64971 , n64972 , n64973 , n64974 , 
 n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , n64981 , n64982 , n64983 , n64984 , 
 n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , n64991 , n64992 , n64993 , n64994 , 
 n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , n65001 , n65002 , n65003 , n65004 , 
 n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , n65011 , n65012 , n65013 , n65014 , 
 n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , n65021 , n65022 , n65023 , n65024 , 
 n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , n65031 , n65032 , n65033 , n65034 , 
 n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , n65041 , n65042 , n65043 , n65044 , 
 n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , n65051 , n65052 , n65053 , n65054 , 
 n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , n65061 , n65062 , n65063 , n65064 , 
 n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , n65071 , n65072 , n65073 , n65074 , 
 n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , n65081 , n65082 , n65083 , n65084 , 
 n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , n65091 , n65092 , n65093 , n65094 , 
 n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , n65101 , n65102 , n65103 , n65104 , 
 n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , n65111 , n65112 , n65113 , n65114 , 
 n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , n65121 , n65122 , n65123 , n65124 , 
 n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , n65131 , n65132 , n65133 , n65134 , 
 n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , n65141 , n65142 , n65143 , n65144 , 
 n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , n65151 , n65152 , n65153 , n65154 , 
 n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , n65161 , n65162 , n65163 , n65164 , 
 n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , n65171 , n65172 , n65173 , n65174 , 
 n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , n65181 , n65182 , n65183 , n65184 , 
 n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , n65191 , n65192 , n65193 , n65194 , 
 n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , n65201 , n65202 , n65203 , n65204 , 
 n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , n65211 , n65212 , n65213 , n65214 , 
 n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , n65221 , n65222 , n65223 , n65224 , 
 n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , n65231 , n65232 , n65233 , n65234 , 
 n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , n65241 , n65242 , n65243 , n65244 , 
 n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , n65251 , n65252 , n65253 , n65254 , 
 n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , n65261 , n65262 , n65263 , n65264 , 
 n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , n65271 , n65272 , n65273 , n65274 , 
 n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , n65281 , n65282 , n65283 , n65284 , 
 n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , n65291 , n65292 , n65293 , n65294 , 
 n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , n65301 , n65302 , n65303 , n65304 , 
 n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , n65311 , n65312 , n65313 , n65314 , 
 n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , n65321 , n65322 , n65323 , n65324 , 
 n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , n65331 , n65332 , n65333 , n65334 , 
 n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , n65341 , n65342 , n65343 , n65344 , 
 n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , n65351 , n65352 , n65353 , n65354 , 
 n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , n65361 , n65362 , n65363 , n65364 , 
 n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , n65371 , n65372 , n65373 , n65374 , 
 n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , n65381 , n65382 , n65383 , n65384 , 
 n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , n65391 , n65392 , n65393 , n65394 , 
 n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , n65401 , n65402 , n65403 , n65404 , 
 n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , n65411 , n65412 , n65413 , n65414 , 
 n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , n65421 , n65422 , n65423 , n65424 , 
 n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , n65431 , n65432 , n65433 , n65434 , 
 n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , n65441 , n65442 , n65443 , n65444 , 
 n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , n65451 , n65452 , n65453 , n65454 , 
 n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , n65461 , n65462 , n65463 , n65464 , 
 n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , n65471 , n65472 , n65473 , n65474 , 
 n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , n65481 , n65482 , n65483 , n65484 , 
 n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , n65491 , n65492 , n65493 , n65494 , 
 n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , n65501 , n65502 , n65503 , n65504 , 
 n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , n65511 , n65512 , n65513 , n65514 , 
 n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , n65521 , n65522 , n65523 , n65524 , 
 n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , n65531 , n65532 , n65533 , n65534 , 
 n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , n65541 , n65542 , n65543 , n65544 , 
 n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , n65551 , n65552 , n65553 , n65554 , 
 n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , n65561 , n65562 , n65563 , n65564 , 
 n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , n65571 , n65572 , n65573 , n65574 , 
 n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , n65581 , n65582 , n65583 , n65584 , 
 n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , n65591 , n65592 , n65593 , n65594 , 
 n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , n65601 , n65602 , n65603 , n65604 , 
 n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , n65611 , n65612 , n65613 , n65614 , 
 n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , n65621 , n65622 , n65623 , n65624 , 
 n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , n65631 , n65632 , n65633 , n65634 , 
 n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , n65641 , n65642 , n65643 , n65644 , 
 n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , 
 n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , n65661 , n65662 , n65663 , n65664 , 
 n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , n65671 , n65672 , n65673 , n65674 , 
 n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , 
 n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , n65691 , n65692 , n65693 , n65694 , 
 n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , n65701 , n65702 , n65703 , n65704 , 
 n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , n65711 , n65712 , n65713 , n65714 , 
 n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , n65721 , n65722 , n65723 , n65724 , 
 n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , n65731 , n65732 , n65733 , n65734 , 
 n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , n65741 , n65742 , n65743 , n65744 , 
 n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , n65751 , n65752 , n65753 , n65754 , 
 n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , n65761 , n65762 , n65763 , n65764 , 
 n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , n65771 , n65772 , n65773 , n65774 , 
 n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , n65781 , n65782 , n65783 , n65784 , 
 n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , n65791 , n65792 , n65793 , n65794 , 
 n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , n65801 , n65802 , n65803 , n65804 , 
 n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , n65811 , n65812 , n65813 , n65814 , 
 n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , n65821 , n65822 , n65823 , n65824 , 
 n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , n65831 , n65832 , n65833 , n65834 , 
 n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , n65841 , n65842 , n65843 , n65844 , 
 n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , n65851 , n65852 , n65853 , n65854 , 
 n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , n65861 , n65862 , n65863 , n65864 , 
 n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , n65871 , n65872 , n65873 , n65874 , 
 n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , n65881 , n65882 , n65883 , n65884 , 
 n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , n65891 , n65892 , n65893 , n65894 , 
 n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , n65901 , n65902 , n65903 , n65904 , 
 n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , n65911 , n65912 , n65913 , n65914 , 
 n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , n65921 , n65922 , n65923 , n65924 , 
 n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , n65931 , n65932 , n65933 , n65934 , 
 n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , n65941 , n65942 , n65943 , n65944 , 
 n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , n65951 , n65952 , n65953 , n65954 , 
 n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , n65961 , n65962 , n65963 , n65964 , 
 n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , n65971 , n65972 , n65973 , n65974 , 
 n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , n65981 , n65982 , n65983 , n65984 , 
 n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , n65991 , n65992 , n65993 , n65994 , 
 n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , n66001 , n66002 , n66003 , n66004 , 
 n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , n66011 , n66012 , n66013 , n66014 , 
 n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , n66021 , n66022 , n66023 , n66024 , 
 n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , n66031 , n66032 , n66033 , n66034 , 
 n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , n66041 , n66042 , n66043 , n66044 , 
 n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , n66051 , n66052 , n66053 , n66054 , 
 n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , n66061 , n66062 , n66063 , n66064 , 
 n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , n66071 , n66072 , n66073 , n66074 , 
 n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , n66081 , n66082 , n66083 , n66084 , 
 n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , n66091 , n66092 , n66093 , n66094 , 
 n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , n66101 , n66102 , n66103 , n66104 , 
 n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , n66111 , n66112 , n66113 , n66114 , 
 n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , n66121 , n66122 , n66123 , n66124 , 
 n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , n66131 , n66132 , n66133 , n66134 , 
 n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , n66141 , n66142 , n66143 , n66144 , 
 n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , n66151 , n66152 , n66153 , n66154 , 
 n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , n66161 , n66162 , n66163 , n66164 , 
 n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , n66171 , n66172 , n66173 , n66174 , 
 n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , n66181 , n66182 , n66183 , n66184 , 
 n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , n66191 , n66192 , n66193 , n66194 , 
 n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , n66201 , n66202 , n66203 , n66204 , 
 n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , n66211 , n66212 , n66213 , n66214 , 
 n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , n66221 , n66222 , n66223 , n66224 , 
 n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , n66231 , n66232 , n66233 , n66234 , 
 n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , n66241 , n66242 , n66243 , n66244 , 
 n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , n66251 , n66252 , n66253 , n66254 , 
 n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , n66261 , n66262 , n66263 , n66264 , 
 n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , n66271 , n66272 , n66273 , n66274 , 
 n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , n66281 , n66282 , n66283 , n66284 , 
 n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , 
 n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , n66301 , n66302 , n66303 , n66304 , 
 n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , n66311 , n66312 , n66313 , n66314 , 
 n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , n66321 , n66322 , n66323 , n66324 , 
 n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , n66331 , n66332 , n66333 , n66334 , 
 n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , n66341 , n66342 , n66343 , n66344 , 
 n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , n66351 , n66352 , n66353 , n66354 , 
 n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , n66361 , n66362 , n66363 , n66364 , 
 n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , n66371 , n66372 , n66373 , n66374 , 
 n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , n66381 , n66382 , n66383 , n66384 , 
 n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , n66391 , n66392 , n66393 , n66394 , 
 n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , n66401 , n66402 , n66403 , n66404 , 
 n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , n66411 , n66412 , n66413 , n66414 , 
 n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , n66421 , n66422 , n66423 , n66424 , 
 n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , n66431 , n66432 , n66433 , n66434 , 
 n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , n66441 , n66442 , n66443 , n66444 , 
 n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , n66451 , n66452 , n66453 , n66454 , 
 n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , n66461 , n66462 , n66463 , n66464 , 
 n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , n66471 , n66472 , n66473 , n66474 , 
 n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , n66481 , n66482 , n66483 , n66484 , 
 n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , n66491 , n66492 , n66493 , n66494 , 
 n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , n66501 , n66502 , n66503 , n66504 , 
 n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , n66511 , n66512 , n66513 , n66514 , 
 n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , n66521 , n66522 , n66523 , n66524 , 
 n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , n66531 , n66532 , n66533 , n66534 , 
 n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , n66541 , n66542 , n66543 , n66544 , 
 n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , n66551 , n66552 , n66553 , n66554 , 
 n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , n66561 , n66562 , n66563 , n66564 , 
 n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , n66571 , n66572 , n66573 , n66574 , 
 n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , n66581 , n66582 , n66583 , n66584 , 
 n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , n66591 , n66592 , n66593 , n66594 , 
 n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , n66601 , n66602 , n66603 , n66604 , 
 n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , n66611 , n66612 , n66613 , n66614 , 
 n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , n66621 , n66622 , n66623 , n66624 , 
 n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , n66631 , n66632 , n66633 , n66634 , 
 n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , n66641 , n66642 , n66643 , n66644 , 
 n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , n66651 , n66652 , n66653 , n66654 , 
 n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , n66661 , n66662 , n66663 , n66664 , 
 n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , 
 n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , n66681 , n66682 , n66683 , n66684 , 
 n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , 
 n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , n66701 , n66702 , n66703 , n66704 , 
 n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , n66711 , n66712 , n66713 , n66714 , 
 n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , n66721 , n66722 , n66723 , n66724 , 
 n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , 
 n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , n66741 , n66742 , n66743 , n66744 , 
 n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , n66751 , n66752 , n66753 , n66754 , 
 n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , n66761 , n66762 , n66763 , n66764 , 
 n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , n66771 , n66772 , n66773 , n66774 , 
 n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , n66781 , n66782 , n66783 , n66784 , 
 n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , n66791 , n66792 , n66793 , n66794 , 
 n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , n66801 , n66802 , n66803 , n66804 , 
 n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , n66811 , n66812 , n66813 , n66814 , 
 n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , n66821 , n66822 , n66823 , n66824 , 
 n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , 
 n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , n66841 , n66842 , n66843 , n66844 , 
 n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , n66851 , n66852 , n66853 , n66854 , 
 n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , n66861 , n66862 , n66863 , n66864 , 
 n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , n66871 , n66872 , n66873 , n66874 , 
 n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , n66881 , n66882 , n66883 , n66884 , 
 n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , n66891 , n66892 , n66893 , n66894 , 
 n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , n66901 , n66902 , n66903 , n66904 , 
 n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , n66911 , n66912 , n66913 , n66914 , 
 n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , n66921 , n66922 , n66923 , n66924 , 
 n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , n66931 , n66932 , n66933 , n66934 , 
 n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , n66941 , n66942 , n66943 , n66944 , 
 n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , n66951 , n66952 , n66953 , n66954 , 
 n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , n66961 , n66962 , n66963 , n66964 , 
 n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , n66971 , n66972 , n66973 , n66974 , 
 n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , n66981 , n66982 , n66983 , n66984 , 
 n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , n66991 , n66992 , n66993 , n66994 , 
 n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , n67001 , n67002 , n67003 , n67004 , 
 n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , n67011 , n67012 , n67013 , n67014 , 
 n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , n67021 , n67022 , n67023 , n67024 , 
 n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , n67031 , n67032 , n67033 , n67034 , 
 n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , n67041 , n67042 , n67043 , n67044 , 
 n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , n67051 , n67052 , n67053 , n67054 , 
 n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , n67061 , n67062 , n67063 , n67064 , 
 n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , n67071 , n67072 , n67073 , n67074 , 
 n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , n67081 , n67082 , n67083 , n67084 , 
 n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , n67091 , n67092 , n67093 , n67094 , 
 n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , n67101 , n67102 , n67103 , n67104 , 
 n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , n67111 , n67112 , n67113 , n67114 , 
 n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , n67121 , n67122 , n67123 , n67124 , 
 n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , n67131 , n67132 , n67133 , n67134 , 
 n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , n67141 , n67142 , n67143 , n67144 , 
 n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , n67151 , n67152 , n67153 , n67154 , 
 n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , n67161 , n67162 , n67163 , n67164 , 
 n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , n67171 , n67172 , n67173 , n67174 , 
 n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , n67181 , n67182 , n67183 , n67184 , 
 n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , n67191 , n67192 , n67193 , n67194 , 
 n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , n67201 , n67202 , n67203 , n67204 , 
 n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , n67211 , n67212 , n67213 , n67214 , 
 n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , n67221 , n67222 , n67223 , n67224 , 
 n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , n67231 , n67232 , n67233 , n67234 , 
 n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , n67241 , n67242 , n67243 , n67244 , 
 n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , n67251 , n67252 , n67253 , n67254 , 
 n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , n67261 , n67262 , n67263 , n67264 , 
 n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , n67271 , n67272 , n67273 , n67274 , 
 n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , n67281 , n67282 , n67283 , n67284 , 
 n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , n67291 , n67292 , n67293 , n67294 , 
 n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , n67301 , n67302 , n67303 , n67304 , 
 n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , 
 n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , n67321 , n67322 , n67323 , n67324 , 
 n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , n67331 , n67332 , n67333 , n67334 , 
 n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , 
 n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , n67351 , n67352 , n67353 , n67354 , 
 n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , n67361 , n67362 , n67363 , n67364 , 
 n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , n67371 , n67372 , n67373 , n67374 , 
 n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , n67381 , n67382 , n67383 , n67384 , 
 n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , n67391 , n67392 , n67393 , n67394 , 
 n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , n67401 , n67402 , n67403 , n67404 , 
 n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , n67411 , n67412 , n67413 , n67414 , 
 n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , 
 n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , n67431 , n67432 , n67433 , n67434 , 
 n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , n67441 , n67442 , n67443 , n67444 , 
 n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , 
 n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , n67461 , n67462 , n67463 , n67464 , 
 n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , 
 n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , 
 n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , n67491 , n67492 , n67493 , n67494 , 
 n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , n67501 , n67502 , n67503 , n67504 , 
 n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , n67511 , n67512 , n67513 , n67514 , 
 n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , n67521 , n67522 , n67523 , n67524 , 
 n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , n67531 , n67532 , n67533 , n67534 , 
 n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , n67541 , n67542 , n67543 , n67544 , 
 n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , n67551 , n67552 , n67553 , n67554 , 
 n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , n67561 , n67562 , n67563 , n67564 , 
 n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , n67571 , n67572 , n67573 , n67574 , 
 n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , n67581 , n67582 , n67583 , n67584 , 
 n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , n67591 , n67592 , n67593 , n67594 , 
 n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , n67601 , n67602 , n67603 , n67604 , 
 n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , 
 n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , n67621 , n67622 , n67623 , n67624 , 
 n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , n67631 , n67632 , n67633 , n67634 , 
 n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , 
 n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , 
 n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , n67661 , n67662 , n67663 , n67664 , 
 n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , n67671 , n67672 , n67673 , n67674 , 
 n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , 
 n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , 
 n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , n67701 , n67702 , n67703 , n67704 , 
 n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , 
 n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , 
 n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , 
 n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , n67741 , n67742 , n67743 , n67744 , 
 n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , n67751 , n67752 , n67753 , n67754 , 
 n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , n67761 , n67762 , n67763 , n67764 , 
 n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , n67771 , n67772 , n67773 , n67774 , 
 n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , n67781 , n67782 , n67783 , n67784 , 
 n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , n67791 , n67792 , n67793 , n67794 , 
 n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , n67801 , n67802 , n67803 , n67804 , 
 n67805 , n67806 , n67807 , n67808 , n67809 , n67810 , n67811 , n67812 , n67813 , n67814 , 
 n67815 , n67816 , n67817 , n67818 , n67819 , n67820 , n67821 , n67822 , n67823 , n67824 , 
 n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , n67831 , n67832 , n67833 , n67834 , 
 n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , n67841 , n67842 , n67843 , n67844 , 
 n67845 , n67846 , n67847 , n67848 , n67849 , n67850 , n67851 , n67852 , n67853 , n67854 , 
 n67855 , n67856 , n67857 , n67858 , n67859 , n67860 , n67861 , n67862 , n67863 , n67864 , 
 n67865 , n67866 , n67867 , n67868 , n67869 , n67870 , n67871 , n67872 , n67873 , n67874 , 
 n67875 , n67876 , n67877 , n67878 , n67879 , n67880 , n67881 , n67882 , n67883 , n67884 , 
 n67885 , n67886 , n67887 , n67888 , n67889 , n67890 , n67891 , n67892 , n67893 , n67894 , 
 n67895 , n67896 , n67897 , n67898 , n67899 , n67900 , n67901 , n67902 , n67903 , n67904 , 
 n67905 , n67906 , n67907 , n67908 , n67909 , n67910 , n67911 , n67912 , n67913 , n67914 , 
 n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , n67921 , n67922 , n67923 , n67924 , 
 n67925 , n67926 , n67927 , n67928 , n67929 , n67930 , n67931 , n67932 , n67933 , n67934 , 
 n67935 , n67936 , n67937 , n67938 , n67939 , n67940 , n67941 , n67942 , n67943 , n67944 , 
 n67945 , n67946 , n67947 , n67948 , n67949 , n67950 , n67951 , n67952 , n67953 , n67954 , 
 n67955 , n67956 , n67957 , n67958 , n67959 , n67960 , n67961 , n67962 , n67963 , n67964 , 
 n67965 , n67966 , n67967 , n67968 , n67969 , n67970 , n67971 , n67972 , n67973 , n67974 , 
 n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , n67981 , n67982 , n67983 , n67984 , 
 n67985 , n67986 , n67987 , n67988 , n67989 , n67990 , n67991 , n67992 , n67993 , n67994 , 
 n67995 , n67996 , n67997 , n67998 , n67999 , n68000 , n68001 , n68002 , n68003 , n68004 , 
 n68005 , n68006 , n68007 , n68008 , n68009 , n68010 , n68011 , n68012 , n68013 , n68014 , 
 n68015 , n68016 , n68017 , n68018 , n68019 , n68020 , n68021 , n68022 , n68023 , n68024 , 
 n68025 , n68026 , n68027 , n68028 , n68029 , n68030 , n68031 , n68032 , n68033 , n68034 , 
 n68035 , n68036 , n68037 , n68038 , n68039 , n68040 , n68041 , n68042 , n68043 , n68044 , 
 n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , n68051 , n68052 , n68053 , n68054 , 
 n68055 , n68056 , n68057 , n68058 , n68059 , n68060 , n68061 , n68062 , n68063 , n68064 , 
 n68065 , n68066 , n68067 , n68068 , n68069 , n68070 , n68071 , n68072 , n68073 , n68074 , 
 n68075 , n68076 , n68077 , n68078 , n68079 , n68080 , n68081 , n68082 , n68083 , n68084 , 
 n68085 , n68086 , n68087 , n68088 , n68089 , n68090 , n68091 , n68092 , n68093 , n68094 , 
 n68095 , n68096 , n68097 , n68098 , n68099 , n68100 , n68101 , n68102 , n68103 , n68104 , 
 n68105 , n68106 , n68107 , n68108 , n68109 , n68110 , n68111 , n68112 , n68113 , n68114 , 
 n68115 , n68116 , n68117 , n68118 , n68119 , n68120 , n68121 , n68122 , n68123 , n68124 , 
 n68125 , n68126 , n68127 , n68128 , n68129 , n68130 , n68131 , n68132 , n68133 , n68134 , 
 n68135 , n68136 , n68137 , n68138 , n68139 , n68140 , n68141 , n68142 , n68143 , n68144 , 
 n68145 , n68146 , n68147 , n68148 , n68149 , n68150 , n68151 , n68152 , n68153 , n68154 , 
 n68155 , n68156 , n68157 , n68158 , n68159 , n68160 , n68161 , n68162 , n68163 , n68164 , 
 n68165 , n68166 , n68167 , n68168 , n68169 , n68170 , n68171 , n68172 , n68173 , n68174 , 
 n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , n68181 , n68182 , n68183 , n68184 , 
 n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , n68191 , n68192 , n68193 , n68194 , 
 n68195 , n68196 , n68197 , n68198 , n68199 , n68200 , n68201 , n68202 , n68203 , n68204 , 
 n68205 , n68206 , n68207 , n68208 , n68209 , n68210 , n68211 , n68212 , n68213 , n68214 , 
 n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , n68221 , n68222 , n68223 , n68224 , 
 n68225 , n68226 , n68227 , n68228 , n68229 , n68230 , n68231 , n68232 , n68233 , n68234 , 
 n68235 , n68236 , n68237 , n68238 , n68239 , n68240 , n68241 , n68242 , n68243 , n68244 , 
 n68245 , n68246 , n68247 , n68248 , n68249 , n68250 , n68251 , n68252 , n68253 , n68254 , 
 n68255 , n68256 , n68257 , n68258 , n68259 , n68260 , n68261 , n68262 , n68263 , n68264 , 
 n68265 , n68266 , n68267 , n68268 , n68269 , n68270 , n68271 , n68272 , n68273 , n68274 , 
 n68275 , n68276 , n68277 , n68278 , n68279 , n68280 , n68281 , n68282 , n68283 , n68284 , 
 n68285 , n68286 , n68287 , n68288 , n68289 , n68290 , n68291 , n68292 , n68293 , n68294 , 
 n68295 , n68296 , n68297 , n68298 , n68299 , n68300 , n68301 , n68302 , n68303 , n68304 , 
 n68305 , n68306 , n68307 , n68308 , n68309 , n68310 , n68311 , n68312 , n68313 , n68314 , 
 n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , n68321 , n68322 , n68323 , n68324 , 
 n68325 , n68326 , n68327 , n68328 , n68329 , n68330 , n68331 , n68332 , n68333 , n68334 , 
 n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , n68341 , n68342 , n68343 , n68344 , 
 n68345 , n68346 , n68347 , n68348 , n68349 , n68350 , n68351 , n68352 , n68353 , n68354 , 
 n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , n68361 , n68362 , n68363 , n68364 , 
 n68365 , n68366 , n68367 , n68368 , n68369 , n68370 , n68371 , n68372 , n68373 , n68374 , 
 n68375 , n68376 , n68377 , n68378 , n68379 , n68380 , n68381 , n68382 , n68383 , n68384 , 
 n68385 , n68386 , n68387 , n68388 , n68389 , n68390 , n68391 , n68392 , n68393 , n68394 , 
 n68395 , n68396 , n68397 , n68398 , n68399 , n68400 , n68401 , n68402 , n68403 , n68404 , 
 n68405 , n68406 , n68407 , n68408 , n68409 , n68410 , n68411 , n68412 , n68413 , n68414 , 
 n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , n68421 , n68422 , n68423 , n68424 , 
 n68425 , n68426 , n68427 , n68428 , n68429 , n68430 , n68431 , n68432 , n68433 , n68434 , 
 n68435 , n68436 , n68437 , n68438 , n68439 , n68440 , n68441 , n68442 , n68443 , n68444 , 
 n68445 , n68446 , n68447 , n68448 , n68449 , n68450 , n68451 , n68452 , n68453 , n68454 , 
 n68455 , n68456 , n68457 , n68458 , n68459 , n68460 , n68461 , n68462 , n68463 , n68464 , 
 n68465 , n68466 , n68467 , n68468 , n68469 , n68470 , n68471 , n68472 , n68473 , n68474 , 
 n68475 , n68476 , n68477 , n68478 , n68479 , n68480 , n68481 , n68482 , n68483 , n68484 , 
 n68485 , n68486 , n68487 , n68488 , n68489 , n68490 , n68491 , n68492 , n68493 , n68494 , 
 n68495 , n68496 , n68497 , n68498 , n68499 , n68500 , n68501 , n68502 , n68503 , n68504 , 
 n68505 , n68506 , n68507 , n68508 , n68509 , n68510 , n68511 , n68512 , n68513 , n68514 , 
 n68515 , n68516 , n68517 , n68518 , n68519 , n68520 , n68521 , n68522 , n68523 , n68524 , 
 n68525 , n68526 , n68527 , n68528 , n68529 , n68530 , n68531 , n68532 , n68533 , n68534 , 
 n68535 , n68536 , n68537 , n68538 , n68539 , n68540 , n68541 , n68542 , n68543 , n68544 , 
 n68545 , n68546 , n68547 , n68548 , n68549 , n68550 , n68551 , n68552 , n68553 , n68554 , 
 n68555 , n68556 , n68557 , n68558 , n68559 , n68560 , n68561 , n68562 , n68563 , n68564 , 
 n68565 , n68566 , n68567 , n68568 , n68569 , n68570 , n68571 , n68572 , n68573 , n68574 , 
 n68575 , n68576 , n68577 , n68578 , n68579 , n68580 , n68581 , n68582 , n68583 , n68584 , 
 n68585 , n68586 , n68587 , n68588 , n68589 , n68590 , n68591 , n68592 , n68593 , n68594 , 
 n68595 , n68596 , n68597 , n68598 , n68599 , n68600 , n68601 , n68602 , n68603 , n68604 , 
 n68605 , n68606 , n68607 , n68608 , n68609 , n68610 , n68611 , n68612 , n68613 , n68614 , 
 n68615 , n68616 , n68617 , n68618 , n68619 , n68620 , n68621 , n68622 , n68623 , n68624 , 
 n68625 , n68626 , n68627 , n68628 , n68629 , n68630 , n68631 , n68632 , n68633 , n68634 , 
 n68635 , n68636 , n68637 , n68638 , n68639 , n68640 , n68641 , n68642 , n68643 , n68644 , 
 n68645 , n68646 , n68647 , n68648 , n68649 , n68650 , n68651 , n68652 , n68653 , n68654 , 
 n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , n68661 , n68662 , n68663 , n68664 , 
 n68665 , n68666 , n68667 , n68668 , n68669 , n68670 , n68671 , n68672 , n68673 , n68674 , 
 n68675 , n68676 , n68677 , n68678 , n68679 , n68680 , n68681 , n68682 , n68683 , n68684 , 
 n68685 , n68686 , n68687 , n68688 , n68689 , n68690 , n68691 , n68692 , n68693 , n68694 , 
 n68695 , n68696 , n68697 , n68698 , n68699 , n68700 , n68701 , n68702 , n68703 , n68704 , 
 n68705 , n68706 , n68707 , n68708 , n68709 , n68710 , n68711 , n68712 , n68713 , n68714 , 
 n68715 , n68716 , n68717 , n68718 , n68719 , n68720 , n68721 , n68722 , n68723 , n68724 , 
 n68725 , n68726 , n68727 , n68728 , n68729 , n68730 , n68731 , n68732 , n68733 , n68734 , 
 n68735 , n68736 , n68737 , n68738 , n68739 , n68740 , n68741 , n68742 , n68743 , n68744 , 
 n68745 , n68746 , n68747 , n68748 , n68749 , n68750 , n68751 , n68752 , n68753 , n68754 , 
 n68755 , n68756 , n68757 , n68758 , n68759 , n68760 , n68761 , n68762 , n68763 , n68764 , 
 n68765 , n68766 , n68767 , n68768 , n68769 , n68770 , n68771 , n68772 , n68773 , n68774 , 
 n68775 , n68776 , n68777 , n68778 , n68779 , n68780 , n68781 , n68782 , n68783 , n68784 , 
 n68785 , n68786 , n68787 , n68788 , n68789 , n68790 , n68791 , n68792 , n68793 , n68794 , 
 n68795 , n68796 , n68797 , n68798 , n68799 , n68800 , n68801 , n68802 , n68803 , n68804 , 
 n68805 , n68806 , n68807 , n68808 , n68809 , n68810 , n68811 , n68812 , n68813 , n68814 , 
 n68815 , n68816 , n68817 , n68818 , n68819 , n68820 , n68821 , n68822 , n68823 , n68824 , 
 n68825 , n68826 , n68827 , n68828 , n68829 , n68830 , n68831 , n68832 , n68833 , n68834 , 
 n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , n68841 , n68842 , n68843 , n68844 , 
 n68845 , n68846 , n68847 , n68848 , n68849 , n68850 , n68851 , n68852 , n68853 , n68854 , 
 n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , n68861 , n68862 , n68863 , n68864 , 
 n68865 , n68866 , n68867 , n68868 , n68869 , n68870 , n68871 , n68872 , n68873 , n68874 , 
 n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , n68881 , n68882 , n68883 , n68884 , 
 n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , n68891 , n68892 , n68893 , n68894 , 
 n68895 , n68896 , n68897 , n68898 , n68899 , n68900 , n68901 , n68902 , n68903 , n68904 , 
 n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , n68911 , n68912 , n68913 , n68914 , 
 n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , n68921 , n68922 , n68923 , n68924 , 
 n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , n68931 , n68932 , n68933 , n68934 , 
 n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , n68941 , n68942 , n68943 , n68944 , 
 n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , 
 n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , n68961 , n68962 , n68963 , n68964 , 
 n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , n68971 , n68972 , n68973 , n68974 , 
 n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , n68981 , n68982 , n68983 , n68984 , 
 n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , n68991 , n68992 , n68993 , n68994 , 
 n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , 
 n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , n69011 , n69012 , n69013 , n69014 , 
 n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , n69021 , n69022 , n69023 , n69024 , 
 n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , n69031 , n69032 , n69033 , n69034 , 
 n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , n69041 , n69042 , n69043 , n69044 , 
 n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , n69051 , n69052 , n69053 , n69054 , 
 n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , n69061 , n69062 , n69063 , n69064 , 
 n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , n69071 , n69072 , n69073 , n69074 , 
 n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , 
 n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , n69091 , n69092 , n69093 , n69094 , 
 n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , n69101 , n69102 , n69103 , n69104 , 
 n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , n69111 , n69112 , n69113 , n69114 , 
 n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , n69121 , n69122 , n69123 , n69124 , 
 n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , n69131 , n69132 , n69133 , n69134 , 
 n69135 , n69136 , n69137 , n69138 , n69139 , n69140 , n69141 , n69142 , n69143 , n69144 , 
 n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , n69151 , n69152 , n69153 , n69154 , 
 n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , n69161 , n69162 , n69163 , n69164 , 
 n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , n69171 , n69172 , n69173 , n69174 , 
 n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , n69181 , n69182 , n69183 , n69184 , 
 n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , n69191 , n69192 , n69193 , n69194 , 
 n69195 , n69196 , n69197 , n69198 , n69199 , n69200 , n69201 , n69202 , n69203 , n69204 , 
 n69205 , n69206 , n69207 , n69208 , n69209 , n69210 , n69211 , n69212 , n69213 , n69214 , 
 n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , n69221 , n69222 , n69223 , n69224 , 
 n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , n69231 , n69232 , n69233 , n69234 , 
 n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , n69241 , n69242 , n69243 , n69244 , 
 n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , 
 n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , n69261 , n69262 , n69263 , n69264 , 
 n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , n69271 , n69272 , n69273 , n69274 , 
 n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , 
 n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , n69291 , n69292 , n69293 , n69294 , 
 n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , n69301 , n69302 , n69303 , n69304 , 
 n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , n69311 , n69312 , n69313 , n69314 , 
 n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , n69321 , n69322 , n69323 , n69324 , 
 n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , n69331 , n69332 , n69333 , n69334 , 
 n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , n69341 , n69342 , n69343 , n69344 , 
 n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , n69351 , n69352 , n69353 , n69354 , 
 n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , n69361 , n69362 , n69363 , n69364 , 
 n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , 
 n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , n69381 , n69382 , n69383 , n69384 , 
 n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , n69391 , n69392 , n69393 , n69394 , 
 n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , n69401 , n69402 , n69403 , n69404 , 
 n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , 
 n69415 , n69416 , n69417 , n69418 , n69419 , n69420 , n69421 , n69422 , n69423 , n69424 , 
 n69425 , n69426 , n69427 , n69428 , n69429 , n69430 , n69431 , n69432 , n69433 , n69434 , 
 n69435 , n69436 , n69437 , n69438 , n69439 , n69440 , n69441 , n69442 , n69443 , n69444 , 
 n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , n69451 , n69452 , n69453 , n69454 , 
 n69455 , n69456 , n69457 , n69458 , n69459 , n69460 , n69461 , n69462 , n69463 , n69464 , 
 n69465 , n69466 , n69467 , n69468 , n69469 , n69470 , n69471 , n69472 , n69473 , n69474 , 
 n69475 , n69476 , n69477 , n69478 , n69479 , n69480 , n69481 , n69482 , n69483 , n69484 , 
 n69485 , n69486 , n69487 , n69488 , n69489 , n69490 , n69491 , n69492 , n69493 , n69494 , 
 n69495 , n69496 , n69497 , n69498 , n69499 , n69500 , n69501 , n69502 , n69503 , n69504 , 
 n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , n69511 , n69512 , n69513 , n69514 , 
 n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , n69521 , n69522 , n69523 , n69524 , 
 n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , n69531 , n69532 , n69533 , n69534 , 
 n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , n69541 , n69542 , n69543 , n69544 , 
 n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , n69551 , n69552 , n69553 , n69554 , 
 n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , n69561 , n69562 , n69563 , n69564 , 
 n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , 
 n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , n69581 , n69582 , n69583 , n69584 , 
 n69585 , n69586 , n69587 , n69588 , n69589 , n69590 , n69591 , n69592 , n69593 , n69594 , 
 n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , n69601 , n69602 , n69603 , n69604 , 
 n69605 , n69606 , n69607 , n69608 , n69609 , n69610 , n69611 , n69612 , n69613 , n69614 , 
 n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , n69621 , n69622 , n69623 , n69624 , 
 n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , n69631 , n69632 , n69633 , n69634 , 
 n69635 , n69636 , n69637 , n69638 , n69639 , n69640 , n69641 , n69642 , n69643 , n69644 , 
 n69645 , n69646 , n69647 , n69648 , n69649 , n69650 , n69651 , n69652 , n69653 , n69654 , 
 n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , n69661 , n69662 , n69663 , n69664 , 
 n69665 , n69666 , n69667 , n69668 , n69669 , n69670 , n69671 , n69672 , n69673 , n69674 , 
 n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , n69681 , n69682 , n69683 , n69684 , 
 n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , n69691 , n69692 , n69693 , n69694 , 
 n69695 , n69696 , n69697 , n69698 , n69699 , n69700 , n69701 , n69702 , n69703 , n69704 , 
 n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , 
 n69715 , n69716 , n69717 , n69718 , n69719 , n69720 , n69721 , n69722 , n69723 , n69724 , 
 n69725 , n69726 , n69727 , n69728 , n69729 , n69730 , n69731 , n69732 , n69733 , n69734 , 
 n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , 
 n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , n69751 , n69752 , n69753 , n69754 , 
 n69755 , n69756 , n69757 , n69758 , n69759 , n69760 , n69761 , n69762 , n69763 , n69764 , 
 n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , n69771 , n69772 , n69773 , n69774 , 
 n69775 , n69776 , n69777 , n69778 , n69779 , n69780 , n69781 , n69782 , n69783 , n69784 , 
 n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , n69791 , n69792 , n69793 , n69794 , 
 n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , n69801 , n69802 , n69803 , n69804 , 
 n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , n69811 , n69812 , n69813 , n69814 , 
 n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , n69821 , n69822 , n69823 , n69824 , 
 n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , n69831 , n69832 , n69833 , n69834 , 
 n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , n69841 , n69842 , n69843 , n69844 , 
 n69845 , n69846 , n69847 , n69848 , n69849 , n69850 , n69851 , n69852 , n69853 , n69854 , 
 n69855 , n69856 , n69857 , n69858 , n69859 , n69860 , n69861 , n69862 , n69863 , n69864 , 
 n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , n69871 , n69872 , n69873 , n69874 , 
 n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , n69881 , n69882 , n69883 , n69884 , 
 n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , n69891 , n69892 , n69893 , n69894 , 
 n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , n69901 , n69902 , n69903 , n69904 , 
 n69905 , n69906 , n69907 , n69908 , n69909 , n69910 , n69911 , n69912 , n69913 , n69914 , 
 n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , n69921 , n69922 , n69923 , n69924 , 
 n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , n69931 , n69932 , n69933 , n69934 , 
 n69935 , n69936 , n69937 , n69938 , n69939 , n69940 , n69941 , n69942 , n69943 , n69944 , 
 n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , n69951 , n69952 , n69953 , n69954 , 
 n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , n69961 , n69962 , n69963 , n69964 , 
 n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , n69971 , n69972 , n69973 , n69974 , 
 n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , n69981 , n69982 , n69983 , n69984 , 
 n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , n69991 , n69992 , n69993 , n69994 , 
 n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , n70001 , n70002 , n70003 , n70004 , 
 n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , n70011 , n70012 , n70013 , n70014 , 
 n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , n70021 , n70022 , n70023 , n70024 , 
 n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , n70031 , n70032 , n70033 , n70034 , 
 n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , n70041 , n70042 , n70043 , n70044 , 
 n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , n70051 , n70052 , n70053 , n70054 , 
 n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , n70061 , n70062 , n70063 , n70064 , 
 n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , n70071 , n70072 , n70073 , n70074 , 
 n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , n70081 , n70082 , n70083 , n70084 , 
 n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , 
 n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , n70101 , n70102 , n70103 , n70104 , 
 n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , n70111 , n70112 , n70113 , n70114 , 
 n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , n70121 , n70122 , n70123 , n70124 , 
 n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , n70131 , n70132 , n70133 , n70134 , 
 n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , 
 n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , n70151 , n70152 , n70153 , n70154 , 
 n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , n70161 , n70162 , n70163 , n70164 , 
 n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , n70171 , n70172 , n70173 , n70174 , 
 n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , n70181 , n70182 , n70183 , n70184 , 
 n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , 
 n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , n70201 , n70202 , n70203 , n70204 , 
 n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , n70211 , n70212 , n70213 , n70214 , 
 n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , n70221 , n70222 , n70223 , n70224 , 
 n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , n70231 , n70232 , n70233 , n70234 , 
 n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , n70241 , n70242 , n70243 , n70244 , 
 n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , n70251 , n70252 , n70253 , n70254 , 
 n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , n70261 , n70262 , n70263 , n70264 , 
 n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , n70271 , n70272 , n70273 , n70274 , 
 n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , 
 n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , n70291 , n70292 , n70293 , n70294 , 
 n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , n70301 , n70302 , n70303 , n70304 , 
 n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , n70311 , n70312 , n70313 , n70314 , 
 n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , n70321 , n70322 , n70323 , n70324 , 
 n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , n70331 , n70332 , n70333 , n70334 , 
 n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , n70341 , n70342 , n70343 , n70344 , 
 n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , n70351 , n70352 , n70353 , n70354 , 
 n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , n70361 , n70362 , n70363 , n70364 , 
 n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , n70371 , n70372 , n70373 , n70374 , 
 n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , n70381 , n70382 , n70383 , n70384 , 
 n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , n70391 , n70392 , n70393 , n70394 , 
 n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , n70401 , n70402 , n70403 , n70404 , 
 n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , n70411 , n70412 , n70413 , n70414 , 
 n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , n70421 , n70422 , n70423 , n70424 , 
 n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , n70431 , n70432 , n70433 , n70434 , 
 n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , n70441 , n70442 , n70443 , n70444 , 
 n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , n70451 , n70452 , n70453 , n70454 , 
 n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , n70461 , n70462 , n70463 , n70464 , 
 n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , n70471 , n70472 , n70473 , n70474 , 
 n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , n70481 , n70482 , n70483 , n70484 , 
 n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , n70491 , n70492 , n70493 , n70494 , 
 n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , n70501 , n70502 , n70503 , n70504 , 
 n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , n70511 , n70512 , n70513 , n70514 , 
 n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , n70521 , n70522 , n70523 , n70524 , 
 n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , n70531 , n70532 , n70533 , n70534 , 
 n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , n70541 , n70542 , n70543 , n70544 , 
 n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , n70551 , n70552 , n70553 , n70554 , 
 n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , n70561 , n70562 , n70563 , n70564 , 
 n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , n70571 , n70572 , n70573 , n70574 , 
 n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , n70581 , n70582 , n70583 , n70584 , 
 n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , n70591 , n70592 , n70593 , n70594 , 
 n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , 
 n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , 
 n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , n70621 , n70622 , n70623 , n70624 , 
 n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , n70631 , n70632 , n70633 , n70634 , 
 n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , n70641 , n70642 , n70643 , n70644 , 
 n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , n70651 , n70652 , n70653 , n70654 , 
 n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , n70661 , n70662 , n70663 , n70664 , 
 n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , n70671 , n70672 , n70673 , n70674 , 
 n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , n70681 , n70682 , n70683 , n70684 , 
 n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , n70691 , n70692 , n70693 , n70694 , 
 n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , n70701 , n70702 , n70703 , n70704 , 
 n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , n70711 , n70712 , n70713 , n70714 , 
 n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , n70721 , n70722 , n70723 , n70724 , 
 n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , n70731 , n70732 , n70733 , n70734 , 
 n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , n70741 , n70742 , n70743 , n70744 , 
 n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , n70751 , n70752 , n70753 , n70754 , 
 n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , n70761 , n70762 , n70763 , n70764 , 
 n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , n70771 , n70772 , n70773 , n70774 , 
 n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , n70781 , n70782 , n70783 , n70784 , 
 n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , n70791 , n70792 , n70793 , n70794 , 
 n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , n70801 , n70802 , n70803 , n70804 , 
 n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , n70811 , n70812 , n70813 , n70814 , 
 n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , n70821 , n70822 , n70823 , n70824 , 
 n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , n70831 , n70832 , n70833 , n70834 , 
 n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , n70841 , n70842 , n70843 , n70844 , 
 n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , n70851 , n70852 , n70853 , n70854 , 
 n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , n70861 , n70862 , n70863 , n70864 , 
 n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , n70871 , n70872 , n70873 , n70874 , 
 n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , n70881 , n70882 , n70883 , n70884 , 
 n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , n70891 , n70892 , n70893 , n70894 , 
 n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , n70901 , n70902 , n70903 , n70904 , 
 n70905 , n70906 , n70907 , n70908 , n70909 , n70910 , n70911 , n70912 , n70913 , n70914 , 
 n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , n70921 , n70922 , n70923 , n70924 , 
 n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , n70931 , n70932 , n70933 , n70934 , 
 n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , n70941 , n70942 , n70943 , n70944 , 
 n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , n70951 , n70952 , n70953 , n70954 , 
 n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , n70961 , n70962 , n70963 , n70964 , 
 n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , n70971 , n70972 , n70973 , n70974 , 
 n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , n70981 , n70982 , n70983 , n70984 , 
 n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , n70991 , n70992 , n70993 , n70994 , 
 n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , n71001 , n71002 , n71003 , n71004 , 
 n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , 
 n71015 , n71016 , n71017 , n71018 , n71019 , n71020 , n71021 , n71022 , n71023 , n71024 , 
 n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , n71031 , n71032 , n71033 , n71034 , 
 n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , n71041 , n71042 , n71043 , n71044 , 
 n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , n71051 , n71052 , n71053 , n71054 , 
 n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , n71061 , n71062 , n71063 , n71064 , 
 n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , n71071 , n71072 , n71073 , n71074 , 
 n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , n71081 , n71082 , n71083 , n71084 , 
 n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , n71091 , n71092 , n71093 , n71094 , 
 n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , n71101 , n71102 , n71103 , n71104 , 
 n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , n71111 , n71112 , n71113 , n71114 , 
 n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , n71121 , n71122 , n71123 , n71124 , 
 n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , n71131 , n71132 , n71133 , n71134 , 
 n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , n71141 , n71142 , n71143 , n71144 , 
 n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , n71151 , n71152 , n71153 , n71154 , 
 n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , n71161 , n71162 , n71163 , n71164 , 
 n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , n71171 , n71172 , n71173 , n71174 , 
 n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , n71181 , n71182 , n71183 , n71184 , 
 n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , n71191 , n71192 , n71193 , n71194 , 
 n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , n71201 , n71202 , n71203 , n71204 , 
 n71205 , n71206 , n71207 , n71208 , n71209 , n71210 , n71211 , n71212 , n71213 , n71214 , 
 n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , n71221 , n71222 , n71223 , n71224 , 
 n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , n71231 , n71232 , n71233 , n71234 , 
 n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , n71241 , n71242 , n71243 , n71244 , 
 n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , n71251 , n71252 , n71253 , n71254 , 
 n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , n71261 , n71262 , n71263 , n71264 , 
 n71265 , n71266 , n71267 , n71268 , n71269 , n71270 , n71271 , n71272 , n71273 , n71274 , 
 n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , n71281 , n71282 , n71283 , n71284 , 
 n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , n71291 , n71292 , n71293 , n71294 , 
 n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , n71301 , n71302 , n71303 , n71304 , 
 n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , n71311 , n71312 , n71313 , n71314 , 
 n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , n71321 , n71322 , n71323 , n71324 , 
 n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , n71331 , n71332 , n71333 , n71334 , 
 n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , n71341 , n71342 , n71343 , n71344 , 
 n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , n71351 , n71352 , n71353 , n71354 , 
 n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , 
 n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , n71371 , n71372 , n71373 , n71374 , 
 n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , n71381 , n71382 , n71383 , n71384 , 
 n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , n71391 , n71392 , n71393 , n71394 , 
 n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , n71401 , n71402 , n71403 , n71404 , 
 n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , n71411 , n71412 , n71413 , n71414 , 
 n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , n71421 , n71422 , n71423 , n71424 , 
 n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , n71431 , n71432 , n71433 , n71434 , 
 n71435 , n71436 , n71437 , n71438 , n71439 , n71440 , n71441 , n71442 , n71443 , n71444 , 
 n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , n71451 , n71452 , n71453 , n71454 , 
 n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , n71461 , n71462 , n71463 , n71464 , 
 n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , n71471 , n71472 , n71473 , n71474 , 
 n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , n71481 , n71482 , n71483 , n71484 , 
 n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , n71491 , n71492 , n71493 , n71494 , 
 n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , n71501 , n71502 , n71503 , n71504 , 
 n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , n71511 , n71512 , n71513 , n71514 , 
 n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , n71521 , n71522 , n71523 , n71524 , 
 n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , n71531 , n71532 , n71533 , n71534 , 
 n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , n71541 , n71542 , n71543 , n71544 , 
 n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , n71551 , n71552 , n71553 , n71554 , 
 n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , n71561 , n71562 , n71563 , n71564 , 
 n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , 
 n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , n71581 , n71582 , n71583 , n71584 , 
 n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , 
 n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , n71601 , n71602 , n71603 , n71604 , 
 n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , n71611 , n71612 , n71613 , n71614 , 
 n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , n71621 , n71622 , n71623 , n71624 , 
 n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , n71631 , n71632 , n71633 , n71634 , 
 n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , n71641 , n71642 , n71643 , n71644 , 
 n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , n71651 , n71652 , n71653 , n71654 , 
 n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , 
 n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , n71671 , n71672 , n71673 , n71674 , 
 n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , n71681 , n71682 , n71683 , n71684 , 
 n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , n71691 , n71692 , n71693 , n71694 , 
 n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , n71701 , n71702 , n71703 , n71704 , 
 n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , n71711 , n71712 , n71713 , n71714 , 
 n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , n71721 , n71722 , n71723 , n71724 , 
 n71725 , n71726 , n71727 , n71728 , n71729 , n71730 , n71731 , n71732 , n71733 , n71734 , 
 n71735 , n71736 , n71737 , n71738 , n71739 , n71740 , n71741 , n71742 , n71743 , n71744 , 
 n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , n71751 , n71752 , n71753 , n71754 , 
 n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , n71761 , n71762 , n71763 , n71764 , 
 n71765 , n71766 , n71767 , n71768 , n71769 , n71770 , n71771 , n71772 , n71773 , n71774 , 
 n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , n71781 , n71782 , n71783 , n71784 , 
 n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , n71791 , n71792 , n71793 , n71794 , 
 n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , n71801 , n71802 , n71803 , n71804 , 
 n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , n71811 , n71812 , n71813 , n71814 , 
 n71815 , n71816 , n71817 , n71818 , n71819 , n71820 , n71821 , n71822 , n71823 , n71824 , 
 n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , n71831 , n71832 , n71833 , n71834 , 
 n71835 , n71836 , n71837 , n71838 , n71839 , n71840 , n71841 , n71842 , n71843 , n71844 , 
 n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , n71851 , n71852 , n71853 , n71854 , 
 n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , n71861 , n71862 , n71863 , n71864 , 
 n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , n71871 , n71872 , n71873 , n71874 , 
 n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , n71881 , n71882 , n71883 , n71884 , 
 n71885 , n71886 , n71887 , n71888 , n71889 , n71890 , n71891 , n71892 , n71893 , n71894 , 
 n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , n71901 , n71902 , n71903 , n71904 , 
 n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , n71911 , n71912 , n71913 , n71914 , 
 n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , 
 n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , n71931 , n71932 , n71933 , n71934 , 
 n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , 
 n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , 
 n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , 
 n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , 
 n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , n71981 , n71982 , n71983 , n71984 , 
 n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , n71991 , n71992 , n71993 , n71994 , 
 n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , n72001 , n72002 , n72003 , n72004 , 
 n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , n72011 , n72012 , n72013 , n72014 , 
 n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , 
 n72025 , n72026 , n72027 , n72028 , n72029 , n72030 , n72031 , n72032 , n72033 , n72034 , 
 n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , n72041 , n72042 , n72043 , n72044 , 
 n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , n72051 , n72052 , n72053 , n72054 , 
 n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , n72061 , n72062 , n72063 , n72064 , 
 n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , n72071 , n72072 , n72073 , n72074 , 
 n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , n72081 , n72082 , n72083 , n72084 , 
 n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , n72091 , n72092 , n72093 , n72094 , 
 n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , n72101 , n72102 , n72103 , n72104 , 
 n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , n72111 , n72112 , n72113 , n72114 , 
 n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , n72121 , n72122 , n72123 , n72124 , 
 n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , n72131 , n72132 , n72133 , n72134 , 
 n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , n72141 , n72142 , n72143 , n72144 , 
 n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , n72151 , n72152 , n72153 , n72154 , 
 n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , n72161 , n72162 , n72163 , n72164 , 
 n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , n72171 , n72172 , n72173 , n72174 , 
 n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , n72181 , n72182 , n72183 , n72184 , 
 n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , n72191 , n72192 , n72193 , n72194 , 
 n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , n72201 , n72202 , n72203 , n72204 , 
 n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , n72211 , n72212 , n72213 , n72214 , 
 n72215 , n72216 , n72217 , n72218 , n72219 , n72220 , n72221 , n72222 , n72223 , n72224 , 
 n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , n72231 , n72232 , n72233 , n72234 , 
 n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , n72241 , n72242 , n72243 , n72244 , 
 n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , n72251 , n72252 , n72253 , n72254 , 
 n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , n72261 , n72262 , n72263 , n72264 , 
 n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , n72271 , n72272 , n72273 , n72274 , 
 n72275 , n72276 , n72277 , n72278 , n72279 , n72280 , n72281 , n72282 , n72283 , n72284 , 
 n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , n72291 , n72292 , n72293 , n72294 , 
 n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , n72301 , n72302 , n72303 , n72304 , 
 n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , n72311 , n72312 , n72313 , n72314 , 
 n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , n72321 , n72322 , n72323 , n72324 , 
 n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , n72331 , n72332 , n72333 , n72334 , 
 n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , n72341 , n72342 , n72343 , n72344 , 
 n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , n72351 , n72352 , n72353 , n72354 , 
 n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , n72361 , n72362 , n72363 , n72364 , 
 n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , n72371 , n72372 , n72373 , n72374 , 
 n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , n72381 , n72382 , n72383 , n72384 , 
 n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , n72391 , n72392 , n72393 , n72394 , 
 n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , n72401 , n72402 , n72403 , n72404 , 
 n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , n72411 , n72412 , n72413 , n72414 , 
 n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , n72421 , n72422 , n72423 , n72424 , 
 n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , n72431 , n72432 , n72433 , n72434 , 
 n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , n72441 , n72442 , n72443 , n72444 , 
 n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , n72451 , n72452 , n72453 , n72454 , 
 n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , n72461 , n72462 , n72463 , n72464 , 
 n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , n72471 , n72472 , n72473 , n72474 , 
 n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , n72481 , n72482 , n72483 , n72484 , 
 n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , n72491 , n72492 , n72493 , n72494 , 
 n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , n72501 , n72502 , n72503 , n72504 , 
 n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , n72511 , n72512 , n72513 , n72514 , 
 n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , n72521 , n72522 , n72523 , n72524 , 
 n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , n72531 , n72532 , n72533 , n72534 , 
 n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , n72541 , n72542 , n72543 , n72544 , 
 n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , n72551 , n72552 , n72553 , n72554 , 
 n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , n72561 , n72562 , n72563 , n72564 , 
 n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , n72571 , n72572 , n72573 , n72574 , 
 n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , 
 n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , n72591 , n72592 , n72593 , n72594 , 
 n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , n72601 , n72602 , n72603 , n72604 , 
 n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , n72611 , n72612 , n72613 , n72614 , 
 n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , n72621 , n72622 , n72623 , n72624 , 
 n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , n72631 , n72632 , n72633 , n72634 , 
 n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , 
 n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , n72651 , n72652 , n72653 , n72654 , 
 n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , n72661 , n72662 , n72663 , n72664 , 
 n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , n72671 , n72672 , n72673 , n72674 , 
 n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , n72681 , n72682 , n72683 , n72684 , 
 n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , n72691 , n72692 , n72693 , n72694 , 
 n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , n72701 , n72702 , n72703 , n72704 , 
 n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , n72711 , n72712 , n72713 , n72714 , 
 n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , n72721 , n72722 , n72723 , n72724 , 
 n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , n72731 , n72732 , n72733 , n72734 , 
 n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , n72741 , n72742 , n72743 , n72744 , 
 n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , n72751 , n72752 , n72753 , n72754 , 
 n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , n72761 , n72762 , n72763 , n72764 , 
 n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , n72771 , n72772 , n72773 , n72774 , 
 n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , n72781 , n72782 , n72783 , n72784 , 
 n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , n72791 , n72792 , n72793 , n72794 , 
 n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , n72801 , n72802 , n72803 , n72804 , 
 n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , n72811 , n72812 , n72813 , n72814 , 
 n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , n72821 , n72822 , n72823 , n72824 , 
 n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , n72831 , n72832 , n72833 , n72834 , 
 n72835 , n72836 , n72837 , n72838 , n72839 , n72840 , n72841 , n72842 , n72843 , n72844 , 
 n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , n72851 , n72852 , n72853 , n72854 , 
 n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , n72861 , n72862 , n72863 , n72864 , 
 n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , n72871 , n72872 , n72873 , n72874 , 
 n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , n72881 , n72882 , n72883 , n72884 , 
 n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , 
 n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , n72901 , n72902 , n72903 , n72904 , 
 n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , n72911 , n72912 , n72913 , n72914 , 
 n72915 , n72916 , n72917 , n72918 , n72919 , n72920 , n72921 , n72922 , n72923 , n72924 , 
 n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , n72931 , n72932 , n72933 , n72934 , 
 n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , n72941 , n72942 , n72943 , n72944 , 
 n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , n72951 , n72952 , n72953 , n72954 , 
 n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , n72961 , n72962 , n72963 , n72964 , 
 n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , n72971 , n72972 , n72973 , n72974 , 
 n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , 
 n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , n72991 , n72992 , n72993 , n72994 , 
 n72995 , n72996 , n72997 , n72998 , n72999 , n73000 , n73001 , n73002 , n73003 , n73004 , 
 n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , n73011 , n73012 , n73013 , n73014 , 
 n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , n73021 , n73022 , n73023 , n73024 , 
 n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , 
 n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , n73041 , n73042 , n73043 , n73044 , 
 n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , 
 n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , n73061 , n73062 , n73063 , n73064 , 
 n73065 , n73066 , n73067 , n73068 , n73069 , n73070 , n73071 , n73072 , n73073 , n73074 , 
 n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , n73081 , n73082 , n73083 , n73084 , 
 n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , n73091 , n73092 , n73093 , n73094 , 
 n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , n73101 , n73102 , n73103 , n73104 , 
 n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , n73111 , n73112 , n73113 , n73114 , 
 n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , n73121 , n73122 , n73123 , n73124 , 
 n73125 , n73126 , n73127 , n73128 , n73129 , n73130 , n73131 , n73132 , n73133 , n73134 , 
 n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , n73141 , n73142 , n73143 , n73144 , 
 n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , n73151 , n73152 , n73153 , n73154 , 
 n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , 
 n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , n73171 , n73172 , n73173 , n73174 , 
 n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , n73181 , n73182 , n73183 , n73184 , 
 n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , n73191 , n73192 , n73193 , n73194 , 
 n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , n73201 , n73202 , n73203 , n73204 , 
 n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , n73211 , n73212 , n73213 , n73214 , 
 n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , n73221 , n73222 , n73223 , n73224 , 
 n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , n73231 , n73232 , n73233 , n73234 , 
 n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , n73241 , n73242 , n73243 , n73244 , 
 n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , n73251 , n73252 , n73253 , n73254 , 
 n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , 
 n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , n73271 , n73272 , n73273 , n73274 , 
 n73275 , n73276 , n73277 , n73278 , n73279 , n73280 , n73281 , n73282 , n73283 , n73284 , 
 n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , n73291 , n73292 , n73293 , n73294 , 
 n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , n73301 , n73302 , n73303 , n73304 , 
 n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , n73311 , n73312 , n73313 , n73314 , 
 n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , n73321 , n73322 , n73323 , n73324 , 
 n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , n73331 , n73332 , n73333 , n73334 , 
 n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , n73341 , n73342 , n73343 , n73344 , 
 n73345 , n73346 , n73347 , n73348 , n73349 , n73350 , n73351 , n73352 , n73353 , n73354 , 
 n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , n73361 , n73362 , n73363 , n73364 , 
 n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , n73371 , n73372 , n73373 , n73374 , 
 n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , n73381 , n73382 , n73383 , n73384 , 
 n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , n73391 , n73392 , n73393 , n73394 , 
 n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , n73401 , n73402 , n73403 , n73404 , 
 n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , n73411 , n73412 , n73413 , n73414 , 
 n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , n73421 , n73422 , n73423 , n73424 , 
 n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , n73431 , n73432 , n73433 , n73434 , 
 n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , n73441 , n73442 , n73443 , n73444 , 
 n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , n73451 , n73452 , n73453 , n73454 , 
 n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , n73461 , n73462 , n73463 , n73464 , 
 n73465 , n73466 , n73467 , n73468 , n73469 , n73470 , n73471 , n73472 , n73473 , n73474 , 
 n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , n73481 , n73482 , n73483 , n73484 , 
 n73485 , n73486 , n73487 , n73488 , n73489 , n73490 , n73491 , n73492 , n73493 , n73494 , 
 n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , n73501 , n73502 , n73503 , n73504 , 
 n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , n73511 , n73512 , n73513 , n73514 , 
 n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , n73521 , n73522 , n73523 , n73524 , 
 n73525 , n73526 , n73527 , n73528 , n73529 , n73530 , n73531 , n73532 , n73533 , n73534 , 
 n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , n73541 , n73542 , n73543 , n73544 , 
 n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , n73551 , n73552 , n73553 , n73554 , 
 n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , n73561 , n73562 , n73563 , n73564 , 
 n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , n73571 , n73572 , n73573 , n73574 , 
 n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , n73581 , n73582 , n73583 , n73584 , 
 n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , n73591 , n73592 , n73593 , n73594 , 
 n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , n73601 , n73602 , n73603 , n73604 , 
 n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , n73611 , n73612 , n73613 , n73614 , 
 n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , n73621 , n73622 , n73623 , n73624 , 
 n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , n73631 , n73632 , n73633 , n73634 , 
 n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , n73641 , n73642 , n73643 , n73644 , 
 n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , n73651 , n73652 , n73653 , n73654 , 
 n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , n73661 , n73662 , n73663 , n73664 , 
 n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , n73671 , n73672 , n73673 , n73674 , 
 n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , n73681 , n73682 , n73683 , n73684 , 
 n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , n73691 , n73692 , n73693 , n73694 , 
 n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , n73701 , n73702 , n73703 , n73704 , 
 n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , n73711 , n73712 , n73713 , n73714 , 
 n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , n73721 , n73722 , n73723 , n73724 , 
 n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , n73731 , n73732 , n73733 , n73734 , 
 n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , n73741 , n73742 , n73743 , n73744 , 
 n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , n73751 , n73752 , n73753 , n73754 , 
 n73755 , n73756 , n73757 , n73758 , n73759 , n73760 , n73761 , n73762 , n73763 , n73764 , 
 n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , n73771 , n73772 , n73773 , n73774 , 
 n73775 , n73776 , n73777 , n73778 , n73779 , n73780 , n73781 , n73782 , n73783 , n73784 , 
 n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , n73791 , n73792 , n73793 , n73794 , 
 n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , n73801 , n73802 , n73803 , n73804 , 
 n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , n73811 , n73812 , n73813 , n73814 , 
 n73815 , n73816 , n73817 , n73818 , n73819 , n73820 , n73821 , n73822 , n73823 , n73824 , 
 n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , n73831 , n73832 , n73833 , n73834 , 
 n73835 , n73836 , n73837 , n73838 , n73839 , n73840 , n73841 , n73842 , n73843 , n73844 , 
 n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , n73851 , n73852 , n73853 , n73854 , 
 n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , n73861 , n73862 , n73863 , n73864 , 
 n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , n73871 , n73872 , n73873 , n73874 , 
 n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , n73881 , n73882 , n73883 , n73884 , 
 n73885 , n73886 , n73887 , n73888 , n73889 , n73890 , n73891 , n73892 , n73893 , n73894 , 
 n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , n73901 , n73902 , n73903 , n73904 , 
 n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , n73911 , n73912 , n73913 , n73914 , 
 n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , n73921 , n73922 , n73923 , n73924 , 
 n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , n73931 , n73932 , n73933 , n73934 , 
 n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , n73941 , n73942 , n73943 , n73944 , 
 n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , n73951 , n73952 , n73953 , n73954 , 
 n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , n73961 , n73962 , n73963 , n73964 , 
 n73965 , n73966 , n73967 , n73968 , n73969 , n73970 , n73971 , n73972 , n73973 , n73974 , 
 n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , n73981 , n73982 , n73983 , n73984 , 
 n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , n73991 , n73992 , n73993 , n73994 , 
 n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , n74001 , n74002 , n74003 , n74004 , 
 n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , n74011 , n74012 , n74013 , n74014 , 
 n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , n74021 , n74022 , n74023 , n74024 , 
 n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , n74031 , n74032 , n74033 , n74034 , 
 n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , n74041 , n74042 , n74043 , n74044 , 
 n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , n74051 , n74052 , n74053 , n74054 , 
 n74055 , n74056 , n74057 , n74058 , n74059 , n74060 , n74061 , n74062 , n74063 , n74064 , 
 n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , n74071 , n74072 , n74073 , n74074 , 
 n74075 , n74076 , n74077 , n74078 , n74079 , n74080 , n74081 , n74082 , n74083 , n74084 , 
 n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , n74091 , n74092 , n74093 , n74094 , 
 n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , n74101 , n74102 , n74103 , n74104 , 
 n74105 , n74106 , n74107 , n74108 , n74109 , n74110 , n74111 , n74112 , n74113 , n74114 , 
 n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , n74121 , n74122 , n74123 , n74124 , 
 n74125 , n74126 , n74127 , n74128 , n74129 , n74130 , n74131 , n74132 , n74133 , n74134 , 
 n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , n74141 , n74142 , n74143 , n74144 , 
 n74145 , n74146 , n74147 , n74148 , n74149 , n74150 , n74151 , n74152 , n74153 , n74154 , 
 n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , n74161 , n74162 , n74163 , n74164 , 
 n74165 , n74166 , n74167 , n74168 , n74169 , n74170 , n74171 , n74172 , n74173 , n74174 , 
 n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , n74181 , n74182 , n74183 , n74184 , 
 n74185 , n74186 , n74187 , n74188 , n74189 , n74190 , n74191 , n74192 , n74193 , n74194 , 
 n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , n74201 , n74202 , n74203 , n74204 , 
 n74205 , n74206 , n74207 , n74208 , n74209 , n74210 , n74211 , n74212 , n74213 , n74214 , 
 n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , n74221 , n74222 , n74223 , n74224 , 
 n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , n74231 , n74232 , n74233 , n74234 , 
 n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , n74241 , n74242 , n74243 , n74244 , 
 n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , 
 n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , n74261 , n74262 , n74263 , n74264 , 
 n74265 , n74266 , n74267 , n74268 , n74269 , n74270 , n74271 , n74272 , n74273 , n74274 , 
 n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , n74281 , n74282 , n74283 , n74284 , 
 n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , n74291 , n74292 , n74293 , n74294 , 
 n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , n74301 , n74302 , n74303 , n74304 , 
 n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , n74311 , n74312 , n74313 , n74314 , 
 n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , n74321 , n74322 , n74323 , n74324 , 
 n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , n74331 , n74332 , n74333 , n74334 , 
 n74335 , n74336 , n74337 , n74338 , n74339 , n74340 , n74341 , n74342 , n74343 , n74344 , 
 n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , n74351 , n74352 , n74353 , n74354 , 
 n74355 , n74356 , n74357 , n74358 , n74359 , n74360 , n74361 , n74362 , n74363 , n74364 , 
 n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , n74371 , n74372 , n74373 , n74374 , 
 n74375 , n74376 , n74377 , n74378 , n74379 , n74380 , n74381 , n74382 , n74383 , n74384 , 
 n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , n74391 , n74392 , n74393 , n74394 , 
 n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , n74401 , n74402 , n74403 , n74404 , 
 n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , n74411 , n74412 , n74413 , n74414 , 
 n74415 , n74416 , n74417 , n74418 , n74419 , n74420 , n74421 , n74422 , n74423 , n74424 , 
 n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , n74431 , n74432 , n74433 , n74434 , 
 n74435 , n74436 , n74437 , n74438 , n74439 , n74440 , n74441 , n74442 , n74443 , n74444 , 
 n74445 , n74446 , n74447 , n74448 , n74449 , n74450 , n74451 , n74452 , n74453 , n74454 , 
 n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , n74461 , n74462 , n74463 , n74464 , 
 n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , n74471 , n74472 , n74473 , n74474 , 
 n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , n74481 , n74482 , n74483 , n74484 , 
 n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , n74491 , n74492 , n74493 , n74494 , 
 n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , n74501 , n74502 , n74503 , n74504 , 
 n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , n74511 , n74512 , n74513 , n74514 , 
 n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , n74521 , n74522 , n74523 , n74524 , 
 n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , n74531 , n74532 , n74533 , n74534 , 
 n74535 , n74536 , n74537 , n74538 , n74539 , n74540 , n74541 , n74542 , n74543 , n74544 , 
 n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , n74551 , n74552 , n74553 , n74554 , 
 n74555 , n74556 , n74557 , n74558 , n74559 , n74560 , n74561 , n74562 , n74563 , n74564 , 
 n74565 , n74566 , n74567 , n74568 , n74569 , n74570 , n74571 , n74572 , n74573 , n74574 , 
 n74575 , n74576 , n74577 , n74578 , n74579 , n74580 , n74581 , n74582 , n74583 , n74584 , 
 n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , n74591 , n74592 , n74593 , n74594 , 
 n74595 , n74596 , n74597 , n74598 , n74599 , n74600 , n74601 , n74602 , n74603 , n74604 , 
 n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , n74611 , n74612 , n74613 , n74614 , 
 n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , n74621 , n74622 , n74623 , n74624 , 
 n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , n74631 , n74632 , n74633 , n74634 , 
 n74635 , n74636 , n74637 , n74638 , n74639 , n74640 , n74641 , n74642 , n74643 , n74644 , 
 n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , n74651 , n74652 , n74653 , n74654 , 
 n74655 , n74656 , n74657 , n74658 , n74659 , n74660 , n74661 , n74662 , n74663 , n74664 , 
 n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , n74671 , n74672 , n74673 , n74674 , 
 n74675 , n74676 , n74677 , n74678 , n74679 , n74680 , n74681 , n74682 , n74683 , n74684 , 
 n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , n74691 , n74692 , n74693 , n74694 , 
 n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , n74701 , n74702 , n74703 , n74704 , 
 n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , n74711 , n74712 , n74713 , n74714 , 
 n74715 , n74716 , n74717 , n74718 , n74719 , n74720 , n74721 , n74722 , n74723 , n74724 , 
 n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , n74731 , n74732 , n74733 , n74734 , 
 n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , n74741 , n74742 , n74743 , n74744 , 
 n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , n74751 , n74752 , n74753 , n74754 , 
 n74755 , n74756 , n74757 , n74758 , n74759 , n74760 , n74761 , n74762 , n74763 , n74764 , 
 n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , n74771 , n74772 , n74773 , n74774 , 
 n74775 , n74776 , n74777 , n74778 , n74779 , n74780 , n74781 , n74782 , n74783 , n74784 , 
 n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , n74791 , n74792 , n74793 , n74794 , 
 n74795 , n74796 , n74797 , n74798 , n74799 , n74800 , n74801 , n74802 , n74803 , n74804 , 
 n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , n74811 , n74812 , n74813 , n74814 , 
 n74815 , n74816 , n74817 , n74818 , n74819 , n74820 , n74821 , n74822 , n74823 , n74824 , 
 n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , n74831 , n74832 , n74833 , n74834 , 
 n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , n74841 , n74842 , n74843 , n74844 , 
 n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , n74851 , n74852 , n74853 , n74854 , 
 n74855 , n74856 , n74857 , n74858 , n74859 , n74860 , n74861 , n74862 , n74863 , n74864 , 
 n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , n74871 , n74872 , n74873 , n74874 , 
 n74875 , n74876 , n74877 , n74878 , n74879 , n74880 , n74881 , n74882 , n74883 , n74884 , 
 n74885 , n74886 , n74887 , n74888 , n74889 , n74890 , n74891 , n74892 , n74893 , n74894 , 
 n74895 , n74896 , n74897 , n74898 , n74899 , n74900 , n74901 , n74902 , n74903 , n74904 , 
 n74905 , n74906 , n74907 , n74908 , n74909 , n74910 , n74911 , n74912 , n74913 , n74914 , 
 n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , n74921 , n74922 , n74923 , n74924 , 
 n74925 , n74926 , n74927 , n74928 , n74929 , n74930 , n74931 , n74932 , n74933 , n74934 , 
 n74935 , n74936 , n74937 , n74938 , n74939 , n74940 , n74941 , n74942 , n74943 , n74944 , 
 n74945 , n74946 , n74947 , n74948 , n74949 , n74950 , n74951 , n74952 , n74953 , n74954 , 
 n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , n74961 , n74962 , n74963 , n74964 , 
 n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , n74971 , n74972 , n74973 , n74974 , 
 n74975 , n74976 , n74977 , n74978 , n74979 , n74980 , n74981 , n74982 , n74983 , n74984 , 
 n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , n74991 , n74992 , n74993 , n74994 , 
 n74995 , n74996 , n74997 , n74998 , n74999 , n75000 , n75001 , n75002 , n75003 , n75004 , 
 n75005 , n75006 , n75007 , n75008 , n75009 , n75010 , n75011 , n75012 , n75013 , n75014 , 
 n75015 , n75016 , n75017 , n75018 , n75019 , n75020 , n75021 , n75022 , n75023 , n75024 , 
 n75025 , n75026 , n75027 , n75028 , n75029 , n75030 , n75031 , n75032 , n75033 , n75034 , 
 n75035 , n75036 , n75037 , n75038 , n75039 , n75040 , n75041 , n75042 , n75043 , n75044 , 
 n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , n75051 , n75052 , n75053 , n75054 , 
 n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , n75061 , n75062 , n75063 , n75064 , 
 n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , n75071 , n75072 , n75073 , n75074 , 
 n75075 , n75076 , n75077 , n75078 , n75079 , n75080 , n75081 , n75082 , n75083 , n75084 , 
 n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , n75091 , n75092 , n75093 , n75094 , 
 n75095 , n75096 , n75097 , n75098 , n75099 , n75100 , n75101 , n75102 , n75103 , n75104 , 
 n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , n75111 , n75112 , n75113 , n75114 , 
 n75115 , n75116 , n75117 , n75118 , n75119 , n75120 , n75121 , n75122 , n75123 , n75124 , 
 n75125 , n75126 , n75127 , n75128 , n75129 , n75130 , n75131 , n75132 , n75133 , n75134 , 
 n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , n75141 , n75142 , n75143 , n75144 , 
 n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , n75151 , n75152 , n75153 , n75154 , 
 n75155 , n75156 , n75157 , n75158 , n75159 , n75160 , n75161 , n75162 , n75163 , n75164 , 
 n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , n75171 , n75172 , n75173 , n75174 , 
 n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , n75181 , n75182 , n75183 , n75184 , 
 n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , n75191 , n75192 , n75193 , n75194 , 
 n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , n75201 , n75202 , n75203 , n75204 , 
 n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , n75211 , n75212 , n75213 , n75214 , 
 n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , n75221 , n75222 , n75223 , n75224 , 
 n75225 , n75226 , n75227 , n75228 , n75229 , n75230 , n75231 , n75232 , n75233 , n75234 , 
 n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , n75241 , n75242 , n75243 , n75244 , 
 n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , n75251 , n75252 , n75253 , n75254 , 
 n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , n75261 , n75262 , n75263 , n75264 , 
 n75265 , n75266 , n75267 , n75268 , n75269 , n75270 , n75271 , n75272 , n75273 , n75274 , 
 n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , n75281 , n75282 , n75283 , n75284 , 
 n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , n75291 , n75292 , n75293 , n75294 , 
 n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , n75301 , n75302 , n75303 , n75304 , 
 n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , n75311 , n75312 , n75313 , n75314 , 
 n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , n75321 , n75322 , n75323 , n75324 , 
 n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , n75331 , n75332 , n75333 , n75334 , 
 n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , n75341 , n75342 , n75343 , n75344 , 
 n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , n75351 , n75352 , n75353 , n75354 , 
 n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , n75361 , n75362 , n75363 , n75364 , 
 n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , n75371 , n75372 , n75373 , n75374 , 
 n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , n75381 , n75382 , n75383 , n75384 , 
 n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , n75391 , n75392 , n75393 , n75394 , 
 n75395 , n75396 , n75397 , n75398 , n75399 , n75400 , n75401 , n75402 , n75403 , n75404 , 
 n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , n75411 , n75412 , n75413 , n75414 , 
 n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , n75421 , n75422 , n75423 , n75424 , 
 n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , n75431 , n75432 , n75433 , n75434 , 
 n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , n75441 , n75442 , n75443 , n75444 , 
 n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , n75451 , n75452 , n75453 , n75454 , 
 n75455 , n75456 , n75457 , n75458 , n75459 , n75460 , n75461 , n75462 , n75463 , n75464 , 
 n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , n75471 , n75472 , n75473 , n75474 , 
 n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , n75481 , n75482 , n75483 , n75484 , 
 n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , n75491 , n75492 , n75493 , n75494 , 
 n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , n75501 , n75502 , n75503 , n75504 , 
 n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , n75511 , n75512 , n75513 , n75514 , 
 n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , n75521 , n75522 , n75523 , n75524 , 
 n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , n75531 , n75532 , n75533 , n75534 , 
 n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , n75541 , n75542 , n75543 , n75544 , 
 n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , n75551 , n75552 , n75553 , n75554 , 
 n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , n75561 , n75562 , n75563 , n75564 , 
 n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , n75571 , n75572 , n75573 , n75574 , 
 n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , n75581 , n75582 , n75583 , n75584 , 
 n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , n75591 , n75592 , n75593 , n75594 , 
 n75595 , n75596 , n75597 , n75598 , n75599 , n75600 , n75601 , n75602 , n75603 , n75604 , 
 n75605 , n75606 , n75607 , n75608 , n75609 , n75610 , n75611 , n75612 , n75613 , n75614 , 
 n75615 , n75616 , n75617 , n75618 , n75619 , n75620 , n75621 , n75622 , n75623 , n75624 , 
 n75625 , n75626 , n75627 , n75628 , n75629 , n75630 , n75631 , n75632 , n75633 , n75634 , 
 n75635 , n75636 , n75637 , n75638 , n75639 , n75640 , n75641 , n75642 , n75643 , n75644 , 
 n75645 , n75646 , n75647 , n75648 , n75649 , n75650 , n75651 , n75652 , n75653 , n75654 , 
 n75655 , n75656 , n75657 , n75658 , n75659 , n75660 , n75661 , n75662 , n75663 , n75664 , 
 n75665 , n75666 , n75667 , n75668 , n75669 , n75670 , n75671 , n75672 , n75673 , n75674 , 
 n75675 , n75676 , n75677 , n75678 , n75679 , n75680 , n75681 , n75682 , n75683 , n75684 , 
 n75685 , n75686 , n75687 , n75688 , n75689 , n75690 , n75691 , n75692 , n75693 , n75694 , 
 n75695 , n75696 , n75697 , n75698 , n75699 , n75700 , n75701 , n75702 , n75703 , n75704 , 
 n75705 , n75706 , n75707 , n75708 , n75709 , n75710 , n75711 , n75712 , n75713 , n75714 , 
 n75715 , n75716 , n75717 , n75718 , n75719 , n75720 , n75721 , n75722 , n75723 , n75724 , 
 n75725 , n75726 , n75727 , n75728 , n75729 , n75730 , n75731 , n75732 , n75733 , n75734 , 
 n75735 , n75736 , n75737 , n75738 , n75739 , n75740 , n75741 , n75742 , n75743 , n75744 , 
 n75745 , n75746 , n75747 , n75748 , n75749 , n75750 , n75751 , n75752 , n75753 , n75754 , 
 n75755 , n75756 , n75757 , n75758 , n75759 , n75760 , n75761 , n75762 , n75763 , n75764 , 
 n75765 , n75766 , n75767 , n75768 , n75769 , n75770 , n75771 , n75772 , n75773 , n75774 , 
 n75775 , n75776 , n75777 , n75778 , n75779 , n75780 , n75781 , n75782 , n75783 , n75784 , 
 n75785 , n75786 , n75787 , n75788 , n75789 , n75790 , n75791 , n75792 , n75793 , n75794 , 
 n75795 , n75796 , n75797 , n75798 , n75799 , n75800 , n75801 , n75802 , n75803 , n75804 , 
 n75805 , n75806 , n75807 , n75808 , n75809 , n75810 , n75811 , n75812 , n75813 , n75814 , 
 n75815 , n75816 , n75817 , n75818 , n75819 , n75820 , n75821 , n75822 , n75823 , n75824 , 
 n75825 , n75826 , n75827 , n75828 , n75829 , n75830 , n75831 , n75832 , n75833 , n75834 , 
 n75835 , n75836 , n75837 , n75838 , n75839 , n75840 , n75841 , n75842 , n75843 , n75844 , 
 n75845 , n75846 , n75847 , n75848 , n75849 , n75850 , n75851 , n75852 , n75853 , n75854 , 
 n75855 , n75856 , n75857 , n75858 , n75859 , n75860 , n75861 , n75862 , n75863 , n75864 , 
 n75865 , n75866 , n75867 , n75868 , n75869 , n75870 , n75871 , n75872 , n75873 , n75874 , 
 n75875 , n75876 , n75877 , n75878 , n75879 , n75880 , n75881 , n75882 , n75883 , n75884 , 
 n75885 , n75886 , n75887 , n75888 , n75889 , n75890 , n75891 , n75892 , n75893 , n75894 , 
 n75895 , n75896 , n75897 , n75898 , n75899 , n75900 , n75901 , n75902 , n75903 , n75904 , 
 n75905 , n75906 , n75907 , n75908 , n75909 , n75910 , n75911 , n75912 , n75913 , n75914 , 
 n75915 , n75916 , n75917 , n75918 , n75919 , n75920 , n75921 , n75922 , n75923 , n75924 , 
 n75925 , n75926 , n75927 , n75928 , n75929 , n75930 , n75931 , n75932 , n75933 , n75934 , 
 n75935 , n75936 , n75937 , n75938 , n75939 , n75940 , n75941 , n75942 , n75943 , n75944 , 
 n75945 , n75946 , n75947 , n75948 , n75949 , n75950 , n75951 , n75952 , n75953 , n75954 , 
 n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , 
 n75965 , n75966 , n75967 , n75968 , n75969 , n75970 , n75971 , n75972 , n75973 , n75974 , 
 n75975 , n75976 , n75977 , n75978 , n75979 , n75980 , n75981 , n75982 , n75983 , n75984 , 
 n75985 , n75986 , n75987 , n75988 , n75989 , n75990 , n75991 , n75992 , n75993 , n75994 , 
 n75995 , n75996 , n75997 , n75998 , n75999 , n76000 , n76001 , n76002 , n76003 , n76004 , 
 n76005 , n76006 , n76007 , n76008 , n76009 , n76010 , n76011 , n76012 , n76013 , n76014 , 
 n76015 , n76016 , n76017 , n76018 , n76019 , n76020 , n76021 , n76022 , n76023 , n76024 , 
 n76025 , n76026 , n76027 , n76028 , n76029 , n76030 , n76031 , n76032 , n76033 , n76034 , 
 n76035 , n76036 , n76037 , n76038 , n76039 , n76040 , n76041 , n76042 , n76043 , n76044 , 
 n76045 , n76046 , n76047 , n76048 , n76049 , n76050 , n76051 , n76052 , n76053 , n76054 , 
 n76055 , n76056 , n76057 , n76058 , n76059 , n76060 , n76061 , n76062 , n76063 , n76064 , 
 n76065 , n76066 , n76067 , n76068 , n76069 , n76070 , n76071 , n76072 , n76073 , n76074 , 
 n76075 , n76076 , n76077 , n76078 , n76079 , n76080 , n76081 , n76082 , n76083 , n76084 , 
 n76085 , n76086 , n76087 , n76088 , n76089 , n76090 , n76091 , n76092 , n76093 , n76094 , 
 n76095 , n76096 , n76097 , n76098 , n76099 , n76100 , n76101 , n76102 , n76103 , n76104 , 
 n76105 , n76106 , n76107 , n76108 , n76109 , n76110 , n76111 , n76112 , n76113 , n76114 , 
 n76115 , n76116 , n76117 , n76118 , n76119 , n76120 , n76121 , n76122 , n76123 , n76124 , 
 n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , 
 n76135 , n76136 , n76137 , n76138 , n76139 , n76140 , n76141 , n76142 , n76143 , n76144 , 
 n76145 , n76146 , n76147 , n76148 , n76149 , n76150 , n76151 , n76152 , n76153 , n76154 , 
 n76155 , n76156 , n76157 , n76158 , n76159 , n76160 , n76161 , n76162 , n76163 , n76164 , 
 n76165 , n76166 , n76167 , n76168 , n76169 , n76170 , n76171 , n76172 , n76173 , n76174 , 
 n76175 , n76176 , n76177 , n76178 , n76179 , n76180 , n76181 , n76182 , n76183 , n76184 , 
 n76185 , n76186 , n76187 , n76188 , n76189 , n76190 , n76191 , n76192 , n76193 , n76194 , 
 n76195 , n76196 , n76197 , n76198 , n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , 
 n76205 , n76206 , n76207 , n76208 , n76209 , n76210 , n76211 , n76212 , n76213 , n76214 , 
 n76215 , n76216 , n76217 , n76218 , n76219 , n76220 , n76221 , n76222 , n76223 , n76224 , 
 n76225 , n76226 , n76227 , n76228 , n76229 , n76230 , n76231 , n76232 , n76233 , n76234 , 
 n76235 , n76236 , n76237 , n76238 , n76239 , n76240 , n76241 , n76242 , n76243 , n76244 , 
 n76245 , n76246 , n76247 , n76248 , n76249 , n76250 , n76251 , n76252 , n76253 , n76254 , 
 n76255 , n76256 , n76257 , n76258 , n76259 , n76260 , n76261 , n76262 , n76263 , n76264 , 
 n76265 , n76266 , n76267 , n76268 , n76269 , n76270 , n76271 , n76272 , n76273 , n76274 , 
 n76275 , n76276 , n76277 , n76278 , n76279 , n76280 , n76281 , n76282 , n76283 , n76284 , 
 n76285 , n76286 , n76287 , n76288 , n76289 , n76290 , n76291 , n76292 , n76293 , n76294 , 
 n76295 , n76296 , n76297 , n76298 , n76299 , n76300 , n76301 , n76302 , n76303 , n76304 , 
 n76305 , n76306 , n76307 , n76308 , n76309 , n76310 , n76311 , n76312 , n76313 , n76314 , 
 n76315 , n76316 , n76317 , n76318 , n76319 , n76320 , n76321 , n76322 , n76323 , n76324 , 
 n76325 , n76326 , n76327 , n76328 , n76329 , n76330 , n76331 , n76332 , n76333 , n76334 , 
 n76335 , n76336 , n76337 , n76338 , n76339 , n76340 , n76341 , n76342 , n76343 , n76344 , 
 n76345 , n76346 , n76347 , n76348 , n76349 , n76350 , n76351 , n76352 , n76353 , n76354 , 
 n76355 , n76356 , n76357 , n76358 , n76359 , n76360 , n76361 , n76362 , n76363 , n76364 , 
 n76365 , n76366 , n76367 , n76368 , n76369 , n76370 , n76371 , n76372 , n76373 , n76374 , 
 n76375 , n76376 , n76377 , n76378 , n76379 , n76380 , n76381 , n76382 , n76383 , n76384 , 
 n76385 , n76386 , n76387 , n76388 , n76389 , n76390 , n76391 , n76392 , n76393 , n76394 , 
 n76395 , n76396 , n76397 , n76398 , n76399 , n76400 , n76401 , n76402 , n76403 , n76404 , 
 n76405 , n76406 , n76407 , n76408 , n76409 , n76410 , n76411 , n76412 , n76413 , n76414 , 
 n76415 , n76416 , n76417 , n76418 , n76419 , n76420 , n76421 , n76422 , n76423 , n76424 , 
 n76425 , n76426 , n76427 , n76428 , n76429 , n76430 , n76431 , n76432 , n76433 , n76434 , 
 n76435 , n76436 , n76437 , n76438 , n76439 , n76440 , n76441 , n76442 , n76443 , n76444 , 
 n76445 , n76446 , n76447 , n76448 , n76449 , n76450 , n76451 , n76452 , n76453 , n76454 , 
 n76455 , n76456 , n76457 , n76458 , n76459 , n76460 , n76461 , n76462 , n76463 , n76464 , 
 n76465 , n76466 , n76467 , n76468 , n76469 , n76470 , n76471 , n76472 , n76473 , n76474 , 
 n76475 , n76476 , n76477 , n76478 , n76479 , n76480 , n76481 , n76482 , n76483 , n76484 , 
 n76485 , n76486 , n76487 , n76488 , n76489 , n76490 , n76491 , n76492 , n76493 , n76494 , 
 n76495 , n76496 , n76497 , n76498 , n76499 , n76500 , n76501 , n76502 , n76503 , n76504 , 
 n76505 , n76506 , n76507 , n76508 , n76509 , n76510 , n76511 , n76512 , n76513 , n76514 , 
 n76515 , n76516 , n76517 , n76518 , n76519 , n76520 , n76521 , n76522 , n76523 , n76524 , 
 n76525 , n76526 , n76527 , n76528 , n76529 , n76530 , n76531 , n76532 , n76533 , n76534 , 
 n76535 , n76536 , n76537 , n76538 , n76539 , n76540 , n76541 , n76542 , n76543 , n76544 , 
 n76545 , n76546 , n76547 , n76548 , n76549 , n76550 , n76551 , n76552 , n76553 , n76554 , 
 n76555 , n76556 , n76557 , n76558 , n76559 , n76560 , n76561 , n76562 , n76563 , n76564 , 
 n76565 , n76566 , n76567 , n76568 , n76569 , n76570 , n76571 , n76572 , n76573 , n76574 , 
 n76575 , n76576 , n76577 , n76578 , n76579 , n76580 , n76581 , n76582 , n76583 , n76584 , 
 n76585 , n76586 , n76587 , n76588 , n76589 , n76590 , n76591 , n76592 , n76593 , n76594 , 
 n76595 , n76596 , n76597 , n76598 , n76599 , n76600 , n76601 , n76602 , n76603 , n76604 , 
 n76605 , n76606 , n76607 , n76608 , n76609 , n76610 , n76611 , n76612 , n76613 , n76614 , 
 n76615 , n76616 , n76617 , n76618 , n76619 , n76620 , n76621 , n76622 , n76623 , n76624 , 
 n76625 , n76626 , n76627 , n76628 , n76629 , n76630 , n76631 , n76632 , n76633 , n76634 , 
 n76635 , n76636 , n76637 , n76638 , n76639 , n76640 , n76641 , n76642 , n76643 , n76644 , 
 n76645 , n76646 , n76647 , n76648 , n76649 , n76650 , n76651 , n76652 , n76653 , n76654 , 
 n76655 , n76656 , n76657 , n76658 , n76659 , n76660 , n76661 , n76662 , n76663 , n76664 , 
 n76665 , n76666 , n76667 , n76668 , n76669 , n76670 , n76671 , n76672 , n76673 , n76674 , 
 n76675 , n76676 , n76677 , n76678 , n76679 , n76680 , n76681 , n76682 , n76683 , n76684 , 
 n76685 , n76686 , n76687 , n76688 , n76689 , n76690 , n76691 , n76692 , n76693 , n76694 , 
 n76695 , n76696 , n76697 , n76698 , n76699 , n76700 , n76701 , n76702 , n76703 , n76704 , 
 n76705 , n76706 , n76707 , n76708 , n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , 
 n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , n76721 , n76722 , n76723 , n76724 , 
 n76725 , n76726 , n76727 , n76728 , n76729 , n76730 , n76731 , n76732 , n76733 , n76734 , 
 n76735 , n76736 , n76737 , n76738 , n76739 , n76740 , n76741 , n76742 , n76743 , n76744 , 
 n76745 , n76746 , n76747 , n76748 , n76749 , n76750 , n76751 , n76752 , n76753 , n76754 , 
 n76755 , n76756 , n76757 , n76758 , n76759 , n76760 , n76761 , n76762 , n76763 , n76764 , 
 n76765 , n76766 , n76767 , n76768 , n76769 , n76770 , n76771 , n76772 , n76773 , n76774 , 
 n76775 , n76776 , n76777 , n76778 , n76779 , n76780 , n76781 , n76782 , n76783 , n76784 , 
 n76785 , n76786 , n76787 , n76788 , n76789 , n76790 , n76791 , n76792 , n76793 , n76794 , 
 n76795 , n76796 , n76797 , n76798 , n76799 , n76800 , n76801 , n76802 , n76803 , n76804 , 
 n76805 , n76806 , n76807 , n76808 , n76809 , n76810 , n76811 , n76812 , n76813 , n76814 , 
 n76815 , n76816 , n76817 , n76818 , n76819 , n76820 , n76821 , n76822 , n76823 , n76824 , 
 n76825 , n76826 , n76827 , n76828 , n76829 , n76830 , n76831 , n76832 , n76833 , n76834 , 
 n76835 , n76836 , n76837 , n76838 , n76839 , n76840 , n76841 , n76842 , n76843 , n76844 , 
 n76845 , n76846 , n76847 , n76848 , n76849 , n76850 , n76851 , n76852 , n76853 , n76854 , 
 n76855 , n76856 , n76857 , n76858 , n76859 , n76860 , n76861 , n76862 , n76863 , n76864 , 
 n76865 , n76866 , n76867 , n76868 , n76869 , n76870 , n76871 , n76872 , n76873 , n76874 , 
 n76875 , n76876 , n76877 , n76878 , n76879 , n76880 , n76881 , n76882 , n76883 , n76884 , 
 n76885 , n76886 , n76887 , n76888 , n76889 , n76890 , n76891 , n76892 , n76893 , n76894 , 
 n76895 , n76896 , n76897 , n76898 , n76899 , n76900 , n76901 , n76902 , n76903 , n76904 , 
 n76905 , n76906 , n76907 , n76908 , n76909 , n76910 , n76911 , n76912 , n76913 , n76914 , 
 n76915 , n76916 , n76917 , n76918 , n76919 , n76920 , n76921 , n76922 , n76923 , n76924 , 
 n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , n76931 , n76932 , n76933 , n76934 , 
 n76935 , n76936 , n76937 , n76938 , n76939 , n76940 , n76941 , n76942 , n76943 , n76944 , 
 n76945 , n76946 , n76947 , n76948 , n76949 , n76950 , n76951 , n76952 , n76953 , n76954 , 
 n76955 , n76956 , n76957 , n76958 , n76959 , n76960 , n76961 , n76962 , n76963 , n76964 , 
 n76965 , n76966 , n76967 , n76968 , n76969 , n76970 , n76971 , n76972 , n76973 , n76974 , 
 n76975 , n76976 , n76977 , n76978 , n76979 , n76980 , n76981 , n76982 , n76983 , n76984 , 
 n76985 , n76986 , n76987 , n76988 , n76989 , n76990 , n76991 , n76992 , n76993 , n76994 , 
 n76995 , n76996 , n76997 , n76998 , n76999 , n77000 , n77001 , n77002 , n77003 , n77004 , 
 n77005 , n77006 , n77007 , n77008 , n77009 , n77010 , n77011 , n77012 , n77013 , n77014 , 
 n77015 , n77016 , n77017 , n77018 , n77019 , n77020 , n77021 , n77022 , n77023 , n77024 , 
 n77025 , n77026 , n77027 , n77028 , n77029 , n77030 , n77031 , n77032 , n77033 , n77034 , 
 n77035 , n77036 , n77037 , n77038 , n77039 , n77040 , n77041 , n77042 , n77043 , n77044 , 
 n77045 , n77046 , n77047 , n77048 , n77049 , n77050 , n77051 , n77052 , n77053 , n77054 , 
 n77055 , n77056 , n77057 , n77058 , n77059 , n77060 , n77061 , n77062 , n77063 , n77064 , 
 n77065 , n77066 , n77067 , n77068 , n77069 , n77070 , n77071 , n77072 , n77073 , n77074 , 
 n77075 , n77076 , n77077 , n77078 , n77079 , n77080 , n77081 , n77082 , n77083 , n77084 , 
 n77085 , n77086 , n77087 , n77088 , n77089 , n77090 , n77091 , n77092 , n77093 , n77094 , 
 n77095 , n77096 , n77097 , n77098 , n77099 , n77100 , n77101 , n77102 , n77103 , n77104 , 
 n77105 , n77106 , n77107 , n77108 , n77109 , n77110 , n77111 , n77112 , n77113 , n77114 , 
 n77115 , n77116 , n77117 , n77118 , n77119 , n77120 , n77121 , n77122 , n77123 , n77124 , 
 n77125 , n77126 , n77127 , n77128 , n77129 , n77130 , n77131 , n77132 , n77133 , n77134 , 
 n77135 , n77136 , n77137 , n77138 , n77139 , n77140 , n77141 , n77142 , n77143 , n77144 , 
 n77145 , n77146 , n77147 , n77148 , n77149 , n77150 , n77151 , n77152 , n77153 , n77154 , 
 n77155 , n77156 , n77157 , n77158 , n77159 , n77160 , n77161 , n77162 , n77163 , n77164 , 
 n77165 , n77166 , n77167 , n77168 , n77169 , n77170 , n77171 , n77172 , n77173 , n77174 , 
 n77175 , n77176 , n77177 , n77178 , n77179 , n77180 , n77181 , n77182 , n77183 , n77184 , 
 n77185 , n77186 , n77187 , n77188 , n77189 , n77190 , n77191 , n77192 , n77193 , n77194 , 
 n77195 , n77196 , n77197 , n77198 , n77199 , n77200 , n77201 , n77202 , n77203 , n77204 , 
 n77205 , n77206 , n77207 , n77208 , n77209 , n77210 , n77211 , n77212 , n77213 , n77214 , 
 n77215 , n77216 , n77217 , n77218 , n77219 , n77220 , n77221 , n77222 , n77223 , n77224 , 
 n77225 , n77226 , n77227 , n77228 , n77229 , n77230 , n77231 , n77232 , n77233 , n77234 , 
 n77235 , n77236 , n77237 , n77238 , n77239 , n77240 , n77241 , n77242 , n77243 , n77244 , 
 n77245 , n77246 , n77247 , n77248 , n77249 , n77250 , n77251 , n77252 , n77253 , n77254 , 
 n77255 , n77256 , n77257 , n77258 , n77259 , n77260 , n77261 , n77262 , n77263 , n77264 , 
 n77265 , n77266 , n77267 , n77268 , n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , 
 n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , n77281 , n77282 , n77283 , n77284 , 
 n77285 , n77286 , n77287 , n77288 , n77289 , n77290 , n77291 , n77292 , n77293 , n77294 , 
 n77295 , n77296 , n77297 , n77298 , n77299 , n77300 , n77301 , n77302 , n77303 , n77304 , 
 n77305 , n77306 , n77307 , n77308 , n77309 , n77310 , n77311 , n77312 , n77313 , n77314 , 
 n77315 , n77316 , n77317 , n77318 , n77319 , n77320 , n77321 , n77322 , n77323 , n77324 , 
 n77325 , n77326 , n77327 , n77328 , n77329 , n77330 , n77331 , n77332 , n77333 , n77334 , 
 n77335 , n77336 , n77337 , n77338 , n77339 , n77340 , n77341 , n77342 , n77343 , n77344 , 
 n77345 , n77346 , n77347 , n77348 , n77349 , n77350 , n77351 , n77352 , n77353 , n77354 , 
 n77355 , n77356 , n77357 , n77358 , n77359 , n77360 , n77361 , n77362 , n77363 , n77364 , 
 n77365 , n77366 , n77367 , n77368 , n77369 , n77370 , n77371 , n77372 , n77373 , n77374 , 
 n77375 , n77376 , n77377 , n77378 , n77379 , n77380 , n77381 , n77382 , n77383 , n77384 , 
 n77385 , n77386 , n77387 , n77388 , n77389 , n77390 , n77391 , n77392 , n77393 , n77394 , 
 n77395 , n77396 , n77397 , n77398 , n77399 , n77400 , n77401 , n77402 , n77403 , n77404 , 
 n77405 , n77406 , n77407 , n77408 , n77409 , n77410 , n77411 , n77412 , n77413 , n77414 , 
 n77415 , n77416 , n77417 , n77418 , n77419 , n77420 , n77421 , n77422 , n77423 , n77424 , 
 n77425 , n77426 , n77427 , n77428 , n77429 , n77430 , n77431 , n77432 , n77433 , n77434 , 
 n77435 , n77436 , n77437 , n77438 , n77439 , n77440 , n77441 , n77442 , n77443 , n77444 , 
 n77445 , n77446 , n77447 , n77448 , n77449 , n77450 , n77451 , n77452 , n77453 , n77454 , 
 n77455 , n77456 , n77457 , n77458 , n77459 , n77460 , n77461 , n77462 , n77463 , n77464 , 
 n77465 , n77466 , n77467 , n77468 , n77469 , n77470 , n77471 , n77472 , n77473 , n77474 , 
 n77475 , n77476 , n77477 , n77478 , n77479 , n77480 , n77481 , n77482 , n77483 , n77484 , 
 n77485 , n77486 , n77487 , n77488 , n77489 , n77490 , n77491 , n77492 , n77493 , n77494 , 
 n77495 , n77496 , n77497 , n77498 , n77499 , n77500 , n77501 , n77502 , n77503 , n77504 , 
 n77505 , n77506 , n77507 , n77508 , n77509 , n77510 , n77511 , n77512 , n77513 , n77514 , 
 n77515 , n77516 , n77517 , n77518 , n77519 , n77520 , n77521 , n77522 , n77523 , n77524 , 
 n77525 , n77526 , n77527 , n77528 , n77529 , n77530 , n77531 , n77532 , n77533 , n77534 , 
 n77535 , n77536 , n77537 , n77538 , n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , 
 n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , n77551 , n77552 , n77553 , n77554 , 
 n77555 , n77556 , n77557 , n77558 , n77559 , n77560 , n77561 , n77562 , n77563 , n77564 , 
 n77565 , n77566 , n77567 , n77568 , n77569 , n77570 , n77571 , n77572 , n77573 , n77574 , 
 n77575 , n77576 , n77577 , n77578 , n77579 , n77580 , n77581 , n77582 , n77583 , n77584 , 
 n77585 , n77586 , n77587 , n77588 , n77589 , n77590 , n77591 , n77592 , n77593 , n77594 , 
 n77595 , n77596 , n77597 , n77598 , n77599 , n77600 , n77601 , n77602 , n77603 , n77604 , 
 n77605 , n77606 , n77607 , n77608 , n77609 , n77610 , n77611 , n77612 , n77613 , n77614 , 
 n77615 , n77616 , n77617 , n77618 , n77619 , n77620 , n77621 , n77622 , n77623 , n77624 , 
 n77625 , n77626 , n77627 , n77628 , n77629 , n77630 , n77631 , n77632 , n77633 , n77634 , 
 n77635 , n77636 , n77637 , n77638 , n77639 , n77640 , n77641 , n77642 , n77643 , n77644 , 
 n77645 , n77646 , n77647 , n77648 , n77649 , n77650 , n77651 , n77652 , n77653 , n77654 , 
 n77655 , n77656 , n77657 , n77658 , n77659 , n77660 , n77661 , n77662 , n77663 , n77664 , 
 n77665 , n77666 , n77667 , n77668 , n77669 , n77670 , n77671 , n77672 , n77673 , n77674 , 
 n77675 , n77676 , n77677 , n77678 , n77679 , n77680 , n77681 , n77682 , n77683 , n77684 , 
 n77685 , n77686 , n77687 , n77688 , n77689 , n77690 , n77691 , n77692 , n77693 , n77694 , 
 n77695 , n77696 , n77697 , n77698 , n77699 , n77700 , n77701 , n77702 , n77703 , n77704 , 
 n77705 , n77706 , n77707 , n77708 , n77709 , n77710 , n77711 , n77712 , n77713 , n77714 , 
 n77715 , n77716 , n77717 , n77718 , n77719 , n77720 , n77721 , n77722 , n77723 , n77724 , 
 n77725 , n77726 , n77727 , n77728 , n77729 , n77730 , n77731 , n77732 , n77733 , n77734 , 
 n77735 , n77736 , n77737 , n77738 , n77739 , n77740 , n77741 , n77742 , n77743 , n77744 , 
 n77745 , n77746 , n77747 , n77748 , n77749 , n77750 , n77751 , n77752 , n77753 , n77754 , 
 n77755 , n77756 , n77757 , n77758 , n77759 , n77760 , n77761 , n77762 , n77763 , n77764 , 
 n77765 , n77766 , n77767 , n77768 , n77769 , n77770 , n77771 , n77772 , n77773 , n77774 , 
 n77775 , n77776 , n77777 , n77778 , n77779 , n77780 , n77781 , n77782 , n77783 , n77784 , 
 n77785 , n77786 , n77787 , n77788 , n77789 , n77790 , n77791 , n77792 , n77793 , n77794 , 
 n77795 , n77796 , n77797 , n77798 , n77799 , n77800 , n77801 , n77802 , n77803 , n77804 , 
 n77805 , n77806 , n77807 , n77808 , n77809 , n77810 , n77811 , n77812 , n77813 , n77814 , 
 n77815 , n77816 , n77817 , n77818 , n77819 , n77820 , n77821 , n77822 , n77823 , n77824 , 
 n77825 , n77826 , n77827 , n77828 , n77829 , n77830 , n77831 , n77832 , n77833 , n77834 , 
 n77835 , n77836 , n77837 , n77838 , n77839 , n77840 , n77841 , n77842 , n77843 , n77844 , 
 n77845 , n77846 , n77847 , n77848 , n77849 , n77850 , n77851 , n77852 , n77853 , n77854 , 
 n77855 , n77856 , n77857 , n77858 , n77859 , n77860 , n77861 , n77862 , n77863 , n77864 , 
 n77865 , n77866 , n77867 , n77868 , n77869 , n77870 , n77871 , n77872 , n77873 , n77874 , 
 n77875 , n77876 , n77877 , n77878 , n77879 , n77880 , n77881 , n77882 , n77883 , n77884 , 
 n77885 , n77886 , n77887 , n77888 , n77889 , n77890 , n77891 , n77892 , n77893 , n77894 , 
 n77895 , n77896 , n77897 , n77898 , n77899 , n77900 , n77901 , n77902 , n77903 , n77904 , 
 n77905 , n77906 , n77907 , n77908 , n77909 , n77910 , n77911 , n77912 , n77913 , n77914 , 
 n77915 , n77916 , n77917 , n77918 , n77919 , n77920 , n77921 , n77922 , n77923 , n77924 , 
 n77925 , n77926 , n77927 , n77928 , n77929 , n77930 , n77931 , n77932 , n77933 , n77934 , 
 n77935 , n77936 , n77937 , n77938 , n77939 , n77940 , n77941 , n77942 , n77943 , n77944 , 
 n77945 , n77946 , n77947 , n77948 , n77949 , n77950 , n77951 , n77952 , n77953 , n77954 , 
 n77955 , n77956 , n77957 , n77958 , n77959 , n77960 , n77961 , n77962 , n77963 , n77964 , 
 n77965 , n77966 , n77967 , n77968 , n77969 , n77970 , n77971 , n77972 , n77973 , n77974 , 
 n77975 , n77976 , n77977 , n77978 , n77979 , n77980 , n77981 , n77982 , n77983 , n77984 , 
 n77985 , n77986 , n77987 , n77988 , n77989 , n77990 , n77991 , n77992 , n77993 , n77994 , 
 n77995 , n77996 , n77997 , n77998 , n77999 , n78000 , n78001 , n78002 , n78003 , n78004 , 
 n78005 , n78006 , n78007 , n78008 , n78009 , n78010 , n78011 , n78012 , n78013 , n78014 , 
 n78015 , n78016 , n78017 , n78018 , n78019 , n78020 , n78021 , n78022 , n78023 , n78024 , 
 n78025 , n78026 , n78027 , n78028 , n78029 , n78030 , n78031 , n78032 , n78033 , n78034 , 
 n78035 , n78036 , n78037 , n78038 , n78039 , n78040 , n78041 , n78042 , n78043 , n78044 , 
 n78045 , n78046 , n78047 , n78048 , n78049 , n78050 , n78051 , n78052 , n78053 , n78054 , 
 n78055 , n78056 , n78057 , n78058 , n78059 , n78060 , n78061 , n78062 , n78063 , n78064 , 
 n78065 , n78066 , n78067 , n78068 , n78069 , n78070 , n78071 , n78072 , n78073 , n78074 , 
 n78075 , n78076 , n78077 , n78078 , n78079 , n78080 , n78081 , n78082 , n78083 , n78084 , 
 n78085 , n78086 , n78087 , n78088 , n78089 , n78090 , n78091 , n78092 , n78093 , n78094 , 
 n78095 , n78096 , n78097 , n78098 , n78099 , n78100 , n78101 , n78102 , n78103 , n78104 , 
 n78105 , n78106 , n78107 , n78108 , n78109 , n78110 , n78111 , n78112 , n78113 , n78114 , 
 n78115 , n78116 , n78117 , n78118 , n78119 , n78120 , n78121 , n78122 , n78123 , n78124 , 
 n78125 , n78126 , n78127 , n78128 , n78129 , n78130 , n78131 , n78132 , n78133 , n78134 , 
 n78135 , n78136 , n78137 , n78138 , n78139 , n78140 , n78141 , n78142 , n78143 , n78144 , 
 n78145 , n78146 , n78147 , n78148 , n78149 , n78150 , n78151 , n78152 , n78153 , n78154 , 
 n78155 , n78156 , n78157 , n78158 , n78159 , n78160 , n78161 , n78162 , n78163 , n78164 , 
 n78165 , n78166 , n78167 , n78168 , n78169 , n78170 , n78171 , n78172 , n78173 , n78174 , 
 n78175 , n78176 , n78177 , n78178 , n78179 , n78180 , n78181 , n78182 , n78183 , n78184 , 
 n78185 , n78186 , n78187 , n78188 , n78189 , n78190 , n78191 , n78192 , n78193 , n78194 , 
 n78195 , n78196 , n78197 , n78198 , n78199 , n78200 , n78201 , n78202 , n78203 , n78204 , 
 n78205 , n78206 , n78207 , n78208 , n78209 , n78210 , n78211 , n78212 , n78213 , n78214 , 
 n78215 , n78216 , n78217 , n78218 , n78219 , n78220 , n78221 , n78222 , n78223 , n78224 , 
 n78225 , n78226 , n78227 , n78228 , n78229 , n78230 , n78231 , n78232 , n78233 , n78234 , 
 n78235 , n78236 , n78237 , n78238 , n78239 , n78240 , n78241 , n78242 , n78243 , n78244 , 
 n78245 , n78246 , n78247 , n78248 , n78249 , n78250 , n78251 , n78252 , n78253 , n78254 , 
 n78255 , n78256 , n78257 , n78258 , n78259 , n78260 , n78261 , n78262 , n78263 , n78264 , 
 n78265 , n78266 , n78267 , n78268 , n78269 , n78270 , n78271 , n78272 , n78273 , n78274 , 
 n78275 , n78276 , n78277 , n78278 , n78279 , n78280 , n78281 , n78282 , n78283 , n78284 , 
 n78285 , n78286 , n78287 , n78288 , n78289 , n78290 , n78291 , n78292 , n78293 , n78294 , 
 n78295 , n78296 , n78297 , n78298 , n78299 , n78300 , n78301 , n78302 , n78303 , n78304 , 
 n78305 , n78306 , n78307 , n78308 , n78309 , n78310 , n78311 , n78312 , n78313 , n78314 , 
 n78315 , n78316 , n78317 , n78318 , n78319 , n78320 , n78321 , n78322 , n78323 , n78324 , 
 n78325 , n78326 , n78327 , n78328 , n78329 , n78330 , n78331 , n78332 , n78333 , n78334 , 
 n78335 , n78336 , n78337 , n78338 , n78339 , n78340 , n78341 , n78342 , n78343 , n78344 , 
 n78345 , n78346 , n78347 , n78348 , n78349 , n78350 , n78351 , n78352 , n78353 , n78354 , 
 n78355 , n78356 , n78357 , n78358 , n78359 , n78360 , n78361 , n78362 , n78363 , n78364 , 
 n78365 , n78366 , n78367 , n78368 , n78369 , n78370 , n78371 , n78372 , n78373 , n78374 , 
 n78375 , n78376 , n78377 , n78378 , n78379 , n78380 , n78381 , n78382 , n78383 , n78384 , 
 n78385 , n78386 , n78387 , n78388 , n78389 , n78390 , n78391 , n78392 , n78393 , n78394 , 
 n78395 , n78396 , n78397 , n78398 , n78399 , n78400 , n78401 , n78402 , n78403 , n78404 , 
 n78405 , n78406 , n78407 , n78408 , n78409 , n78410 , n78411 , n78412 , n78413 , n78414 , 
 n78415 , n78416 , n78417 , n78418 , n78419 , n78420 , n78421 , n78422 , n78423 , n78424 , 
 n78425 , n78426 , n78427 , n78428 , n78429 , n78430 , n78431 , n78432 , n78433 , n78434 , 
 n78435 , n78436 , n78437 , n78438 , n78439 , n78440 , n78441 , n78442 , n78443 , n78444 , 
 n78445 , n78446 , n78447 , n78448 , n78449 , n78450 , n78451 , n78452 , n78453 , n78454 , 
 n78455 , n78456 , n78457 , n78458 , n78459 , n78460 , n78461 , n78462 , n78463 , n78464 , 
 n78465 , n78466 , n78467 , n78468 , n78469 , n78470 , n78471 , n78472 , n78473 , n78474 , 
 n78475 , n78476 , n78477 , n78478 , n78479 , n78480 , n78481 , n78482 , n78483 , n78484 , 
 n78485 , n78486 , n78487 , n78488 , n78489 , n78490 , n78491 , n78492 , n78493 , n78494 , 
 n78495 , n78496 , n78497 , n78498 , n78499 , n78500 , n78501 , n78502 , n78503 , n78504 , 
 n78505 , n78506 , n78507 , n78508 , n78509 , n78510 , n78511 , n78512 , n78513 , n78514 , 
 n78515 , n78516 , n78517 , n78518 , n78519 , n78520 , n78521 , n78522 , n78523 , n78524 , 
 n78525 , n78526 , n78527 , n78528 , n78529 , n78530 , n78531 , n78532 , n78533 , n78534 , 
 n78535 , n78536 , n78537 , n78538 , n78539 , n78540 , n78541 , n78542 , n78543 , n78544 , 
 n78545 , n78546 , n78547 , n78548 , n78549 , n78550 , n78551 , n78552 , n78553 , n78554 , 
 n78555 , n78556 , n78557 , n78558 , n78559 , n78560 , n78561 , n78562 , n78563 , n78564 , 
 n78565 , n78566 , n78567 , n78568 , n78569 , n78570 , n78571 , n78572 , n78573 , n78574 , 
 n78575 , n78576 , n78577 , n78578 , n78579 , n78580 , n78581 , n78582 , n78583 , n78584 , 
 n78585 , n78586 , n78587 , n78588 , n78589 , n78590 , n78591 , n78592 , n78593 , n78594 , 
 n78595 , n78596 , n78597 , n78598 , n78599 , n78600 , n78601 , n78602 , n78603 , n78604 , 
 n78605 , n78606 , n78607 , n78608 , n78609 , n78610 , n78611 , n78612 , n78613 , n78614 , 
 n78615 , n78616 , n78617 , n78618 , n78619 , n78620 , n78621 , n78622 , n78623 , n78624 , 
 n78625 , n78626 , n78627 , n78628 , n78629 , n78630 , n78631 , n78632 , n78633 , n78634 , 
 n78635 , n78636 , n78637 , n78638 , n78639 , n78640 , n78641 , n78642 , n78643 , n78644 , 
 n78645 , n78646 , n78647 , n78648 , n78649 , n78650 , n78651 , n78652 , n78653 , n78654 , 
 n78655 , n78656 , n78657 , n78658 , n78659 , n78660 , n78661 , n78662 , n78663 , n78664 , 
 n78665 , n78666 , n78667 , n78668 , n78669 , n78670 , n78671 , n78672 , n78673 , n78674 , 
 n78675 , n78676 , n78677 , n78678 , n78679 , n78680 , n78681 , n78682 , n78683 , n78684 , 
 n78685 , n78686 , n78687 , n78688 , n78689 , n78690 , n78691 , n78692 , n78693 , n78694 , 
 n78695 , n78696 , n78697 , n78698 , n78699 , n78700 , n78701 , n78702 , n78703 , n78704 , 
 n78705 , n78706 , n78707 , n78708 , n78709 , n78710 , n78711 , n78712 , n78713 , n78714 , 
 n78715 , n78716 , n78717 , n78718 , n78719 , n78720 , n78721 , n78722 , n78723 , n78724 , 
 n78725 , n78726 , n78727 , n78728 , n78729 , n78730 , n78731 , n78732 , n78733 , n78734 , 
 n78735 , n78736 , n78737 , n78738 , n78739 , n78740 , n78741 , n78742 , n78743 , n78744 , 
 n78745 , n78746 , n78747 , n78748 , n78749 , n78750 , n78751 , n78752 , n78753 , n78754 , 
 n78755 , n78756 , n78757 , n78758 , n78759 , n78760 , n78761 , n78762 , n78763 , n78764 , 
 n78765 , n78766 , n78767 , n78768 , n78769 , n78770 , n78771 , n78772 , n78773 , n78774 , 
 n78775 , n78776 , n78777 , n78778 , n78779 , n78780 , n78781 , n78782 , n78783 , n78784 , 
 n78785 , n78786 , n78787 , n78788 , n78789 , n78790 , n78791 , n78792 , n78793 , n78794 , 
 n78795 , n78796 , n78797 , n78798 , n78799 , n78800 , n78801 , n78802 , n78803 , n78804 , 
 n78805 , n78806 , n78807 , n78808 , n78809 , n78810 , n78811 , n78812 , n78813 , n78814 , 
 n78815 , n78816 , n78817 , n78818 , n78819 , n78820 , n78821 , n78822 , n78823 , n78824 , 
 n78825 , n78826 , n78827 , n78828 , n78829 , n78830 , n78831 , n78832 , n78833 , n78834 , 
 n78835 , n78836 , n78837 , n78838 , n78839 , n78840 , n78841 , n78842 , n78843 , n78844 , 
 n78845 , n78846 , n78847 , n78848 , n78849 , n78850 , n78851 , n78852 , n78853 , n78854 , 
 n78855 , n78856 , n78857 , n78858 , n78859 , n78860 , n78861 , n78862 , n78863 , n78864 , 
 n78865 , n78866 , n78867 , n78868 , n78869 , n78870 , n78871 , n78872 , n78873 , n78874 , 
 n78875 , n78876 , n78877 , n78878 , n78879 , n78880 , n78881 , n78882 , n78883 , n78884 , 
 n78885 , n78886 , n78887 , n78888 , n78889 , n78890 , n78891 , n78892 , n78893 , n78894 , 
 n78895 , n78896 , n78897 , n78898 , n78899 , n78900 , n78901 , n78902 , n78903 , n78904 , 
 n78905 , n78906 , n78907 , n78908 , n78909 , n78910 , n78911 , n78912 , n78913 , n78914 , 
 n78915 , n78916 , n78917 , n78918 , n78919 , n78920 , n78921 , n78922 , n78923 , n78924 , 
 n78925 , n78926 , n78927 , n78928 , n78929 , n78930 , n78931 , n78932 , n78933 , n78934 , 
 n78935 , n78936 , n78937 , n78938 , n78939 , n78940 , n78941 , n78942 , n78943 , n78944 , 
 n78945 , n78946 , n78947 , n78948 , n78949 , n78950 , n78951 , n78952 , n78953 , n78954 , 
 n78955 , n78956 , n78957 , n78958 , n78959 , n78960 , n78961 , n78962 , n78963 , n78964 , 
 n78965 , n78966 , n78967 , n78968 , n78969 , n78970 , n78971 , n78972 , n78973 , n78974 , 
 n78975 , n78976 , n78977 , n78978 , n78979 , n78980 , n78981 , n78982 , n78983 , n78984 , 
 n78985 , n78986 , n78987 , n78988 , n78989 , n78990 , n78991 , n78992 , n78993 , n78994 , 
 n78995 , n78996 , n78997 , n78998 , n78999 , n79000 , n79001 , n79002 , n79003 , n79004 , 
 n79005 , n79006 , n79007 , n79008 , n79009 , n79010 , n79011 , n79012 , n79013 , n79014 , 
 n79015 , n79016 , n79017 , n79018 , n79019 , n79020 , n79021 , n79022 , n79023 , n79024 , 
 n79025 , n79026 , n79027 , n79028 , n79029 , n79030 , n79031 , n79032 , n79033 , n79034 , 
 n79035 , n79036 , n79037 , n79038 , n79039 , n79040 , n79041 , n79042 , n79043 , n79044 , 
 n79045 , n79046 , n79047 , n79048 , n79049 , n79050 , n79051 , n79052 , n79053 , n79054 , 
 n79055 , n79056 , n79057 , n79058 , n79059 , n79060 , n79061 , n79062 , n79063 , n79064 , 
 n79065 , n79066 , n79067 , n79068 , n79069 , n79070 , n79071 , n79072 , n79073 , n79074 , 
 n79075 , n79076 , n79077 , n79078 , n79079 , n79080 , n79081 , n79082 , n79083 , n79084 , 
 n79085 , n79086 , n79087 , n79088 , n79089 , n79090 , n79091 , n79092 , n79093 , n79094 , 
 n79095 , n79096 , n79097 , n79098 , n79099 , n79100 , n79101 , n79102 , n79103 , n79104 , 
 n79105 , n79106 , n79107 , n79108 , n79109 , n79110 , n79111 , n79112 , n79113 , n79114 , 
 n79115 , n79116 , n79117 , n79118 , n79119 , n79120 , n79121 , n79122 , n79123 , n79124 , 
 n79125 , n79126 , n79127 , n79128 , n79129 , n79130 , n79131 , n79132 , n79133 , n79134 , 
 n79135 , n79136 , n79137 , n79138 , n79139 , n79140 , n79141 , n79142 , n79143 , n79144 , 
 n79145 , n79146 , n79147 , n79148 , n79149 , n79150 , n79151 , n79152 , n79153 , n79154 , 
 n79155 , n79156 , n79157 , n79158 , n79159 , n79160 , n79161 , n79162 , n79163 , n79164 , 
 n79165 , n79166 , n79167 , n79168 , n79169 , n79170 , n79171 , n79172 , n79173 , n79174 , 
 n79175 , n79176 , n79177 , n79178 , n79179 , n79180 , n79181 , n79182 , n79183 , n79184 , 
 n79185 , n79186 , n79187 , n79188 , n79189 , n79190 , n79191 , n79192 , n79193 , n79194 , 
 n79195 , n79196 , n79197 , n79198 , n79199 , n79200 , n79201 , n79202 , n79203 , n79204 , 
 n79205 , n79206 , n79207 , n79208 , n79209 , n79210 , n79211 , n79212 , n79213 , n79214 , 
 n79215 , n79216 , n79217 , n79218 , n79219 , n79220 , n79221 , n79222 , n79223 , n79224 , 
 n79225 , n79226 , n79227 , n79228 , n79229 , n79230 , n79231 , n79232 , n79233 , n79234 , 
 n79235 , n79236 , n79237 , n79238 , n79239 , n79240 , n79241 , n79242 , n79243 , n79244 , 
 n79245 , n79246 , n79247 , n79248 , n79249 , n79250 , n79251 , n79252 , n79253 , n79254 , 
 n79255 , n79256 , n79257 , n79258 , n79259 , n79260 , n79261 , n79262 , n79263 , n79264 , 
 n79265 , n79266 , n79267 , n79268 , n79269 , n79270 , n79271 , n79272 , n79273 , n79274 , 
 n79275 , n79276 , n79277 , n79278 , n79279 , n79280 , n79281 , n79282 , n79283 , n79284 , 
 n79285 , n79286 , n79287 , n79288 , n79289 , n79290 , n79291 , n79292 , n79293 , n79294 , 
 n79295 , n79296 , n79297 , n79298 , n79299 , n79300 , n79301 , n79302 , n79303 , n79304 , 
 n79305 , n79306 , n79307 , n79308 , n79309 , n79310 , n79311 , n79312 , n79313 , n79314 , 
 n79315 , n79316 , n79317 , n79318 , n79319 , n79320 , n79321 , n79322 , n79323 , n79324 , 
 n79325 , n79326 , n79327 , n79328 , n79329 , n79330 , n79331 , n79332 , n79333 , n79334 , 
 n79335 , n79336 , n79337 , n79338 , n79339 , n79340 , n79341 , n79342 , n79343 , n79344 , 
 n79345 , n79346 , n79347 , n79348 , n79349 , n79350 , n79351 , n79352 , n79353 , n79354 , 
 n79355 , n79356 , n79357 , n79358 , n79359 , n79360 , n79361 , n79362 , n79363 , n79364 , 
 n79365 , n79366 , n79367 , n79368 , n79369 , n79370 , n79371 , n79372 , n79373 , n79374 , 
 n79375 , n79376 , n79377 , n79378 , n79379 , n79380 , n79381 , n79382 , n79383 , n79384 , 
 n79385 , n79386 , n79387 , n79388 , n79389 , n79390 , n79391 , n79392 , n79393 , n79394 , 
 n79395 , n79396 , n79397 , n79398 , n79399 , n79400 , n79401 , n79402 , n79403 , n79404 , 
 n79405 , n79406 , n79407 , n79408 , n79409 , n79410 , n79411 , n79412 , n79413 , n79414 , 
 n79415 , n79416 , n79417 , n79418 , n79419 , n79420 , n79421 , n79422 , n79423 , n79424 , 
 n79425 , n79426 , n79427 , n79428 , n79429 , n79430 , n79431 , n79432 , n79433 , n79434 , 
 n79435 , n79436 , n79437 , n79438 , n79439 , n79440 , n79441 , n79442 , n79443 , n79444 , 
 n79445 , n79446 , n79447 , n79448 , n79449 , n79450 , n79451 , n79452 , n79453 , n79454 , 
 n79455 , n79456 , n79457 , n79458 , n79459 , n79460 , n79461 , n79462 , n79463 , n79464 , 
 n79465 , n79466 , n79467 , n79468 , n79469 , n79470 , n79471 , n79472 , n79473 , n79474 , 
 n79475 , n79476 , n79477 , n79478 , n79479 , n79480 , n79481 , n79482 , n79483 , n79484 , 
 n79485 , n79486 , n79487 , n79488 , n79489 , n79490 , n79491 , n79492 , n79493 , n79494 , 
 n79495 , n79496 , n79497 , n79498 , n79499 , n79500 , n79501 , n79502 , n79503 , n79504 , 
 n79505 , n79506 , n79507 , n79508 , n79509 , n79510 , n79511 , n79512 , n79513 , n79514 , 
 n79515 , n79516 , n79517 , n79518 , n79519 , n79520 , n79521 , n79522 , n79523 , n79524 , 
 n79525 , n79526 , n79527 , n79528 , n79529 , n79530 , n79531 , n79532 , n79533 , n79534 , 
 n79535 , n79536 , n79537 , n79538 , n79539 , n79540 , n79541 , n79542 , n79543 , n79544 , 
 n79545 , n79546 , n79547 , n79548 , n79549 , n79550 , n79551 , n79552 , n79553 , n79554 , 
 n79555 , n79556 , n79557 , n79558 , n79559 , n79560 , n79561 , n79562 , n79563 , n79564 , 
 n79565 , n79566 , n79567 , n79568 , n79569 , n79570 , n79571 , n79572 , n79573 , n79574 , 
 n79575 , n79576 , n79577 , n79578 , n79579 , n79580 , n79581 , n79582 , n79583 , n79584 , 
 n79585 , n79586 , n79587 , n79588 , n79589 , n79590 , n79591 , n79592 , n79593 , n79594 , 
 n79595 , n79596 , n79597 , n79598 , n79599 , n79600 , n79601 , n79602 , n79603 , n79604 , 
 n79605 , n79606 , n79607 , n79608 , n79609 , n79610 , n79611 , n79612 , n79613 , n79614 , 
 n79615 , n79616 , n79617 , n79618 , n79619 , n79620 , n79621 , n79622 , n79623 , n79624 , 
 n79625 , n79626 , n79627 , n79628 , n79629 , n79630 , n79631 , n79632 , n79633 , n79634 , 
 n79635 , n79636 , n79637 , n79638 , n79639 , n79640 , n79641 , n79642 , n79643 , n79644 , 
 n79645 , n79646 , n79647 , n79648 , n79649 , n79650 , n79651 , n79652 , n79653 , n79654 , 
 n79655 , n79656 , n79657 , n79658 , n79659 , n79660 , n79661 , n79662 , n79663 , n79664 , 
 n79665 , n79666 , n79667 , n79668 , n79669 , n79670 , n79671 , n79672 , n79673 , n79674 , 
 n79675 , n79676 , n79677 , n79678 , n79679 , n79680 , n79681 , n79682 , n79683 , n79684 , 
 n79685 , n79686 , n79687 , n79688 , n79689 , n79690 , n79691 , n79692 , n79693 , n79694 , 
 n79695 , n79696 , n79697 , n79698 , n79699 , n79700 , n79701 , n79702 , n79703 , n79704 , 
 n79705 , n79706 , n79707 , n79708 , n79709 , n79710 , n79711 , n79712 , n79713 , n79714 , 
 n79715 , n79716 , n79717 , n79718 , n79719 , n79720 , n79721 , n79722 , n79723 , n79724 , 
 n79725 , n79726 , n79727 , n79728 , n79729 , n79730 , n79731 , n79732 , n79733 , n79734 , 
 n79735 , n79736 , n79737 , n79738 , n79739 , n79740 , n79741 , n79742 , n79743 , n79744 , 
 n79745 , n79746 , n79747 , n79748 , n79749 , n79750 , n79751 , n79752 , n79753 , n79754 , 
 n79755 , n79756 , n79757 , n79758 , n79759 , n79760 , n79761 , n79762 , n79763 , n79764 , 
 n79765 , n79766 , n79767 , n79768 , n79769 , n79770 , n79771 , n79772 , n79773 , n79774 , 
 n79775 , n79776 , n79777 , n79778 , n79779 , n79780 , n79781 , n79782 , n79783 , n79784 , 
 n79785 , n79786 , n79787 , n79788 , n79789 , n79790 , n79791 , n79792 , n79793 , n79794 , 
 n79795 , n79796 , n79797 , n79798 , n79799 , n79800 , n79801 , n79802 , n79803 , n79804 , 
 n79805 , n79806 , n79807 , n79808 , n79809 , n79810 , n79811 , n79812 , n79813 , n79814 , 
 n79815 , n79816 , n79817 , n79818 , n79819 , n79820 , n79821 , n79822 , n79823 , n79824 , 
 n79825 , n79826 , n79827 , n79828 , n79829 , n79830 , n79831 , n79832 , n79833 , n79834 , 
 n79835 , n79836 , n79837 , n79838 , n79839 , n79840 , n79841 , n79842 , n79843 , n79844 , 
 n79845 , n79846 , n79847 , n79848 , n79849 , n79850 , n79851 , n79852 , n79853 , n79854 , 
 n79855 , n79856 , n79857 , n79858 , n79859 , n79860 , n79861 , n79862 , n79863 , n79864 , 
 n79865 , n79866 , n79867 , n79868 , n79869 , n79870 , n79871 , n79872 , n79873 , n79874 , 
 n79875 , n79876 , n79877 , n79878 , n79879 , n79880 , n79881 , n79882 , n79883 , n79884 , 
 n79885 , n79886 , n79887 , n79888 , n79889 , n79890 , n79891 , n79892 , n79893 , n79894 , 
 n79895 , n79896 , n79897 , n79898 , n79899 , n79900 , n79901 , n79902 , n79903 , n79904 , 
 n79905 , n79906 , n79907 , n79908 , n79909 , n79910 , n79911 , n79912 , n79913 , n79914 , 
 n79915 , n79916 , n79917 , n79918 , n79919 , n79920 , n79921 , n79922 , n79923 , n79924 , 
 n79925 , n79926 , n79927 , n79928 , n79929 , n79930 , n79931 , n79932 , n79933 , n79934 , 
 n79935 , n79936 , n79937 , n79938 , n79939 , n79940 , n79941 , n79942 , n79943 , n79944 , 
 n79945 , n79946 , n79947 , n79948 , n79949 , n79950 , n79951 , n79952 , n79953 , n79954 , 
 n79955 , n79956 , n79957 , n79958 , n79959 , n79960 , n79961 , n79962 , n79963 , n79964 , 
 n79965 , n79966 , n79967 , n79968 , n79969 , n79970 , n79971 , n79972 , n79973 , n79974 , 
 n79975 , n79976 , n79977 , n79978 , n79979 , n79980 , n79981 , n79982 , n79983 , n79984 , 
 n79985 , n79986 , n79987 , n79988 , n79989 , n79990 , n79991 , n79992 , n79993 , n79994 , 
 n79995 , n79996 , n79997 , n79998 , n79999 , n80000 , n80001 , n80002 , n80003 , n80004 , 
 n80005 , n80006 , n80007 , n80008 , n80009 , n80010 , n80011 , n80012 , n80013 , n80014 , 
 n80015 , n80016 , n80017 , n80018 , n80019 , n80020 , n80021 , n80022 , n80023 , n80024 , 
 n80025 , n80026 , n80027 , n80028 , n80029 , n80030 , n80031 , n80032 , n80033 , n80034 , 
 n80035 , n80036 , n80037 , n80038 , n80039 , n80040 , n80041 , n80042 , n80043 , n80044 , 
 n80045 , n80046 , n80047 , n80048 , n80049 , n80050 , n80051 , n80052 , n80053 , n80054 , 
 n80055 , n80056 , n80057 , n80058 , n80059 , n80060 , n80061 , n80062 , n80063 , n80064 , 
 n80065 , n80066 , n80067 , n80068 , n80069 , n80070 , n80071 , n80072 , n80073 , n80074 , 
 n80075 , n80076 , n80077 , n80078 , n80079 , n80080 , n80081 , n80082 , n80083 , n80084 , 
 n80085 , n80086 , n80087 , n80088 , n80089 , n80090 , n80091 , n80092 , n80093 , n80094 , 
 n80095 , n80096 , n80097 , n80098 , n80099 , n80100 , n80101 , n80102 , n80103 , n80104 , 
 n80105 , n80106 , n80107 , n80108 , n80109 , n80110 , n80111 , n80112 , n80113 , n80114 , 
 n80115 , n80116 , n80117 , n80118 , n80119 , n80120 , n80121 , n80122 , n80123 , n80124 , 
 n80125 , n80126 , n80127 , n80128 , n80129 , n80130 , n80131 , n80132 , n80133 , n80134 , 
 n80135 , n80136 , n80137 , n80138 , n80139 , n80140 , n80141 , n80142 , n80143 , n80144 , 
 n80145 , n80146 , n80147 , n80148 , n80149 , n80150 , n80151 , n80152 , n80153 , n80154 , 
 n80155 , n80156 , n80157 , n80158 , n80159 , n80160 , n80161 , n80162 , n80163 , n80164 , 
 n80165 , n80166 , n80167 , n80168 , n80169 , n80170 , n80171 , n80172 , n80173 , n80174 , 
 n80175 , n80176 , n80177 , n80178 , n80179 , n80180 , n80181 , n80182 , n80183 , n80184 , 
 n80185 , n80186 , n80187 , n80188 , n80189 , n80190 , n80191 , n80192 , n80193 , n80194 , 
 n80195 , n80196 , n80197 , n80198 , n80199 , n80200 , n80201 , n80202 , n80203 , n80204 , 
 n80205 , n80206 , n80207 , n80208 , n80209 , n80210 , n80211 , n80212 , n80213 , n80214 , 
 n80215 , n80216 , n80217 , n80218 , n80219 , n80220 , n80221 , n80222 , n80223 , n80224 , 
 n80225 , n80226 , n80227 , n80228 , n80229 , n80230 , n80231 , n80232 , n80233 , n80234 , 
 n80235 , n80236 , n80237 , n80238 , n80239 , n80240 , n80241 , n80242 , n80243 , n80244 , 
 n80245 , n80246 , n80247 , n80248 , n80249 , n80250 , n80251 , n80252 , n80253 , n80254 , 
 n80255 , n80256 , n80257 , n80258 , n80259 , n80260 , n80261 , n80262 , n80263 , n80264 , 
 n80265 , n80266 , n80267 , n80268 , n80269 , n80270 , n80271 , n80272 , n80273 , n80274 , 
 n80275 , n80276 , n80277 , n80278 , n80279 , n80280 , n80281 , n80282 , n80283 , n80284 , 
 n80285 , n80286 , n80287 , n80288 , n80289 , n80290 , n80291 , n80292 , n80293 , n80294 , 
 n80295 , n80296 , n80297 , n80298 , n80299 , n80300 , n80301 , n80302 , n80303 , n80304 , 
 n80305 , n80306 , n80307 , n80308 , n80309 , n80310 , n80311 , n80312 , n80313 , n80314 , 
 n80315 , n80316 , n80317 , n80318 , n80319 , n80320 , n80321 , n80322 , n80323 , n80324 , 
 n80325 , n80326 , n80327 , n80328 , n80329 , n80330 , n80331 , n80332 , n80333 , n80334 , 
 n80335 , n80336 , n80337 , n80338 , n80339 , n80340 , n80341 , n80342 , n80343 , n80344 , 
 n80345 , n80346 , n80347 , n80348 , n80349 , n80350 , n80351 , n80352 , n80353 , n80354 , 
 n80355 , n80356 , n80357 , n80358 , n80359 , n80360 , n80361 , n80362 , n80363 , n80364 , 
 n80365 , n80366 , n80367 , n80368 , n80369 , n80370 , n80371 , n80372 , n80373 , n80374 , 
 n80375 , n80376 , n80377 , n80378 , n80379 , n80380 , n80381 , n80382 , n80383 , n80384 , 
 n80385 , n80386 , n80387 , n80388 , n80389 , n80390 , n80391 , n80392 , n80393 , n80394 , 
 n80395 , n80396 , n80397 , n80398 , n80399 , n80400 , n80401 , n80402 , n80403 , n80404 , 
 n80405 , n80406 , n80407 , n80408 , n80409 , n80410 , n80411 , n80412 , n80413 , n80414 , 
 n80415 , n80416 , n80417 , n80418 , n80419 , n80420 , n80421 , n80422 , n80423 , n80424 , 
 n80425 , n80426 , n80427 , n80428 , n80429 , n80430 , n80431 , n80432 , n80433 , n80434 , 
 n80435 , n80436 , n80437 , n80438 , n80439 , n80440 , n80441 , n80442 , n80443 , n80444 , 
 n80445 , n80446 , n80447 , n80448 , n80449 , n80450 , n80451 , n80452 , n80453 , n80454 , 
 n80455 , n80456 , n80457 , n80458 , n80459 , n80460 , n80461 , n80462 , n80463 , n80464 , 
 n80465 , n80466 , n80467 , n80468 , n80469 , n80470 , n80471 , n80472 , n80473 , n80474 , 
 n80475 , n80476 , n80477 , n80478 , n80479 , n80480 , n80481 , n80482 , n80483 , n80484 , 
 n80485 , n80486 , n80487 , n80488 , n80489 , n80490 , n80491 , n80492 , n80493 , n80494 , 
 n80495 , n80496 , n80497 , n80498 , n80499 , n80500 , n80501 , n80502 , n80503 , n80504 , 
 n80505 , n80506 , n80507 , n80508 , n80509 , n80510 , n80511 , n80512 , n80513 , n80514 , 
 n80515 , n80516 , n80517 , n80518 , n80519 , n80520 , n80521 , n80522 , n80523 , n80524 , 
 n80525 , n80526 , n80527 , n80528 , n80529 , n80530 , n80531 , n80532 , n80533 , n80534 , 
 n80535 , n80536 , n80537 , n80538 , n80539 , n80540 , n80541 , n80542 , n80543 , n80544 , 
 n80545 , n80546 , n80547 , n80548 , n80549 , n80550 , n80551 , n80552 , n80553 , n80554 , 
 n80555 , n80556 , n80557 , n80558 , n80559 , n80560 , n80561 , n80562 , n80563 , n80564 , 
 n80565 , n80566 , n80567 , n80568 , n80569 , n80570 , n80571 , n80572 , n80573 , n80574 , 
 n80575 , n80576 , n80577 , n80578 , n80579 , n80580 , n80581 , n80582 , n80583 , n80584 , 
 n80585 , n80586 , n80587 , n80588 , n80589 , n80590 , n80591 , n80592 , n80593 , n80594 , 
 n80595 , n80596 , n80597 , n80598 , n80599 , n80600 , n80601 , n80602 , n80603 , n80604 , 
 n80605 , n80606 , n80607 , n80608 , n80609 , n80610 , n80611 , n80612 , n80613 , n80614 , 
 n80615 , n80616 , n80617 , n80618 , n80619 , n80620 , n80621 , n80622 , n80623 , n80624 , 
 n80625 , n80626 , n80627 , n80628 , n80629 , n80630 , n80631 , n80632 , n80633 , n80634 , 
 n80635 , n80636 , n80637 , n80638 , n80639 , n80640 , n80641 , n80642 , n80643 , n80644 , 
 n80645 , n80646 , n80647 , n80648 , n80649 , n80650 , n80651 , n80652 , n80653 , n80654 , 
 n80655 , n80656 , n80657 , n80658 , n80659 , n80660 , n80661 , n80662 , n80663 , n80664 , 
 n80665 , n80666 , n80667 , n80668 , n80669 , n80670 , n80671 , n80672 , n80673 , n80674 , 
 n80675 , n80676 , n80677 , n80678 , n80679 , n80680 , n80681 , n80682 , n80683 , n80684 , 
 n80685 , n80686 , n80687 , n80688 , n80689 , n80690 , n80691 , n80692 , n80693 , n80694 , 
 n80695 , n80696 , n80697 , n80698 , n80699 , n80700 , n80701 , n80702 , n80703 , n80704 , 
 n80705 , n80706 , n80707 , n80708 , n80709 , n80710 , n80711 , n80712 , n80713 , n80714 , 
 n80715 , n80716 , n80717 , n80718 , n80719 , n80720 , n80721 , n80722 , n80723 , n80724 , 
 n80725 , n80726 , n80727 , n80728 , n80729 , n80730 , n80731 , n80732 , n80733 , n80734 , 
 n80735 , n80736 , n80737 , n80738 , n80739 , n80740 , n80741 , n80742 , n80743 , n80744 , 
 n80745 , n80746 , n80747 , n80748 , n80749 , n80750 , n80751 , n80752 , n80753 , n80754 , 
 n80755 , n80756 , n80757 , n80758 , n80759 , n80760 , n80761 , n80762 , n80763 , n80764 , 
 n80765 , n80766 , n80767 , n80768 , n80769 , n80770 , n80771 , n80772 , n80773 , n80774 , 
 n80775 , n80776 , n80777 , n80778 , n80779 , n80780 , n80781 , n80782 , n80783 , n80784 , 
 n80785 , n80786 , n80787 , n80788 , n80789 , n80790 , n80791 , n80792 , n80793 , n80794 , 
 n80795 , n80796 , n80797 , n80798 , n80799 , n80800 , n80801 , n80802 , n80803 , n80804 , 
 n80805 , n80806 , n80807 , n80808 , n80809 , n80810 , n80811 , n80812 , n80813 , n80814 , 
 n80815 , n80816 , n80817 , n80818 , n80819 , n80820 , n80821 , n80822 , n80823 , n80824 , 
 n80825 , n80826 , n80827 , n80828 , n80829 , n80830 , n80831 , n80832 , n80833 , n80834 , 
 n80835 , n80836 , n80837 , n80838 , n80839 , n80840 , n80841 , n80842 , n80843 , n80844 , 
 n80845 , n80846 , n80847 , n80848 , n80849 , n80850 , n80851 , n80852 , n80853 , n80854 , 
 n80855 , n80856 , n80857 , n80858 , n80859 , n80860 , n80861 , n80862 , n80863 , n80864 , 
 n80865 , n80866 , n80867 , n80868 , n80869 , n80870 , n80871 , n80872 , n80873 , n80874 , 
 n80875 , n80876 , n80877 , n80878 , n80879 , n80880 , n80881 , n80882 , n80883 , n80884 , 
 n80885 , n80886 , n80887 , n80888 , n80889 , n80890 , n80891 , n80892 , n80893 , n80894 , 
 n80895 , n80896 , n80897 , n80898 , n80899 , n80900 , n80901 , n80902 , n80903 , n80904 , 
 n80905 , n80906 , n80907 , n80908 , n80909 , n80910 , n80911 , n80912 , n80913 , n80914 , 
 n80915 , n80916 , n80917 , n80918 , n80919 , n80920 , n80921 , n80922 , n80923 , n80924 , 
 n80925 , n80926 , n80927 , n80928 , n80929 , n80930 , n80931 , n80932 , n80933 , n80934 , 
 n80935 , n80936 , n80937 , n80938 , n80939 , n80940 , n80941 , n80942 , n80943 , n80944 , 
 n80945 , n80946 , n80947 , n80948 , n80949 , n80950 , n80951 , n80952 , n80953 , n80954 , 
 n80955 , n80956 , n80957 , n80958 , n80959 , n80960 , n80961 , n80962 , n80963 , n80964 , 
 n80965 , n80966 , n80967 , n80968 , n80969 , n80970 , n80971 , n80972 , n80973 , n80974 , 
 n80975 , n80976 , n80977 , n80978 , n80979 , n80980 , n80981 , n80982 , n80983 , n80984 , 
 n80985 , n80986 , n80987 , n80988 , n80989 , n80990 , n80991 , n80992 , n80993 , n80994 , 
 n80995 , n80996 , n80997 , n80998 , n80999 , n81000 , n81001 , n81002 , n81003 , n81004 , 
 n81005 , n81006 , n81007 , n81008 , n81009 , n81010 , n81011 , n81012 , n81013 , n81014 , 
 n81015 , n81016 , n81017 , n81018 , n81019 , n81020 , n81021 , n81022 , n81023 , n81024 , 
 n81025 , n81026 , n81027 , n81028 , n81029 , n81030 , n81031 , n81032 , n81033 , n81034 , 
 n81035 , n81036 , n81037 , n81038 , n81039 , n81040 , n81041 , n81042 , n81043 , n81044 , 
 n81045 , n81046 , n81047 , n81048 , n81049 , n81050 , n81051 , n81052 , n81053 , n81054 , 
 n81055 , n81056 , n81057 , n81058 , n81059 , n81060 , n81061 , n81062 , n81063 , n81064 , 
 n81065 , n81066 , n81067 , n81068 , n81069 , n81070 , n81071 , n81072 , n81073 , n81074 , 
 n81075 , n81076 , n81077 , n81078 , n81079 , n81080 , n81081 , n81082 , n81083 , n81084 , 
 n81085 , n81086 , n81087 , n81088 , n81089 , n81090 , n81091 , n81092 , n81093 , n81094 , 
 n81095 , n81096 , n81097 , n81098 , n81099 , n81100 , n81101 , n81102 , n81103 , n81104 , 
 n81105 , n81106 , n81107 , n81108 , n81109 , n81110 , n81111 , n81112 , n81113 , n81114 , 
 n81115 , n81116 , n81117 , n81118 , n81119 , n81120 , n81121 , n81122 , n81123 , n81124 , 
 n81125 , n81126 , n81127 , n81128 , n81129 , n81130 , n81131 , n81132 , n81133 , n81134 , 
 n81135 , n81136 , n81137 , n81138 , n81139 , n81140 , n81141 , n81142 , n81143 , n81144 , 
 n81145 , n81146 , n81147 , n81148 , n81149 , n81150 , n81151 , n81152 , n81153 , n81154 , 
 n81155 , n81156 , n81157 , n81158 , n81159 , n81160 , n81161 , n81162 , n81163 , n81164 , 
 n81165 , n81166 , n81167 , n81168 , n81169 , n81170 , n81171 , n81172 , n81173 , n81174 , 
 n81175 , n81176 , n81177 , n81178 , n81179 , n81180 , n81181 , n81182 , n81183 , n81184 , 
 n81185 , n81186 , n81187 , n81188 , n81189 , n81190 , n81191 , n81192 , n81193 , n81194 , 
 n81195 , n81196 , n81197 , n81198 , n81199 , n81200 , n81201 , n81202 , n81203 , n81204 , 
 n81205 , n81206 , n81207 , n81208 , n81209 , n81210 , n81211 , n81212 , n81213 , n81214 , 
 n81215 , n81216 , n81217 , n81218 , n81219 , n81220 , n81221 , n81222 , n81223 , n81224 , 
 n81225 , n81226 , n81227 , n81228 , n81229 , n81230 , n81231 , n81232 , n81233 , n81234 , 
 n81235 , n81236 , n81237 , n81238 , n81239 , n81240 , n81241 , n81242 , n81243 , n81244 , 
 n81245 , n81246 , n81247 , n81248 , n81249 , n81250 , n81251 , n81252 , n81253 , n81254 , 
 n81255 , n81256 , n81257 , n81258 , n81259 , n81260 , n81261 , n81262 , n81263 , n81264 , 
 n81265 , n81266 , n81267 , n81268 , n81269 , n81270 , n81271 , n81272 , n81273 , n81274 , 
 n81275 , n81276 , n81277 , n81278 , n81279 , n81280 , n81281 , n81282 , n81283 , n81284 , 
 n81285 , n81286 , n81287 , n81288 , n81289 , n81290 , n81291 , n81292 , n81293 , n81294 , 
 n81295 , n81296 , n81297 , n81298 , n81299 , n81300 , n81301 , n81302 , n81303 , n81304 , 
 n81305 , n81306 , n81307 , n81308 , n81309 , n81310 , n81311 , n81312 , n81313 , n81314 , 
 n81315 , n81316 , n81317 , n81318 , n81319 , n81320 , n81321 , n81322 , n81323 , n81324 , 
 n81325 , n81326 , n81327 , n81328 , n81329 , n81330 , n81331 , n81332 , n81333 , n81334 , 
 n81335 , n81336 , n81337 , n81338 , n81339 , n81340 , n81341 , n81342 , n81343 , n81344 , 
 n81345 , n81346 , n81347 , n81348 , n81349 , n81350 , n81351 , n81352 , n81353 , n81354 , 
 n81355 , n81356 , n81357 , n81358 , n81359 , n81360 , n81361 , n81362 , n81363 , n81364 , 
 n81365 , n81366 , n81367 , n81368 , n81369 , n81370 , n81371 , n81372 , n81373 , n81374 , 
 n81375 , n81376 , n81377 , n81378 , n81379 , n81380 , n81381 , n81382 , n81383 , n81384 , 
 n81385 , n81386 , n81387 , n81388 , n81389 , n81390 , n81391 , n81392 , n81393 , n81394 , 
 n81395 , n81396 , n81397 , n81398 , n81399 , n81400 , n81401 , n81402 , n81403 , n81404 , 
 n81405 , n81406 , n81407 , n81408 , n81409 , n81410 , n81411 , n81412 , n81413 , n81414 , 
 n81415 , n81416 , n81417 , n81418 , n81419 , n81420 , n81421 , n81422 , n81423 , n81424 , 
 n81425 , n81426 , n81427 , n81428 , n81429 , n81430 , n81431 , n81432 , n81433 , n81434 , 
 n81435 , n81436 , n81437 , n81438 , n81439 , n81440 , n81441 , n81442 , n81443 , n81444 , 
 n81445 , n81446 , n81447 , n81448 , n81449 , n81450 , n81451 , n81452 , n81453 , n81454 , 
 n81455 , n81456 , n81457 , n81458 , n81459 , n81460 , n81461 , n81462 , n81463 , n81464 , 
 n81465 , n81466 , n81467 , n81468 , n81469 , n81470 , n81471 , n81472 , n81473 , n81474 , 
 n81475 , n81476 , n81477 , n81478 , n81479 , n81480 , n81481 , n81482 , n81483 , n81484 , 
 n81485 , n81486 , n81487 , n81488 , n81489 , n81490 , n81491 , n81492 , n81493 , n81494 , 
 n81495 , n81496 , n81497 , n81498 , n81499 , n81500 , n81501 , n81502 , n81503 , n81504 , 
 n81505 , n81506 , n81507 , n81508 , n81509 , n81510 , n81511 , n81512 , n81513 , n81514 , 
 n81515 , n81516 , n81517 , n81518 , n81519 , n81520 , n81521 , n81522 , n81523 , n81524 , 
 n81525 , n81526 , n81527 , n81528 , n81529 , n81530 , n81531 , n81532 , n81533 , n81534 , 
 n81535 , n81536 , n81537 , n81538 , n81539 , n81540 , n81541 , n81542 , n81543 , n81544 , 
 n81545 , n81546 , n81547 , n81548 , n81549 , n81550 , n81551 , n81552 , n81553 , n81554 , 
 n81555 , n81556 , n81557 , n81558 , n81559 , n81560 , n81561 , n81562 , n81563 , n81564 , 
 n81565 , n81566 , n81567 , n81568 , n81569 , n81570 , n81571 , n81572 , n81573 , n81574 , 
 n81575 , n81576 , n81577 , n81578 , n81579 , n81580 , n81581 , n81582 , n81583 , n81584 , 
 n81585 , n81586 , n81587 , n81588 , n81589 , n81590 , n81591 , n81592 , n81593 , n81594 , 
 n81595 , n81596 , n81597 , n81598 , n81599 , n81600 , n81601 , n81602 , n81603 , n81604 , 
 n81605 , n81606 , n81607 , n81608 , n81609 , n81610 , n81611 , n81612 , n81613 , n81614 , 
 n81615 , n81616 , n81617 , n81618 , n81619 , n81620 , n81621 , n81622 , n81623 , n81624 , 
 n81625 , n81626 , n81627 , n81628 , n81629 , n81630 , n81631 , n81632 , n81633 , n81634 , 
 n81635 , n81636 , n81637 , n81638 , n81639 , n81640 , n81641 , n81642 , n81643 , n81644 , 
 n81645 , n81646 , n81647 , n81648 , n81649 , n81650 , n81651 , n81652 , n81653 , n81654 , 
 n81655 , n81656 , n81657 , n81658 , n81659 , n81660 , n81661 , n81662 , n81663 , n81664 , 
 n81665 , n81666 , n81667 , n81668 , n81669 , n81670 , n81671 , n81672 , n81673 , n81674 , 
 n81675 , n81676 , n81677 , n81678 , n81679 , n81680 , n81681 , n81682 , n81683 , n81684 , 
 n81685 , n81686 , n81687 , n81688 , n81689 , n81690 , n81691 , n81692 , n81693 , n81694 , 
 n81695 , n81696 , n81697 , n81698 , n81699 , n81700 , n81701 , n81702 , n81703 , n81704 , 
 n81705 , n81706 , n81707 , n81708 , n81709 , n81710 , n81711 , n81712 , n81713 , n81714 , 
 n81715 , n81716 , n81717 , n81718 , n81719 , n81720 , n81721 , n81722 , n81723 , n81724 , 
 n81725 , n81726 , n81727 , n81728 , n81729 , n81730 , n81731 , n81732 , n81733 , n81734 , 
 n81735 , n81736 , n81737 , n81738 , n81739 , n81740 , n81741 , n81742 , n81743 , n81744 , 
 n81745 , n81746 , n81747 , n81748 , n81749 , n81750 , n81751 , n81752 , n81753 , n81754 , 
 n81755 , n81756 , n81757 , n81758 , n81759 , n81760 , n81761 , n81762 , n81763 , n81764 , 
 n81765 , n81766 , n81767 , n81768 , n81769 , n81770 , n81771 , n81772 , n81773 , n81774 , 
 n81775 , n81776 , n81777 , n81778 , n81779 , n81780 , n81781 , n81782 , n81783 , n81784 , 
 n81785 , n81786 , n81787 , n81788 , n81789 , n81790 , n81791 , n81792 , n81793 , n81794 , 
 n81795 , n81796 , n81797 , n81798 , n81799 , n81800 , n81801 , n81802 , n81803 , n81804 , 
 n81805 , n81806 , n81807 , n81808 , n81809 , n81810 , n81811 , n81812 , n81813 , n81814 , 
 n81815 , n81816 , n81817 , n81818 , n81819 , n81820 , n81821 , n81822 , n81823 , n81824 , 
 n81825 , n81826 , n81827 , n81828 , n81829 , n81830 , n81831 , n81832 , n81833 , n81834 , 
 n81835 , n81836 , n81837 , n81838 , n81839 , n81840 , n81841 , n81842 , n81843 , n81844 , 
 n81845 , n81846 , n81847 , n81848 , n81849 , n81850 , n81851 , n81852 , n81853 , n81854 , 
 n81855 , n81856 , n81857 , n81858 , n81859 , n81860 , n81861 , n81862 , n81863 , n81864 , 
 n81865 , n81866 , n81867 , n81868 , n81869 , n81870 , n81871 , n81872 , n81873 , n81874 , 
 n81875 , n81876 , n81877 , n81878 , n81879 , n81880 , n81881 , n81882 , n81883 , n81884 , 
 n81885 , n81886 , n81887 , n81888 , n81889 , n81890 , n81891 , n81892 , n81893 , n81894 , 
 n81895 , n81896 , n81897 , n81898 , n81899 , n81900 , n81901 , n81902 , n81903 , n81904 , 
 n81905 , n81906 , n81907 , n81908 , n81909 , n81910 , n81911 , n81912 , n81913 , n81914 , 
 n81915 , n81916 , n81917 , n81918 , n81919 , n81920 , n81921 , n81922 , n81923 , n81924 , 
 n81925 , n81926 , n81927 , n81928 , n81929 , n81930 , n81931 , n81932 , n81933 , n81934 , 
 n81935 , n81936 , n81937 , n81938 , n81939 , n81940 , n81941 , n81942 , n81943 , n81944 , 
 n81945 , n81946 , n81947 , n81948 , n81949 , n81950 , n81951 , n81952 , n81953 , n81954 , 
 n81955 , n81956 , n81957 , n81958 , n81959 , n81960 , n81961 , n81962 , n81963 , n81964 , 
 n81965 , n81966 , n81967 , n81968 , n81969 , n81970 , n81971 , n81972 , n81973 , n81974 , 
 n81975 , n81976 , n81977 , n81978 , n81979 , n81980 , n81981 , n81982 , n81983 , n81984 , 
 n81985 , n81986 , n81987 , n81988 , n81989 , n81990 , n81991 , n81992 , n81993 , n81994 , 
 n81995 , n81996 , n81997 , n81998 , n81999 , n82000 , n82001 , n82002 , n82003 , n82004 , 
 n82005 , n82006 , n82007 , n82008 , n82009 , n82010 , n82011 , n82012 , n82013 , n82014 , 
 n82015 , n82016 , n82017 , n82018 , n82019 , n82020 , n82021 , n82022 , n82023 , n82024 , 
 n82025 , n82026 , n82027 , n82028 , n82029 , n82030 , n82031 , n82032 , n82033 , n82034 , 
 n82035 , n82036 , n82037 , n82038 , n82039 , n82040 , n82041 , n82042 , n82043 , n82044 , 
 n82045 , n82046 , n82047 , n82048 , n82049 , n82050 , n82051 , n82052 , n82053 , n82054 , 
 n82055 , n82056 , n82057 , n82058 , n82059 , n82060 , n82061 , n82062 , n82063 , n82064 , 
 n82065 , n82066 , n82067 , n82068 , n82069 , n82070 , n82071 , n82072 , n82073 , n82074 , 
 n82075 , n82076 , n82077 , n82078 , n82079 , n82080 , n82081 , n82082 , n82083 , n82084 , 
 n82085 , n82086 , n82087 , n82088 , n82089 , n82090 , n82091 , n82092 , n82093 , n82094 , 
 n82095 , n82096 , n82097 , n82098 , n82099 , n82100 , n82101 , n82102 , n82103 , n82104 , 
 n82105 , n82106 , n82107 , n82108 , n82109 , n82110 , n82111 , n82112 , n82113 , n82114 , 
 n82115 , n82116 , n82117 , n82118 , n82119 , n82120 , n82121 , n82122 , n82123 , n82124 , 
 n82125 , n82126 , n82127 , n82128 , n82129 , n82130 , n82131 , n82132 , n82133 , n82134 , 
 n82135 , n82136 , n82137 , n82138 , n82139 , n82140 , n82141 , n82142 , n82143 , n82144 , 
 n82145 , n82146 , n82147 , n82148 , n82149 , n82150 , n82151 , n82152 , n82153 , n82154 , 
 n82155 , n82156 , n82157 , n82158 , n82159 , n82160 , n82161 , n82162 , n82163 , n82164 , 
 n82165 , n82166 , n82167 , n82168 , n82169 , n82170 , n82171 , n82172 , n82173 , n82174 , 
 n82175 , n82176 , n82177 , n82178 , n82179 , n82180 , n82181 , n82182 , n82183 , n82184 , 
 n82185 , n82186 , n82187 , n82188 , n82189 , n82190 , n82191 , n82192 , n82193 , n82194 , 
 n82195 , n82196 , n82197 , n82198 , n82199 , n82200 , n82201 , n82202 , n82203 , n82204 , 
 n82205 , n82206 , n82207 , n82208 , n82209 , n82210 , n82211 , n82212 , n82213 , n82214 , 
 n82215 , n82216 , n82217 , n82218 , n82219 , n82220 , n82221 , n82222 , n82223 , n82224 , 
 n82225 , n82226 , n82227 , n82228 , n82229 , n82230 , n82231 , n82232 , n82233 , n82234 , 
 n82235 , n82236 , n82237 , n82238 , n82239 , n82240 , n82241 , n82242 , n82243 , n82244 , 
 n82245 , n82246 , n82247 , n82248 , n82249 , n82250 , n82251 , n82252 , n82253 , n82254 , 
 n82255 , n82256 , n82257 , n82258 , n82259 , n82260 , n82261 , n82262 , n82263 , n82264 , 
 n82265 , n82266 , n82267 , n82268 , n82269 , n82270 , n82271 , n82272 , n82273 , n82274 , 
 n82275 , n82276 , n82277 , n82278 , n82279 , n82280 , n82281 , n82282 , n82283 , n82284 , 
 n82285 , n82286 , n82287 , n82288 , n82289 , n82290 , n82291 , n82292 , n82293 , n82294 , 
 n82295 , n82296 , n82297 , n82298 , n82299 , n82300 , n82301 , n82302 , n82303 , n82304 , 
 n82305 , n82306 , n82307 , n82308 , n82309 , n82310 , n82311 , n82312 , n82313 , n82314 , 
 n82315 , n82316 , n82317 , n82318 , n82319 , n82320 , n82321 , n82322 , n82323 , n82324 , 
 n82325 , n82326 , n82327 , n82328 , n82329 , n82330 , n82331 , n82332 , n82333 , n82334 , 
 n82335 , n82336 , n82337 , n82338 , n82339 , n82340 , n82341 , n82342 , n82343 , n82344 , 
 n82345 , n82346 , n82347 , n82348 , n82349 , n82350 , n82351 , n82352 , n82353 , n82354 , 
 n82355 , n82356 , n82357 , n82358 , n82359 , n82360 , n82361 , n82362 , n82363 , n82364 , 
 n82365 , n82366 , n82367 , n82368 , n82369 , n82370 , n82371 , n82372 , n82373 , n82374 , 
 n82375 , n82376 , n82377 , n82378 , n82379 , n82380 , n82381 , n82382 , n82383 , n82384 , 
 n82385 , n82386 , n82387 , n82388 , n82389 , n82390 , n82391 , n82392 , n82393 , n82394 , 
 n82395 , n82396 , n82397 , n82398 , n82399 , n82400 , n82401 , n82402 , n82403 , n82404 , 
 n82405 , n82406 , n82407 , n82408 , n82409 , n82410 , n82411 , n82412 , n82413 , n82414 , 
 n82415 , n82416 , n82417 , n82418 , n82419 , n82420 , n82421 , n82422 , n82423 , n82424 , 
 n82425 , n82426 , n82427 , n82428 , n82429 , n82430 , n82431 , n82432 , n82433 , n82434 , 
 n82435 , n82436 , n82437 , n82438 , n82439 , n82440 , n82441 , n82442 , n82443 , n82444 , 
 n82445 , n82446 , n82447 , n82448 , n82449 , n82450 , n82451 , n82452 , n82453 , n82454 , 
 n82455 , n82456 , n82457 , n82458 , n82459 , n82460 , n82461 , n82462 , n82463 , n82464 , 
 n82465 , n82466 , n82467 , n82468 , n82469 , n82470 , n82471 , n82472 , n82473 , n82474 , 
 n82475 , n82476 , n82477 , n82478 , n82479 , n82480 , n82481 , n82482 , n82483 , n82484 , 
 n82485 , n82486 , n82487 , n82488 , n82489 , n82490 , n82491 , n82492 , n82493 , n82494 , 
 n82495 , n82496 , n82497 , n82498 , n82499 , n82500 , n82501 , n82502 , n82503 , n82504 , 
 n82505 , n82506 , n82507 , n82508 , n82509 , n82510 , n82511 , n82512 , n82513 , n82514 , 
 n82515 , n82516 , n82517 , n82518 , n82519 , n82520 , n82521 , n82522 , n82523 , n82524 , 
 n82525 , n82526 , n82527 , n82528 , n82529 , n82530 , n82531 , n82532 , n82533 , n82534 , 
 n82535 , n82536 , n82537 , n82538 , n82539 , n82540 , n82541 , n82542 , n82543 , n82544 , 
 n82545 , n82546 , n82547 , n82548 , n82549 , n82550 , n82551 , n82552 , n82553 , n82554 , 
 n82555 , n82556 , n82557 , n82558 , n82559 , n82560 , n82561 , n82562 , n82563 , n82564 , 
 n82565 , n82566 , n82567 , n82568 , n82569 , n82570 , n82571 , n82572 , n82573 , n82574 , 
 n82575 , n82576 , n82577 , n82578 , n82579 , n82580 , n82581 , n82582 , n82583 , n82584 , 
 n82585 , n82586 , n82587 , n82588 , n82589 , n82590 , n82591 , n82592 , n82593 , n82594 , 
 n82595 , n82596 , n82597 , n82598 , n82599 , n82600 , n82601 , n82602 , n82603 , n82604 , 
 n82605 , n82606 , n82607 , n82608 , n82609 , n82610 , n82611 , n82612 , n82613 , n82614 , 
 n82615 , n82616 , n82617 , n82618 , n82619 , n82620 , n82621 , n82622 , n82623 , n82624 , 
 n82625 , n82626 , n82627 , n82628 , n82629 , n82630 , n82631 , n82632 , n82633 , n82634 , 
 n82635 , n82636 , n82637 , n82638 , n82639 , n82640 , n82641 , n82642 , n82643 , n82644 , 
 n82645 , n82646 , n82647 , n82648 , n82649 , n82650 , n82651 , n82652 , n82653 , n82654 , 
 n82655 , n82656 , n82657 , n82658 , n82659 , n82660 , n82661 , n82662 , n82663 , n82664 , 
 n82665 , n82666 , n82667 , n82668 , n82669 , n82670 , n82671 , n82672 , n82673 , n82674 , 
 n82675 , n82676 , n82677 , n82678 , n82679 , n82680 , n82681 , n82682 , n82683 , n82684 , 
 n82685 , n82686 , n82687 , n82688 , n82689 , n82690 , n82691 , n82692 , n82693 , n82694 , 
 n82695 , n82696 , n82697 , n82698 , n82699 , n82700 , n82701 , n82702 , n82703 , n82704 , 
 n82705 , n82706 , n82707 , n82708 , n82709 , n82710 , n82711 , n82712 , n82713 , n82714 , 
 n82715 , n82716 , n82717 , n82718 , n82719 , n82720 , n82721 , n82722 , n82723 , n82724 , 
 n82725 , n82726 , n82727 , n82728 , n82729 , n82730 , n82731 , n82732 , n82733 , n82734 , 
 n82735 , n82736 , n82737 , n82738 , n82739 , n82740 , n82741 , n82742 , n82743 , n82744 , 
 n82745 , n82746 , n82747 , n82748 , n82749 , n82750 , n82751 , n82752 , n82753 , n82754 , 
 n82755 , n82756 , n82757 , n82758 , n82759 , n82760 , n82761 , n82762 , n82763 , n82764 , 
 n82765 , n82766 , n82767 , n82768 , n82769 , n82770 , n82771 , n82772 , n82773 , n82774 , 
 n82775 , n82776 , n82777 , n82778 , n82779 , n82780 , n82781 , n82782 , n82783 , n82784 , 
 n82785 , n82786 , n82787 , n82788 , n82789 , n82790 , n82791 , n82792 , n82793 , n82794 , 
 n82795 , n82796 , n82797 , n82798 , n82799 , n82800 , n82801 , n82802 , n82803 , n82804 , 
 n82805 , n82806 , n82807 , n82808 , n82809 , n82810 , n82811 , n82812 , n82813 , n82814 , 
 n82815 , n82816 , n82817 , n82818 , n82819 , n82820 , n82821 , n82822 , n82823 , n82824 , 
 n82825 , n82826 , n82827 , n82828 , n82829 , n82830 , n82831 , n82832 , n82833 , n82834 , 
 n82835 , n82836 , n82837 , n82838 , n82839 , n82840 , n82841 , n82842 , n82843 , n82844 , 
 n82845 , n82846 , n82847 , n82848 , n82849 , n82850 , n82851 , n82852 , n82853 , n82854 , 
 n82855 , n82856 , n82857 , n82858 , n82859 , n82860 , n82861 , n82862 , n82863 , n82864 , 
 n82865 , n82866 , n82867 , n82868 , n82869 , n82870 , n82871 , n82872 , n82873 , n82874 , 
 n82875 , n82876 , n82877 , n82878 , n82879 , n82880 , n82881 , n82882 , n82883 , n82884 , 
 n82885 , n82886 , n82887 , n82888 , n82889 , n82890 , n82891 , n82892 , n82893 , n82894 , 
 n82895 , n82896 , n82897 , n82898 , n82899 , n82900 , n82901 , n82902 , n82903 , n82904 , 
 n82905 , n82906 , n82907 , n82908 , n82909 , n82910 , n82911 , n82912 , n82913 , n82914 , 
 n82915 , n82916 , n82917 , n82918 , n82919 , n82920 , n82921 , n82922 , n82923 , n82924 , 
 n82925 , n82926 , n82927 , n82928 , n82929 , n82930 , n82931 , n82932 , n82933 , n82934 , 
 n82935 , n82936 , n82937 , n82938 , n82939 , n82940 , n82941 , n82942 , n82943 , n82944 , 
 n82945 , n82946 , n82947 , n82948 , n82949 , n82950 , n82951 , n82952 , n82953 , n82954 , 
 n82955 , n82956 , n82957 , n82958 , n82959 , n82960 , n82961 , n82962 , n82963 , n82964 , 
 n82965 , n82966 , n82967 , n82968 , n82969 , n82970 , n82971 , n82972 , n82973 , n82974 , 
 n82975 , n82976 , n82977 , n82978 , n82979 , n82980 , n82981 , n82982 , n82983 , n82984 , 
 n82985 , n82986 , n82987 , n82988 , n82989 , n82990 , n82991 , n82992 , n82993 , n82994 , 
 n82995 , n82996 , n82997 , n82998 , n82999 , n83000 , n83001 , n83002 , n83003 , n83004 , 
 n83005 , n83006 , n83007 , n83008 , n83009 , n83010 , n83011 , n83012 , n83013 , n83014 , 
 n83015 , n83016 , n83017 , n83018 , n83019 , n83020 , n83021 , n83022 , n83023 , n83024 , 
 n83025 , n83026 , n83027 , n83028 , n83029 , n83030 , n83031 , n83032 , n83033 , n83034 , 
 n83035 , n83036 , n83037 , n83038 , n83039 , n83040 , n83041 , n83042 , n83043 , n83044 , 
 n83045 , n83046 , n83047 , n83048 , n83049 , n83050 , n83051 , n83052 , n83053 , n83054 , 
 n83055 , n83056 , n83057 , n83058 , n83059 , n83060 , n83061 , n83062 , n83063 , n83064 , 
 n83065 , n83066 , n83067 , n83068 , n83069 , n83070 , n83071 , n83072 , n83073 , n83074 , 
 n83075 , n83076 , n83077 , n83078 , n83079 , n83080 , n83081 , n83082 , n83083 , n83084 , 
 n83085 , n83086 , n83087 , n83088 , n83089 , n83090 , n83091 , n83092 , n83093 , n83094 , 
 n83095 , n83096 , n83097 , n83098 , n83099 , n83100 , n83101 , n83102 , n83103 , n83104 , 
 n83105 , n83106 , n83107 , n83108 , n83109 , n83110 , n83111 , n83112 , n83113 , n83114 , 
 n83115 , n83116 , n83117 , n83118 , n83119 , n83120 , n83121 , n83122 , n83123 , n83124 , 
 n83125 , n83126 , n83127 , n83128 , n83129 , n83130 , n83131 , n83132 , n83133 , n83134 , 
 n83135 , n83136 , n83137 , n83138 , n83139 , n83140 , n83141 , n83142 , n83143 , n83144 , 
 n83145 , n83146 , n83147 , n83148 , n83149 , n83150 , n83151 , n83152 , n83153 , n83154 , 
 n83155 , n83156 , n83157 , n83158 , n83159 , n83160 , n83161 , n83162 , n83163 , n83164 , 
 n83165 , n83166 , n83167 , n83168 , n83169 , n83170 , n83171 , n83172 , n83173 , n83174 , 
 n83175 , n83176 , n83177 , n83178 , n83179 , n83180 , n83181 , n83182 , n83183 , n83184 , 
 n83185 , n83186 , n83187 , n83188 , n83189 , n83190 , n83191 , n83192 , n83193 , n83194 , 
 n83195 , n83196 , n83197 , n83198 , n83199 , n83200 , n83201 , n83202 , n83203 , n83204 , 
 n83205 , n83206 , n83207 , n83208 , n83209 , n83210 , n83211 , n83212 , n83213 , n83214 , 
 n83215 , n83216 , n83217 , n83218 , n83219 , n83220 , n83221 , n83222 , n83223 , n83224 , 
 n83225 , n83226 , n83227 , n83228 , n83229 , n83230 , n83231 , n83232 , n83233 , n83234 , 
 n83235 , n83236 , n83237 , n83238 , n83239 , n83240 , n83241 , n83242 , n83243 , n83244 , 
 n83245 , n83246 , n83247 , n83248 , n83249 , n83250 , n83251 , n83252 , n83253 , n83254 , 
 n83255 , n83256 , n83257 , n83258 , n83259 , n83260 , n83261 , n83262 , n83263 , n83264 , 
 n83265 , n83266 , n83267 , n83268 , n83269 , n83270 , n83271 , n83272 , n83273 , n83274 , 
 n83275 , n83276 , n83277 , n83278 , n83279 , n83280 , n83281 , n83282 , n83283 , n83284 , 
 n83285 , n83286 , n83287 , n83288 , n83289 , n83290 , n83291 , n83292 , n83293 , n83294 , 
 n83295 , n83296 , n83297 , n83298 , n83299 , n83300 , n83301 , n83302 , n83303 , n83304 , 
 n83305 , n83306 , n83307 , n83308 , n83309 , n83310 , n83311 , n83312 , n83313 , n83314 , 
 n83315 , n83316 , n83317 , n83318 , n83319 , n83320 , n83321 , n83322 , n83323 , n83324 , 
 n83325 , n83326 , n83327 , n83328 , n83329 , n83330 , n83331 , n83332 , n83333 , n83334 , 
 n83335 , n83336 , n83337 , n83338 , n83339 , n83340 , n83341 , n83342 , n83343 , n83344 , 
 n83345 , n83346 , n83347 , n83348 , n83349 , n83350 , n83351 , n83352 , n83353 , n83354 , 
 n83355 , n83356 , n83357 , n83358 , n83359 , n83360 , n83361 , n83362 , n83363 , n83364 , 
 n83365 , n83366 , n83367 , n83368 , n83369 , n83370 , n83371 , n83372 , n83373 , n83374 , 
 n83375 , n83376 , n83377 , n83378 , n83379 , n83380 , n83381 , n83382 , n83383 , n83384 , 
 n83385 , n83386 , n83387 , n83388 , n83389 , n83390 , n83391 , n83392 , n83393 , n83394 , 
 n83395 , n83396 , n83397 , n83398 , n83399 , n83400 , n83401 , n83402 , n83403 , n83404 , 
 n83405 , n83406 , n83407 , n83408 , n83409 , n83410 , n83411 , n83412 , n83413 , n83414 , 
 n83415 , n83416 , n83417 , n83418 , n83419 , n83420 , n83421 , n83422 , n83423 , n83424 , 
 n83425 , n83426 , n83427 , n83428 , n83429 , n83430 , n83431 , n83432 , n83433 , n83434 , 
 n83435 , n83436 , n83437 , n83438 , n83439 , n83440 , n83441 , n83442 , n83443 , n83444 , 
 n83445 , n83446 , n83447 , n83448 , n83449 , n83450 , n83451 , n83452 , n83453 , n83454 , 
 n83455 , n83456 , n83457 , n83458 , n83459 , n83460 , n83461 , n83462 , n83463 , n83464 , 
 n83465 , n83466 , n83467 , n83468 , n83469 , n83470 , n83471 , n83472 , n83473 , n83474 , 
 n83475 , n83476 , n83477 , n83478 , n83479 , n83480 , n83481 , n83482 , n83483 , n83484 , 
 n83485 , n83486 , n83487 , n83488 , n83489 , n83490 , n83491 , n83492 , n83493 , n83494 , 
 n83495 , n83496 , n83497 , n83498 , n83499 , n83500 , n83501 , n83502 , n83503 , n83504 , 
 n83505 , n83506 , n83507 , n83508 , n83509 , n83510 , n83511 , n83512 , n83513 , n83514 , 
 n83515 , n83516 , n83517 , n83518 , n83519 , n83520 , n83521 , n83522 , n83523 , n83524 , 
 n83525 , n83526 , n83527 , n83528 , n83529 , n83530 , n83531 , n83532 , n83533 , n83534 , 
 n83535 , n83536 , n83537 , n83538 , n83539 , n83540 , n83541 , n83542 , n83543 , n83544 , 
 n83545 , n83546 , n83547 , n83548 , n83549 , n83550 , n83551 , n83552 , n83553 , n83554 , 
 n83555 , n83556 , n83557 , n83558 , n83559 , n83560 , n83561 , n83562 , n83563 , n83564 , 
 n83565 , n83566 , n83567 , n83568 , n83569 , n83570 , n83571 , n83572 , n83573 , n83574 , 
 n83575 , n83576 , n83577 , n83578 , n83579 , n83580 , n83581 , n83582 , n83583 , n83584 , 
 n83585 , n83586 , n83587 , n83588 , n83589 , n83590 , n83591 , n83592 , n83593 , n83594 , 
 n83595 , n83596 , n83597 , n83598 , n83599 , n83600 , n83601 , n83602 , n83603 , n83604 , 
 n83605 , n83606 , n83607 , n83608 , n83609 , n83610 , n83611 , n83612 , n83613 , n83614 , 
 n83615 , n83616 , n83617 , n83618 , n83619 , n83620 , n83621 , n83622 , n83623 , n83624 , 
 n83625 , n83626 , n83627 , n83628 , n83629 , n83630 , n83631 , n83632 , n83633 , n83634 , 
 n83635 , n83636 , n83637 , n83638 , n83639 , n83640 , n83641 , n83642 , n83643 , n83644 , 
 n83645 , n83646 , n83647 , n83648 , n83649 , n83650 , n83651 , n83652 , n83653 , n83654 , 
 n83655 , n83656 , n83657 , n83658 , n83659 , n83660 , n83661 , n83662 , n83663 , n83664 , 
 n83665 , n83666 , n83667 , n83668 , n83669 , n83670 , n83671 , n83672 , n83673 , n83674 , 
 n83675 , n83676 , n83677 , n83678 , n83679 , n83680 , n83681 , n83682 , n83683 , n83684 , 
 n83685 , n83686 , n83687 , n83688 , n83689 , n83690 , n83691 , n83692 , n83693 , n83694 , 
 n83695 , n83696 , n83697 , n83698 , n83699 , n83700 , n83701 , n83702 , n83703 , n83704 , 
 n83705 , n83706 , n83707 , n83708 , n83709 , n83710 , n83711 , n83712 , n83713 , n83714 , 
 n83715 , n83716 , n83717 , n83718 , n83719 , n83720 , n83721 , n83722 , n83723 , n83724 , 
 n83725 , n83726 , n83727 , n83728 , n83729 , n83730 , n83731 , n83732 , n83733 , n83734 , 
 n83735 , n83736 , n83737 , n83738 , n83739 , n83740 , n83741 , n83742 , n83743 , n83744 , 
 n83745 , n83746 , n83747 , n83748 , n83749 , n83750 , n83751 , n83752 , n83753 , n83754 , 
 n83755 , n83756 , n83757 , n83758 , n83759 , n83760 , n83761 , n83762 , n83763 , n83764 , 
 n83765 , n83766 , n83767 , n83768 , n83769 , n83770 , n83771 , n83772 , n83773 , n83774 , 
 n83775 , n83776 , n83777 , n83778 , n83779 , n83780 , n83781 , n83782 , n83783 , n83784 , 
 n83785 , n83786 , n83787 , n83788 , n83789 , n83790 , n83791 , n83792 , n83793 , n83794 , 
 n83795 , n83796 , n83797 , n83798 , n83799 , n83800 , n83801 , n83802 , n83803 , n83804 , 
 n83805 , n83806 , n83807 , n83808 , n83809 , n83810 , n83811 , n83812 , n83813 , n83814 , 
 n83815 , n83816 , n83817 , n83818 , n83819 , n83820 , n83821 , n83822 , n83823 , n83824 , 
 n83825 , n83826 , n83827 , n83828 , n83829 , n83830 , n83831 , n83832 , n83833 , n83834 , 
 n83835 , n83836 , n83837 , n83838 , n83839 , n83840 , n83841 , n83842 , n83843 , n83844 , 
 n83845 , n83846 , n83847 , n83848 , n83849 , n83850 , n83851 , n83852 , n83853 , n83854 , 
 n83855 , n83856 , n83857 , n83858 , n83859 , n83860 , n83861 , n83862 , n83863 , n83864 , 
 n83865 , n83866 , n83867 , n83868 , n83869 , n83870 , n83871 , n83872 , n83873 , n83874 , 
 n83875 , n83876 , n83877 , n83878 , n83879 , n83880 , n83881 , n83882 , n83883 , n83884 , 
 n83885 , n83886 , n83887 , n83888 , n83889 , n83890 , n83891 , n83892 , n83893 , n83894 , 
 n83895 , n83896 , n83897 , n83898 , n83899 , n83900 , n83901 , n83902 , n83903 , n83904 , 
 n83905 , n83906 , n83907 , n83908 , n83909 , n83910 , n83911 , n83912 , n83913 , n83914 , 
 n83915 , n83916 , n83917 , n83918 , n83919 , n83920 , n83921 , n83922 , n83923 , n83924 , 
 n83925 , n83926 , n83927 , n83928 , n83929 , n83930 , n83931 , n83932 , n83933 , n83934 , 
 n83935 , n83936 , n83937 , n83938 , n83939 , n83940 , n83941 , n83942 , n83943 , n83944 , 
 n83945 , n83946 , n83947 , n83948 , n83949 , n83950 , n83951 , n83952 , n83953 , n83954 , 
 n83955 , n83956 , n83957 , n83958 , n83959 , n83960 , n83961 , n83962 , n83963 , n83964 , 
 n83965 , n83966 , n83967 , n83968 , n83969 , n83970 , n83971 , n83972 , n83973 , n83974 , 
 n83975 , n83976 , n83977 , n83978 , n83979 , n83980 , n83981 , n83982 , n83983 , n83984 , 
 n83985 , n83986 , n83987 , n83988 , n83989 , n83990 , n83991 , n83992 , n83993 , n83994 , 
 n83995 , n83996 , n83997 , n83998 , n83999 , n84000 , n84001 , n84002 , n84003 , n84004 , 
 n84005 , n84006 , n84007 , n84008 , n84009 , n84010 , n84011 , n84012 , n84013 , n84014 , 
 n84015 , n84016 , n84017 , n84018 , n84019 , n84020 , n84021 , n84022 , n84023 , n84024 , 
 n84025 , n84026 , n84027 , n84028 , n84029 , n84030 , n84031 , n84032 , n84033 , n84034 , 
 n84035 , n84036 , n84037 , n84038 , n84039 , n84040 , n84041 , n84042 , n84043 , n84044 , 
 n84045 , n84046 , n84047 , n84048 , n84049 , n84050 , n84051 , n84052 , n84053 , n84054 , 
 n84055 , n84056 , n84057 , n84058 , n84059 , n84060 , n84061 , n84062 , n84063 , n84064 , 
 n84065 , n84066 , n84067 , n84068 , n84069 , n84070 , n84071 , n84072 , n84073 , n84074 , 
 n84075 , n84076 , n84077 , n84078 , n84079 , n84080 , n84081 , n84082 , n84083 , n84084 , 
 n84085 , n84086 , n84087 , n84088 , n84089 , n84090 , n84091 , n84092 , n84093 , n84094 , 
 n84095 , n84096 , n84097 , n84098 , n84099 , n84100 , n84101 , n84102 , n84103 , n84104 , 
 n84105 , n84106 , n84107 , n84108 , n84109 , n84110 , n84111 , n84112 , n84113 , n84114 , 
 n84115 , n84116 , n84117 , n84118 , n84119 , n84120 , n84121 , n84122 , n84123 , n84124 , 
 n84125 , n84126 , n84127 , n84128 , n84129 , n84130 , n84131 , n84132 , n84133 , n84134 , 
 n84135 , n84136 , n84137 , n84138 , n84139 , n84140 , n84141 , n84142 , n84143 , n84144 , 
 n84145 , n84146 , n84147 , n84148 , n84149 , n84150 , n84151 , n84152 , n84153 , n84154 , 
 n84155 , n84156 , n84157 , n84158 , n84159 , n84160 , n84161 , n84162 , n84163 , n84164 , 
 n84165 , n84166 , n84167 , n84168 , n84169 , n84170 , n84171 , n84172 , n84173 , n84174 , 
 n84175 , n84176 , n84177 , n84178 , n84179 , n84180 , n84181 , n84182 , n84183 , n84184 , 
 n84185 , n84186 , n84187 , n84188 , n84189 , n84190 , n84191 , n84192 , n84193 , n84194 , 
 n84195 , n84196 , n84197 , n84198 , n84199 , n84200 , n84201 , n84202 , n84203 , n84204 , 
 n84205 , n84206 , n84207 , n84208 , n84209 , n84210 , n84211 , n84212 , n84213 , n84214 , 
 n84215 , n84216 , n84217 , n84218 , n84219 , n84220 , n84221 , n84222 , n84223 , n84224 , 
 n84225 , n84226 , n84227 , n84228 , n84229 , n84230 , n84231 , n84232 , n84233 , n84234 , 
 n84235 , n84236 , n84237 , n84238 , n84239 , n84240 , n84241 , n84242 , n84243 , n84244 , 
 n84245 , n84246 , n84247 , n84248 , n84249 , n84250 , n84251 , n84252 , n84253 , n84254 , 
 n84255 , n84256 , n84257 , n84258 , n84259 , n84260 , n84261 , n84262 , n84263 , n84264 , 
 n84265 , n84266 , n84267 , n84268 , n84269 , n84270 , n84271 , n84272 , n84273 , n84274 , 
 n84275 , n84276 , n84277 , n84278 , n84279 , n84280 , n84281 , n84282 , n84283 , n84284 , 
 n84285 , n84286 , n84287 , n84288 , n84289 , n84290 , n84291 , n84292 , n84293 , n84294 , 
 n84295 , n84296 , n84297 , n84298 , n84299 , n84300 , n84301 , n84302 , n84303 , n84304 , 
 n84305 , n84306 , n84307 , n84308 , n84309 , n84310 , n84311 , n84312 , n84313 , n84314 , 
 n84315 , n84316 , n84317 , n84318 , n84319 , n84320 , n84321 , n84322 , n84323 , n84324 , 
 n84325 , n84326 , n84327 , n84328 , n84329 , n84330 , n84331 , n84332 , n84333 , n84334 , 
 n84335 , n84336 , n84337 , n84338 , n84339 , n84340 , n84341 , n84342 , n84343 , n84344 , 
 n84345 , n84346 , n84347 , n84348 , n84349 , n84350 , n84351 , n84352 , n84353 , n84354 , 
 n84355 , n84356 , n84357 , n84358 , n84359 , n84360 , n84361 , n84362 , n84363 , n84364 , 
 n84365 , n84366 , n84367 , n84368 , n84369 , n84370 , n84371 , n84372 , n84373 , n84374 , 
 n84375 , n84376 , n84377 , n84378 , n84379 , n84380 , n84381 , n84382 , n84383 , n84384 , 
 n84385 , n84386 , n84387 , n84388 , n84389 , n84390 , n84391 , n84392 , n84393 , n84394 , 
 n84395 , n84396 , n84397 , n84398 , n84399 , n84400 , n84401 , n84402 , n84403 , n84404 , 
 n84405 , n84406 , n84407 , n84408 , n84409 , n84410 , n84411 , n84412 , n84413 , n84414 , 
 n84415 , n84416 , n84417 , n84418 , n84419 , n84420 , n84421 , n84422 , n84423 , n84424 , 
 n84425 , n84426 , n84427 , n84428 , n84429 , n84430 , n84431 , n84432 , n84433 , n84434 , 
 n84435 , n84436 , n84437 , n84438 , n84439 , n84440 , n84441 , n84442 , n84443 , n84444 , 
 n84445 , n84446 , n84447 , n84448 , n84449 , n84450 , n84451 , n84452 , n84453 , n84454 , 
 n84455 , n84456 , n84457 , n84458 , n84459 , n84460 , n84461 , n84462 , n84463 , n84464 , 
 n84465 , n84466 , n84467 , n84468 , n84469 , n84470 , n84471 , n84472 , n84473 , n84474 , 
 n84475 , n84476 , n84477 , n84478 , n84479 , n84480 , n84481 , n84482 , n84483 , n84484 , 
 n84485 , n84486 , n84487 , n84488 , n84489 , n84490 , n84491 , n84492 , n84493 , n84494 , 
 n84495 , n84496 , n84497 , n84498 , n84499 , n84500 , n84501 , n84502 , n84503 , n84504 , 
 n84505 , n84506 , n84507 , n84508 , n84509 , n84510 , n84511 , n84512 , n84513 , n84514 , 
 n84515 , n84516 , n84517 , n84518 , n84519 , n84520 , n84521 , n84522 , n84523 , n84524 , 
 n84525 , n84526 , n84527 , n84528 , n84529 , n84530 , n84531 , n84532 , n84533 , n84534 , 
 n84535 , n84536 , n84537 , n84538 , n84539 , n84540 , n84541 , n84542 , n84543 , n84544 , 
 n84545 , n84546 , n84547 , n84548 , n84549 , n84550 , n84551 , n84552 , n84553 , n84554 , 
 n84555 , n84556 , n84557 , n84558 , n84559 , n84560 , n84561 , n84562 , n84563 , n84564 , 
 n84565 , n84566 , n84567 , n84568 , n84569 , n84570 , n84571 , n84572 , n84573 , n84574 , 
 n84575 , n84576 , n84577 , n84578 , n84579 , n84580 , n84581 , n84582 , n84583 , n84584 , 
 n84585 , n84586 , n84587 , n84588 , n84589 , n84590 , n84591 , n84592 , n84593 , n84594 , 
 n84595 , n84596 , n84597 , n84598 , n84599 , n84600 , n84601 , n84602 , n84603 , n84604 , 
 n84605 , n84606 , n84607 , n84608 , n84609 , n84610 , n84611 , n84612 , n84613 , n84614 , 
 n84615 , n84616 , n84617 , n84618 , n84619 , n84620 , n84621 , n84622 , n84623 , n84624 , 
 n84625 , n84626 , n84627 , n84628 , n84629 , n84630 , n84631 , n84632 , n84633 , n84634 , 
 n84635 , n84636 , n84637 , n84638 , n84639 , n84640 , n84641 , n84642 , n84643 , n84644 , 
 n84645 , n84646 , n84647 , n84648 , n84649 , n84650 , n84651 , n84652 , n84653 , n84654 , 
 n84655 , n84656 , n84657 , n84658 , n84659 , n84660 , n84661 , n84662 , n84663 , n84664 , 
 n84665 , n84666 , n84667 , n84668 , n84669 , n84670 , n84671 , n84672 , n84673 , n84674 , 
 n84675 , n84676 , n84677 , n84678 , n84679 , n84680 , n84681 , n84682 , n84683 , n84684 , 
 n84685 , n84686 , n84687 , n84688 , n84689 , n84690 , n84691 , n84692 , n84693 , n84694 , 
 n84695 , n84696 , n84697 , n84698 , n84699 , n84700 , n84701 , n84702 , n84703 , n84704 , 
 n84705 , n84706 , n84707 , n84708 , n84709 , n84710 , n84711 , n84712 , n84713 , n84714 , 
 n84715 , n84716 , n84717 , n84718 , n84719 , n84720 , n84721 , n84722 , n84723 , n84724 , 
 n84725 , n84726 , n84727 , n84728 , n84729 , n84730 , n84731 , n84732 , n84733 , n84734 , 
 n84735 , n84736 , n84737 , n84738 , n84739 , n84740 , n84741 , n84742 , n84743 , n84744 , 
 n84745 , n84746 , n84747 , n84748 , n84749 , n84750 , n84751 , n84752 , n84753 , n84754 , 
 n84755 , n84756 , n84757 , n84758 , n84759 , n84760 , n84761 , n84762 , n84763 , n84764 , 
 n84765 , n84766 , n84767 , n84768 , n84769 , n84770 , n84771 , n84772 , n84773 , n84774 , 
 n84775 , n84776 , n84777 , n84778 , n84779 , n84780 , n84781 , n84782 , n84783 , n84784 , 
 n84785 , n84786 , n84787 , n84788 , n84789 , n84790 , n84791 , n84792 , n84793 , n84794 , 
 n84795 , n84796 , n84797 , n84798 , n84799 , n84800 , n84801 , n84802 , n84803 , n84804 , 
 n84805 , n84806 , n84807 , n84808 , n84809 , n84810 , n84811 , n84812 , n84813 , n84814 , 
 n84815 , n84816 , n84817 , n84818 , n84819 , n84820 , n84821 , n84822 , n84823 , n84824 , 
 n84825 , n84826 , n84827 , n84828 , n84829 , n84830 , n84831 , n84832 , n84833 , n84834 , 
 n84835 , n84836 , n84837 , n84838 , n84839 , n84840 , n84841 , n84842 , n84843 , n84844 , 
 n84845 , n84846 , n84847 , n84848 , n84849 , n84850 , n84851 , n84852 , n84853 , n84854 , 
 n84855 , n84856 , n84857 , n84858 , n84859 , n84860 , n84861 , n84862 , n84863 , n84864 , 
 n84865 , n84866 , n84867 , n84868 , n84869 , n84870 , n84871 , n84872 , n84873 , n84874 , 
 n84875 , n84876 , n84877 , n84878 , n84879 , n84880 , n84881 , n84882 , n84883 , n84884 , 
 n84885 , n84886 , n84887 , n84888 , n84889 , n84890 , n84891 , n84892 , n84893 , n84894 , 
 n84895 , n84896 , n84897 , n84898 , n84899 , n84900 , n84901 , n84902 , n84903 , n84904 , 
 n84905 , n84906 , n84907 , n84908 , n84909 , n84910 , n84911 , n84912 , n84913 , n84914 , 
 n84915 , n84916 , n84917 , n84918 , n84919 , n84920 , n84921 , n84922 , n84923 , n84924 , 
 n84925 , n84926 , n84927 , n84928 , n84929 , n84930 , n84931 , n84932 , n84933 , n84934 , 
 n84935 , n84936 , n84937 , n84938 , n84939 , n84940 , n84941 , n84942 , n84943 , n84944 , 
 n84945 , n84946 , n84947 , n84948 , n84949 , n84950 , n84951 , n84952 , n84953 , n84954 , 
 n84955 , n84956 , n84957 , n84958 , n84959 , n84960 , n84961 , n84962 , n84963 , n84964 , 
 n84965 , n84966 , n84967 , n84968 , n84969 , n84970 , n84971 , n84972 , n84973 , n84974 , 
 n84975 , n84976 , n84977 , n84978 , n84979 , n84980 , n84981 , n84982 , n84983 , n84984 , 
 n84985 , n84986 , n84987 , n84988 , n84989 , n84990 , n84991 , n84992 , n84993 , n84994 , 
 n84995 , n84996 , n84997 , n84998 , n84999 , n85000 , n85001 , n85002 , n85003 , n85004 , 
 n85005 , n85006 , n85007 , n85008 , n85009 , n85010 , n85011 , n85012 , n85013 , n85014 , 
 n85015 , n85016 , n85017 , n85018 , n85019 , n85020 , n85021 , n85022 , n85023 , n85024 , 
 n85025 , n85026 , n85027 , n85028 , n85029 , n85030 , n85031 , n85032 , n85033 , n85034 , 
 n85035 , n85036 , n85037 , n85038 , n85039 , n85040 , n85041 , n85042 , n85043 , n85044 , 
 n85045 , n85046 , n85047 , n85048 , n85049 , n85050 , n85051 , n85052 , n85053 , n85054 , 
 n85055 , n85056 , n85057 , n85058 , n85059 , n85060 , n85061 , n85062 , n85063 , n85064 , 
 n85065 , n85066 , n85067 , n85068 , n85069 , n85070 , n85071 , n85072 , n85073 , n85074 , 
 n85075 , n85076 , n85077 , n85078 , n85079 , n85080 , n85081 , n85082 , n85083 , n85084 , 
 n85085 , n85086 , n85087 , n85088 , n85089 , n85090 , n85091 , n85092 , n85093 , n85094 , 
 n85095 , n85096 , n85097 , n85098 , n85099 , n85100 , n85101 , n85102 , n85103 , n85104 , 
 n85105 , n85106 , n85107 , n85108 , n85109 , n85110 , n85111 , n85112 , n85113 , n85114 , 
 n85115 , n85116 , n85117 , n85118 , n85119 , n85120 , n85121 , n85122 , n85123 , n85124 , 
 n85125 , n85126 , n85127 , n85128 , n85129 , n85130 , n85131 , n85132 , n85133 , n85134 , 
 n85135 , n85136 , n85137 , n85138 , n85139 , n85140 , n85141 , n85142 , n85143 , n85144 , 
 n85145 , n85146 , n85147 , n85148 , n85149 , n85150 , n85151 , n85152 , n85153 , n85154 , 
 n85155 , n85156 , n85157 , n85158 , n85159 , n85160 , n85161 , n85162 , n85163 , n85164 , 
 n85165 , n85166 , n85167 , n85168 , n85169 , n85170 , n85171 , n85172 , n85173 , n85174 , 
 n85175 , n85176 , n85177 , n85178 , n85179 , n85180 , n85181 , n85182 , n85183 , n85184 , 
 n85185 , n85186 , n85187 , n85188 , n85189 , n85190 , n85191 , n85192 , n85193 , n85194 , 
 n85195 , n85196 , n85197 , n85198 , n85199 , n85200 , n85201 , n85202 , n85203 , n85204 , 
 n85205 , n85206 , n85207 , n85208 , n85209 , n85210 , n85211 , n85212 , n85213 , n85214 , 
 n85215 , n85216 , n85217 , n85218 , n85219 , n85220 , n85221 , n85222 , n85223 , n85224 , 
 n85225 , n85226 , n85227 , n85228 , n85229 , n85230 , n85231 , n85232 , n85233 , n85234 , 
 n85235 , n85236 , n85237 , n85238 , n85239 , n85240 , n85241 , n85242 , n85243 , n85244 , 
 n85245 , n85246 , n85247 , n85248 , n85249 , n85250 , n85251 , n85252 , n85253 , n85254 , 
 n85255 , n85256 , n85257 , n85258 , n85259 , n85260 , n85261 , n85262 , n85263 , n85264 , 
 n85265 , n85266 , n85267 , n85268 , n85269 , n85270 , n85271 , n85272 , n85273 , n85274 , 
 n85275 , n85276 , n85277 , n85278 , n85279 , n85280 , n85281 , n85282 , n85283 , n85284 , 
 n85285 , n85286 , n85287 , n85288 , n85289 , n85290 , n85291 , n85292 , n85293 , n85294 , 
 n85295 , n85296 , n85297 , n85298 , n85299 , n85300 , n85301 , n85302 , n85303 , n85304 , 
 n85305 , n85306 , n85307 , n85308 , n85309 , n85310 , n85311 , n85312 , n85313 , n85314 , 
 n85315 , n85316 , n85317 , n85318 , n85319 , n85320 , n85321 , n85322 , n85323 , n85324 , 
 n85325 , n85326 , n85327 , n85328 , n85329 , n85330 , n85331 , n85332 , n85333 , n85334 , 
 n85335 , n85336 , n85337 , n85338 , n85339 , n85340 , n85341 , n85342 , n85343 , n85344 , 
 n85345 , n85346 , n85347 , n85348 , n85349 , n85350 , n85351 , n85352 , n85353 , n85354 , 
 n85355 , n85356 , n85357 , n85358 , n85359 , n85360 , n85361 , n85362 , n85363 , n85364 , 
 n85365 , n85366 , n85367 , n85368 , n85369 , n85370 , n85371 , n85372 , n85373 , n85374 , 
 n85375 , n85376 , n85377 , n85378 , n85379 , n85380 , n85381 , n85382 , n85383 , n85384 , 
 n85385 , n85386 , n85387 , n85388 , n85389 , n85390 , n85391 , n85392 , n85393 , n85394 , 
 n85395 , n85396 , n85397 , n85398 , n85399 , n85400 , n85401 , n85402 , n85403 , n85404 , 
 n85405 , n85406 , n85407 , n85408 , n85409 , n85410 , n85411 , n85412 , n85413 , n85414 , 
 n85415 , n85416 , n85417 , n85418 , n85419 , n85420 , n85421 , n85422 , n85423 , n85424 , 
 n85425 , n85426 , n85427 , n85428 , n85429 , n85430 , n85431 , n85432 , n85433 , n85434 , 
 n85435 , n85436 , n85437 , n85438 , n85439 , n85440 , n85441 , n85442 , n85443 , n85444 , 
 n85445 , n85446 , n85447 , n85448 , n85449 , n85450 , n85451 , n85452 , n85453 , n85454 , 
 n85455 , n85456 , n85457 , n85458 , n85459 , n85460 , n85461 , n85462 , n85463 , n85464 , 
 n85465 , n85466 , n85467 , n85468 , n85469 , n85470 , n85471 , n85472 , n85473 , n85474 , 
 n85475 , n85476 , n85477 , n85478 , n85479 , n85480 , n85481 , n85482 , n85483 , n85484 , 
 n85485 , n85486 , n85487 , n85488 , n85489 , n85490 , n85491 , n85492 , n85493 , n85494 , 
 n85495 , n85496 , n85497 , n85498 , n85499 , n85500 , n85501 , n85502 , n85503 , n85504 , 
 n85505 , n85506 , n85507 , n85508 , n85509 , n85510 , n85511 , n85512 , n85513 , n85514 , 
 n85515 , n85516 , n85517 , n85518 , n85519 , n85520 , n85521 , n85522 , n85523 , n85524 , 
 n85525 , n85526 , n85527 , n85528 , n85529 , n85530 , n85531 , n85532 , n85533 , n85534 , 
 n85535 , n85536 , n85537 , n85538 , n85539 , n85540 , n85541 , n85542 , n85543 , n85544 , 
 n85545 , n85546 , n85547 , n85548 , n85549 , n85550 , n85551 , n85552 , n85553 , n85554 , 
 n85555 , n85556 , n85557 , n85558 , n85559 , n85560 , n85561 , n85562 , n85563 , n85564 , 
 n85565 , n85566 , n85567 , n85568 , n85569 , n85570 , n85571 , n85572 , n85573 , n85574 , 
 n85575 , n85576 , n85577 , n85578 , n85579 , n85580 , n85581 , n85582 , n85583 , n85584 , 
 n85585 , n85586 , n85587 , n85588 , n85589 , n85590 , n85591 , n85592 , n85593 , n85594 , 
 n85595 , n85596 , n85597 , n85598 , n85599 , n85600 , n85601 , n85602 , n85603 , n85604 , 
 n85605 , n85606 , n85607 , n85608 , n85609 , n85610 , n85611 , n85612 , n85613 , n85614 , 
 n85615 , n85616 , n85617 , n85618 , n85619 , n85620 , n85621 , n85622 , n85623 , n85624 , 
 n85625 , n85626 , n85627 , n85628 , n85629 , n85630 , n85631 , n85632 , n85633 , n85634 , 
 n85635 , n85636 , n85637 , n85638 , n85639 , n85640 , n85641 , n85642 , n85643 , n85644 , 
 n85645 , n85646 , n85647 , n85648 , n85649 , n85650 , n85651 , n85652 , n85653 , n85654 , 
 n85655 , n85656 , n85657 , n85658 , n85659 , n85660 , n85661 , n85662 , n85663 , n85664 , 
 n85665 , n85666 , n85667 , n85668 , n85669 , n85670 , n85671 , n85672 , n85673 , n85674 , 
 n85675 , n85676 , n85677 , n85678 , n85679 , n85680 , n85681 , n85682 , n85683 , n85684 , 
 n85685 , n85686 , n85687 , n85688 , n85689 , n85690 , n85691 , n85692 , n85693 , n85694 , 
 n85695 , n85696 , n85697 , n85698 , n85699 , n85700 , n85701 , n85702 , n85703 , n85704 , 
 n85705 , n85706 , n85707 , n85708 , n85709 , n85710 , n85711 , n85712 , n85713 , n85714 , 
 n85715 , n85716 , n85717 , n85718 , n85719 , n85720 , n85721 , n85722 , n85723 , n85724 , 
 n85725 , n85726 , n85727 , n85728 , n85729 , n85730 , n85731 , n85732 , n85733 , n85734 , 
 n85735 , n85736 , n85737 , n85738 , n85739 , n85740 , n85741 , n85742 , n85743 , n85744 , 
 n85745 , n85746 , n85747 , n85748 , n85749 , n85750 , n85751 , n85752 , n85753 , n85754 , 
 n85755 , n85756 , n85757 , n85758 , n85759 , n85760 , n85761 , n85762 , n85763 , n85764 , 
 n85765 , n85766 , n85767 , n85768 , n85769 , n85770 , n85771 , n85772 , n85773 , n85774 , 
 n85775 , n85776 , n85777 , n85778 , n85779 , n85780 , n85781 , n85782 , n85783 , n85784 , 
 n85785 , n85786 , n85787 , n85788 , n85789 , n85790 , n85791 , n85792 , n85793 , n85794 , 
 n85795 , n85796 , n85797 , n85798 , n85799 , n85800 , n85801 , n85802 , n85803 , n85804 , 
 n85805 , n85806 , n85807 , n85808 , n85809 , n85810 , n85811 , n85812 , n85813 , n85814 , 
 n85815 , n85816 , n85817 , n85818 , n85819 , n85820 , n85821 , n85822 , n85823 , n85824 , 
 n85825 , n85826 , n85827 , n85828 , n85829 , n85830 , n85831 , n85832 , n85833 , n85834 , 
 n85835 , n85836 , n85837 , n85838 , n85839 , n85840 , n85841 , n85842 , n85843 , n85844 , 
 n85845 , n85846 , n85847 , n85848 , n85849 , n85850 , n85851 , n85852 , n85853 , n85854 , 
 n85855 , n85856 , n85857 , n85858 , n85859 , n85860 , n85861 , n85862 , n85863 , n85864 , 
 n85865 , n85866 , n85867 , n85868 , n85869 , n85870 , n85871 , n85872 , n85873 , n85874 , 
 n85875 , n85876 , n85877 , n85878 , n85879 , n85880 , n85881 , n85882 , n85883 , n85884 , 
 n85885 , n85886 , n85887 , n85888 , n85889 , n85890 , n85891 , n85892 , n85893 , n85894 , 
 n85895 , n85896 , n85897 , n85898 , n85899 , n85900 , n85901 , n85902 , n85903 , n85904 , 
 n85905 , n85906 , n85907 , n85908 , n85909 , n85910 , n85911 , n85912 , n85913 , n85914 , 
 n85915 , n85916 , n85917 , n85918 , n85919 , n85920 , n85921 , n85922 , n85923 , n85924 , 
 n85925 , n85926 , n85927 , n85928 , n85929 , n85930 , n85931 , n85932 , n85933 , n85934 , 
 n85935 , n85936 , n85937 , n85938 , n85939 , n85940 , n85941 , n85942 , n85943 , n85944 , 
 n85945 , n85946 , n85947 , n85948 , n85949 , n85950 , n85951 , n85952 , n85953 , n85954 , 
 n85955 , n85956 , n85957 , n85958 , n85959 , n85960 , n85961 , n85962 , n85963 , n85964 , 
 n85965 , n85966 , n85967 , n85968 , n85969 , n85970 , n85971 , n85972 , n85973 , n85974 , 
 n85975 , n85976 , n85977 , n85978 , n85979 , n85980 , n85981 , n85982 , n85983 , n85984 , 
 n85985 , n85986 , n85987 , n85988 , n85989 , n85990 , n85991 , n85992 , n85993 , n85994 , 
 n85995 , n85996 , n85997 , n85998 , n85999 , n86000 , n86001 , n86002 , n86003 , n86004 , 
 n86005 , n86006 , n86007 , n86008 , n86009 , n86010 , n86011 , n86012 , n86013 , n86014 , 
 n86015 , n86016 , n86017 , n86018 , n86019 , n86020 , n86021 , n86022 , n86023 , n86024 , 
 n86025 , n86026 , n86027 , n86028 , n86029 , n86030 , n86031 , n86032 , n86033 , n86034 , 
 n86035 , n86036 , n86037 , n86038 , n86039 , n86040 , n86041 , n86042 , n86043 , n86044 , 
 n86045 , n86046 , n86047 , n86048 , n86049 , n86050 , n86051 , n86052 , n86053 , n86054 , 
 n86055 , n86056 , n86057 , n86058 , n86059 , n86060 , n86061 , n86062 , n86063 , n86064 , 
 n86065 , n86066 , n86067 , n86068 , n86069 , n86070 , n86071 , n86072 , n86073 , n86074 , 
 n86075 , n86076 , n86077 , n86078 , n86079 , n86080 , n86081 , n86082 , n86083 , n86084 , 
 n86085 , n86086 , n86087 , n86088 , n86089 , n86090 , n86091 , n86092 , n86093 , n86094 , 
 n86095 , n86096 , n86097 , n86098 , n86099 , n86100 , n86101 , n86102 , n86103 , n86104 , 
 n86105 , n86106 , n86107 , n86108 , n86109 , n86110 , n86111 , n86112 , n86113 , n86114 , 
 n86115 , n86116 , n86117 , n86118 , n86119 , n86120 , n86121 , n86122 , n86123 , n86124 , 
 n86125 , n86126 , n86127 , n86128 , n86129 , n86130 , n86131 , n86132 , n86133 , n86134 , 
 n86135 , n86136 , n86137 , n86138 , n86139 , n86140 , n86141 , n86142 , n86143 , n86144 , 
 n86145 , n86146 , n86147 , n86148 , n86149 , n86150 , n86151 , n86152 , n86153 , n86154 , 
 n86155 , n86156 , n86157 , n86158 , n86159 , n86160 , n86161 , n86162 , n86163 , n86164 , 
 n86165 , n86166 , n86167 , n86168 , n86169 , n86170 , n86171 , n86172 , n86173 , n86174 , 
 n86175 , n86176 , n86177 , n86178 , n86179 , n86180 , n86181 , n86182 , n86183 , n86184 , 
 n86185 , n86186 , n86187 , n86188 , n86189 , n86190 , n86191 , n86192 , n86193 , n86194 , 
 n86195 , n86196 , n86197 , n86198 , n86199 , n86200 , n86201 , n86202 , n86203 , n86204 , 
 n86205 , n86206 , n86207 , n86208 , n86209 , n86210 , n86211 , n86212 , n86213 , n86214 , 
 n86215 , n86216 , n86217 , n86218 , n86219 , n86220 , n86221 , n86222 , n86223 , n86224 , 
 n86225 , n86226 , n86227 , n86228 , n86229 , n86230 , n86231 , n86232 , n86233 , n86234 , 
 n86235 , n86236 , n86237 , n86238 , n86239 , n86240 , n86241 , n86242 , n86243 , n86244 , 
 n86245 , n86246 , n86247 , n86248 , n86249 , n86250 , n86251 , n86252 , n86253 , n86254 , 
 n86255 , n86256 , n86257 , n86258 , n86259 , n86260 , n86261 , n86262 , n86263 , n86264 , 
 n86265 , n86266 , n86267 , n86268 , n86269 , n86270 , n86271 , n86272 , n86273 , n86274 , 
 n86275 , n86276 , n86277 , n86278 , n86279 , n86280 , n86281 , n86282 , n86283 , n86284 , 
 n86285 , n86286 , n86287 , n86288 , n86289 , n86290 , n86291 , n86292 , n86293 , n86294 , 
 n86295 , n86296 , n86297 , n86298 , n86299 , n86300 , n86301 , n86302 , n86303 , n86304 , 
 n86305 , n86306 , n86307 , n86308 , n86309 , n86310 , n86311 , n86312 , n86313 , n86314 , 
 n86315 , n86316 , n86317 , n86318 , n86319 , n86320 , n86321 , n86322 , n86323 , n86324 , 
 n86325 , n86326 , n86327 , n86328 , n86329 , n86330 , n86331 , n86332 , n86333 , n86334 , 
 n86335 , n86336 , n86337 , n86338 , n86339 , n86340 , n86341 , n86342 , n86343 , n86344 , 
 n86345 , n86346 , n86347 , n86348 , n86349 , n86350 , n86351 , n86352 , n86353 , n86354 , 
 n86355 , n86356 , n86357 , n86358 , n86359 , n86360 , n86361 , n86362 , n86363 , n86364 , 
 n86365 , n86366 , n86367 , n86368 , n86369 , n86370 , n86371 , n86372 , n86373 , n86374 , 
 n86375 , n86376 , n86377 , n86378 , n86379 , n86380 , n86381 , n86382 , n86383 , n86384 , 
 n86385 , n86386 , n86387 , n86388 , n86389 , n86390 , n86391 , n86392 , n86393 , n86394 , 
 n86395 , n86396 , n86397 , n86398 , n86399 , n86400 , n86401 , n86402 , n86403 , n86404 , 
 n86405 , n86406 , n86407 , n86408 , n86409 , n86410 , n86411 , n86412 , n86413 , n86414 , 
 n86415 , n86416 , n86417 , n86418 , n86419 , n86420 , n86421 , n86422 , n86423 , n86424 , 
 n86425 , n86426 , n86427 , n86428 , n86429 , n86430 , n86431 , n86432 , n86433 , n86434 , 
 n86435 , n86436 , n86437 , n86438 , n86439 , n86440 , n86441 , n86442 , n86443 , n86444 , 
 n86445 , n86446 , n86447 , n86448 , n86449 , n86450 , n86451 , n86452 , n86453 , n86454 , 
 n86455 , n86456 , n86457 , n86458 , n86459 , n86460 , n86461 , n86462 , n86463 , n86464 , 
 n86465 , n86466 , n86467 , n86468 , n86469 , n86470 , n86471 , n86472 , n86473 , n86474 , 
 n86475 , n86476 , n86477 , n86478 , n86479 , n86480 , n86481 , n86482 , n86483 , n86484 , 
 n86485 , n86486 , n86487 , n86488 , n86489 , n86490 , n86491 , n86492 , n86493 , n86494 , 
 n86495 , n86496 , n86497 , n86498 , n86499 , n86500 , n86501 , n86502 , n86503 , n86504 , 
 n86505 , n86506 , n86507 , n86508 , n86509 , n86510 , n86511 , n86512 , n86513 , n86514 , 
 n86515 , n86516 , n86517 , n86518 , n86519 , n86520 , n86521 , n86522 , n86523 , n86524 , 
 n86525 , n86526 , n86527 , n86528 , n86529 , n86530 , n86531 , n86532 , n86533 , n86534 , 
 n86535 , n86536 , n86537 , n86538 , n86539 , n86540 , n86541 , n86542 , n86543 , n86544 , 
 n86545 , n86546 , n86547 , n86548 , n86549 , n86550 , n86551 , n86552 , n86553 , n86554 , 
 n86555 , n86556 , n86557 , n86558 , n86559 , n86560 , n86561 , n86562 , n86563 , n86564 , 
 n86565 , n86566 , n86567 , n86568 , n86569 , n86570 , n86571 , n86572 , n86573 , n86574 , 
 n86575 , n86576 , n86577 , n86578 , n86579 , n86580 , n86581 , n86582 , n86583 , n86584 , 
 n86585 , n86586 , n86587 , n86588 , n86589 , n86590 , n86591 , n86592 , n86593 , n86594 , 
 n86595 , n86596 , n86597 , n86598 , n86599 , n86600 , n86601 , n86602 , n86603 , n86604 , 
 n86605 , n86606 , n86607 , n86608 , n86609 , n86610 , n86611 , n86612 , n86613 , n86614 , 
 n86615 , n86616 , n86617 , n86618 , n86619 , n86620 , n86621 , n86622 , n86623 , n86624 , 
 n86625 , n86626 , n86627 , n86628 , n86629 , n86630 , n86631 , n86632 , n86633 , n86634 , 
 n86635 , n86636 , n86637 , n86638 , n86639 , n86640 , n86641 , n86642 , n86643 , n86644 , 
 n86645 , n86646 , n86647 , n86648 , n86649 , n86650 , n86651 , n86652 , n86653 , n86654 , 
 n86655 , n86656 , n86657 , n86658 , n86659 , n86660 , n86661 , n86662 , n86663 , n86664 , 
 n86665 , n86666 , n86667 , n86668 , n86669 , n86670 , n86671 , n86672 , n86673 , n86674 , 
 n86675 , n86676 , n86677 , n86678 , n86679 , n86680 , n86681 , n86682 , n86683 , n86684 , 
 n86685 , n86686 , n86687 , n86688 , n86689 , n86690 , n86691 , n86692 , n86693 , n86694 , 
 n86695 , n86696 , n86697 , n86698 , n86699 , n86700 , n86701 , n86702 , n86703 , n86704 , 
 n86705 , n86706 , n86707 , n86708 , n86709 , n86710 , n86711 , n86712 , n86713 , n86714 , 
 n86715 , n86716 , n86717 , n86718 , n86719 , n86720 , n86721 , n86722 , n86723 , n86724 , 
 n86725 , n86726 , n86727 , n86728 , n86729 , n86730 , n86731 , n86732 , n86733 , n86734 , 
 n86735 , n86736 , n86737 , n86738 , n86739 , n86740 , n86741 , n86742 , n86743 , n86744 , 
 n86745 , n86746 , n86747 , n86748 , n86749 , n86750 , n86751 , n86752 , n86753 , n86754 , 
 n86755 , n86756 , n86757 , n86758 , n86759 , n86760 , n86761 , n86762 , n86763 , n86764 , 
 n86765 , n86766 , n86767 , n86768 , n86769 , n86770 , n86771 , n86772 , n86773 , n86774 , 
 n86775 , n86776 , n86777 , n86778 , n86779 , n86780 , n86781 , n86782 , n86783 , n86784 , 
 n86785 , n86786 , n86787 , n86788 , n86789 , n86790 , n86791 , n86792 , n86793 , n86794 , 
 n86795 , n86796 , n86797 , n86798 , n86799 , n86800 , n86801 , n86802 , n86803 , n86804 , 
 n86805 , n86806 , n86807 , n86808 , n86809 , n86810 , n86811 , n86812 , n86813 , n86814 , 
 n86815 , n86816 , n86817 , n86818 , n86819 , n86820 , n86821 , n86822 , n86823 , n86824 , 
 n86825 , n86826 , n86827 , n86828 , n86829 , n86830 , n86831 , n86832 , n86833 , n86834 , 
 n86835 , n86836 , n86837 , n86838 , n86839 , n86840 , n86841 , n86842 , n86843 , n86844 , 
 n86845 , n86846 , n86847 , n86848 , n86849 , n86850 , n86851 , n86852 , n86853 , n86854 , 
 n86855 , n86856 , n86857 , n86858 , n86859 , n86860 , n86861 , n86862 , n86863 , n86864 , 
 n86865 , n86866 , n86867 , n86868 , n86869 , n86870 , n86871 , n86872 , n86873 , n86874 , 
 n86875 , n86876 , n86877 , n86878 , n86879 , n86880 , n86881 , n86882 , n86883 , n86884 , 
 n86885 , n86886 , n86887 , n86888 , n86889 , n86890 , n86891 , n86892 , n86893 , n86894 , 
 n86895 , n86896 , n86897 , n86898 , n86899 , n86900 , n86901 , n86902 , n86903 , n86904 , 
 n86905 , n86906 , n86907 , n86908 , n86909 , n86910 , n86911 , n86912 , n86913 , n86914 , 
 n86915 , n86916 , n86917 , n86918 , n86919 , n86920 , n86921 , n86922 , n86923 , n86924 , 
 n86925 , n86926 , n86927 , n86928 , n86929 , n86930 , n86931 , n86932 , n86933 , n86934 , 
 n86935 , n86936 , n86937 , n86938 , n86939 , n86940 , n86941 , n86942 , n86943 , n86944 , 
 n86945 , n86946 , n86947 , n86948 , n86949 , n86950 , n86951 , n86952 , n86953 , n86954 , 
 n86955 , n86956 , n86957 , n86958 , n86959 , n86960 , n86961 , n86962 , n86963 , n86964 , 
 n86965 , n86966 , n86967 , n86968 , n86969 , n86970 , n86971 , n86972 , n86973 , n86974 , 
 n86975 , n86976 , n86977 , n86978 , n86979 , n86980 , n86981 , n86982 , n86983 , n86984 , 
 n86985 , n86986 , n86987 , n86988 , n86989 , n86990 , n86991 , n86992 , n86993 , n86994 , 
 n86995 , n86996 , n86997 , n86998 , n86999 , n87000 , n87001 , n87002 , n87003 , n87004 , 
 n87005 , n87006 , n87007 , n87008 , n87009 , n87010 , n87011 , n87012 , n87013 , n87014 , 
 n87015 , n87016 , n87017 , n87018 , n87019 , n87020 , n87021 , n87022 , n87023 , n87024 , 
 n87025 , n87026 , n87027 , n87028 , n87029 , n87030 , n87031 , n87032 , n87033 , n87034 , 
 n87035 , n87036 , n87037 , n87038 , n87039 , n87040 , n87041 , n87042 , n87043 , n87044 , 
 n87045 , n87046 , n87047 , n87048 , n87049 , n87050 , n87051 , n87052 , n87053 , n87054 , 
 n87055 , n87056 , n87057 , n87058 , n87059 , n87060 , n87061 , n87062 , n87063 , n87064 , 
 n87065 , n87066 , n87067 , n87068 , n87069 , n87070 , n87071 , n87072 , n87073 , n87074 , 
 n87075 , n87076 , n87077 , n87078 , n87079 , n87080 , n87081 , n87082 , n87083 , n87084 , 
 n87085 , n87086 , n87087 , n87088 , n87089 , n87090 , n87091 , n87092 , n87093 , n87094 , 
 n87095 , n87096 , n87097 , n87098 , n87099 , n87100 , n87101 , n87102 , n87103 , n87104 , 
 n87105 , n87106 , n87107 , n87108 , n87109 , n87110 , n87111 , n87112 , n87113 , n87114 , 
 n87115 , n87116 , n87117 , n87118 , n87119 , n87120 , n87121 , n87122 , n87123 , n87124 , 
 n87125 , n87126 , n87127 , n87128 , n87129 , n87130 , n87131 , n87132 , n87133 , n87134 , 
 n87135 , n87136 , n87137 , n87138 , n87139 , n87140 , n87141 , n87142 , n87143 , n87144 , 
 n87145 , n87146 , n87147 , n87148 , n87149 , n87150 , n87151 , n87152 , n87153 , n87154 , 
 n87155 , n87156 , n87157 , n87158 , n87159 , n87160 , n87161 , n87162 , n87163 , n87164 , 
 n87165 , n87166 , n87167 , n87168 , n87169 , n87170 , n87171 , n87172 , n87173 , n87174 , 
 n87175 , n87176 , n87177 , n87178 , n87179 , n87180 , n87181 , n87182 , n87183 , n87184 , 
 n87185 , n87186 , n87187 , n87188 , n87189 , n87190 , n87191 , n87192 , n87193 , n87194 , 
 n87195 , n87196 , n87197 , n87198 , n87199 , n87200 , n87201 , n87202 , n87203 , n87204 , 
 n87205 , n87206 , n87207 , n87208 , n87209 , n87210 , n87211 , n87212 , n87213 , n87214 , 
 n87215 , n87216 , n87217 , n87218 , n87219 , n87220 , n87221 , n87222 , n87223 , n87224 , 
 n87225 , n87226 , n87227 , n87228 , n87229 , n87230 , n87231 , n87232 , n87233 , n87234 , 
 n87235 , n87236 , n87237 , n87238 , n87239 , n87240 , n87241 , n87242 , n87243 , n87244 , 
 n87245 , n87246 , n87247 , n87248 , n87249 , n87250 , n87251 , n87252 , n87253 , n87254 , 
 n87255 , n87256 , n87257 , n87258 , n87259 , n87260 , n87261 , n87262 , n87263 , n87264 , 
 n87265 , n87266 , n87267 , n87268 , n87269 , n87270 , n87271 , n87272 , n87273 , n87274 , 
 n87275 , n87276 , n87277 , n87278 , n87279 , n87280 , n87281 , n87282 , n87283 , n87284 , 
 n87285 , n87286 , n87287 , n87288 , n87289 , n87290 , n87291 , n87292 , n87293 , n87294 , 
 n87295 , n87296 , n87297 , n87298 , n87299 , n87300 , n87301 , n87302 , n87303 , n87304 , 
 n87305 , n87306 , n87307 , n87308 , n87309 , n87310 , n87311 , n87312 , n87313 , n87314 , 
 n87315 , n87316 , n87317 , n87318 , n87319 , n87320 , n87321 , n87322 , n87323 , n87324 , 
 n87325 , n87326 , n87327 , n87328 , n87329 , n87330 , n87331 , n87332 , n87333 , n87334 , 
 n87335 , n87336 , n87337 , n87338 , n87339 , n87340 , n87341 , n87342 , n87343 , n87344 , 
 n87345 , n87346 , n87347 , n87348 , n87349 , n87350 , n87351 , n87352 , n87353 , n87354 , 
 n87355 , n87356 , n87357 , n87358 , n87359 , n87360 , n87361 , n87362 , n87363 , n87364 , 
 n87365 , n87366 , n87367 , n87368 , n87369 , n87370 , n87371 , n87372 , n87373 , n87374 , 
 n87375 , n87376 , n87377 , n87378 , n87379 , n87380 , n87381 , n87382 , n87383 , n87384 , 
 n87385 , n87386 , n87387 , n87388 , n87389 , n87390 , n87391 , n87392 , n87393 , n87394 , 
 n87395 , n87396 , n87397 , n87398 , n87399 , n87400 , n87401 , n87402 , n87403 , n87404 , 
 n87405 , n87406 , n87407 , n87408 , n87409 , n87410 , n87411 , n87412 , n87413 , n87414 , 
 n87415 , n87416 , n87417 , n87418 , n87419 , n87420 , n87421 , n87422 , n87423 , n87424 , 
 n87425 , n87426 , n87427 , n87428 , n87429 , n87430 , n87431 , n87432 , n87433 , n87434 , 
 n87435 , n87436 , n87437 , n87438 , n87439 , n87440 , n87441 , n87442 , n87443 , n87444 , 
 n87445 , n87446 , n87447 , n87448 , n87449 , n87450 , n87451 , n87452 , n87453 , n87454 , 
 n87455 , n87456 , n87457 , n87458 , n87459 , n87460 , n87461 , n87462 , n87463 , n87464 , 
 n87465 , n87466 , n87467 , n87468 , n87469 , n87470 , n87471 , n87472 , n87473 , n87474 , 
 n87475 , n87476 , n87477 , n87478 , n87479 , n87480 , n87481 , n87482 , n87483 , n87484 , 
 n87485 , n87486 , n87487 , n87488 , n87489 , n87490 , n87491 , n87492 , n87493 , n87494 , 
 n87495 , n87496 , n87497 , n87498 , n87499 , n87500 , n87501 , n87502 , n87503 , n87504 , 
 n87505 , n87506 , n87507 , n87508 , n87509 , n87510 , n87511 , n87512 , n87513 , n87514 , 
 n87515 , n87516 , n87517 , n87518 , n87519 , n87520 , n87521 , n87522 , n87523 , n87524 , 
 n87525 , n87526 , n87527 , n87528 , n87529 , n87530 , n87531 , n87532 , n87533 , n87534 , 
 n87535 , n87536 , n87537 , n87538 , n87539 , n87540 , n87541 , n87542 , n87543 , n87544 , 
 n87545 , n87546 , n87547 , n87548 , n87549 , n87550 , n87551 , n87552 , n87553 , n87554 , 
 n87555 , n87556 , n87557 , n87558 , n87559 , n87560 , n87561 , n87562 , n87563 , n87564 , 
 n87565 , n87566 , n87567 , n87568 , n87569 , n87570 , n87571 , n87572 , n87573 , n87574 , 
 n87575 , n87576 , n87577 , n87578 , n87579 , n87580 , n87581 , n87582 , n87583 , n87584 , 
 n87585 , n87586 , n87587 , n87588 , n87589 , n87590 , n87591 , n87592 , n87593 , n87594 , 
 n87595 , n87596 , n87597 , n87598 , n87599 , n87600 , n87601 , n87602 , n87603 , n87604 , 
 n87605 , n87606 , n87607 , n87608 , n87609 , n87610 , n87611 , n87612 , n87613 , n87614 , 
 n87615 , n87616 , n87617 , n87618 , n87619 , n87620 , n87621 , n87622 , n87623 , n87624 , 
 n87625 , n87626 , n87627 , n87628 , n87629 , n87630 , n87631 , n87632 , n87633 , n87634 , 
 n87635 , n87636 , n87637 , n87638 , n87639 , n87640 , n87641 , n87642 , n87643 , n87644 , 
 n87645 , n87646 , n87647 , n87648 , n87649 , n87650 , n87651 , n87652 , n87653 , n87654 , 
 n87655 , n87656 , n87657 , n87658 , n87659 , n87660 , n87661 , n87662 , n87663 , n87664 , 
 n87665 , n87666 , n87667 , n87668 , n87669 , n87670 , n87671 , n87672 , n87673 , n87674 , 
 n87675 , n87676 , n87677 , n87678 , n87679 , n87680 , n87681 , n87682 , n87683 , n87684 , 
 n87685 , n87686 , n87687 , n87688 , n87689 , n87690 , n87691 , n87692 , n87693 , n87694 , 
 n87695 , n87696 , n87697 , n87698 , n87699 , n87700 , n87701 , n87702 , n87703 , n87704 , 
 n87705 , n87706 , n87707 , n87708 , n87709 , n87710 , n87711 , n87712 , n87713 , n87714 , 
 n87715 , n87716 , n87717 , n87718 , n87719 , n87720 , n87721 , n87722 , n87723 , n87724 , 
 n87725 , n87726 , n87727 , n87728 , n87729 , n87730 , n87731 , n87732 , n87733 , n87734 , 
 n87735 , n87736 , n87737 , n87738 , n87739 , n87740 , n87741 , n87742 , n87743 , n87744 , 
 n87745 , n87746 , n87747 , n87748 , n87749 , n87750 , n87751 , n87752 , n87753 , n87754 , 
 n87755 , n87756 , n87757 , n87758 , n87759 , n87760 , n87761 , n87762 , n87763 , n87764 , 
 n87765 , n87766 , n87767 , n87768 , n87769 , n87770 , n87771 , n87772 , n87773 , n87774 , 
 n87775 , n87776 , n87777 , n87778 , n87779 , n87780 , n87781 , n87782 , n87783 , n87784 , 
 n87785 , n87786 , n87787 , n87788 , n87789 , n87790 , n87791 , n87792 , n87793 , n87794 , 
 n87795 , n87796 , n87797 , n87798 , n87799 , n87800 , n87801 , n87802 , n87803 , n87804 , 
 n87805 , n87806 , n87807 , n87808 , n87809 , n87810 , n87811 , n87812 , n87813 , n87814 , 
 n87815 , n87816 , n87817 , n87818 , n87819 , n87820 , n87821 , n87822 , n87823 , n87824 , 
 n87825 , n87826 , n87827 , n87828 , n87829 , n87830 , n87831 , n87832 , n87833 , n87834 , 
 n87835 , n87836 , n87837 , n87838 , n87839 , n87840 , n87841 , n87842 , n87843 , n87844 , 
 n87845 , n87846 , n87847 , n87848 , n87849 , n87850 , n87851 , n87852 , n87853 , n87854 , 
 n87855 , n87856 , n87857 , n87858 , n87859 , n87860 , n87861 , n87862 , n87863 , n87864 , 
 n87865 , n87866 , n87867 , n87868 , n87869 , n87870 , n87871 , n87872 , n87873 , n87874 , 
 n87875 , n87876 , n87877 , n87878 , n87879 , n87880 , n87881 , n87882 , n87883 , n87884 , 
 n87885 , n87886 , n87887 , n87888 , n87889 , n87890 , n87891 , n87892 , n87893 , n87894 , 
 n87895 , n87896 , n87897 , n87898 , n87899 , n87900 , n87901 , n87902 , n87903 , n87904 , 
 n87905 , n87906 , n87907 , n87908 , n87909 , n87910 , n87911 , n87912 , n87913 , n87914 , 
 n87915 , n87916 , n87917 , n87918 , n87919 , n87920 , n87921 , n87922 , n87923 , n87924 , 
 n87925 , n87926 , n87927 , n87928 , n87929 , n87930 , n87931 , n87932 , n87933 , n87934 , 
 n87935 , n87936 , n87937 , n87938 , n87939 , n87940 , n87941 , n87942 , n87943 , n87944 , 
 n87945 , n87946 , n87947 , n87948 , n87949 , n87950 , n87951 , n87952 , n87953 , n87954 , 
 n87955 , n87956 , n87957 , n87958 , n87959 , n87960 , n87961 , n87962 , n87963 , n87964 , 
 n87965 , n87966 , n87967 , n87968 , n87969 , n87970 , n87971 , n87972 , n87973 , n87974 , 
 n87975 , n87976 , n87977 , n87978 , n87979 , n87980 , n87981 , n87982 , n87983 , n87984 , 
 n87985 , n87986 , n87987 , n87988 , n87989 , n87990 , n87991 , n87992 , n87993 , n87994 , 
 n87995 , n87996 , n87997 , n87998 , n87999 , n88000 , n88001 , n88002 , n88003 , n88004 , 
 n88005 , n88006 , n88007 , n88008 , n88009 , n88010 , n88011 , n88012 , n88013 , n88014 , 
 n88015 , n88016 , n88017 , n88018 , n88019 , n88020 , n88021 , n88022 , n88023 , n88024 , 
 n88025 , n88026 , n88027 , n88028 , n88029 , n88030 , n88031 , n88032 , n88033 , n88034 , 
 n88035 , n88036 , n88037 , n88038 , n88039 , n88040 , n88041 , n88042 , n88043 , n88044 , 
 n88045 , n88046 , n88047 , n88048 , n88049 , n88050 , n88051 , n88052 , n88053 , n88054 , 
 n88055 , n88056 , n88057 , n88058 , n88059 , n88060 , n88061 , n88062 , n88063 , n88064 , 
 n88065 , n88066 , n88067 , n88068 , n88069 , n88070 , n88071 , n88072 , n88073 , n88074 , 
 n88075 , n88076 , n88077 , n88078 , n88079 , n88080 , n88081 , n88082 , n88083 , n88084 , 
 n88085 , n88086 , n88087 , n88088 , n88089 , n88090 , n88091 , n88092 , n88093 , n88094 , 
 n88095 , n88096 , n88097 , n88098 , n88099 , n88100 , n88101 , n88102 , n88103 , n88104 , 
 n88105 , n88106 , n88107 , n88108 , n88109 , n88110 , n88111 , n88112 , n88113 , n88114 , 
 n88115 , n88116 , n88117 , n88118 , n88119 , n88120 , n88121 , n88122 , n88123 , n88124 , 
 n88125 , n88126 , n88127 , n88128 , n88129 , n88130 , n88131 , n88132 , n88133 , n88134 , 
 n88135 , n88136 , n88137 , n88138 , n88139 , n88140 , n88141 , n88142 , n88143 , n88144 , 
 n88145 , n88146 , n88147 , n88148 , n88149 , n88150 , n88151 , n88152 , n88153 , n88154 , 
 n88155 , n88156 , n88157 , n88158 , n88159 , n88160 , n88161 , n88162 , n88163 , n88164 , 
 n88165 , n88166 , n88167 , n88168 , n88169 , n88170 , n88171 , n88172 , n88173 , n88174 , 
 n88175 , n88176 , n88177 , n88178 , n88179 , n88180 , n88181 , n88182 , n88183 , n88184 , 
 n88185 , n88186 , n88187 , n88188 , n88189 , n88190 , n88191 , n88192 , n88193 , n88194 , 
 n88195 , n88196 , n88197 , n88198 , n88199 , n88200 , n88201 , n88202 , n88203 , n88204 , 
 n88205 , n88206 , n88207 , n88208 , n88209 , n88210 , n88211 , n88212 , n88213 , n88214 , 
 n88215 , n88216 , n88217 , n88218 , n88219 , n88220 , n88221 , n88222 , n88223 , n88224 , 
 n88225 , n88226 , n88227 , n88228 , n88229 , n88230 , n88231 , n88232 , n88233 , n88234 , 
 n88235 , n88236 , n88237 , n88238 , n88239 , n88240 , n88241 , n88242 , n88243 , n88244 , 
 n88245 , n88246 , n88247 , n88248 , n88249 , n88250 , n88251 , n88252 , n88253 , n88254 , 
 n88255 , n88256 , n88257 , n88258 , n88259 , n88260 , n88261 , n88262 , n88263 , n88264 , 
 n88265 , n88266 , n88267 , n88268 , n88269 , n88270 , n88271 , n88272 , n88273 , n88274 , 
 n88275 , n88276 , n88277 , n88278 , n88279 , n88280 , n88281 , n88282 , n88283 , n88284 , 
 n88285 , n88286 , n88287 , n88288 , n88289 , n88290 , n88291 , n88292 , n88293 , n88294 , 
 n88295 , n88296 , n88297 , n88298 , n88299 , n88300 , n88301 , n88302 , n88303 , n88304 , 
 n88305 , n88306 , n88307 , n88308 , n88309 , n88310 , n88311 , n88312 , n88313 , n88314 , 
 n88315 , n88316 , n88317 , n88318 , n88319 , n88320 , n88321 , n88322 , n88323 , n88324 , 
 n88325 , n88326 , n88327 , n88328 , n88329 , n88330 , n88331 , n88332 , n88333 , n88334 , 
 n88335 , n88336 , n88337 , n88338 , n88339 , n88340 , n88341 , n88342 , n88343 , n88344 , 
 n88345 , n88346 , n88347 , n88348 , n88349 , n88350 , n88351 , n88352 , n88353 , n88354 , 
 n88355 , n88356 , n88357 , n88358 , n88359 , n88360 , n88361 , n88362 , n88363 , n88364 , 
 n88365 , n88366 , n88367 , n88368 , n88369 , n88370 , n88371 , n88372 , n88373 , n88374 , 
 n88375 , n88376 , n88377 , n88378 , n88379 , n88380 , n88381 , n88382 , n88383 , n88384 , 
 n88385 , n88386 , n88387 , n88388 , n88389 , n88390 , n88391 , n88392 , n88393 , n88394 , 
 n88395 , n88396 , n88397 , n88398 , n88399 , n88400 , n88401 , n88402 , n88403 , n88404 , 
 n88405 , n88406 , n88407 , n88408 , n88409 , n88410 , n88411 , n88412 , n88413 , n88414 , 
 n88415 , n88416 , n88417 , n88418 , n88419 , n88420 , n88421 , n88422 , n88423 , n88424 , 
 n88425 , n88426 , n88427 , n88428 , n88429 , n88430 , n88431 , n88432 , n88433 , n88434 , 
 n88435 , n88436 , n88437 , n88438 , n88439 , n88440 , n88441 , n88442 , n88443 , n88444 , 
 n88445 , n88446 , n88447 , n88448 , n88449 , n88450 , n88451 , n88452 , n88453 , n88454 , 
 n88455 , n88456 , n88457 , n88458 , n88459 , n88460 , n88461 , n88462 , n88463 , n88464 , 
 n88465 , n88466 , n88467 , n88468 , n88469 , n88470 , n88471 , n88472 , n88473 , n88474 , 
 n88475 , n88476 , n88477 , n88478 , n88479 , n88480 , n88481 , n88482 , n88483 , n88484 , 
 n88485 , n88486 , n88487 , n88488 , n88489 , n88490 , n88491 , n88492 , n88493 , n88494 , 
 n88495 , n88496 , n88497 , n88498 , n88499 , n88500 , n88501 , n88502 , n88503 , n88504 , 
 n88505 , n88506 , n88507 , n88508 , n88509 , n88510 , n88511 , n88512 , n88513 , n88514 , 
 n88515 , n88516 , n88517 , n88518 , n88519 , n88520 , n88521 , n88522 , n88523 , n88524 , 
 n88525 , n88526 , n88527 , n88528 , n88529 , n88530 , n88531 , n88532 , n88533 , n88534 , 
 n88535 , n88536 , n88537 , n88538 , n88539 , n88540 , n88541 , n88542 , n88543 , n88544 , 
 n88545 , n88546 , n88547 , n88548 , n88549 , n88550 , n88551 , n88552 , n88553 , n88554 , 
 n88555 , n88556 , n88557 , n88558 , n88559 , n88560 , n88561 , n88562 , n88563 , n88564 , 
 n88565 , n88566 , n88567 , n88568 , n88569 , n88570 , n88571 , n88572 , n88573 , n88574 , 
 n88575 , n88576 , n88577 , n88578 , n88579 , n88580 , n88581 , n88582 , n88583 , n88584 , 
 n88585 , n88586 , n88587 , n88588 , n88589 , n88590 , n88591 , n88592 , n88593 , n88594 , 
 n88595 , n88596 , n88597 , n88598 , n88599 , n88600 , n88601 , n88602 , n88603 , n88604 , 
 n88605 , n88606 , n88607 , n88608 , n88609 , n88610 , n88611 , n88612 , n88613 , n88614 , 
 n88615 , n88616 , n88617 , n88618 , n88619 , n88620 , n88621 , n88622 , n88623 , n88624 , 
 n88625 , n88626 , n88627 , n88628 , n88629 , n88630 , n88631 , n88632 , n88633 , n88634 , 
 n88635 , n88636 , n88637 , n88638 , n88639 , n88640 , n88641 , n88642 , n88643 , n88644 , 
 n88645 , n88646 , n88647 , n88648 , n88649 , n88650 , n88651 , n88652 , n88653 , n88654 , 
 n88655 , n88656 , n88657 , n88658 , n88659 , n88660 , n88661 , n88662 , n88663 , n88664 , 
 n88665 , n88666 , n88667 , n88668 , n88669 , n88670 , n88671 , n88672 , n88673 , n88674 , 
 n88675 , n88676 , n88677 , n88678 , n88679 , n88680 , n88681 , n88682 , n88683 , n88684 , 
 n88685 , n88686 , n88687 , n88688 , n88689 , n88690 , n88691 , n88692 , n88693 , n88694 , 
 n88695 , n88696 , n88697 , n88698 , n88699 , n88700 , n88701 , n88702 , n88703 , n88704 , 
 n88705 , n88706 , n88707 , n88708 , n88709 , n88710 , n88711 , n88712 , n88713 , n88714 , 
 n88715 , n88716 , n88717 , n88718 , n88719 , n88720 , n88721 , n88722 , n88723 , n88724 , 
 n88725 , n88726 , n88727 , n88728 , n88729 , n88730 , n88731 , n88732 , n88733 , n88734 , 
 n88735 , n88736 , n88737 , n88738 , n88739 , n88740 , n88741 , n88742 , n88743 , n88744 , 
 n88745 , n88746 , n88747 , n88748 , n88749 , n88750 , n88751 , n88752 , n88753 , n88754 , 
 n88755 , n88756 , n88757 , n88758 , n88759 , n88760 , n88761 , n88762 , n88763 , n88764 , 
 n88765 , n88766 , n88767 , n88768 , n88769 , n88770 , n88771 , n88772 , n88773 , n88774 , 
 n88775 , n88776 , n88777 , n88778 , n88779 , n88780 , n88781 , n88782 , n88783 , n88784 , 
 n88785 , n88786 , n88787 , n88788 , n88789 , n88790 , n88791 , n88792 , n88793 , n88794 , 
 n88795 , n88796 , n88797 , n88798 , n88799 , n88800 , n88801 , n88802 , n88803 , n88804 , 
 n88805 , n88806 , n88807 , n88808 , n88809 , n88810 , n88811 , n88812 , n88813 , n88814 , 
 n88815 , n88816 , n88817 , n88818 , n88819 , n88820 , n88821 , n88822 , n88823 , n88824 , 
 n88825 , n88826 , n88827 , n88828 , n88829 , n88830 , n88831 , n88832 , n88833 , n88834 , 
 n88835 , n88836 , n88837 , n88838 , n88839 , n88840 , n88841 , n88842 , n88843 , n88844 , 
 n88845 , n88846 , n88847 , n88848 , n88849 , n88850 , n88851 , n88852 , n88853 , n88854 , 
 n88855 , n88856 , n88857 , n88858 , n88859 , n88860 , n88861 , n88862 , n88863 , n88864 , 
 n88865 , n88866 , n88867 , n88868 , n88869 , n88870 , n88871 , n88872 , n88873 , n88874 , 
 n88875 , n88876 , n88877 , n88878 , n88879 , n88880 , n88881 , n88882 , n88883 , n88884 , 
 n88885 , n88886 , n88887 , n88888 , n88889 , n88890 , n88891 , n88892 , n88893 , n88894 , 
 n88895 , n88896 , n88897 , n88898 , n88899 , n88900 , n88901 , n88902 , n88903 , n88904 , 
 n88905 , n88906 , n88907 , n88908 , n88909 , n88910 , n88911 , n88912 , n88913 , n88914 , 
 n88915 , n88916 , n88917 , n88918 , n88919 , n88920 , n88921 , n88922 , n88923 , n88924 , 
 n88925 , n88926 , n88927 , n88928 , n88929 , n88930 , n88931 , n88932 , n88933 , n88934 , 
 n88935 , n88936 , n88937 , n88938 , n88939 , n88940 , n88941 , n88942 , n88943 , n88944 , 
 n88945 , n88946 , n88947 , n88948 , n88949 , n88950 , n88951 , n88952 , n88953 , n88954 , 
 n88955 , n88956 , n88957 , n88958 , n88959 , n88960 , n88961 , n88962 , n88963 , n88964 , 
 n88965 , n88966 , n88967 , n88968 , n88969 , n88970 , n88971 , n88972 , n88973 , n88974 , 
 n88975 , n88976 , n88977 , n88978 , n88979 , n88980 , n88981 , n88982 , n88983 , n88984 , 
 n88985 , n88986 , n88987 , n88988 , n88989 , n88990 , n88991 , n88992 , n88993 , n88994 , 
 n88995 , n88996 , n88997 , n88998 , n88999 , n89000 , n89001 , n89002 , n89003 , n89004 , 
 n89005 , n89006 , n89007 , n89008 , n89009 , n89010 , n89011 , n89012 , n89013 , n89014 , 
 n89015 , n89016 , n89017 , n89018 , n89019 , n89020 , n89021 , n89022 , n89023 , n89024 , 
 n89025 , n89026 , n89027 , n89028 , n89029 , n89030 , n89031 , n89032 , n89033 , n89034 , 
 n89035 , n89036 , n89037 , n89038 , n89039 , n89040 , n89041 , n89042 , n89043 , n89044 , 
 n89045 , n89046 , n89047 , n89048 , n89049 , n89050 , n89051 , n89052 , n89053 , n89054 , 
 n89055 , n89056 , n89057 , n89058 , n89059 , n89060 , n89061 , n89062 , n89063 , n89064 , 
 n89065 , n89066 , n89067 , n89068 , n89069 , n89070 , n89071 , n89072 , n89073 , n89074 , 
 n89075 , n89076 , n89077 , n89078 , n89079 , n89080 , n89081 , n89082 , n89083 , n89084 , 
 n89085 , n89086 , n89087 , n89088 , n89089 , n89090 , n89091 , n89092 , n89093 , n89094 , 
 n89095 , n89096 , n89097 , n89098 , n89099 , n89100 , n89101 , n89102 , n89103 , n89104 , 
 n89105 , n89106 , n89107 , n89108 , n89109 , n89110 , n89111 , n89112 , n89113 , n89114 , 
 n89115 , n89116 , n89117 , n89118 , n89119 , n89120 , n89121 , n89122 , n89123 , n89124 , 
 n89125 , n89126 , n89127 , n89128 , n89129 , n89130 , n89131 , n89132 , n89133 , n89134 , 
 n89135 , n89136 , n89137 , n89138 , n89139 , n89140 , n89141 , n89142 , n89143 , n89144 , 
 n89145 , n89146 , n89147 , n89148 , n89149 , n89150 , n89151 , n89152 , n89153 , n89154 , 
 n89155 , n89156 , n89157 , n89158 , n89159 , n89160 , n89161 , n89162 , n89163 , n89164 , 
 n89165 , n89166 , n89167 , n89168 , n89169 , n89170 , n89171 , n89172 , n89173 , n89174 , 
 n89175 , n89176 , n89177 , n89178 , n89179 , n89180 , n89181 , n89182 , n89183 , n89184 , 
 n89185 , n89186 , n89187 , n89188 , n89189 , n89190 , n89191 , n89192 , n89193 , n89194 , 
 n89195 , n89196 , n89197 , n89198 , n89199 , n89200 , n89201 , n89202 , n89203 , n89204 , 
 n89205 , n89206 , n89207 , n89208 , n89209 , n89210 , n89211 , n89212 , n89213 , n89214 , 
 n89215 , n89216 , n89217 , n89218 , n89219 , n89220 , n89221 , n89222 , n89223 , n89224 , 
 n89225 , n89226 , n89227 , n89228 , n89229 , n89230 , n89231 , n89232 , n89233 , n89234 , 
 n89235 , n89236 , n89237 , n89238 , n89239 , n89240 , n89241 , n89242 , n89243 , n89244 , 
 n89245 , n89246 , n89247 , n89248 , n89249 , n89250 , n89251 , n89252 , n89253 , n89254 , 
 n89255 , n89256 , n89257 , n89258 , n89259 , n89260 , n89261 , n89262 , n89263 , n89264 , 
 n89265 , n89266 , n89267 , n89268 , n89269 , n89270 , n89271 , n89272 , n89273 , n89274 , 
 n89275 , n89276 , n89277 , n89278 , n89279 , n89280 , n89281 , n89282 , n89283 , n89284 , 
 n89285 , n89286 , n89287 , n89288 , n89289 , n89290 , n89291 , n89292 , n89293 , n89294 , 
 n89295 , n89296 , n89297 , n89298 , n89299 , n89300 , n89301 , n89302 , n89303 , n89304 , 
 n89305 , n89306 , n89307 , n89308 , n89309 , n89310 , n89311 , n89312 , n89313 , n89314 , 
 n89315 , n89316 , n89317 , n89318 , n89319 , n89320 , n89321 , n89322 , n89323 , n89324 , 
 n89325 , n89326 , n89327 , n89328 , n89329 , n89330 , n89331 , n89332 , n89333 , n89334 , 
 n89335 , n89336 , n89337 , n89338 , n89339 , n89340 , n89341 , n89342 , n89343 , n89344 , 
 n89345 , n89346 , n89347 , n89348 , n89349 , n89350 , n89351 , n89352 , n89353 , n89354 , 
 n89355 , n89356 , n89357 , n89358 , n89359 , n89360 , n89361 , n89362 , n89363 , n89364 , 
 n89365 , n89366 , n89367 , n89368 , n89369 , n89370 , n89371 , n89372 , n89373 , n89374 , 
 n89375 , n89376 , n89377 , n89378 , n89379 , n89380 , n89381 , n89382 , n89383 , n89384 , 
 n89385 , n89386 , n89387 , n89388 , n89389 , n89390 , n89391 , n89392 , n89393 , n89394 , 
 n89395 , n89396 , n89397 , n89398 , n89399 , n89400 , n89401 , n89402 , n89403 , n89404 , 
 n89405 , n89406 , n89407 , n89408 , n89409 , n89410 , n89411 , n89412 , n89413 , n89414 , 
 n89415 , n89416 , n89417 , n89418 , n89419 , n89420 , n89421 , n89422 , n89423 , n89424 , 
 n89425 , n89426 , n89427 , n89428 , n89429 , n89430 , n89431 , n89432 , n89433 , n89434 , 
 n89435 , n89436 , n89437 , n89438 , n89439 , n89440 , n89441 , n89442 , n89443 , n89444 , 
 n89445 , n89446 , n89447 , n89448 , n89449 , n89450 , n89451 , n89452 , n89453 , n89454 , 
 n89455 , n89456 , n89457 , n89458 , n89459 , n89460 , n89461 , n89462 , n89463 , n89464 , 
 n89465 , n89466 , n89467 , n89468 , n89469 , n89470 , n89471 , n89472 , n89473 , n89474 , 
 n89475 , n89476 , n89477 , n89478 , n89479 , n89480 , n89481 , n89482 , n89483 , n89484 , 
 n89485 , n89486 , n89487 , n89488 , n89489 , n89490 , n89491 , n89492 , n89493 , n89494 , 
 n89495 , n89496 , n89497 , n89498 , n89499 , n89500 , n89501 , n89502 , n89503 , n89504 , 
 n89505 , n89506 , n89507 , n89508 , n89509 , n89510 , n89511 , n89512 , n89513 , n89514 , 
 n89515 , n89516 , n89517 , n89518 , n89519 , n89520 , n89521 , n89522 , n89523 , n89524 , 
 n89525 , n89526 , n89527 , n89528 , n89529 , n89530 , n89531 , n89532 , n89533 , n89534 , 
 n89535 , n89536 , n89537 , n89538 , n89539 , n89540 , n89541 , n89542 , n89543 , n89544 , 
 n89545 , n89546 , n89547 , n89548 , n89549 , n89550 , n89551 , n89552 , n89553 , n89554 , 
 n89555 , n89556 , n89557 , n89558 , n89559 , n89560 , n89561 , n89562 , n89563 , n89564 , 
 n89565 , n89566 , n89567 , n89568 , n89569 , n89570 , n89571 , n89572 , n89573 , n89574 , 
 n89575 , n89576 , n89577 , n89578 , n89579 , n89580 , n89581 , n89582 , n89583 , n89584 , 
 n89585 , n89586 , n89587 , n89588 , n89589 , n89590 , n89591 , n89592 , n89593 , n89594 , 
 n89595 , n89596 , n89597 , n89598 , n89599 , n89600 , n89601 , n89602 , n89603 , n89604 , 
 n89605 , n89606 , n89607 , n89608 , n89609 , n89610 , n89611 , n89612 , n89613 , n89614 , 
 n89615 , n89616 , n89617 , n89618 , n89619 , n89620 , n89621 , n89622 , n89623 , n89624 , 
 n89625 , n89626 , n89627 , n89628 , n89629 , n89630 , n89631 , n89632 , n89633 , n89634 , 
 n89635 , n89636 , n89637 , n89638 , n89639 , n89640 , n89641 , n89642 , n89643 , n89644 , 
 n89645 , n89646 , n89647 , n89648 , n89649 , n89650 , n89651 , n89652 , n89653 , n89654 , 
 n89655 , n89656 , n89657 , n89658 , n89659 , n89660 , n89661 , n89662 , n89663 , n89664 , 
 n89665 , n89666 , n89667 , n89668 , n89669 , n89670 , n89671 , n89672 , n89673 , n89674 , 
 n89675 , n89676 , n89677 , n89678 , n89679 , n89680 , n89681 , n89682 , n89683 , n89684 , 
 n89685 , n89686 , n89687 , n89688 , n89689 , n89690 , n89691 , n89692 , n89693 , n89694 , 
 n89695 , n89696 , n89697 , n89698 , n89699 , n89700 , n89701 , n89702 , n89703 , n89704 , 
 n89705 , n89706 , n89707 , n89708 , n89709 , n89710 , n89711 , n89712 , n89713 , n89714 , 
 n89715 , n89716 , n89717 , n89718 , n89719 , n89720 , n89721 , n89722 , n89723 , n89724 , 
 n89725 , n89726 , n89727 , n89728 , n89729 , n89730 , n89731 , n89732 , n89733 , n89734 , 
 n89735 , n89736 , n89737 , n89738 , n89739 , n89740 , n89741 , n89742 , n89743 , n89744 , 
 n89745 , n89746 , n89747 , n89748 , n89749 , n89750 , n89751 , n89752 , n89753 , n89754 , 
 n89755 , n89756 , n89757 , n89758 , n89759 , n89760 , n89761 , n89762 , n89763 , n89764 , 
 n89765 , n89766 , n89767 , n89768 , n89769 , n89770 , n89771 , n89772 , n89773 , n89774 , 
 n89775 , n89776 , n89777 , n89778 , n89779 , n89780 , n89781 , n89782 , n89783 , n89784 , 
 n89785 , n89786 , n89787 , n89788 , n89789 , n89790 , n89791 , n89792 , n89793 , n89794 , 
 n89795 , n89796 , n89797 , n89798 , n89799 , n89800 , n89801 , n89802 , n89803 , n89804 , 
 n89805 , n89806 , n89807 , n89808 , n89809 , n89810 , n89811 , n89812 , n89813 , n89814 , 
 n89815 , n89816 , n89817 , n89818 , n89819 , n89820 , n89821 , n89822 , n89823 , n89824 , 
 n89825 , n89826 , n89827 , n89828 , n89829 , n89830 , n89831 , n89832 , n89833 , n89834 , 
 n89835 , n89836 , n89837 , n89838 , n89839 , n89840 , n89841 , n89842 , n89843 , n89844 , 
 n89845 , n89846 , n89847 , n89848 , n89849 , n89850 , n89851 , n89852 , n89853 , n89854 , 
 n89855 , n89856 , n89857 , n89858 , n89859 , n89860 , n89861 , n89862 , n89863 , n89864 , 
 n89865 , n89866 , n89867 , n89868 , n89869 , n89870 , n89871 , n89872 , n89873 , n89874 , 
 n89875 , n89876 , n89877 , n89878 , n89879 , n89880 , n89881 , n89882 , n89883 , n89884 , 
 n89885 , n89886 , n89887 , n89888 , n89889 , n89890 , n89891 , n89892 , n89893 , n89894 , 
 n89895 , n89896 , n89897 , n89898 , n89899 , n89900 , n89901 , n89902 , n89903 , n89904 , 
 n89905 , n89906 , n89907 , n89908 , n89909 , n89910 , n89911 , n89912 , n89913 , n89914 , 
 n89915 , n89916 , n89917 , n89918 , n89919 , n89920 , n89921 , n89922 , n89923 , n89924 , 
 n89925 , n89926 , n89927 , n89928 , n89929 , n89930 , n89931 , n89932 , n89933 , n89934 , 
 n89935 , n89936 , n89937 , n89938 , n89939 , n89940 , n89941 , n89942 , n89943 , n89944 , 
 n89945 , n89946 , n89947 , n89948 , n89949 , n89950 , n89951 , n89952 , n89953 , n89954 , 
 n89955 , n89956 , n89957 , n89958 , n89959 , n89960 , n89961 , n89962 , n89963 , n89964 , 
 n89965 , n89966 , n89967 , n89968 , n89969 , n89970 , n89971 , n89972 , n89973 , n89974 , 
 n89975 , n89976 , n89977 , n89978 , n89979 , n89980 , n89981 , n89982 , n89983 , n89984 , 
 n89985 , n89986 , n89987 , n89988 , n89989 , n89990 , n89991 , n89992 , n89993 , n89994 , 
 n89995 , n89996 , n89997 , n89998 , n89999 , n90000 , n90001 , n90002 , n90003 , n90004 , 
 n90005 , n90006 , n90007 , n90008 , n90009 , n90010 , n90011 , n90012 , n90013 , n90014 , 
 n90015 , n90016 , n90017 , n90018 , n90019 , n90020 , n90021 , n90022 , n90023 , n90024 , 
 n90025 , n90026 , n90027 , n90028 , n90029 , n90030 , n90031 , n90032 , n90033 , n90034 , 
 n90035 , n90036 , n90037 , n90038 , n90039 , n90040 , n90041 , n90042 , n90043 , n90044 , 
 n90045 , n90046 , n90047 , n90048 , n90049 , n90050 , n90051 , n90052 , n90053 , n90054 , 
 n90055 , n90056 , n90057 , n90058 , n90059 , n90060 , n90061 , n90062 , n90063 , n90064 , 
 n90065 , n90066 , n90067 , n90068 , n90069 , n90070 , n90071 , n90072 , n90073 , n90074 , 
 n90075 , n90076 , n90077 , n90078 , n90079 , n90080 , n90081 , n90082 , n90083 , n90084 , 
 n90085 , n90086 , n90087 , n90088 , n90089 , n90090 , n90091 , n90092 , n90093 , n90094 , 
 n90095 , n90096 , n90097 , n90098 , n90099 , n90100 , n90101 , n90102 , n90103 , n90104 , 
 n90105 , n90106 , n90107 , n90108 , n90109 , n90110 , n90111 , n90112 , n90113 , n90114 , 
 n90115 , n90116 , n90117 , n90118 , n90119 , n90120 , n90121 , n90122 , n90123 , n90124 , 
 n90125 , n90126 , n90127 , n90128 , n90129 , n90130 , n90131 , n90132 , n90133 , n90134 , 
 n90135 , n90136 , n90137 , n90138 , n90139 , n90140 , n90141 , n90142 , n90143 , n90144 , 
 n90145 , n90146 , n90147 , n90148 , n90149 , n90150 , n90151 , n90152 , n90153 , n90154 , 
 n90155 , n90156 , n90157 , n90158 , n90159 , n90160 , n90161 , n90162 , n90163 , n90164 , 
 n90165 , n90166 , n90167 , n90168 , n90169 , n90170 , n90171 , n90172 , n90173 , n90174 , 
 n90175 , n90176 , n90177 , n90178 , n90179 , n90180 , n90181 , n90182 , n90183 , n90184 , 
 n90185 , n90186 , n90187 , n90188 , n90189 , n90190 , n90191 , n90192 , n90193 , n90194 , 
 n90195 , n90196 , n90197 , n90198 , n90199 , n90200 , n90201 , n90202 , n90203 , n90204 , 
 n90205 , n90206 , n90207 , n90208 , n90209 , n90210 , n90211 , n90212 , n90213 , n90214 , 
 n90215 , n90216 , n90217 , n90218 , n90219 , n90220 , n90221 , n90222 , n90223 , n90224 , 
 n90225 , n90226 , n90227 , n90228 , n90229 , n90230 , n90231 , n90232 , n90233 , n90234 , 
 n90235 , n90236 , n90237 , n90238 , n90239 , n90240 , n90241 , n90242 , n90243 , n90244 , 
 n90245 , n90246 , n90247 , n90248 , n90249 , n90250 , n90251 , n90252 , n90253 , n90254 , 
 n90255 , n90256 , n90257 , n90258 , n90259 , n90260 , n90261 , n90262 , n90263 , n90264 , 
 n90265 , n90266 , n90267 , n90268 , n90269 , n90270 , n90271 , n90272 , n90273 , n90274 , 
 n90275 , n90276 , n90277 , n90278 , n90279 , n90280 , n90281 , n90282 , n90283 , n90284 , 
 n90285 , n90286 , n90287 , n90288 , n90289 , n90290 , n90291 , n90292 , n90293 , n90294 , 
 n90295 , n90296 , n90297 , n90298 , n90299 , n90300 , n90301 , n90302 , n90303 , n90304 , 
 n90305 , n90306 , n90307 , n90308 , n90309 , n90310 , n90311 , n90312 , n90313 , n90314 , 
 n90315 , n90316 , n90317 , n90318 , n90319 , n90320 , n90321 , n90322 , n90323 , n90324 , 
 n90325 , n90326 , n90327 , n90328 , n90329 , n90330 , n90331 , n90332 , n90333 , n90334 , 
 n90335 , n90336 , n90337 , n90338 , n90339 , n90340 , n90341 , n90342 , n90343 , n90344 , 
 n90345 , n90346 , n90347 , n90348 , n90349 , n90350 , n90351 , n90352 , n90353 , n90354 , 
 n90355 , n90356 , n90357 , n90358 , n90359 , n90360 , n90361 , n90362 , n90363 , n90364 , 
 n90365 , n90366 , n90367 , n90368 , n90369 , n90370 , n90371 , n90372 , n90373 , n90374 , 
 n90375 , n90376 , n90377 , n90378 , n90379 , n90380 , n90381 , n90382 , n90383 , n90384 , 
 n90385 , n90386 , n90387 , n90388 , n90389 , n90390 , n90391 , n90392 , n90393 , n90394 , 
 n90395 , n90396 , n90397 , n90398 , n90399 , n90400 , n90401 , n90402 , n90403 , n90404 , 
 n90405 , n90406 , n90407 , n90408 , n90409 , n90410 , n90411 , n90412 , n90413 , n90414 , 
 n90415 , n90416 , n90417 , n90418 , n90419 , n90420 , n90421 , n90422 , n90423 , n90424 , 
 n90425 , n90426 , n90427 , n90428 , n90429 , n90430 , n90431 , n90432 , n90433 , n90434 , 
 n90435 , n90436 , n90437 , n90438 , n90439 , n90440 , n90441 , n90442 , n90443 , n90444 , 
 n90445 , n90446 , n90447 , n90448 , n90449 , n90450 , n90451 , n90452 , n90453 , n90454 , 
 n90455 , n90456 , n90457 , n90458 , n90459 , n90460 , n90461 , n90462 , n90463 , n90464 , 
 n90465 , n90466 , n90467 , n90468 , n90469 , n90470 , n90471 , n90472 , n90473 , n90474 , 
 n90475 , n90476 , n90477 , n90478 , n90479 , n90480 , n90481 , n90482 , n90483 , n90484 , 
 n90485 , n90486 , n90487 , n90488 , n90489 , n90490 , n90491 , n90492 , n90493 , n90494 , 
 n90495 , n90496 , n90497 , n90498 , n90499 , n90500 , n90501 , n90502 , n90503 , n90504 , 
 n90505 , n90506 , n90507 , n90508 , n90509 , n90510 , n90511 , n90512 , n90513 , n90514 , 
 n90515 , n90516 , n90517 , n90518 , n90519 , n90520 , n90521 , n90522 , n90523 , n90524 , 
 n90525 , n90526 , n90527 , n90528 , n90529 , n90530 , n90531 , n90532 , n90533 , n90534 , 
 n90535 , n90536 , n90537 , n90538 , n90539 , n90540 , n90541 , n90542 , n90543 , n90544 , 
 n90545 , n90546 , n90547 , n90548 , n90549 , n90550 , n90551 , n90552 , n90553 , n90554 , 
 n90555 , n90556 , n90557 , n90558 , n90559 , n90560 , n90561 , n90562 , n90563 , n90564 , 
 n90565 , n90566 , n90567 , n90568 , n90569 , n90570 , n90571 , n90572 , n90573 , n90574 , 
 n90575 , n90576 , n90577 , n90578 , n90579 , n90580 , n90581 , n90582 , n90583 , n90584 , 
 n90585 , n90586 , n90587 , n90588 , n90589 , n90590 , n90591 , n90592 , n90593 , n90594 , 
 n90595 , n90596 , n90597 , n90598 , n90599 , n90600 , n90601 , n90602 , n90603 , n90604 , 
 n90605 , n90606 , n90607 , n90608 , n90609 , n90610 , n90611 , n90612 , n90613 , n90614 , 
 n90615 , n90616 , n90617 , n90618 , n90619 , n90620 , n90621 , n90622 , n90623 , n90624 , 
 n90625 , n90626 , n90627 , n90628 , n90629 , n90630 , n90631 , n90632 , n90633 , n90634 , 
 n90635 , n90636 , n90637 , n90638 , n90639 , n90640 , n90641 , n90642 , n90643 , n90644 , 
 n90645 , n90646 , n90647 , n90648 , n90649 , n90650 , n90651 , n90652 , n90653 , n90654 , 
 n90655 , n90656 , n90657 , n90658 , n90659 , n90660 , n90661 , n90662 , n90663 , n90664 , 
 n90665 , n90666 , n90667 , n90668 , n90669 , n90670 , n90671 , n90672 , n90673 , n90674 , 
 n90675 , n90676 , n90677 , n90678 , n90679 , n90680 , n90681 , n90682 , n90683 , n90684 , 
 n90685 , n90686 , n90687 , n90688 , n90689 , n90690 , n90691 , n90692 , n90693 , n90694 , 
 n90695 , n90696 , n90697 , n90698 , n90699 , n90700 , n90701 , n90702 , n90703 , n90704 , 
 n90705 , n90706 , n90707 , n90708 , n90709 , n90710 , n90711 , n90712 , n90713 , n90714 , 
 n90715 , n90716 , n90717 , n90718 , n90719 , n90720 , n90721 , n90722 , n90723 , n90724 , 
 n90725 , n90726 , n90727 , n90728 , n90729 , n90730 , n90731 , n90732 , n90733 , n90734 , 
 n90735 , n90736 , n90737 , n90738 , n90739 , n90740 , n90741 , n90742 , n90743 , n90744 , 
 n90745 , n90746 , n90747 , n90748 , n90749 , n90750 , n90751 , n90752 , n90753 , n90754 , 
 n90755 , n90756 , n90757 , n90758 , n90759 , n90760 , n90761 , n90762 , n90763 , n90764 , 
 n90765 , n90766 , n90767 , n90768 , n90769 , n90770 , n90771 , n90772 , n90773 , n90774 , 
 n90775 , n90776 , n90777 , n90778 , n90779 , n90780 , n90781 , n90782 , n90783 , n90784 , 
 n90785 , n90786 , n90787 , n90788 , n90789 , n90790 , n90791 , n90792 , n90793 , n90794 , 
 n90795 , n90796 , n90797 , n90798 , n90799 , n90800 , n90801 , n90802 , n90803 , n90804 , 
 n90805 , n90806 , n90807 , n90808 , n90809 , n90810 , n90811 , n90812 , n90813 , n90814 , 
 n90815 , n90816 , n90817 , n90818 , n90819 , n90820 , n90821 , n90822 , n90823 , n90824 , 
 n90825 , n90826 , n90827 , n90828 , n90829 , n90830 , n90831 , n90832 , n90833 , n90834 , 
 n90835 , n90836 , n90837 , n90838 , n90839 , n90840 , n90841 , n90842 , n90843 , n90844 , 
 n90845 , n90846 , n90847 , n90848 , n90849 , n90850 , n90851 , n90852 , n90853 , n90854 , 
 n90855 , n90856 , n90857 , n90858 , n90859 , n90860 , n90861 , n90862 , n90863 , n90864 , 
 n90865 , n90866 , n90867 , n90868 , n90869 , n90870 , n90871 , n90872 , n90873 , n90874 , 
 n90875 , n90876 , n90877 , n90878 , n90879 , n90880 , n90881 , n90882 , n90883 , n90884 , 
 n90885 , n90886 , n90887 , n90888 , n90889 , n90890 , n90891 , n90892 , n90893 , n90894 , 
 n90895 , n90896 , n90897 , n90898 , n90899 , n90900 , n90901 , n90902 , n90903 , n90904 , 
 n90905 , n90906 , n90907 , n90908 , n90909 , n90910 , n90911 , n90912 , n90913 , n90914 , 
 n90915 , n90916 , n90917 , n90918 , n90919 , n90920 , n90921 , n90922 , n90923 , n90924 , 
 n90925 , n90926 , n90927 , n90928 , n90929 , n90930 , n90931 , n90932 , n90933 , n90934 , 
 n90935 , n90936 , n90937 , n90938 , n90939 , n90940 , n90941 , n90942 , n90943 , n90944 , 
 n90945 , n90946 , n90947 , n90948 , n90949 , n90950 , n90951 , n90952 , n90953 , n90954 , 
 n90955 , n90956 , n90957 , n90958 , n90959 , n90960 , n90961 , n90962 , n90963 , n90964 , 
 n90965 , n90966 , n90967 , n90968 , n90969 , n90970 , n90971 , n90972 , n90973 , n90974 , 
 n90975 , n90976 , n90977 , n90978 , n90979 , n90980 , n90981 , n90982 , n90983 , n90984 , 
 n90985 , n90986 , n90987 , n90988 , n90989 , n90990 , n90991 , n90992 , n90993 , n90994 , 
 n90995 , n90996 , n90997 , n90998 , n90999 , n91000 , n91001 , n91002 , n91003 , n91004 , 
 n91005 , n91006 , n91007 , n91008 , n91009 , n91010 , n91011 , n91012 , n91013 , n91014 , 
 n91015 , n91016 , n91017 , n91018 , n91019 , n91020 , n91021 , n91022 , n91023 , n91024 , 
 n91025 , n91026 , n91027 , n91028 , n91029 , n91030 , n91031 , n91032 , n91033 , n91034 , 
 n91035 , n91036 , n91037 , n91038 , n91039 , n91040 , n91041 , n91042 , n91043 , n91044 , 
 n91045 , n91046 , n91047 , n91048 , n91049 , n91050 , n91051 , n91052 , n91053 , n91054 , 
 n91055 , n91056 , n91057 , n91058 , n91059 , n91060 , n91061 , n91062 , n91063 , n91064 , 
 n91065 , n91066 , n91067 , n91068 , n91069 , n91070 , n91071 , n91072 , n91073 , n91074 , 
 n91075 , n91076 , n91077 , n91078 , n91079 , n91080 , n91081 , n91082 , n91083 , n91084 , 
 n91085 , n91086 , n91087 , n91088 , n91089 , n91090 , n91091 , n91092 , n91093 , n91094 , 
 n91095 , n91096 , n91097 , n91098 , n91099 , n91100 , n91101 , n91102 , n91103 , n91104 , 
 n91105 , n91106 , n91107 , n91108 , n91109 , n91110 , n91111 , n91112 , n91113 , n91114 , 
 n91115 , n91116 , n91117 , n91118 , n91119 , n91120 , n91121 , n91122 , n91123 , n91124 , 
 n91125 , n91126 , n91127 , n91128 , n91129 , n91130 , n91131 , n91132 , n91133 , n91134 , 
 n91135 , n91136 , n91137 , n91138 , n91139 , n91140 , n91141 , n91142 , n91143 , n91144 , 
 n91145 , n91146 , n91147 , n91148 , n91149 , n91150 , n91151 , n91152 , n91153 , n91154 , 
 n91155 , n91156 , n91157 , n91158 , n91159 , n91160 , n91161 , n91162 , n91163 , n91164 , 
 n91165 , n91166 , n91167 , n91168 , n91169 , n91170 , n91171 , n91172 , n91173 , n91174 , 
 n91175 , n91176 , n91177 , n91178 , n91179 , n91180 , n91181 , n91182 , n91183 , n91184 , 
 n91185 , n91186 , n91187 , n91188 , n91189 , n91190 , n91191 , n91192 , n91193 , n91194 , 
 n91195 , n91196 , n91197 , n91198 , n91199 , n91200 , n91201 , n91202 , n91203 , n91204 , 
 n91205 , n91206 , n91207 , n91208 , n91209 , n91210 , n91211 , n91212 , n91213 , n91214 , 
 n91215 , n91216 , n91217 , n91218 , n91219 , n91220 , n91221 , n91222 , n91223 , n91224 , 
 n91225 , n91226 , n91227 , n91228 , n91229 , n91230 , n91231 , n91232 , n91233 , n91234 , 
 n91235 , n91236 , n91237 , n91238 , n91239 , n91240 , n91241 , n91242 , n91243 , n91244 , 
 n91245 , n91246 , n91247 , n91248 , n91249 , n91250 , n91251 , n91252 , n91253 , n91254 , 
 n91255 , n91256 , n91257 , n91258 , n91259 , n91260 , n91261 , n91262 , n91263 , n91264 , 
 n91265 , n91266 , n91267 , n91268 , n91269 , n91270 , n91271 , n91272 , n91273 , n91274 , 
 n91275 , n91276 , n91277 , n91278 , n91279 , n91280 , n91281 , n91282 , n91283 , n91284 , 
 n91285 , n91286 , n91287 , n91288 , n91289 , n91290 , n91291 , n91292 , n91293 , n91294 , 
 n91295 , n91296 , n91297 , n91298 , n91299 , n91300 , n91301 , n91302 , n91303 , n91304 , 
 n91305 , n91306 , n91307 , n91308 , n91309 , n91310 , n91311 , n91312 , n91313 , n91314 , 
 n91315 , n91316 , n91317 , n91318 , n91319 , n91320 , n91321 , n91322 , n91323 , n91324 , 
 n91325 , n91326 , n91327 , n91328 , n91329 , n91330 , n91331 , n91332 , n91333 , n91334 , 
 n91335 , n91336 , n91337 , n91338 , n91339 , n91340 , n91341 , n91342 , n91343 , n91344 , 
 n91345 , n91346 , n91347 , n91348 , n91349 , n91350 , n91351 , n91352 , n91353 , n91354 , 
 n91355 , n91356 , n91357 , n91358 , n91359 , n91360 , n91361 , n91362 , n91363 , n91364 , 
 n91365 , n91366 , n91367 , n91368 , n91369 , n91370 , n91371 , n91372 , n91373 , n91374 , 
 n91375 , n91376 , n91377 , n91378 , n91379 , n91380 , n91381 , n91382 , n91383 , n91384 , 
 n91385 , n91386 , n91387 , n91388 , n91389 , n91390 , n91391 , n91392 , n91393 , n91394 , 
 n91395 , n91396 , n91397 , n91398 , n91399 , n91400 , n91401 , n91402 , n91403 , n91404 , 
 n91405 , n91406 , n91407 , n91408 , n91409 , n91410 , n91411 , n91412 , n91413 , n91414 , 
 n91415 , n91416 , n91417 , n91418 , n91419 , n91420 , n91421 , n91422 , n91423 , n91424 , 
 n91425 , n91426 , n91427 , n91428 , n91429 , n91430 , n91431 , n91432 , n91433 , n91434 , 
 n91435 , n91436 , n91437 , n91438 , n91439 , n91440 , n91441 , n91442 , n91443 , n91444 , 
 n91445 , n91446 , n91447 , n91448 , n91449 , n91450 , n91451 , n91452 , n91453 , n91454 , 
 n91455 , n91456 , n91457 , n91458 , n91459 , n91460 , n91461 , n91462 , n91463 , n91464 , 
 n91465 , n91466 , n91467 , n91468 , n91469 , n91470 , n91471 , n91472 , n91473 , n91474 , 
 n91475 , n91476 , n91477 , n91478 , n91479 , n91480 , n91481 , n91482 , n91483 , n91484 , 
 n91485 , n91486 , n91487 , n91488 , n91489 , n91490 , n91491 , n91492 , n91493 , n91494 , 
 n91495 , n91496 , n91497 , n91498 , n91499 , n91500 , n91501 , n91502 , n91503 , n91504 , 
 n91505 , n91506 , n91507 , n91508 , n91509 , n91510 , n91511 , n91512 , n91513 , n91514 , 
 n91515 , n91516 , n91517 , n91518 , n91519 , n91520 , n91521 , n91522 , n91523 , n91524 , 
 n91525 , n91526 , n91527 , n91528 , n91529 , n91530 , n91531 , n91532 , n91533 , n91534 , 
 n91535 , n91536 , n91537 , n91538 , n91539 , n91540 , n91541 , n91542 , n91543 , n91544 , 
 n91545 , n91546 , n91547 , n91548 , n91549 , n91550 , n91551 , n91552 , n91553 , n91554 , 
 n91555 , n91556 , n91557 , n91558 , n91559 , n91560 , n91561 , n91562 , n91563 , n91564 , 
 n91565 , n91566 , n91567 , n91568 , n91569 , n91570 , n91571 , n91572 , n91573 , n91574 , 
 n91575 , n91576 , n91577 , n91578 , n91579 , n91580 , n91581 , n91582 , n91583 , n91584 , 
 n91585 , n91586 , n91587 , n91588 , n91589 , n91590 , n91591 , n91592 , n91593 , n91594 , 
 n91595 , n91596 , n91597 , n91598 , n91599 , n91600 , n91601 , n91602 , n91603 , n91604 , 
 n91605 , n91606 , n91607 , n91608 , n91609 , n91610 , n91611 , n91612 , n91613 , n91614 , 
 n91615 , n91616 , n91617 , n91618 , n91619 , n91620 , n91621 , n91622 , n91623 , n91624 , 
 n91625 , n91626 , n91627 , n91628 , n91629 , n91630 , n91631 , n91632 , n91633 , n91634 , 
 n91635 , n91636 , n91637 , n91638 , n91639 , n91640 , n91641 , n91642 , n91643 , n91644 , 
 n91645 , n91646 , n91647 , n91648 , n91649 , n91650 , n91651 , n91652 , n91653 , n91654 , 
 n91655 , n91656 , n91657 , n91658 , n91659 , n91660 , n91661 , n91662 , n91663 , n91664 , 
 n91665 , n91666 , n91667 , n91668 , n91669 , n91670 , n91671 , n91672 , n91673 , n91674 , 
 n91675 , n91676 , n91677 , n91678 , n91679 , n91680 , n91681 , n91682 , n91683 , n91684 , 
 n91685 , n91686 , n91687 , n91688 , n91689 , n91690 , n91691 , n91692 , n91693 , n91694 , 
 n91695 , n91696 , n91697 , n91698 , n91699 , n91700 , n91701 , n91702 , n91703 , n91704 , 
 n91705 , n91706 , n91707 , n91708 , n91709 , n91710 , n91711 , n91712 , n91713 , n91714 , 
 n91715 , n91716 , n91717 , n91718 , n91719 , n91720 , n91721 , n91722 , n91723 , n91724 , 
 n91725 , n91726 , n91727 , n91728 , n91729 , n91730 , n91731 , n91732 , n91733 , n91734 , 
 n91735 , n91736 , n91737 , n91738 , n91739 , n91740 , n91741 , n91742 , n91743 , n91744 , 
 n91745 , n91746 , n91747 , n91748 , n91749 , n91750 , n91751 , n91752 , n91753 , n91754 , 
 n91755 , n91756 , n91757 , n91758 , n91759 , n91760 , n91761 , n91762 , n91763 , n91764 , 
 n91765 , n91766 , n91767 , n91768 , n91769 , n91770 , n91771 , n91772 , n91773 , n91774 , 
 n91775 , n91776 , n91777 , n91778 , n91779 , n91780 , n91781 , n91782 , n91783 , n91784 , 
 n91785 , n91786 , n91787 , n91788 , n91789 , n91790 , n91791 , n91792 , n91793 , n91794 , 
 n91795 , n91796 , n91797 , n91798 , n91799 , n91800 , n91801 , n91802 , n91803 , n91804 , 
 n91805 , n91806 , n91807 , n91808 , n91809 , n91810 , n91811 , n91812 , n91813 , n91814 , 
 n91815 , n91816 , n91817 , n91818 , n91819 , n91820 , n91821 , n91822 , n91823 , n91824 , 
 n91825 , n91826 , n91827 , n91828 , n91829 , n91830 , n91831 , n91832 , n91833 , n91834 , 
 n91835 , n91836 , n91837 , n91838 , n91839 , n91840 , n91841 , n91842 , n91843 , n91844 , 
 n91845 , n91846 , n91847 , n91848 , n91849 , n91850 , n91851 , n91852 , n91853 , n91854 , 
 n91855 , n91856 , n91857 , n91858 , n91859 , n91860 , n91861 , n91862 , n91863 , n91864 , 
 n91865 , n91866 , n91867 , n91868 , n91869 , n91870 , n91871 , n91872 , n91873 , n91874 , 
 n91875 , n91876 , n91877 , n91878 , n91879 , n91880 , n91881 , n91882 , n91883 , n91884 , 
 n91885 , n91886 , n91887 , n91888 , n91889 , n91890 , n91891 , n91892 , n91893 , n91894 , 
 n91895 , n91896 , n91897 , n91898 , n91899 , n91900 , n91901 , n91902 , n91903 , n91904 , 
 n91905 , n91906 , n91907 , n91908 , n91909 , n91910 , n91911 , n91912 , n91913 , n91914 , 
 n91915 , n91916 , n91917 , n91918 , n91919 , n91920 , n91921 , n91922 , n91923 , n91924 , 
 n91925 , n91926 , n91927 , n91928 , n91929 , n91930 , n91931 , n91932 , n91933 , n91934 , 
 n91935 , n91936 , n91937 , n91938 , n91939 , n91940 , n91941 , n91942 , n91943 , n91944 , 
 n91945 , n91946 , n91947 , n91948 , n91949 , n91950 , n91951 , n91952 , n91953 , n91954 , 
 n91955 , n91956 , n91957 , n91958 , n91959 , n91960 , n91961 , n91962 , n91963 , n91964 , 
 n91965 , n91966 , n91967 , n91968 , n91969 , n91970 , n91971 , n91972 , n91973 , n91974 , 
 n91975 , n91976 , n91977 , n91978 , n91979 , n91980 , n91981 , n91982 , n91983 , n91984 , 
 n91985 , n91986 , n91987 , n91988 , n91989 , n91990 , n91991 , n91992 , n91993 , n91994 , 
 n91995 , n91996 , n91997 , n91998 , n91999 , n92000 , n92001 , n92002 , n92003 , n92004 , 
 n92005 , n92006 , n92007 , n92008 , n92009 , n92010 , n92011 , n92012 , n92013 , n92014 , 
 n92015 , n92016 , n92017 , n92018 , n92019 , n92020 , n92021 , n92022 , n92023 , n92024 , 
 n92025 , n92026 , n92027 , n92028 , n92029 , n92030 , n92031 , n92032 , n92033 , n92034 , 
 n92035 , n92036 , n92037 , n92038 , n92039 , n92040 , n92041 , n92042 , n92043 , n92044 , 
 n92045 , n92046 , n92047 , n92048 , n92049 , n92050 , n92051 , n92052 , n92053 , n92054 , 
 n92055 , n92056 , n92057 , n92058 , n92059 , n92060 , n92061 , n92062 , n92063 , n92064 , 
 n92065 , n92066 , n92067 , n92068 , n92069 , n92070 , n92071 , n92072 , n92073 , n92074 , 
 n92075 , n92076 , n92077 , n92078 , n92079 , n92080 , n92081 , n92082 , n92083 , n92084 , 
 n92085 , n92086 , n92087 , n92088 , n92089 , n92090 , n92091 , n92092 , n92093 , n92094 , 
 n92095 , n92096 , n92097 , n92098 , n92099 , n92100 , n92101 , n92102 , n92103 , n92104 , 
 n92105 , n92106 , n92107 , n92108 , n92109 , n92110 , n92111 , n92112 , n92113 , n92114 , 
 n92115 , n92116 , n92117 , n92118 , n92119 , n92120 , n92121 , n92122 , n92123 , n92124 , 
 n92125 , n92126 , n92127 , n92128 , n92129 , n92130 , n92131 , n92132 , n92133 , n92134 , 
 n92135 , n92136 , n92137 , n92138 , n92139 , n92140 , n92141 , n92142 , n92143 , n92144 , 
 n92145 , n92146 , n92147 , n92148 , n92149 , n92150 , n92151 , n92152 , n92153 , n92154 , 
 n92155 , n92156 , n92157 , n92158 , n92159 , n92160 , n92161 , n92162 , n92163 , n92164 , 
 n92165 , n92166 , n92167 , n92168 , n92169 , n92170 , n92171 , n92172 , n92173 , n92174 , 
 n92175 , n92176 , n92177 , n92178 , n92179 , n92180 , n92181 , n92182 , n92183 , n92184 , 
 n92185 , n92186 , n92187 , n92188 , n92189 , n92190 , n92191 , n92192 , n92193 , n92194 , 
 n92195 , n92196 , n92197 , n92198 , n92199 , n92200 , n92201 , n92202 , n92203 , n92204 , 
 n92205 , n92206 , n92207 , n92208 , n92209 , n92210 , n92211 , n92212 , n92213 , n92214 , 
 n92215 , n92216 , n92217 , n92218 , n92219 , n92220 , n92221 , n92222 , n92223 , n92224 , 
 n92225 , n92226 , n92227 , n92228 , n92229 , n92230 , n92231 , n92232 , n92233 , n92234 , 
 n92235 , n92236 , n92237 , n92238 , n92239 , n92240 , n92241 , n92242 , n92243 , n92244 , 
 n92245 , n92246 , n92247 , n92248 , n92249 , n92250 , n92251 , n92252 , n92253 , n92254 , 
 n92255 , n92256 , n92257 , n92258 , n92259 , n92260 , n92261 , n92262 , n92263 , n92264 , 
 n92265 , n92266 , n92267 , n92268 , n92269 , n92270 , n92271 , n92272 , n92273 , n92274 , 
 n92275 , n92276 , n92277 , n92278 , n92279 , n92280 , n92281 , n92282 , n92283 , n92284 , 
 n92285 , n92286 , n92287 , n92288 , n92289 , n92290 , n92291 , n92292 , n92293 , n92294 , 
 n92295 , n92296 , n92297 , n92298 , n92299 , n92300 , n92301 , n92302 , n92303 , n92304 , 
 n92305 , n92306 , n92307 , n92308 , n92309 , n92310 , n92311 , n92312 , n92313 , n92314 , 
 n92315 , n92316 , n92317 , n92318 , n92319 , n92320 , n92321 , n92322 , n92323 , n92324 , 
 n92325 , n92326 , n92327 , n92328 , n92329 , n92330 , n92331 , n92332 , n92333 , n92334 , 
 n92335 , n92336 , n92337 , n92338 , n92339 , n92340 , n92341 , n92342 , n92343 , n92344 , 
 n92345 , n92346 , n92347 , n92348 , n92349 , n92350 , n92351 , n92352 , n92353 , n92354 , 
 n92355 , n92356 , n92357 , n92358 , n92359 , n92360 , n92361 , n92362 , n92363 , n92364 , 
 n92365 , n92366 , n92367 , n92368 , n92369 , n92370 , n92371 , n92372 , n92373 , n92374 , 
 n92375 , n92376 , n92377 , n92378 , n92379 , n92380 , n92381 , n92382 , n92383 , n92384 , 
 n92385 , n92386 , n92387 , n92388 , n92389 , n92390 , n92391 , n92392 , n92393 , n92394 , 
 n92395 , n92396 , n92397 , n92398 , n92399 , n92400 , n92401 , n92402 , n92403 , n92404 , 
 n92405 , n92406 , n92407 , n92408 , n92409 , n92410 , n92411 , n92412 , n92413 , n92414 , 
 n92415 , n92416 , n92417 , n92418 , n92419 , n92420 , n92421 , n92422 , n92423 , n92424 , 
 n92425 , n92426 , n92427 , n92428 , n92429 , n92430 , n92431 , n92432 , n92433 , n92434 , 
 n92435 , n92436 , n92437 , n92438 , n92439 , n92440 , n92441 , n92442 , n92443 , n92444 , 
 n92445 , n92446 , n92447 , n92448 , n92449 , n92450 , n92451 , n92452 , n92453 , n92454 , 
 n92455 , n92456 , n92457 , n92458 , n92459 , n92460 , n92461 , n92462 , n92463 , n92464 , 
 n92465 , n92466 , n92467 , n92468 , n92469 , n92470 , n92471 , n92472 , n92473 , n92474 , 
 n92475 , n92476 , n92477 , n92478 , n92479 , n92480 , n92481 , n92482 , n92483 , n92484 , 
 n92485 , n92486 , n92487 , n92488 , n92489 , n92490 , n92491 , n92492 , n92493 , n92494 , 
 n92495 , n92496 , n92497 , n92498 , n92499 , n92500 , n92501 , n92502 , n92503 , n92504 , 
 n92505 , n92506 , n92507 , n92508 , n92509 , n92510 , n92511 , n92512 , n92513 , n92514 , 
 n92515 , n92516 , n92517 , n92518 , n92519 , n92520 , n92521 , n92522 , n92523 , n92524 , 
 n92525 , n92526 , n92527 , n92528 , n92529 , n92530 , n92531 , n92532 , n92533 , n92534 , 
 n92535 , n92536 , n92537 , n92538 , n92539 , n92540 , n92541 , n92542 , n92543 , n92544 , 
 n92545 , n92546 , n92547 , n92548 , n92549 , n92550 , n92551 , n92552 , n92553 , n92554 , 
 n92555 , n92556 , n92557 , n92558 , n92559 , n92560 , n92561 , n92562 , n92563 , n92564 , 
 n92565 , n92566 , n92567 , n92568 , n92569 , n92570 , n92571 , n92572 , n92573 , n92574 , 
 n92575 , n92576 , n92577 , n92578 , n92579 , n92580 , n92581 , n92582 , n92583 , n92584 , 
 n92585 , n92586 , n92587 , n92588 , n92589 , n92590 , n92591 , n92592 , n92593 , n92594 , 
 n92595 , n92596 , n92597 , n92598 , n92599 , n92600 , n92601 , n92602 , n92603 , n92604 , 
 n92605 , n92606 , n92607 , n92608 , n92609 , n92610 , n92611 , n92612 , n92613 , n92614 , 
 n92615 , n92616 , n92617 , n92618 , n92619 , n92620 , n92621 , n92622 , n92623 , n92624 , 
 n92625 , n92626 , n92627 , n92628 , n92629 , n92630 , n92631 , n92632 , n92633 , n92634 , 
 n92635 , n92636 , n92637 , n92638 , n92639 , n92640 , n92641 , n92642 , n92643 , n92644 , 
 n92645 , n92646 , n92647 , n92648 , n92649 , n92650 , n92651 , n92652 , n92653 , n92654 , 
 n92655 , n92656 , n92657 , n92658 , n92659 , n92660 , n92661 , n92662 , n92663 , n92664 , 
 n92665 , n92666 , n92667 , n92668 , n92669 , n92670 , n92671 , n92672 , n92673 , n92674 , 
 n92675 , n92676 , n92677 , n92678 , n92679 , n92680 , n92681 , n92682 , n92683 , n92684 , 
 n92685 , n92686 , n92687 , n92688 , n92689 , n92690 , n92691 , n92692 , n92693 , n92694 , 
 n92695 , n92696 , n92697 , n92698 , n92699 , n92700 , n92701 , n92702 , n92703 , n92704 , 
 n92705 , n92706 , n92707 , n92708 , n92709 , n92710 , n92711 , n92712 , n92713 , n92714 , 
 n92715 , n92716 , n92717 , n92718 , n92719 , n92720 , n92721 , n92722 , n92723 , n92724 , 
 n92725 , n92726 , n92727 , n92728 , n92729 , n92730 , n92731 , n92732 , n92733 , n92734 , 
 n92735 , n92736 , n92737 , n92738 , n92739 , n92740 , n92741 , n92742 , n92743 , n92744 , 
 n92745 , n92746 , n92747 , n92748 , n92749 , n92750 , n92751 , n92752 , n92753 , n92754 , 
 n92755 , n92756 , n92757 , n92758 , n92759 , n92760 , n92761 , n92762 , n92763 , n92764 , 
 n92765 , n92766 , n92767 , n92768 , n92769 , n92770 , n92771 , n92772 , n92773 , n92774 , 
 n92775 , n92776 , n92777 , n92778 , n92779 , n92780 , n92781 , n92782 , n92783 , n92784 , 
 n92785 , n92786 , n92787 , n92788 , n92789 , n92790 , n92791 , n92792 , n92793 , n92794 , 
 n92795 , n92796 , n92797 , n92798 , n92799 , n92800 , n92801 , n92802 , n92803 , n92804 , 
 n92805 , n92806 , n92807 , n92808 , n92809 , n92810 , n92811 , n92812 , n92813 , n92814 , 
 n92815 , n92816 , n92817 , n92818 , n92819 , n92820 , n92821 , n92822 , n92823 , n92824 , 
 n92825 , n92826 , n92827 , n92828 , n92829 , n92830 , n92831 , n92832 , n92833 , n92834 , 
 n92835 , n92836 , n92837 , n92838 , n92839 , n92840 , n92841 , n92842 , n92843 , n92844 , 
 n92845 , n92846 , n92847 , n92848 , n92849 , n92850 , n92851 , n92852 , n92853 , n92854 , 
 n92855 , n92856 , n92857 , n92858 , n92859 , n92860 , n92861 , n92862 , n92863 , n92864 , 
 n92865 , n92866 , n92867 , n92868 , n92869 , n92870 , n92871 , n92872 , n92873 , n92874 , 
 n92875 , n92876 , n92877 , n92878 , n92879 , n92880 , n92881 , n92882 , n92883 , n92884 , 
 n92885 , n92886 , n92887 , n92888 , n92889 , n92890 , n92891 , n92892 , n92893 , n92894 , 
 n92895 , n92896 , n92897 , n92898 , n92899 , n92900 , n92901 , n92902 , n92903 , n92904 , 
 n92905 , n92906 , n92907 , n92908 , n92909 , n92910 , n92911 , n92912 , n92913 , n92914 , 
 n92915 , n92916 , n92917 , n92918 , n92919 , n92920 , n92921 , n92922 , n92923 , n92924 , 
 n92925 , n92926 , n92927 , n92928 , n92929 , n92930 , n92931 , n92932 , n92933 , n92934 , 
 n92935 , n92936 , n92937 , n92938 , n92939 , n92940 , n92941 , n92942 , n92943 , n92944 , 
 n92945 , n92946 , n92947 , n92948 , n92949 , n92950 , n92951 , n92952 , n92953 , n92954 , 
 n92955 , n92956 , n92957 , n92958 , n92959 , n92960 , n92961 , n92962 , n92963 , n92964 , 
 n92965 , n92966 , n92967 , n92968 , n92969 , n92970 , n92971 , n92972 , n92973 , n92974 , 
 n92975 , n92976 , n92977 , n92978 , n92979 , n92980 , n92981 , n92982 , n92983 , n92984 , 
 n92985 , n92986 , n92987 , n92988 , n92989 , n92990 , n92991 , n92992 , n92993 , n92994 , 
 n92995 , n92996 , n92997 , n92998 , n92999 , n93000 , n93001 , n93002 , n93003 , n93004 , 
 n93005 , n93006 , n93007 , n93008 , n93009 , n93010 , n93011 , n93012 , n93013 , n93014 , 
 n93015 , n93016 , n93017 , n93018 , n93019 , n93020 , n93021 , n93022 , n93023 , n93024 , 
 n93025 , n93026 , n93027 , n93028 , n93029 , n93030 , n93031 , n93032 , n93033 , n93034 , 
 n93035 , n93036 , n93037 , n93038 , n93039 , n93040 , n93041 , n93042 , n93043 , n93044 , 
 n93045 , n93046 , n93047 , n93048 , n93049 , n93050 , n93051 , n93052 , n93053 , n93054 , 
 n93055 , n93056 , n93057 , n93058 , n93059 , n93060 , n93061 , n93062 , n93063 , n93064 , 
 n93065 , n93066 , n93067 , n93068 , n93069 , n93070 , n93071 , n93072 , n93073 , n93074 , 
 n93075 , n93076 , n93077 , n93078 , n93079 , n93080 , n93081 , n93082 , n93083 , n93084 , 
 n93085 , n93086 , n93087 , n93088 , n93089 , n93090 , n93091 , n93092 , n93093 , n93094 , 
 n93095 , n93096 , n93097 , n93098 , n93099 , n93100 , n93101 , n93102 , n93103 , n93104 , 
 n93105 , n93106 , n93107 , n93108 , n93109 , n93110 , n93111 , n93112 , n93113 , n93114 , 
 n93115 , n93116 , n93117 , n93118 , n93119 , n93120 , n93121 , n93122 , n93123 , n93124 , 
 n93125 , n93126 , n93127 , n93128 , n93129 , n93130 , n93131 , n93132 , n93133 , n93134 , 
 n93135 , n93136 , n93137 , n93138 , n93139 , n93140 , n93141 , n93142 , n93143 , n93144 , 
 n93145 , n93146 , n93147 , n93148 , n93149 , n93150 , n93151 , n93152 , n93153 , n93154 , 
 n93155 , n93156 , n93157 , n93158 , n93159 , n93160 , n93161 , n93162 , n93163 , n93164 , 
 n93165 , n93166 , n93167 , n93168 , n93169 , n93170 , n93171 , n93172 , n93173 , n93174 , 
 n93175 , n93176 , n93177 , n93178 , n93179 , n93180 , n93181 , n93182 , n93183 , n93184 , 
 n93185 , n93186 , n93187 , n93188 , n93189 , n93190 , n93191 , n93192 , n93193 , n93194 , 
 n93195 , n93196 , n93197 , n93198 , n93199 , n93200 , n93201 , n93202 , n93203 , n93204 , 
 n93205 , n93206 , n93207 , n93208 , n93209 , n93210 , n93211 , n93212 , n93213 , n93214 , 
 n93215 , n93216 , n93217 , n93218 , n93219 , n93220 , n93221 , n93222 , n93223 , n93224 , 
 n93225 , n93226 , n93227 , n93228 , n93229 , n93230 , n93231 , n93232 , n93233 , n93234 , 
 n93235 , n93236 , n93237 , n93238 , n93239 , n93240 , n93241 , n93242 , n93243 , n93244 , 
 n93245 , n93246 , n93247 , n93248 , n93249 , n93250 , n93251 , n93252 , n93253 , n93254 , 
 n93255 , n93256 , n93257 , n93258 , n93259 , n93260 , n93261 , n93262 , n93263 , n93264 , 
 n93265 , n93266 , n93267 , n93268 , n93269 , n93270 , n93271 , n93272 , n93273 , n93274 , 
 n93275 , n93276 , n93277 , n93278 , n93279 , n93280 , n93281 , n93282 , n93283 , n93284 , 
 n93285 , n93286 , n93287 , n93288 , n93289 , n93290 , n93291 , n93292 , n93293 , n93294 , 
 n93295 , n93296 , n93297 , n93298 , n93299 , n93300 , n93301 , n93302 , n93303 , n93304 , 
 n93305 , n93306 , n93307 , n93308 , n93309 , n93310 , n93311 , n93312 , n93313 , n93314 , 
 n93315 , n93316 , n93317 , n93318 , n93319 , n93320 , n93321 , n93322 , n93323 , n93324 , 
 n93325 , n93326 , n93327 , n93328 , n93329 , n93330 , n93331 , n93332 , n93333 , n93334 , 
 n93335 , n93336 , n93337 , n93338 , n93339 , n93340 , n93341 , n93342 , n93343 , n93344 , 
 n93345 , n93346 , n93347 , n93348 , n93349 , n93350 , n93351 , n93352 , n93353 , n93354 , 
 n93355 , n93356 , n93357 , n93358 , n93359 , n93360 , n93361 , n93362 , n93363 , n93364 , 
 n93365 , n93366 , n93367 , n93368 , n93369 , n93370 , n93371 , n93372 , n93373 , n93374 , 
 n93375 , n93376 , n93377 , n93378 , n93379 , n93380 , n93381 , n93382 , n93383 , n93384 , 
 n93385 , n93386 , n93387 , n93388 , n93389 , n93390 , n93391 , n93392 , n93393 , n93394 , 
 n93395 , n93396 , n93397 , n93398 , n93399 , n93400 , n93401 , n93402 , n93403 , n93404 , 
 n93405 , n93406 , n93407 , n93408 , n93409 , n93410 , n93411 , n93412 , n93413 , n93414 , 
 n93415 , n93416 , n93417 , n93418 , n93419 , n93420 , n93421 , n93422 , n93423 , n93424 , 
 n93425 , n93426 , n93427 , n93428 , n93429 , n93430 , n93431 , n93432 , n93433 , n93434 , 
 n93435 , n93436 , n93437 , n93438 , n93439 , n93440 , n93441 , n93442 , n93443 , n93444 , 
 n93445 , n93446 , n93447 , n93448 , n93449 , n93450 , n93451 , n93452 , n93453 , n93454 , 
 n93455 , n93456 , n93457 , n93458 , n93459 , n93460 , n93461 , n93462 , n93463 , n93464 , 
 n93465 , n93466 , n93467 , n93468 , n93469 , n93470 , n93471 , n93472 , n93473 , n93474 , 
 n93475 , n93476 , n93477 , n93478 , n93479 , n93480 , n93481 , n93482 , n93483 , n93484 , 
 n93485 , n93486 , n93487 , n93488 , n93489 , n93490 , n93491 , n93492 , n93493 , n93494 , 
 n93495 , n93496 , n93497 , n93498 , n93499 , n93500 , n93501 , n93502 , n93503 , n93504 , 
 n93505 , n93506 , n93507 , n93508 , n93509 , n93510 , n93511 , n93512 , n93513 , n93514 , 
 n93515 , n93516 , n93517 , n93518 , n93519 , n93520 , n93521 , n93522 , n93523 , n93524 , 
 n93525 , n93526 , n93527 , n93528 , n93529 , n93530 , n93531 , n93532 , n93533 , n93534 , 
 n93535 , n93536 , n93537 , n93538 , n93539 , n93540 , n93541 , n93542 , n93543 , n93544 , 
 n93545 , n93546 , n93547 , n93548 , n93549 , n93550 , n93551 , n93552 , n93553 , n93554 , 
 n93555 , n93556 , n93557 , n93558 , n93559 , n93560 , n93561 , n93562 , n93563 , n93564 , 
 n93565 , n93566 , n93567 , n93568 , n93569 , n93570 , n93571 , n93572 , n93573 , n93574 , 
 n93575 , n93576 , n93577 , n93578 , n93579 , n93580 , n93581 , n93582 , n93583 , n93584 , 
 n93585 , n93586 , n93587 , n93588 , n93589 , n93590 , n93591 , n93592 , n93593 , n93594 , 
 n93595 , n93596 , n93597 , n93598 , n93599 , n93600 , n93601 , n93602 , n93603 , n93604 , 
 n93605 , n93606 , n93607 , n93608 , n93609 , n93610 , n93611 , n93612 , n93613 , n93614 , 
 n93615 , n93616 , n93617 , n93618 , n93619 , n93620 , n93621 , n93622 , n93623 , n93624 , 
 n93625 , n93626 , n93627 , n93628 , n93629 , n93630 , n93631 , n93632 , n93633 , n93634 , 
 n93635 , n93636 , n93637 , n93638 , n93639 , n93640 , n93641 , n93642 , n93643 , n93644 , 
 n93645 , n93646 , n93647 , n93648 , n93649 , n93650 , n93651 , n93652 , n93653 , n93654 , 
 n93655 , n93656 , n93657 , n93658 , n93659 , n93660 , n93661 , n93662 , n93663 , n93664 , 
 n93665 , n93666 , n93667 , n93668 , n93669 , n93670 , n93671 , n93672 , n93673 , n93674 , 
 n93675 , n93676 , n93677 , n93678 , n93679 , n93680 , n93681 , n93682 , n93683 , n93684 , 
 n93685 , n93686 , n93687 , n93688 , n93689 , n93690 , n93691 , n93692 , n93693 , n93694 , 
 n93695 , n93696 , n93697 , n93698 , n93699 , n93700 , n93701 , n93702 , n93703 , n93704 , 
 n93705 , n93706 , n93707 , n93708 , n93709 , n93710 , n93711 , n93712 , n93713 , n93714 , 
 n93715 , n93716 , n93717 , n93718 , n93719 , n93720 , n93721 , n93722 , n93723 , n93724 , 
 n93725 , n93726 , n93727 , n93728 , n93729 , n93730 , n93731 , n93732 , n93733 , n93734 , 
 n93735 , n93736 , n93737 , n93738 , n93739 , n93740 , n93741 , n93742 , n93743 , n93744 , 
 n93745 , n93746 , n93747 , n93748 , n93749 , n93750 , n93751 , n93752 , n93753 , n93754 , 
 n93755 , n93756 , n93757 , n93758 , n93759 , n93760 , n93761 , n93762 , n93763 , n93764 , 
 n93765 , n93766 , n93767 , n93768 , n93769 , n93770 , n93771 , n93772 , n93773 , n93774 , 
 n93775 , n93776 , n93777 , n93778 , n93779 , n93780 , n93781 , n93782 , n93783 , n93784 , 
 n93785 , n93786 , n93787 , n93788 , n93789 , n93790 , n93791 , n93792 , n93793 , n93794 , 
 n93795 , n93796 , n93797 , n93798 , n93799 , n93800 , n93801 , n93802 , n93803 , n93804 , 
 n93805 , n93806 , n93807 , n93808 , n93809 , n93810 , n93811 , n93812 , n93813 , n93814 , 
 n93815 , n93816 , n93817 , n93818 , n93819 , n93820 , n93821 , n93822 , n93823 , n93824 , 
 n93825 , n93826 , n93827 , n93828 , n93829 , n93830 , n93831 , n93832 , n93833 , n93834 , 
 n93835 , n93836 , n93837 , n93838 , n93839 , n93840 , n93841 , n93842 , n93843 , n93844 , 
 n93845 , n93846 , n93847 , n93848 , n93849 , n93850 , n93851 , n93852 , n93853 , n93854 , 
 n93855 , n93856 , n93857 , n93858 , n93859 , n93860 , n93861 , n93862 , n93863 , n93864 , 
 n93865 , n93866 , n93867 , n93868 , n93869 , n93870 , n93871 , n93872 , n93873 , n93874 , 
 n93875 , n93876 , n93877 , n93878 , n93879 , n93880 , n93881 , n93882 , n93883 , n93884 , 
 n93885 , n93886 , n93887 , n93888 , n93889 , n93890 , n93891 , n93892 , n93893 , n93894 , 
 n93895 , n93896 , n93897 , n93898 , n93899 , n93900 , n93901 , n93902 , n93903 , n93904 , 
 n93905 , n93906 , n93907 , n93908 , n93909 , n93910 , n93911 , n93912 , n93913 , n93914 , 
 n93915 , n93916 , n93917 , n93918 , n93919 , n93920 , n93921 , n93922 , n93923 , n93924 , 
 n93925 , n93926 , n93927 , n93928 , n93929 , n93930 , n93931 , n93932 , n93933 , n93934 , 
 n93935 , n93936 , n93937 , n93938 , n93939 , n93940 , n93941 , n93942 , n93943 , n93944 , 
 n93945 , n93946 , n93947 , n93948 , n93949 , n93950 , n93951 , n93952 , n93953 , n93954 , 
 n93955 , n93956 , n93957 , n93958 , n93959 , n93960 , n93961 , n93962 , n93963 , n93964 , 
 n93965 , n93966 , n93967 , n93968 , n93969 , n93970 , n93971 , n93972 , n93973 , n93974 , 
 n93975 , n93976 , n93977 , n93978 , n93979 , n93980 , n93981 , n93982 , n93983 , n93984 , 
 n93985 , n93986 , n93987 , n93988 , n93989 , n93990 , n93991 , n93992 , n93993 , n93994 , 
 n93995 , n93996 , n93997 , n93998 , n93999 , n94000 , n94001 , n94002 , n94003 , n94004 , 
 n94005 , n94006 , n94007 , n94008 , n94009 , n94010 , n94011 , n94012 , n94013 , n94014 , 
 n94015 , n94016 , n94017 , n94018 , n94019 , n94020 , n94021 , n94022 , n94023 , n94024 , 
 n94025 , n94026 , n94027 , n94028 , n94029 , n94030 , n94031 , n94032 , n94033 , n94034 , 
 n94035 , n94036 , n94037 , n94038 , n94039 , n94040 , n94041 , n94042 , n94043 , n94044 , 
 n94045 , n94046 , n94047 , n94048 , n94049 , n94050 , n94051 , n94052 , n94053 , n94054 , 
 n94055 , n94056 , n94057 , n94058 , n94059 , n94060 , n94061 , n94062 , n94063 , n94064 , 
 n94065 , n94066 , n94067 , n94068 , n94069 , n94070 , n94071 , n94072 , n94073 , n94074 , 
 n94075 , n94076 , n94077 , n94078 , n94079 , n94080 , n94081 , n94082 , n94083 , n94084 , 
 n94085 , n94086 , n94087 , n94088 , n94089 , n94090 , n94091 , n94092 , n94093 , n94094 , 
 n94095 , n94096 , n94097 , n94098 , n94099 , n94100 , n94101 , n94102 , n94103 , n94104 , 
 n94105 , n94106 , n94107 , n94108 , n94109 , n94110 , n94111 , n94112 , n94113 , n94114 , 
 n94115 , n94116 , n94117 , n94118 , n94119 , n94120 , n94121 , n94122 , n94123 , n94124 , 
 n94125 , n94126 , n94127 , n94128 , n94129 , n94130 , n94131 , n94132 , n94133 , n94134 , 
 n94135 , n94136 , n94137 , n94138 , n94139 , n94140 , n94141 , n94142 , n94143 , n94144 , 
 n94145 , n94146 , n94147 , n94148 , n94149 , n94150 , n94151 , n94152 , n94153 , n94154 , 
 n94155 , n94156 , n94157 , n94158 , n94159 , n94160 , n94161 , n94162 , n94163 , n94164 , 
 n94165 , n94166 , n94167 , n94168 , n94169 , n94170 , n94171 , n94172 , n94173 , n94174 , 
 n94175 , n94176 , n94177 , n94178 , n94179 , n94180 , n94181 , n94182 , n94183 , n94184 , 
 n94185 , n94186 , n94187 , n94188 , n94189 , n94190 , n94191 , n94192 , n94193 , n94194 , 
 n94195 , n94196 , n94197 , n94198 , n94199 , n94200 , n94201 , n94202 , n94203 , n94204 , 
 n94205 , n94206 , n94207 , n94208 , n94209 , n94210 , n94211 , n94212 , n94213 , n94214 , 
 n94215 , n94216 , n94217 , n94218 , n94219 , n94220 , n94221 , n94222 , n94223 , n94224 , 
 n94225 , n94226 , n94227 , n94228 , n94229 , n94230 , n94231 , n94232 , n94233 , n94234 , 
 n94235 , n94236 , n94237 , n94238 , n94239 , n94240 , n94241 , n94242 , n94243 , n94244 , 
 n94245 , n94246 , n94247 , n94248 , n94249 , n94250 , n94251 , n94252 , n94253 , n94254 , 
 n94255 , n94256 , n94257 , n94258 , n94259 , n94260 , n94261 , n94262 , n94263 , n94264 , 
 n94265 , n94266 , n94267 , n94268 , n94269 , n94270 , n94271 , n94272 , n94273 , n94274 , 
 n94275 , n94276 , n94277 , n94278 , n94279 , n94280 , n94281 , n94282 , n94283 , n94284 , 
 n94285 , n94286 , n94287 , n94288 , n94289 , n94290 , n94291 , n94292 , n94293 , n94294 , 
 n94295 , n94296 , n94297 , n94298 , n94299 , n94300 , n94301 , n94302 , n94303 , n94304 , 
 n94305 , n94306 , n94307 , n94308 , n94309 , n94310 , n94311 , n94312 , n94313 , n94314 , 
 n94315 , n94316 , n94317 , n94318 , n94319 , n94320 , n94321 , n94322 , n94323 , n94324 , 
 n94325 , n94326 , n94327 , n94328 , n94329 , n94330 , n94331 , n94332 , n94333 , n94334 , 
 n94335 , n94336 , n94337 , n94338 , n94339 , n94340 , n94341 , n94342 , n94343 , n94344 , 
 n94345 , n94346 , n94347 , n94348 , n94349 , n94350 , n94351 , n94352 , n94353 , n94354 , 
 n94355 , n94356 , n94357 , n94358 , n94359 , n94360 , n94361 , n94362 , n94363 , n94364 , 
 n94365 , n94366 , n94367 , n94368 , n94369 , n94370 , n94371 , n94372 , n94373 , n94374 , 
 n94375 , n94376 , n94377 , n94378 , n94379 , n94380 , n94381 , n94382 , n94383 , n94384 , 
 n94385 , n94386 , n94387 , n94388 , n94389 , n94390 , n94391 , n94392 , n94393 , n94394 , 
 n94395 , n94396 , n94397 , n94398 , n94399 , n94400 , n94401 , n94402 , n94403 , n94404 , 
 n94405 , n94406 , n94407 , n94408 , n94409 , n94410 , n94411 , n94412 , n94413 , n94414 , 
 n94415 , n94416 , n94417 , n94418 , n94419 , n94420 , n94421 , n94422 , n94423 , n94424 , 
 n94425 , n94426 , n94427 , n94428 , n94429 , n94430 , n94431 , n94432 , n94433 , n94434 , 
 n94435 , n94436 , n94437 , n94438 , n94439 , n94440 , n94441 , n94442 , n94443 , n94444 , 
 n94445 , n94446 , n94447 , n94448 , n94449 , n94450 , n94451 , n94452 , n94453 , n94454 , 
 n94455 , n94456 , n94457 , n94458 , n94459 , n94460 , n94461 , n94462 , n94463 , n94464 , 
 n94465 , n94466 , n94467 , n94468 , n94469 , n94470 , n94471 , n94472 , n94473 , n94474 , 
 n94475 , n94476 , n94477 , n94478 , n94479 , n94480 , n94481 , n94482 , n94483 , n94484 , 
 n94485 , n94486 , n94487 , n94488 , n94489 , n94490 , n94491 , n94492 , n94493 , n94494 , 
 n94495 , n94496 , n94497 , n94498 , n94499 , n94500 , n94501 , n94502 , n94503 , n94504 , 
 n94505 , n94506 , n94507 , n94508 , n94509 , n94510 , n94511 , n94512 , n94513 , n94514 , 
 n94515 , n94516 , n94517 , n94518 , n94519 , n94520 , n94521 , n94522 , n94523 , n94524 , 
 n94525 , n94526 , n94527 , n94528 , n94529 , n94530 , n94531 , n94532 , n94533 , n94534 , 
 n94535 , n94536 , n94537 , n94538 , n94539 , n94540 , n94541 , n94542 , n94543 , n94544 , 
 n94545 , n94546 , n94547 , n94548 , n94549 , n94550 , n94551 , n94552 , n94553 , n94554 , 
 n94555 , n94556 , n94557 , n94558 , n94559 , n94560 , n94561 , n94562 , n94563 , n94564 , 
 n94565 , n94566 , n94567 , n94568 , n94569 , n94570 , n94571 , n94572 , n94573 , n94574 , 
 n94575 , n94576 , n94577 , n94578 , n94579 , n94580 , n94581 , n94582 , n94583 , n94584 , 
 n94585 , n94586 , n94587 , n94588 , n94589 , n94590 , n94591 , n94592 , n94593 , n94594 , 
 n94595 , n94596 , n94597 , n94598 , n94599 , n94600 , n94601 , n94602 , n94603 , n94604 , 
 n94605 , n94606 , n94607 , n94608 , n94609 , n94610 , n94611 , n94612 , n94613 , n94614 , 
 n94615 , n94616 , n94617 , n94618 , n94619 , n94620 , n94621 , n94622 , n94623 , n94624 , 
 n94625 , n94626 , n94627 , n94628 , n94629 , n94630 , n94631 , n94632 , n94633 , n94634 , 
 n94635 , n94636 , n94637 , n94638 , n94639 , n94640 , n94641 , n94642 , n94643 , n94644 , 
 n94645 , n94646 , n94647 , n94648 , n94649 , n94650 , n94651 , n94652 , n94653 , n94654 , 
 n94655 , n94656 , n94657 , n94658 , n94659 , n94660 , n94661 , n94662 , n94663 , n94664 , 
 n94665 , n94666 , n94667 , n94668 , n94669 , n94670 , n94671 , n94672 , n94673 , n94674 , 
 n94675 , n94676 , n94677 , n94678 , n94679 , n94680 , n94681 , n94682 , n94683 , n94684 , 
 n94685 , n94686 , n94687 , n94688 , n94689 , n94690 , n94691 , n94692 , n94693 , n94694 , 
 n94695 , n94696 , n94697 , n94698 , n94699 , n94700 , n94701 , n94702 , n94703 , n94704 , 
 n94705 , n94706 , n94707 , n94708 , n94709 , n94710 , n94711 , n94712 , n94713 , n94714 , 
 n94715 , n94716 , n94717 , n94718 , n94719 , n94720 , n94721 , n94722 , n94723 , n94724 , 
 n94725 , n94726 , n94727 , n94728 , n94729 , n94730 , n94731 , n94732 , n94733 , n94734 , 
 n94735 , n94736 , n94737 , n94738 , n94739 , n94740 , n94741 , n94742 , n94743 , n94744 , 
 n94745 , n94746 , n94747 , n94748 , n94749 , n94750 , n94751 , n94752 , n94753 , n94754 , 
 n94755 , n94756 , n94757 , n94758 , n94759 , n94760 , n94761 , n94762 , n94763 , n94764 , 
 n94765 , n94766 , n94767 , n94768 , n94769 , n94770 , n94771 , n94772 , n94773 , n94774 , 
 n94775 , n94776 , n94777 , n94778 , n94779 , n94780 , n94781 , n94782 , n94783 , n94784 , 
 n94785 , n94786 , n94787 , n94788 , n94789 , n94790 , n94791 , n94792 , n94793 , n94794 , 
 n94795 , n94796 , n94797 , n94798 , n94799 , n94800 , n94801 , n94802 , n94803 , n94804 , 
 n94805 , n94806 , n94807 , n94808 , n94809 , n94810 , n94811 , n94812 , n94813 , n94814 , 
 n94815 , n94816 , n94817 , n94818 , n94819 , n94820 , n94821 , n94822 , n94823 , n94824 , 
 n94825 , n94826 , n94827 , n94828 , n94829 , n94830 , n94831 , n94832 , n94833 , n94834 , 
 n94835 , n94836 , n94837 , n94838 , n94839 , n94840 , n94841 , n94842 , n94843 , n94844 , 
 n94845 , n94846 , n94847 , n94848 , n94849 , n94850 , n94851 , n94852 , n94853 , n94854 , 
 n94855 , n94856 , n94857 , n94858 , n94859 , n94860 , n94861 , n94862 , n94863 , n94864 , 
 n94865 , n94866 , n94867 , n94868 , n94869 , n94870 , n94871 , n94872 , n94873 , n94874 , 
 n94875 , n94876 , n94877 , n94878 , n94879 , n94880 , n94881 , n94882 , n94883 , n94884 , 
 n94885 , n94886 , n94887 , n94888 , n94889 , n94890 , n94891 , n94892 , n94893 , n94894 , 
 n94895 , n94896 , n94897 , n94898 , n94899 , n94900 , n94901 , n94902 , n94903 , n94904 , 
 n94905 , n94906 , n94907 , n94908 , n94909 , n94910 , n94911 , n94912 , n94913 , n94914 , 
 n94915 , n94916 , n94917 , n94918 , n94919 , n94920 , n94921 , n94922 , n94923 , n94924 , 
 n94925 , n94926 , n94927 , n94928 , n94929 , n94930 , n94931 , n94932 , n94933 , n94934 , 
 n94935 , n94936 , n94937 , n94938 , n94939 , n94940 , n94941 , n94942 , n94943 , n94944 , 
 n94945 , n94946 , n94947 , n94948 , n94949 , n94950 , n94951 , n94952 , n94953 , n94954 , 
 n94955 , n94956 , n94957 , n94958 , n94959 , n94960 , n94961 , n94962 , n94963 , n94964 , 
 n94965 , n94966 , n94967 , n94968 , n94969 , n94970 , n94971 , n94972 , n94973 , n94974 , 
 n94975 , n94976 , n94977 , n94978 , n94979 , n94980 , n94981 , n94982 , n94983 , n94984 , 
 n94985 , n94986 , n94987 , n94988 , n94989 , n94990 , n94991 , n94992 , n94993 , n94994 , 
 n94995 , n94996 , n94997 , n94998 , n94999 , n95000 , n95001 , n95002 , n95003 , n95004 , 
 n95005 , n95006 , n95007 , n95008 , n95009 , n95010 , n95011 , n95012 , n95013 , n95014 , 
 n95015 , n95016 , n95017 , n95018 , n95019 , n95020 , n95021 , n95022 , n95023 , n95024 , 
 n95025 , n95026 , n95027 , n95028 , n95029 , n95030 , n95031 , n95032 , n95033 , n95034 , 
 n95035 , n95036 , n95037 , n95038 , n95039 , n95040 , n95041 , n95042 , n95043 , n95044 , 
 n95045 , n95046 , n95047 , n95048 , n95049 , n95050 , n95051 , n95052 , n95053 , n95054 , 
 C0n , C0 , C1n , C1 ;
buf ( n544 , n0 );
buf ( n545 , n1 );
buf ( n546 , n2 );
buf ( n547 , n3 );
buf ( n548 , n4 );
buf ( n549 , n5 );
buf ( n550 , n6 );
buf ( n551 , n7 );
buf ( n552 , n8 );
buf ( n553 , n9 );
buf ( n554 , n10 );
buf ( n555 , n11 );
buf ( n556 , n12 );
buf ( n557 , n13 );
buf ( n558 , n14 );
buf ( n559 , n15 );
buf ( n560 , n16 );
buf ( n561 , n17 );
buf ( n562 , n18 );
buf ( n563 , n19 );
buf ( n564 , n20 );
buf ( n565 , n21 );
buf ( n566 , n22 );
buf ( n567 , n23 );
buf ( n568 , n24 );
buf ( n569 , n25 );
buf ( n570 , n26 );
buf ( n571 , n27 );
buf ( n572 , n28 );
buf ( n573 , n29 );
buf ( n574 , n30 );
buf ( n575 , n31 );
buf ( n576 , n32 );
buf ( n577 , n33 );
buf ( n578 , n34 );
buf ( n579 , n35 );
buf ( n580 , n36 );
buf ( n581 , n37 );
buf ( n582 , n38 );
buf ( n583 , n39 );
buf ( n584 , n40 );
buf ( n585 , n41 );
buf ( n586 , n42 );
buf ( n587 , n43 );
buf ( n588 , n44 );
buf ( n589 , n45 );
buf ( n590 , n46 );
buf ( n591 , n47 );
buf ( n592 , n48 );
buf ( n593 , n49 );
buf ( n594 , n50 );
buf ( n595 , n51 );
buf ( n596 , n52 );
buf ( n597 , n53 );
buf ( n598 , n54 );
buf ( n599 , n55 );
buf ( n600 , n56 );
buf ( n601 , n57 );
buf ( n602 , n58 );
buf ( n603 , n59 );
buf ( n604 , n60 );
buf ( n605 , n61 );
buf ( n606 , n62 );
buf ( n607 , n63 );
buf ( n608 , n64 );
buf ( n609 , n65 );
buf ( n610 , n66 );
buf ( n611 , n67 );
buf ( n612 , n68 );
buf ( n613 , n69 );
buf ( n614 , n70 );
buf ( n615 , n71 );
buf ( n616 , n72 );
buf ( n617 , n73 );
buf ( n618 , n74 );
buf ( n619 , n75 );
buf ( n620 , n76 );
buf ( n621 , n77 );
buf ( n622 , n78 );
buf ( n623 , n79 );
buf ( n80 , n624 );
buf ( n81 , n625 );
buf ( n82 , n626 );
buf ( n83 , n627 );
buf ( n84 , n628 );
buf ( n85 , n629 );
buf ( n86 , n630 );
buf ( n87 , n631 );
buf ( n88 , n632 );
buf ( n89 , n633 );
buf ( n90 , n634 );
buf ( n91 , n635 );
buf ( n92 , n636 );
buf ( n93 , n637 );
buf ( n94 , n638 );
buf ( n95 , n639 );
buf ( n96 , n640 );
buf ( n97 , n641 );
buf ( n98 , n642 );
buf ( n99 , n643 );
buf ( n100 , n644 );
buf ( n101 , n645 );
buf ( n102 , n646 );
buf ( n103 , n647 );
buf ( n104 , n648 );
buf ( n105 , n649 );
buf ( n106 , n650 );
buf ( n107 , n651 );
buf ( n108 , n652 );
buf ( n109 , n653 );
buf ( n110 , n654 );
buf ( n111 , n655 );
buf ( n112 , n656 );
buf ( n113 , n657 );
buf ( n114 , n658 );
buf ( n115 , n659 );
buf ( n116 , n660 );
buf ( n117 , n661 );
buf ( n118 , n662 );
buf ( n119 , n663 );
buf ( n120 , n664 );
buf ( n121 , n665 );
buf ( n122 , n666 );
buf ( n123 , n667 );
buf ( n124 , n668 );
buf ( n125 , n669 );
buf ( n126 , n670 );
buf ( n127 , n671 );
buf ( n128 , n672 );
buf ( n129 , n673 );
buf ( n130 , n674 );
buf ( n131 , n675 );
buf ( n132 , n676 );
buf ( n133 , n677 );
buf ( n134 , n678 );
buf ( n135 , n679 );
buf ( n136 , n680 );
buf ( n137 , n681 );
buf ( n138 , n682 );
buf ( n139 , n683 );
buf ( n140 , n684 );
buf ( n141 , n685 );
buf ( n142 , n686 );
buf ( n143 , n687 );
buf ( n144 , n688 );
buf ( n145 , n689 );
buf ( n146 , n690 );
buf ( n147 , n691 );
buf ( n148 , n692 );
buf ( n149 , n693 );
buf ( n150 , n694 );
buf ( n151 , n695 );
buf ( n152 , n696 );
buf ( n153 , n697 );
buf ( n154 , n698 );
buf ( n155 , n699 );
buf ( n156 , n700 );
buf ( n157 , n701 );
buf ( n158 , n702 );
buf ( n159 , n703 );
buf ( n160 , n704 );
buf ( n161 , n705 );
buf ( n162 , n706 );
buf ( n163 , n707 );
buf ( n164 , n708 );
buf ( n165 , n709 );
buf ( n166 , n710 );
buf ( n167 , n711 );
buf ( n168 , n712 );
buf ( n169 , n713 );
buf ( n170 , n714 );
buf ( n171 , n715 );
buf ( n172 , n716 );
buf ( n173 , n717 );
buf ( n174 , n718 );
buf ( n175 , n719 );
buf ( n176 , n720 );
buf ( n177 , n721 );
buf ( n178 , n722 );
buf ( n179 , n723 );
buf ( n180 , n724 );
buf ( n181 , n725 );
buf ( n182 , n726 );
buf ( n183 , n727 );
buf ( n184 , n728 );
buf ( n185 , n729 );
buf ( n186 , n730 );
buf ( n187 , n731 );
buf ( n188 , n732 );
buf ( n189 , n733 );
buf ( n190 , n734 );
buf ( n191 , n735 );
buf ( n192 , n736 );
buf ( n193 , n737 );
buf ( n194 , n738 );
buf ( n195 , n739 );
buf ( n196 , n740 );
buf ( n197 , n741 );
buf ( n198 , n742 );
buf ( n199 , n743 );
buf ( n200 , n744 );
buf ( n201 , n745 );
buf ( n202 , n746 );
buf ( n203 , n747 );
buf ( n204 , n748 );
buf ( n205 , n749 );
buf ( n206 , n750 );
buf ( n207 , n751 );
buf ( n208 , n752 );
buf ( n209 , n753 );
buf ( n210 , n754 );
buf ( n211 , n755 );
buf ( n212 , n756 );
buf ( n213 , n757 );
buf ( n214 , n758 );
buf ( n215 , n759 );
buf ( n216 , n760 );
buf ( n217 , n761 );
buf ( n218 , n762 );
buf ( n219 , n763 );
buf ( n220 , n764 );
buf ( n221 , n765 );
buf ( n222 , n766 );
buf ( n223 , n767 );
buf ( n224 , n768 );
buf ( n225 , n769 );
buf ( n226 , n770 );
buf ( n227 , n771 );
buf ( n228 , n772 );
buf ( n229 , n773 );
buf ( n230 , n774 );
buf ( n231 , n775 );
buf ( n232 , n776 );
buf ( n233 , n777 );
buf ( n234 , n778 );
buf ( n235 , n779 );
buf ( n236 , n780 );
buf ( n237 , n781 );
buf ( n238 , n782 );
buf ( n239 , n783 );
buf ( n240 , n784 );
buf ( n241 , n785 );
buf ( n242 , n786 );
buf ( n243 , n787 );
buf ( n244 , n788 );
buf ( n245 , n789 );
buf ( n246 , n790 );
buf ( n247 , n791 );
buf ( n248 , n792 );
buf ( n249 , n793 );
buf ( n250 , n794 );
buf ( n251 , n795 );
buf ( n252 , n796 );
buf ( n253 , n797 );
buf ( n254 , n798 );
buf ( n255 , n799 );
buf ( n256 , n800 );
buf ( n257 , n801 );
buf ( n258 , n802 );
buf ( n259 , n803 );
buf ( n260 , n804 );
buf ( n261 , n805 );
buf ( n262 , n806 );
buf ( n263 , n807 );
buf ( n264 , n808 );
buf ( n265 , n809 );
buf ( n266 , n810 );
buf ( n267 , n811 );
buf ( n268 , n812 );
buf ( n269 , n813 );
buf ( n270 , n814 );
buf ( n271 , n815 );
buf ( n624 , n25691 );
buf ( n625 , n25709 );
buf ( n626 , n25712 );
buf ( n627 , n25715 );
buf ( n628 , n25718 );
buf ( n629 , n25721 );
buf ( n630 , n25724 );
buf ( n631 , n25727 );
buf ( n632 , n25730 );
buf ( n633 , n25733 );
buf ( n634 , n25736 );
buf ( n635 , n25739 );
buf ( n636 , n25742 );
buf ( n637 , n25745 );
buf ( n638 , n25759 );
buf ( n639 , n25773 );
buf ( n640 , n25787 );
buf ( n641 , n25795 );
buf ( n642 , n25803 );
buf ( n643 , n95036 );
buf ( n644 , n95051 );
buf ( n645 , n25815 );
buf ( n646 , n25823 );
buf ( n647 , n25826 );
buf ( n648 , n25874 );
buf ( n649 , n95038 );
buf ( n650 , n95054 );
buf ( n651 , n25834 );
buf ( n652 , n25837 );
buf ( n653 , n25856 );
buf ( n654 , n25858 );
buf ( n655 , n1531 );
buf ( n656 , n30241 );
buf ( n657 , n30259 );
buf ( n658 , n30262 );
buf ( n659 , n30265 );
buf ( n660 , n30268 );
buf ( n661 , n30271 );
buf ( n662 , n95032 );
buf ( n663 , n95035 );
buf ( n664 , n30490 );
buf ( n665 , n30486 );
buf ( n666 , n30482 );
buf ( n667 , n30478 );
buf ( n668 , n30470 );
buf ( n669 , n30466 );
buf ( n670 , n30289 );
buf ( n671 , n30301 );
buf ( n672 , n30319 );
buf ( n673 , n30333 );
buf ( n674 , n30347 );
buf ( n675 , n95017 );
buf ( n676 , n30359 );
buf ( n677 , n30362 );
buf ( n678 , n30370 );
buf ( n679 , n30378 );
buf ( n680 , n30386 );
buf ( n681 , n30398 );
buf ( n682 , n30401 );
buf ( n683 , n30404 );
buf ( n684 , n30407 );
buf ( n685 , n30410 );
buf ( n686 , n95020 );
buf ( n687 , n1542 );
buf ( n688 , n94902 );
buf ( n689 , n94902 );
buf ( n690 , n94902 );
buf ( n691 , n94902 );
buf ( n692 , n94902 );
buf ( n693 , n94902 );
buf ( n694 , n94902 );
buf ( n695 , n94902 );
buf ( n696 , n94902 );
buf ( n697 , n94902 );
buf ( n698 , n94902 );
buf ( n699 , n94902 );
buf ( n700 , n94902 );
buf ( n701 , n94902 );
buf ( n702 , n94902 );
buf ( n703 , n94902 );
buf ( n704 , n94902 );
buf ( n705 , n94902 );
buf ( n706 , n94902 );
buf ( n707 , n94902 );
buf ( n708 , n94902 );
buf ( n709 , n94902 );
buf ( n710 , n94902 );
buf ( n711 , n94902 );
buf ( n712 , n94902 );
buf ( n713 , n94902 );
buf ( n714 , n94902 );
buf ( n715 , n94902 );
buf ( n716 , n94838 );
buf ( n717 , n94853 );
buf ( n718 , n95050 );
buf ( n719 , n93173 );
buf ( n720 , n94780 );
buf ( n721 , n93208 );
buf ( n722 , n93284 );
buf ( n723 , n93234 );
buf ( n724 , n93393 );
buf ( n725 , n94973 );
buf ( n726 , n93309 );
buf ( n727 , n93265 );
buf ( n728 , n93408 );
buf ( n729 , n93434 );
buf ( n730 , n93464 );
buf ( n731 , n93381 );
buf ( n732 , n93969 );
buf ( n733 , n93495 );
buf ( n734 , n93359 );
buf ( n735 , n93521 );
buf ( n736 , n93551 );
buf ( n737 , n93577 );
buf ( n738 , n94878 );
buf ( n739 , n94865 );
buf ( n740 , n93986 );
buf ( n741 , n93605 );
buf ( n742 , n93627 );
buf ( n743 , n93654 );
buf ( n744 , n94001 );
buf ( n745 , n94799 );
buf ( n746 , n94997 );
buf ( n747 , n93820 );
buf ( n748 , n94704 );
buf ( n749 , n93722 );
buf ( n750 , n93777 );
buf ( n751 , n93795 );
buf ( n752 , n94040 );
buf ( n753 , n93928 );
buf ( n754 , n94027 );
buf ( n755 , n93952 );
buf ( n756 , n94102 );
buf ( n757 , n94899 );
buf ( n758 , n93888 );
buf ( n759 , n93865 );
buf ( n760 , n94090 );
buf ( n761 , n94156 );
buf ( n762 , n94129 );
buf ( n763 , n94813 );
buf ( n764 , n94941 );
buf ( n765 , n94803 );
buf ( n766 , n94075 );
buf ( n767 , n94908 );
buf ( n768 , n94916 );
buf ( n769 , n94738 );
buf ( n770 , n94210 );
buf ( n771 , n94233 );
buf ( n772 , n94742 );
buf ( n773 , n94274 );
buf ( n774 , n94289 );
buf ( n775 , n94315 );
buf ( n776 , n94949 );
buf ( n777 , n94991 );
buf ( n778 , n94346 );
buf ( n779 , n94960 );
buf ( n780 , n94721 );
buf ( n781 , n94372 );
buf ( n782 , n94709 );
buf ( n783 , n94952 );
buf ( n784 , n94717 );
buf ( n785 , n94936 );
buf ( n786 , n94424 );
buf ( n787 , n94439 );
buf ( n788 , n94461 );
buf ( n789 , n95004 );
buf ( n790 , n94888 );
buf ( n791 , n95000 );
buf ( n792 , n94464 );
buf ( n793 , n94478 );
buf ( n794 , n94492 );
buf ( n795 , n94510 );
buf ( n796 , n94746 );
buf ( n797 , n94921 );
buf ( n798 , n94926 );
buf ( n799 , n95029 );
buf ( n800 , n94538 );
buf ( n801 , n94771 );
buf ( n802 , n94555 );
buf ( n803 , n94558 );
buf ( n804 , n94572 );
buf ( n805 , n95011 );
buf ( n806 , n94590 );
buf ( n807 , n94612 );
buf ( n808 , n94615 );
buf ( n809 , n94617 );
buf ( n810 , n94619 );
buf ( n811 , n94629 );
buf ( n812 , n94632 );
buf ( n813 , n94642 );
buf ( n814 , n94692 );
buf ( n815 , n94696 );
buf ( n816 , n598 );
not ( n817 , n816 );
buf ( n818 , n817 );
or ( n819 , n818 , n597 );
buf ( n820 , n597 );
not ( n821 , n820 );
buf ( n822 , n821 );
or ( n823 , n822 , n598 );
nand ( n824 , n819 , n823 );
buf ( n825 , n824 );
buf ( n826 , n825 );
not ( n827 , n826 );
buf ( n828 , n596 );
not ( n829 , n828 );
buf ( n830 , n559 );
buf ( n831 , n570 );
xor ( n832 , n830 , n831 );
buf ( n833 , n832 );
buf ( n834 , n833 );
not ( n835 , n834 );
buf ( n836 , n571 );
buf ( n837 , n572 );
xor ( n838 , n836 , n837 );
buf ( n839 , n838 );
buf ( n840 , n839 );
not ( n841 , n840 );
buf ( n842 , n841 );
buf ( n843 , n842 );
xor ( n844 , n571 , n570 );
buf ( n845 , n844 );
nand ( n846 , n843 , n845 );
buf ( n847 , n846 );
buf ( n848 , n847 );
not ( n849 , n848 );
buf ( n850 , n849 );
buf ( n851 , n850 );
not ( n852 , n851 );
or ( n853 , n835 , n852 );
buf ( n854 , n842 );
not ( n855 , n854 );
buf ( n856 , n855 );
buf ( n857 , n856 );
buf ( n858 , n558 );
buf ( n859 , n570 );
xor ( n860 , n858 , n859 );
buf ( n861 , n860 );
buf ( n862 , n861 );
nand ( n863 , n857 , n862 );
buf ( n864 , n863 );
buf ( n865 , n864 );
nand ( n866 , n853 , n865 );
buf ( n867 , n866 );
buf ( n868 , n557 );
buf ( n869 , n572 );
xor ( n870 , n868 , n869 );
buf ( n871 , n870 );
buf ( n872 , n871 );
not ( n873 , n872 );
not ( n874 , n572 );
nand ( n875 , n874 , n573 );
not ( n876 , n875 );
not ( n877 , n573 );
nand ( n878 , n877 , n572 );
not ( n879 , n878 );
or ( n880 , n876 , n879 );
xor ( n881 , n573 , n574 );
not ( n882 , n881 );
nand ( n883 , n880 , n882 );
not ( n884 , n883 );
buf ( n885 , n884 );
not ( n886 , n885 );
or ( n887 , n873 , n886 );
buf ( n888 , n881 );
buf ( n889 , n888 );
buf ( n890 , n556 );
buf ( n891 , n572 );
xor ( n892 , n890 , n891 );
buf ( n893 , n892 );
buf ( n894 , n893 );
nand ( n895 , n889 , n894 );
buf ( n896 , n895 );
buf ( n897 , n896 );
nand ( n898 , n887 , n897 );
buf ( n899 , n898 );
xor ( n900 , n867 , n899 );
buf ( n901 , n574 );
not ( n902 , n901 );
buf ( n903 , n575 );
nor ( n904 , n902 , n903 );
buf ( n905 , n904 );
not ( n906 , n905 );
buf ( n907 , n555 );
buf ( n908 , n574 );
xor ( n909 , n907 , n908 );
buf ( n910 , n909 );
not ( n911 , n910 );
or ( n912 , n906 , n911 );
buf ( n913 , n554 );
buf ( n914 , n574 );
xor ( n915 , n913 , n914 );
buf ( n916 , n915 );
buf ( n917 , n916 );
buf ( n918 , n575 );
nand ( n919 , n917 , n918 );
buf ( n920 , n919 );
nand ( n921 , n912 , n920 );
or ( n922 , n559 , n571 );
nand ( n923 , n922 , n572 );
buf ( n924 , n559 );
buf ( n925 , n571 );
nand ( n926 , n924 , n925 );
buf ( n927 , n926 );
nand ( n928 , n923 , n927 , n570 );
not ( n929 , n928 );
and ( n930 , n921 , n929 );
not ( n931 , n921 );
and ( n932 , n931 , n928 );
nor ( n933 , n930 , n932 );
xor ( n934 , n900 , n933 );
buf ( n935 , n934 );
buf ( n936 , n905 );
not ( n937 , n936 );
buf ( n938 , n557 );
buf ( n939 , n574 );
xor ( n940 , n938 , n939 );
buf ( n941 , n940 );
buf ( n942 , n941 );
not ( n943 , n942 );
or ( n944 , n937 , n943 );
buf ( n945 , n556 );
buf ( n946 , n574 );
xor ( n947 , n945 , n946 );
buf ( n948 , n947 );
buf ( n949 , n948 );
buf ( n950 , n575 );
nand ( n951 , n949 , n950 );
buf ( n952 , n951 );
buf ( n953 , n952 );
nand ( n954 , n944 , n953 );
buf ( n955 , n954 );
buf ( n956 , n955 );
buf ( n957 , n559 );
buf ( n958 , n573 );
or ( n959 , n957 , n958 );
buf ( n960 , n574 );
nand ( n961 , n959 , n960 );
buf ( n962 , n961 );
buf ( n963 , n962 );
buf ( n964 , n559 );
buf ( n965 , n573 );
nand ( n966 , n964 , n965 );
buf ( n967 , n966 );
buf ( n968 , n967 );
buf ( n969 , n572 );
nand ( n970 , n963 , n968 , n969 );
buf ( n971 , n970 );
buf ( n972 , n971 );
not ( n973 , n972 );
buf ( n974 , n973 );
buf ( n975 , n974 );
and ( n976 , n956 , n975 );
buf ( n977 , n976 );
buf ( n978 , n977 );
xor ( n979 , n590 , n557 );
buf ( n980 , n979 );
not ( n981 , n980 );
not ( n982 , n591 );
nand ( n983 , n982 , n590 );
not ( n984 , n983 );
buf ( n985 , n984 );
not ( n986 , n985 );
or ( n987 , n981 , n986 );
and ( n988 , n556 , n590 );
not ( n989 , n556 );
not ( n990 , n590 );
and ( n991 , n989 , n990 );
nor ( n992 , n988 , n991 );
buf ( n993 , n992 );
buf ( n994 , n591 );
nand ( n995 , n993 , n994 );
buf ( n996 , n995 );
buf ( n997 , n996 );
nand ( n998 , n987 , n997 );
buf ( n999 , n998 );
buf ( n1000 , n999 );
buf ( n1001 , n559 );
buf ( n1002 , n589 );
or ( n1003 , n1001 , n1002 );
buf ( n1004 , n590 );
nand ( n1005 , n1003 , n1004 );
buf ( n1006 , n1005 );
buf ( n1007 , n1006 );
buf ( n1008 , n559 );
buf ( n1009 , n589 );
nand ( n1010 , n1008 , n1009 );
buf ( n1011 , n1010 );
buf ( n1012 , n1011 );
buf ( n1013 , n588 );
nand ( n1014 , n1007 , n1012 , n1013 );
buf ( n1015 , n1014 );
buf ( n1016 , n1015 );
not ( n1017 , n1016 );
buf ( n1018 , n1017 );
buf ( n1019 , n1018 );
and ( n1020 , n1000 , n1019 );
buf ( n1021 , n1020 );
buf ( n1022 , n1021 );
xor ( n1023 , n978 , n1022 );
not ( n1024 , n590 );
nor ( n1025 , n1024 , n591 );
not ( n1026 , n1025 );
not ( n1027 , n992 );
or ( n1028 , n1026 , n1027 );
and ( n1029 , n590 , n555 );
not ( n1030 , n590 );
not ( n1031 , n555 );
and ( n1032 , n1030 , n1031 );
nor ( n1033 , n1029 , n1032 );
nand ( n1034 , n1033 , n591 );
nand ( n1035 , n1028 , n1034 );
xor ( n1036 , n587 , n588 );
buf ( n1037 , n1036 );
buf ( n1038 , n559 );
and ( n1039 , n1037 , n1038 );
buf ( n1040 , n1039 );
xor ( n1041 , n1035 , n1040 );
not ( n1042 , n590 );
nand ( n1043 , n1042 , n589 );
buf ( n1044 , n1043 );
buf ( n1045 , n589 );
not ( n1046 , n1045 );
buf ( n1047 , n590 );
nand ( n1048 , n1046 , n1047 );
buf ( n1049 , n1048 );
buf ( n1050 , n1049 );
buf ( n1051 , n588 );
buf ( n1052 , n589 );
xor ( n1053 , n1051 , n1052 );
buf ( n1054 , n1053 );
buf ( n1055 , n1054 );
and ( n1056 , n1044 , n1050 , n1055 );
buf ( n1057 , n1056 );
buf ( n1058 , n1057 );
buf ( n1059 , n1058 );
buf ( n1060 , n1059 );
buf ( n1061 , n1060 );
not ( n1062 , n1061 );
buf ( n1063 , n1062 );
buf ( n1064 , n1063 );
buf ( n1065 , n558 );
buf ( n1066 , n588 );
xnor ( n1067 , n1065 , n1066 );
buf ( n1068 , n1067 );
buf ( n1069 , n1068 );
or ( n1070 , n1064 , n1069 );
xor ( n1071 , n589 , n590 );
buf ( n1072 , n1071 );
buf ( n1073 , n1072 );
buf ( n1074 , n1073 );
buf ( n1075 , n1074 );
buf ( n1076 , n557 );
buf ( n1077 , n588 );
xor ( n1078 , n1076 , n1077 );
buf ( n1079 , n1078 );
buf ( n1080 , n1079 );
nand ( n1081 , n1075 , n1080 );
buf ( n1082 , n1081 );
buf ( n1083 , n1082 );
nand ( n1084 , n1070 , n1083 );
buf ( n1085 , n1084 );
xor ( n1086 , n1041 , n1085 );
buf ( n1087 , n1086 );
and ( n1088 , n1023 , n1087 );
and ( n1089 , n978 , n1022 );
or ( n1090 , n1088 , n1089 );
buf ( n1091 , n1090 );
buf ( n1092 , n1091 );
xor ( n1093 , n935 , n1092 );
xor ( n1094 , n1035 , n1040 );
and ( n1095 , n1094 , n1085 );
and ( n1096 , n1035 , n1040 );
or ( n1097 , n1095 , n1096 );
buf ( n1098 , n1097 );
buf ( n1099 , n856 );
buf ( n1100 , n559 );
and ( n1101 , n1099 , n1100 );
buf ( n1102 , n1101 );
buf ( n1103 , n1102 );
buf ( n1104 , n948 );
not ( n1105 , n1104 );
buf ( n1106 , n574 );
not ( n1107 , n1106 );
buf ( n1108 , n575 );
nor ( n1109 , n1107 , n1108 );
buf ( n1110 , n1109 );
buf ( n1111 , n1110 );
not ( n1112 , n1111 );
or ( n1113 , n1105 , n1112 );
buf ( n1114 , n910 );
buf ( n1115 , n575 );
nand ( n1116 , n1114 , n1115 );
buf ( n1117 , n1116 );
buf ( n1118 , n1117 );
nand ( n1119 , n1113 , n1118 );
buf ( n1120 , n1119 );
buf ( n1121 , n1120 );
xor ( n1122 , n1103 , n1121 );
buf ( n1123 , n558 );
buf ( n1124 , n572 );
xor ( n1125 , n1123 , n1124 );
buf ( n1126 , n1125 );
buf ( n1127 , n1126 );
not ( n1128 , n1127 );
buf ( n1129 , n884 );
not ( n1130 , n1129 );
or ( n1131 , n1128 , n1130 );
buf ( n1132 , n888 );
buf ( n1133 , n871 );
nand ( n1134 , n1132 , n1133 );
buf ( n1135 , n1134 );
buf ( n1136 , n1135 );
nand ( n1137 , n1131 , n1136 );
buf ( n1138 , n1137 );
buf ( n1139 , n1138 );
and ( n1140 , n1122 , n1139 );
and ( n1141 , n1103 , n1121 );
or ( n1142 , n1140 , n1141 );
buf ( n1143 , n1142 );
buf ( n1144 , n1143 );
xor ( n1145 , n1098 , n1144 );
buf ( n1146 , n1079 );
not ( n1147 , n1146 );
buf ( n1148 , n1060 );
not ( n1149 , n1148 );
or ( n1150 , n1147 , n1149 );
buf ( n1151 , n1071 );
buf ( n1152 , n556 );
buf ( n1153 , n588 );
xor ( n1154 , n1152 , n1153 );
buf ( n1155 , n1154 );
buf ( n1156 , n1155 );
nand ( n1157 , n1151 , n1156 );
buf ( n1158 , n1157 );
buf ( n1159 , n1158 );
nand ( n1160 , n1150 , n1159 );
buf ( n1161 , n1160 );
buf ( n1162 , n1161 );
buf ( n1163 , n559 );
buf ( n1164 , n586 );
xor ( n1165 , n1163 , n1164 );
buf ( n1166 , n1165 );
buf ( n1167 , n1166 );
not ( n1168 , n1167 );
xor ( n1169 , n587 , n588 );
not ( n1170 , n1169 );
not ( n1171 , n586 );
not ( n1172 , n587 );
and ( n1173 , n1171 , n1172 );
and ( n1174 , n586 , n587 );
nor ( n1175 , n1173 , n1174 );
nand ( n1176 , n1170 , n1175 );
not ( n1177 , n1176 );
buf ( n1178 , n1177 );
not ( n1179 , n1178 );
or ( n1180 , n1168 , n1179 );
buf ( n1181 , n1036 );
buf ( n1182 , n558 );
buf ( n1183 , n586 );
xor ( n1184 , n1182 , n1183 );
buf ( n1185 , n1184 );
buf ( n1186 , n1185 );
nand ( n1187 , n1181 , n1186 );
buf ( n1188 , n1187 );
buf ( n1189 , n1188 );
nand ( n1190 , n1180 , n1189 );
buf ( n1191 , n1190 );
buf ( n1192 , n1191 );
xor ( n1193 , n1162 , n1192 );
buf ( n1194 , n1033 );
not ( n1195 , n1194 );
buf ( n1196 , n984 );
not ( n1197 , n1196 );
or ( n1198 , n1195 , n1197 );
and ( n1199 , n554 , n590 );
not ( n1200 , n554 );
buf ( n1201 , n590 );
not ( n1202 , n1201 );
buf ( n1203 , n1202 );
and ( n1204 , n1200 , n1203 );
nor ( n1205 , n1199 , n1204 );
buf ( n1206 , n1205 );
buf ( n1207 , n591 );
nand ( n1208 , n1206 , n1207 );
buf ( n1209 , n1208 );
buf ( n1210 , n1209 );
nand ( n1211 , n1198 , n1210 );
buf ( n1212 , n1211 );
or ( n1213 , n559 , n587 );
nand ( n1214 , n1213 , n588 );
nand ( n1215 , n559 , n587 );
and ( n1216 , n1214 , n1215 , n586 );
and ( n1217 , n1212 , n1216 );
not ( n1218 , n1212 );
not ( n1219 , n1216 );
and ( n1220 , n1218 , n1219 );
nor ( n1221 , n1217 , n1220 );
buf ( n1222 , n1221 );
xor ( n1223 , n1193 , n1222 );
buf ( n1224 , n1223 );
buf ( n1225 , n1224 );
xor ( n1226 , n1145 , n1225 );
buf ( n1227 , n1226 );
buf ( n1228 , n1227 );
xor ( n1229 , n1093 , n1228 );
buf ( n1230 , n1229 );
buf ( n1231 , n1230 );
not ( n1232 , n1231 );
xor ( n1233 , n1103 , n1121 );
xor ( n1234 , n1233 , n1139 );
buf ( n1235 , n1234 );
buf ( n1236 , n1235 );
buf ( n1237 , n559 );
buf ( n1238 , n572 );
xor ( n1239 , n1237 , n1238 );
buf ( n1240 , n1239 );
buf ( n1241 , n1240 );
not ( n1242 , n1241 );
not ( n1243 , n883 );
buf ( n1244 , n1243 );
not ( n1245 , n1244 );
or ( n1246 , n1242 , n1245 );
buf ( n1247 , n888 );
buf ( n1248 , n1126 );
nand ( n1249 , n1247 , n1248 );
buf ( n1250 , n1249 );
buf ( n1251 , n1250 );
nand ( n1252 , n1246 , n1251 );
buf ( n1253 , n1252 );
buf ( n1254 , n1253 );
buf ( n1255 , n559 );
buf ( n1256 , n588 );
xor ( n1257 , n1255 , n1256 );
buf ( n1258 , n1257 );
buf ( n1259 , n1258 );
not ( n1260 , n1259 );
buf ( n1261 , n1060 );
buf ( n1262 , n1261 );
buf ( n1263 , n1262 );
buf ( n1264 , n1263 );
not ( n1265 , n1264 );
or ( n1266 , n1260 , n1265 );
buf ( n1267 , n1068 );
not ( n1268 , n1267 );
buf ( n1269 , n1074 );
nand ( n1270 , n1268 , n1269 );
buf ( n1271 , n1270 );
buf ( n1272 , n1271 );
nand ( n1273 , n1266 , n1272 );
buf ( n1274 , n1273 );
buf ( n1275 , n1274 );
xor ( n1276 , n1254 , n1275 );
xnor ( n1277 , n1015 , n999 );
buf ( n1278 , n1277 );
and ( n1279 , n1276 , n1278 );
and ( n1280 , n1254 , n1275 );
or ( n1281 , n1279 , n1280 );
buf ( n1282 , n1281 );
buf ( n1283 , n1282 );
xor ( n1284 , n1236 , n1283 );
xor ( n1285 , n978 , n1022 );
xor ( n1286 , n1285 , n1087 );
buf ( n1287 , n1286 );
buf ( n1288 , n1287 );
and ( n1289 , n1284 , n1288 );
and ( n1290 , n1236 , n1283 );
or ( n1291 , n1289 , n1290 );
buf ( n1292 , n1291 );
buf ( n1293 , n1292 );
not ( n1294 , n1293 );
buf ( n1295 , n1294 );
buf ( n1296 , n1295 );
nand ( n1297 , n1232 , n1296 );
buf ( n1298 , n1297 );
buf ( n1299 , n1298 );
buf ( n1300 , n1230 );
buf ( n1301 , n1292 );
nand ( n1302 , n1300 , n1301 );
buf ( n1303 , n1302 );
buf ( n1304 , n1303 );
nand ( n1305 , n1299 , n1304 );
buf ( n1306 , n1305 );
xor ( n1307 , n590 , n558 );
buf ( n1308 , n1307 );
not ( n1309 , n1308 );
buf ( n1310 , n984 );
not ( n1311 , n1310 );
or ( n1312 , n1309 , n1311 );
buf ( n1313 , n979 );
buf ( n1314 , n591 );
nand ( n1315 , n1313 , n1314 );
buf ( n1316 , n1315 );
buf ( n1317 , n1316 );
nand ( n1318 , n1312 , n1317 );
buf ( n1319 , n1318 );
buf ( n1320 , n1319 );
buf ( n1321 , n888 );
buf ( n1322 , n559 );
and ( n1323 , n1321 , n1322 );
buf ( n1324 , n1323 );
buf ( n1325 , n1324 );
nand ( n1326 , n1320 , n1325 );
buf ( n1327 , n1326 );
buf ( n1328 , n1327 );
buf ( n1329 , n955 );
buf ( n1330 , n974 );
and ( n1331 , n1329 , n1330 );
not ( n1332 , n1329 );
buf ( n1333 , n971 );
and ( n1334 , n1332 , n1333 );
nor ( n1335 , n1331 , n1334 );
buf ( n1336 , n1335 );
buf ( n1337 , n1336 );
not ( n1338 , n1337 );
buf ( n1339 , n1338 );
buf ( n1340 , n1339 );
nand ( n1341 , n1328 , n1340 );
buf ( n1342 , n1341 );
buf ( n1343 , n1342 );
not ( n1344 , n1343 );
xor ( n1345 , n1254 , n1275 );
xor ( n1346 , n1345 , n1278 );
buf ( n1347 , n1346 );
buf ( n1348 , n1347 );
not ( n1349 , n1348 );
or ( n1350 , n1344 , n1349 );
buf ( n1351 , n1339 );
not ( n1352 , n1351 );
buf ( n1353 , n1327 );
not ( n1354 , n1353 );
buf ( n1355 , n1354 );
buf ( n1356 , n1355 );
nand ( n1357 , n1352 , n1356 );
buf ( n1358 , n1357 );
buf ( n1359 , n1358 );
nand ( n1360 , n1350 , n1359 );
buf ( n1361 , n1360 );
buf ( n1362 , n1361 );
xor ( n1363 , n1236 , n1283 );
xor ( n1364 , n1363 , n1288 );
buf ( n1365 , n1364 );
buf ( n1366 , n1365 );
nor ( n1367 , n1362 , n1366 );
buf ( n1368 , n1367 );
buf ( n1369 , n1368 );
not ( n1370 , n1369 );
buf ( n1371 , n1370 );
buf ( n1372 , n1371 );
not ( n1373 , n1372 );
not ( n1374 , n1347 );
buf ( n1375 , n1355 );
not ( n1376 , n1375 );
buf ( n1377 , n1339 );
not ( n1378 , n1377 );
and ( n1379 , n1376 , n1378 );
buf ( n1380 , n1355 );
buf ( n1381 , n1339 );
and ( n1382 , n1380 , n1381 );
nor ( n1383 , n1379 , n1382 );
buf ( n1384 , n1383 );
not ( n1385 , n1384 );
nand ( n1386 , n1374 , n1385 );
not ( n1387 , n1386 );
nand ( n1388 , n1347 , n1384 );
not ( n1389 , n1388 );
or ( n1390 , n1387 , n1389 );
buf ( n1391 , n558 );
buf ( n1392 , n574 );
xor ( n1393 , n1391 , n1392 );
buf ( n1394 , n1393 );
buf ( n1395 , n1394 );
not ( n1396 , n1395 );
buf ( n1397 , n905 );
not ( n1398 , n1397 );
or ( n1399 , n1396 , n1398 );
buf ( n1400 , n575 );
buf ( n1401 , n941 );
nand ( n1402 , n1400 , n1401 );
buf ( n1403 , n1402 );
buf ( n1404 , n1403 );
nand ( n1405 , n1399 , n1404 );
buf ( n1406 , n1405 );
buf ( n1407 , n1406 );
buf ( n1408 , n1407 );
buf ( n1409 , n1074 );
buf ( n1410 , n559 );
and ( n1411 , n1409 , n1410 );
buf ( n1412 , n1411 );
buf ( n1413 , n1412 );
buf ( n1414 , n1413 );
buf ( n1415 , n1414 );
buf ( n1416 , n1415 );
or ( n1417 , n1408 , n1416 );
buf ( n1418 , n1417 );
buf ( n1419 , n1418 );
not ( n1420 , n1419 );
buf ( n1421 , n1324 );
buf ( n1422 , n1319 );
xnor ( n1423 , n1421 , n1422 );
buf ( n1424 , n1423 );
buf ( n1425 , n1424 );
not ( n1426 , n1425 );
buf ( n1427 , n1426 );
buf ( n1428 , n1427 );
not ( n1429 , n1428 );
or ( n1430 , n1420 , n1429 );
buf ( n1431 , n1415 );
buf ( n1432 , n1407 );
nand ( n1433 , n1431 , n1432 );
buf ( n1434 , n1433 );
buf ( n1435 , n1434 );
nand ( n1436 , n1430 , n1435 );
buf ( n1437 , n1436 );
nand ( n1438 , n1390 , n1437 );
buf ( n1439 , n1438 );
not ( n1440 , n1439 );
buf ( n1441 , n1440 );
not ( n1442 , n1441 );
xor ( n1443 , n1406 , n1412 );
buf ( n1444 , n1443 );
not ( n1445 , n1444 );
buf ( n1446 , n1445 );
buf ( n1447 , n1446 );
not ( n1448 , n1447 );
buf ( n1449 , n1427 );
not ( n1450 , n1449 );
or ( n1451 , n1448 , n1450 );
buf ( n1452 , n1443 );
buf ( n1453 , n1424 );
nand ( n1454 , n1452 , n1453 );
buf ( n1455 , n1454 );
buf ( n1456 , n1455 );
nand ( n1457 , n1451 , n1456 );
buf ( n1458 , n1457 );
buf ( n1459 , n1458 );
buf ( n1460 , n559 );
buf ( n1461 , n591 );
nand ( n1462 , n1460 , n1461 );
buf ( n1463 , n1462 );
buf ( n1464 , n1463 );
buf ( n1465 , n590 );
and ( n1466 , n1464 , n1465 );
buf ( n1467 , n1466 );
buf ( n1468 , n1467 );
buf ( n1469 , n1468 );
buf ( n1470 , n1469 );
buf ( n1471 , n1470 );
buf ( n1472 , n559 );
buf ( n1473 , n575 );
nand ( n1474 , n1472 , n1473 );
buf ( n1475 , n1474 );
buf ( n1476 , n1475 );
buf ( n1477 , n574 );
and ( n1478 , n1476 , n1477 );
buf ( n1479 , n1478 );
buf ( n1480 , n1479 );
buf ( n1481 , n1480 );
buf ( n1482 , n1481 );
buf ( n1483 , n1482 );
or ( n1484 , n1471 , n1483 );
buf ( n1485 , n1484 );
buf ( n1486 , n1485 );
not ( n1487 , n1486 );
buf ( n1488 , n559 );
not ( n1489 , n1488 );
buf ( n1490 , n1489 );
buf ( n1491 , n1490 );
not ( n1492 , n1491 );
buf ( n1493 , n984 );
not ( n1494 , n1493 );
or ( n1495 , n1492 , n1494 );
buf ( n1496 , n591 );
buf ( n1497 , n1307 );
nand ( n1498 , n1496 , n1497 );
buf ( n1499 , n1498 );
buf ( n1500 , n1499 );
nand ( n1501 , n1495 , n1500 );
buf ( n1502 , n1501 );
buf ( n1503 , n1502 );
not ( n1504 , n1503 );
or ( n1505 , n1487 , n1504 );
buf ( n1506 , n1482 );
buf ( n1507 , n1470 );
nand ( n1508 , n1506 , n1507 );
buf ( n1509 , n1508 );
buf ( n1510 , n1509 );
nand ( n1511 , n1505 , n1510 );
buf ( n1512 , n1511 );
buf ( n1513 , n1512 );
nand ( n1514 , n1459 , n1513 );
buf ( n1515 , n1514 );
not ( n1516 , n1515 );
buf ( n1517 , n1458 );
not ( n1518 , n1517 );
buf ( n1519 , n1518 );
buf ( n1520 , n1519 );
buf ( n1521 , n1512 );
not ( n1522 , n1521 );
buf ( n1523 , n1522 );
buf ( n1524 , n1523 );
nand ( n1525 , n1520 , n1524 );
buf ( n1526 , n1525 );
buf ( n1527 , n1526 );
buf ( n1528 , n559 );
buf ( n1529 , n575 );
and ( n1530 , n1528 , n1529 );
buf ( n1531 , n1530 );
buf ( n1532 , n1531 );
not ( n1533 , n1532 );
buf ( n1534 , n1533 );
buf ( n1535 , n1534 );
buf ( n1536 , n559 );
buf ( n1537 , n591 );
and ( n1538 , n1536 , n1537 );
buf ( n1539 , n1538 );
buf ( n1540 , n1539 );
not ( n1541 , n1540 );
buf ( n1542 , n1541 );
buf ( n1543 , n1542 );
nor ( n1544 , n1535 , n1543 );
buf ( n1545 , n1544 );
buf ( n1546 , n1545 );
buf ( n1547 , n1490 );
not ( n1548 , n1547 );
buf ( n1549 , n905 );
not ( n1550 , n1549 );
or ( n1551 , n1548 , n1550 );
buf ( n1552 , n1394 );
buf ( n1553 , n575 );
nand ( n1554 , n1552 , n1553 );
buf ( n1555 , n1554 );
buf ( n1556 , n1555 );
nand ( n1557 , n1551 , n1556 );
buf ( n1558 , n1557 );
buf ( n1559 , n1558 );
xor ( n1560 , n1546 , n1559 );
buf ( n1561 , n1467 );
buf ( n1562 , n1479 );
xnor ( n1563 , n1561 , n1562 );
buf ( n1564 , n1563 );
xnor ( n1565 , n1502 , n1564 );
buf ( n1566 , n1565 );
and ( n1567 , n1560 , n1566 );
and ( n1568 , n1546 , n1559 );
or ( n1569 , n1567 , n1568 );
buf ( n1570 , n1569 );
buf ( n1571 , n1570 );
nand ( n1572 , n1527 , n1571 );
buf ( n1573 , n1572 );
not ( n1574 , n1573 );
or ( n1575 , n1516 , n1574 );
not ( n1576 , n1437 );
nand ( n1577 , n1347 , n1576 , n1385 );
not ( n1578 , n1577 );
and ( n1579 , n1374 , n1576 , n1384 );
nor ( n1580 , n1578 , n1579 );
nand ( n1581 , n1575 , n1580 );
nand ( n1582 , n1442 , n1581 );
buf ( n1583 , n1582 );
not ( n1584 , n1583 );
or ( n1585 , n1373 , n1584 );
buf ( n1586 , n1365 );
buf ( n1587 , n1361 );
nand ( n1588 , n1586 , n1587 );
buf ( n1589 , n1588 );
buf ( n1590 , n1589 );
nand ( n1591 , n1585 , n1590 );
buf ( n1592 , n1591 );
xor ( n1593 , n1306 , n1592 );
xor ( n1594 , n557 , n558 );
not ( n1595 , n1594 );
not ( n1596 , n1595 );
not ( n1597 , n1596 );
not ( n1598 , n556 );
not ( n1599 , n573 );
not ( n1600 , n589 );
or ( n1601 , n1599 , n1600 );
nor ( n1602 , n574 , n590 );
nor ( n1603 , n573 , n589 );
nor ( n1604 , n1602 , n1603 );
nand ( n1605 , n574 , n590 );
nand ( n1606 , n575 , n591 );
nand ( n1607 , n1605 , n1606 );
nand ( n1608 , n1604 , n1607 );
nand ( n1609 , n1601 , n1608 );
nand ( n1610 , n572 , n588 );
not ( n1611 , n1610 );
nor ( n1612 , n572 , n588 );
nor ( n1613 , n1611 , n1612 );
and ( n1614 , n1609 , n1613 );
not ( n1615 , n1609 );
not ( n1616 , n588 );
nand ( n1617 , n874 , n1616 );
nand ( n1618 , n1617 , n1610 );
and ( n1619 , n1615 , n1618 );
nor ( n1620 , n1614 , n1619 );
not ( n1621 , n1620 );
not ( n1622 , n1621 );
or ( n1623 , n1598 , n1622 );
buf ( n1624 , n1620 );
not ( n1625 , n556 );
nand ( n1626 , n1624 , n1625 );
nand ( n1627 , n1623 , n1626 );
not ( n1628 , n1627 );
or ( n1629 , n1597 , n1628 );
not ( n1630 , n556 );
nand ( n1631 , n575 , n591 );
not ( n1632 , n1631 );
not ( n1633 , n1632 );
not ( n1634 , n574 );
not ( n1635 , n590 );
nand ( n1636 , n1634 , n1635 );
not ( n1637 , n1636 );
or ( n1638 , n1633 , n1637 );
nand ( n1639 , n574 , n590 );
nand ( n1640 , n1638 , n1639 );
and ( n1641 , n573 , n589 );
not ( n1642 , n573 );
not ( n1643 , n589 );
and ( n1644 , n1642 , n1643 );
nor ( n1645 , n1641 , n1644 );
not ( n1646 , n1645 );
and ( n1647 , n1640 , n1646 );
not ( n1648 , n1640 );
and ( n1649 , n1648 , n1645 );
nor ( n1650 , n1647 , n1649 );
not ( n1651 , n1650 );
not ( n1652 , n1651 );
not ( n1653 , n1652 );
or ( n1654 , n1630 , n1653 );
nand ( n1655 , n1625 , n1651 );
nand ( n1656 , n1654 , n1655 );
xor ( n1657 , n556 , n557 );
nand ( n1658 , n1595 , n1657 );
not ( n1659 , n1658 );
nand ( n1660 , n1656 , n1659 );
nand ( n1661 , n1629 , n1660 );
or ( n1662 , n555 , n556 );
xor ( n1663 , n591 , n575 );
buf ( n1664 , n1663 );
nand ( n1665 , n1662 , n1664 );
nand ( n1666 , n555 , n556 );
and ( n1667 , n1665 , n1666 , n554 );
xor ( n1668 , n556 , n555 );
not ( n1669 , n1668 );
not ( n1670 , n554 );
xor ( n1671 , n574 , n590 );
nand ( n1672 , n575 , n591 );
and ( n1673 , n1671 , n1672 );
not ( n1674 , n1671 );
and ( n1675 , n575 , n591 );
and ( n1676 , n1674 , n1675 );
nor ( n1677 , n1673 , n1676 );
not ( n1678 , n1677 );
or ( n1679 , n1670 , n1678 );
not ( n1680 , n1677 );
not ( n1681 , n554 );
nand ( n1682 , n1680 , n1681 );
nand ( n1683 , n1679 , n1682 );
not ( n1684 , n1683 );
or ( n1685 , n1669 , n1684 );
not ( n1686 , n554 );
not ( n1687 , n1664 );
not ( n1688 , n1687 );
or ( n1689 , n1686 , n1688 );
nand ( n1690 , n1664 , n1681 );
nand ( n1691 , n1689 , n1690 );
xor ( n1692 , n554 , n555 );
not ( n1693 , n1692 );
nor ( n1694 , n1693 , n1668 );
nand ( n1695 , n1691 , n1694 );
nand ( n1696 , n1685 , n1695 );
xor ( n1697 , n1667 , n1696 );
xor ( n1698 , n1661 , n1697 );
not ( n1699 , n558 );
not ( n1700 , n573 );
not ( n1701 , n589 );
and ( n1702 , n1700 , n1701 );
nor ( n1703 , n1702 , n1612 );
not ( n1704 , n1703 );
not ( n1705 , n574 );
not ( n1706 , n590 );
or ( n1707 , n1705 , n1706 );
nor ( n1708 , n574 , n590 );
nand ( n1709 , n575 , n591 );
or ( n1710 , n1708 , n1709 );
nand ( n1711 , n1707 , n1710 );
not ( n1712 , n1711 );
or ( n1713 , n1704 , n1712 );
nor ( n1714 , n572 , n588 );
nand ( n1715 , n573 , n589 );
or ( n1716 , n1714 , n1715 );
nand ( n1717 , n572 , n588 );
nand ( n1718 , n1716 , n1717 );
not ( n1719 , n1718 );
nand ( n1720 , n1713 , n1719 );
not ( n1721 , n571 );
not ( n1722 , n587 );
and ( n1723 , n1721 , n1722 );
nand ( n1724 , n587 , n571 );
not ( n1725 , n1724 );
nor ( n1726 , n1723 , n1725 );
and ( n1727 , n1720 , n1726 );
not ( n1728 , n1720 );
not ( n1729 , n1726 );
and ( n1730 , n1728 , n1729 );
nor ( n1731 , n1727 , n1730 );
buf ( n1732 , n1731 );
not ( n1733 , n1732 );
not ( n1734 , n1733 );
or ( n1735 , n1699 , n1734 );
not ( n1736 , n558 );
nand ( n1737 , n1732 , n1736 );
nand ( n1738 , n1735 , n1737 );
nor ( n1739 , n1736 , n559 );
buf ( n1740 , n1739 );
nand ( n1741 , n1738 , n1740 );
not ( n1742 , n558 );
nand ( n1743 , n1742 , n559 );
not ( n1744 , n1743 );
or ( n1745 , n587 , n571 );
not ( n1746 , n1745 );
not ( n1747 , n1703 );
nor ( n1748 , n574 , n590 );
nand ( n1749 , n575 , n591 );
or ( n1750 , n1748 , n1749 );
nand ( n1751 , n1750 , n1639 );
not ( n1752 , n1751 );
or ( n1753 , n1747 , n1752 );
nand ( n1754 , n1753 , n1719 );
not ( n1755 , n1754 );
or ( n1756 , n1746 , n1755 );
nand ( n1757 , n1756 , n1724 );
nand ( n1758 , n570 , n586 );
not ( n1759 , n1758 );
nor ( n1760 , n570 , n586 );
nor ( n1761 , n1759 , n1760 );
and ( n1762 , n1757 , n1761 );
not ( n1763 , n1757 );
not ( n1764 , n570 );
not ( n1765 , n1764 );
not ( n1766 , n586 );
not ( n1767 , n1766 );
or ( n1768 , n1765 , n1767 );
nand ( n1769 , n1768 , n1758 );
and ( n1770 , n1763 , n1769 );
nor ( n1771 , n1762 , n1770 );
buf ( n1772 , n1771 );
nand ( n1773 , n1744 , n1772 );
nand ( n1774 , n558 , n559 );
not ( n1775 , n1774 );
not ( n1776 , n1772 );
nand ( n1777 , n1775 , n1776 );
nand ( n1778 , n1741 , n1773 , n1777 );
xor ( n1779 , n1698 , n1778 );
and ( n1780 , n1664 , n1668 );
not ( n1781 , n1594 );
not ( n1782 , n1656 );
or ( n1783 , n1781 , n1782 );
and ( n1784 , n556 , n1677 );
not ( n1785 , n556 );
nand ( n1786 , n575 , n591 );
and ( n1787 , n1671 , n1786 );
not ( n1788 , n1671 );
and ( n1789 , n1788 , n1675 );
nor ( n1790 , n1787 , n1789 );
not ( n1791 , n1790 );
and ( n1792 , n1785 , n1791 );
or ( n1793 , n1784 , n1792 );
nand ( n1794 , n1793 , n1659 );
nand ( n1795 , n1783 , n1794 );
xor ( n1796 , n1780 , n1795 );
or ( n1797 , n557 , n558 );
xor ( n1798 , n591 , n575 );
nand ( n1799 , n1797 , n1798 );
nand ( n1800 , n557 , n558 );
and ( n1801 , n1799 , n1800 , n556 );
not ( n1802 , n1594 );
not ( n1803 , n1793 );
or ( n1804 , n1802 , n1803 );
and ( n1805 , n556 , n1664 );
not ( n1806 , n556 );
not ( n1807 , n1798 );
and ( n1808 , n1806 , n1807 );
nor ( n1809 , n1805 , n1808 );
and ( n1810 , n1595 , n1657 );
nand ( n1811 , n1809 , n1810 );
nand ( n1812 , n1804 , n1811 );
and ( n1813 , n1801 , n1812 );
and ( n1814 , n1796 , n1813 );
and ( n1815 , n1780 , n1795 );
or ( n1816 , n1814 , n1815 );
not ( n1817 , n1816 );
and ( n1818 , n1779 , n1817 );
not ( n1819 , n1779 );
and ( n1820 , n1819 , n1816 );
nor ( n1821 , n1818 , n1820 );
xor ( n1822 , n1780 , n1795 );
xor ( n1823 , n1822 , n1813 );
not ( n1824 , n559 );
not ( n1825 , n1738 );
or ( n1826 , n1824 , n1825 );
and ( n1827 , n558 , n1624 );
not ( n1828 , n558 );
and ( n1829 , n1828 , n1621 );
nor ( n1830 , n1827 , n1829 );
nand ( n1831 , n1830 , n1739 );
nand ( n1832 , n1826 , n1831 );
nor ( n1833 , n1823 , n1832 );
not ( n1834 , n559 );
not ( n1835 , n1830 );
or ( n1836 , n1834 , n1835 );
not ( n1837 , n1650 );
not ( n1838 , n1837 );
nand ( n1839 , n1838 , n558 );
not ( n1840 , n1839 );
not ( n1841 , n558 );
nand ( n1842 , n1841 , n1651 );
not ( n1843 , n1842 );
or ( n1844 , n1840 , n1843 );
nand ( n1845 , n1844 , n1740 );
nand ( n1846 , n1836 , n1845 );
xor ( n1847 , n1801 , n1812 );
xor ( n1848 , n1846 , n1847 );
not ( n1849 , n559 );
nand ( n1850 , n1839 , n1842 );
not ( n1851 , n1850 );
or ( n1852 , n1849 , n1851 );
not ( n1853 , n558 );
not ( n1854 , n1790 );
not ( n1855 , n1854 );
not ( n1856 , n1855 );
or ( n1857 , n1853 , n1856 );
not ( n1858 , n558 );
nand ( n1859 , n1858 , n1680 );
nand ( n1860 , n1857 , n1859 );
nand ( n1861 , n1860 , n1740 );
nand ( n1862 , n1852 , n1861 );
not ( n1863 , n1862 );
and ( n1864 , n1664 , n1594 );
not ( n1865 , n1864 );
or ( n1866 , n1863 , n1865 );
nor ( n1867 , n1862 , n1864 );
not ( n1868 , n559 );
not ( n1869 , n1860 );
or ( n1870 , n1868 , n1869 );
nand ( n1871 , n1687 , n1740 );
nand ( n1872 , n1870 , n1871 );
not ( n1873 , n559 );
not ( n1874 , n1664 );
or ( n1875 , n1873 , n1874 );
nand ( n1876 , n1875 , n558 );
not ( n1877 , n1876 );
nand ( n1878 , n1872 , n1877 );
or ( n1879 , n1867 , n1878 );
nand ( n1880 , n1866 , n1879 );
and ( n1881 , n1848 , n1880 );
and ( n1882 , n1846 , n1847 );
or ( n1883 , n1881 , n1882 );
not ( n1884 , n1883 );
or ( n1885 , n1833 , n1884 );
nand ( n1886 , n1823 , n1832 );
nand ( n1887 , n1885 , n1886 );
buf ( n1888 , n1887 );
not ( n1889 , n1888 );
and ( n1890 , n1821 , n1889 );
not ( n1891 , n1821 );
and ( n1892 , n1891 , n1888 );
nor ( n1893 , n1890 , n1892 );
nand ( n1894 , n1593 , n1893 );
buf ( n1895 , n1580 );
buf ( n1896 , n1438 );
nand ( n1897 , n1895 , n1896 );
buf ( n1898 , n1897 );
buf ( n1899 , n1898 );
buf ( n1900 , n1573 );
buf ( n1901 , n1515 );
nand ( n1902 , n1900 , n1901 );
buf ( n1903 , n1902 );
buf ( n1904 , n1903 );
not ( n1905 , n1904 );
buf ( n1906 , n1905 );
buf ( n1907 , n1906 );
and ( n1908 , n1899 , n1907 );
not ( n1909 , n1899 );
buf ( n1910 , n1903 );
and ( n1911 , n1909 , n1910 );
nor ( n1912 , n1908 , n1911 );
buf ( n1913 , n1912 );
xor ( n1914 , n1846 , n1847 );
xor ( n1915 , n1914 , n1880 );
not ( n1916 , n1915 );
nand ( n1917 , n1916 , n1913 );
buf ( n1918 , n1582 );
not ( n1919 , n1918 );
buf ( n1920 , n1919 );
buf ( n1921 , n1920 );
buf ( n1922 , n1365 );
buf ( n1923 , n1361 );
nor ( n1924 , n1922 , n1923 );
buf ( n1925 , n1924 );
buf ( n1926 , n1925 );
not ( n1927 , n1926 );
buf ( n1928 , n1927 );
buf ( n1929 , n1928 );
buf ( n1930 , n1589 );
nand ( n1931 , n1929 , n1930 );
buf ( n1932 , n1931 );
buf ( n1933 , n1932 );
and ( n1934 , n1921 , n1933 );
not ( n1935 , n1921 );
buf ( n1936 , n1932 );
not ( n1937 , n1936 );
buf ( n1938 , n1937 );
buf ( n1939 , n1938 );
and ( n1940 , n1935 , n1939 );
nor ( n1941 , n1934 , n1940 );
buf ( n1942 , n1941 );
not ( n1943 , n1942 );
not ( n1944 , n1833 );
nand ( n1945 , n1944 , n1886 );
and ( n1946 , n1945 , n1884 );
not ( n1947 , n1945 );
and ( n1948 , n1947 , n1883 );
nor ( n1949 , n1946 , n1948 );
nand ( n1950 , n1943 , n1949 );
and ( n1951 , n1894 , C1 , n1950 );
not ( n1952 , n1949 );
nand ( n1953 , n1952 , n1942 );
not ( n1954 , n1953 );
not ( n1955 , n1954 );
not ( n1956 , n1894 );
or ( n1957 , n1955 , n1956 );
not ( n1958 , n1593 );
not ( n1959 , n1893 );
nand ( n1960 , n1958 , n1959 );
nand ( n1961 , n1957 , n1960 );
nor ( n1962 , n1951 , n1961 );
not ( n1963 , n1962 );
xor ( n1964 , n1098 , n1144 );
and ( n1965 , n1964 , n1225 );
and ( n1966 , n1098 , n1144 );
or ( n1967 , n1965 , n1966 );
buf ( n1968 , n1967 );
buf ( n1969 , n861 );
not ( n1970 , n1969 );
buf ( n1971 , n847 );
not ( n1972 , n1971 );
buf ( n1973 , n1972 );
buf ( n1974 , n1973 );
not ( n1975 , n1974 );
or ( n1976 , n1970 , n1975 );
buf ( n1977 , n842 );
not ( n1978 , n1977 );
buf ( n1979 , n1978 );
buf ( n1980 , n1979 );
buf ( n1981 , n1980 );
buf ( n1982 , n1981 );
buf ( n1983 , n1982 );
buf ( n1984 , n557 );
buf ( n1985 , n570 );
xor ( n1986 , n1984 , n1985 );
buf ( n1987 , n1986 );
buf ( n1988 , n1987 );
nand ( n1989 , n1983 , n1988 );
buf ( n1990 , n1989 );
buf ( n1991 , n1990 );
nand ( n1992 , n1976 , n1991 );
buf ( n1993 , n1992 );
buf ( n1994 , n1993 );
buf ( n1995 , n921 );
buf ( n1996 , n929 );
and ( n1997 , n1995 , n1996 );
buf ( n1998 , n1997 );
buf ( n1999 , n1998 );
xor ( n2000 , n1994 , n1999 );
xor ( n2001 , n569 , n570 );
buf ( n2002 , n2001 );
buf ( n2003 , n559 );
and ( n2004 , n2002 , n2003 );
buf ( n2005 , n2004 );
not ( n2006 , n905 );
not ( n2007 , n916 );
or ( n2008 , n2006 , n2007 );
buf ( n2009 , n553 );
buf ( n2010 , n574 );
xor ( n2011 , n2009 , n2010 );
buf ( n2012 , n2011 );
buf ( n2013 , n2012 );
buf ( n2014 , n575 );
nand ( n2015 , n2013 , n2014 );
buf ( n2016 , n2015 );
nand ( n2017 , n2008 , n2016 );
xor ( n2018 , n2005 , n2017 );
buf ( n2019 , n893 );
not ( n2020 , n2019 );
buf ( n2021 , n884 );
not ( n2022 , n2021 );
or ( n2023 , n2020 , n2022 );
buf ( n2024 , n888 );
buf ( n2025 , n555 );
buf ( n2026 , n572 );
xor ( n2027 , n2025 , n2026 );
buf ( n2028 , n2027 );
buf ( n2029 , n2028 );
nand ( n2030 , n2024 , n2029 );
buf ( n2031 , n2030 );
buf ( n2032 , n2031 );
nand ( n2033 , n2023 , n2032 );
buf ( n2034 , n2033 );
xor ( n2035 , n2018 , n2034 );
buf ( n2036 , n2035 );
xor ( n2037 , n2000 , n2036 );
buf ( n2038 , n2037 );
not ( n2039 , n2038 );
and ( n2040 , n1968 , n2039 );
not ( n2041 , n1968 );
and ( n2042 , n2041 , n2038 );
nor ( n2043 , n2040 , n2042 );
buf ( n2044 , n899 );
not ( n2045 , n2044 );
buf ( n2046 , n933 );
not ( n2047 , n2046 );
or ( n2048 , n2045 , n2047 );
buf ( n2049 , n899 );
buf ( n2050 , n933 );
or ( n2051 , n2049 , n2050 );
buf ( n2052 , n867 );
nand ( n2053 , n2051 , n2052 );
buf ( n2054 , n2053 );
buf ( n2055 , n2054 );
nand ( n2056 , n2048 , n2055 );
buf ( n2057 , n2056 );
xor ( n2058 , n1162 , n1192 );
and ( n2059 , n2058 , n1222 );
and ( n2060 , n1162 , n1192 );
or ( n2061 , n2059 , n2060 );
buf ( n2062 , n2061 );
not ( n2063 , n2062 );
xor ( n2064 , n2057 , n2063 );
buf ( n2065 , n1185 );
not ( n2066 , n2065 );
buf ( n2067 , n1177 );
not ( n2068 , n2067 );
or ( n2069 , n2066 , n2068 );
buf ( n2070 , n1036 );
buf ( n2071 , n557 );
buf ( n2072 , n586 );
xor ( n2073 , n2071 , n2072 );
buf ( n2074 , n2073 );
buf ( n2075 , n2074 );
nand ( n2076 , n2070 , n2075 );
buf ( n2077 , n2076 );
buf ( n2078 , n2077 );
nand ( n2079 , n2069 , n2078 );
buf ( n2080 , n2079 );
buf ( n2081 , n2080 );
not ( n2082 , n2081 );
buf ( n2083 , n2082 );
buf ( n2084 , n1212 );
buf ( n2085 , n1216 );
and ( n2086 , n2084 , n2085 );
buf ( n2087 , n2086 );
not ( n2088 , n2087 );
xor ( n2089 , n2083 , n2088 );
buf ( n2090 , n2089 );
not ( n2091 , n2090 );
buf ( n2092 , n2091 );
not ( n2093 , n2092 );
buf ( n2094 , n1205 );
not ( n2095 , n2094 );
buf ( n2096 , n984 );
not ( n2097 , n2096 );
or ( n2098 , n2095 , n2097 );
and ( n2099 , n553 , n590 );
not ( n2100 , n553 );
buf ( n2101 , n590 );
not ( n2102 , n2101 );
buf ( n2103 , n2102 );
and ( n2104 , n2100 , n2103 );
nor ( n2105 , n2099 , n2104 );
nand ( n2106 , n2105 , n591 );
buf ( n2107 , n2106 );
nand ( n2108 , n2098 , n2107 );
buf ( n2109 , n2108 );
buf ( n2110 , n2109 );
not ( n2111 , n2110 );
buf ( n2112 , n1490 );
not ( n2113 , n2112 );
buf ( n2114 , n585 );
buf ( n2115 , n586 );
xor ( n2116 , n2114 , n2115 );
buf ( n2117 , n2116 );
buf ( n2118 , n2117 );
not ( n2119 , n2118 );
buf ( n2120 , n2119 );
buf ( n2121 , n2120 );
not ( n2122 , n2121 );
buf ( n2123 , n2122 );
buf ( n2124 , n2123 );
nand ( n2125 , n2113 , n2124 );
buf ( n2126 , n2125 );
buf ( n2127 , n2126 );
not ( n2128 , n2127 );
and ( n2129 , n2111 , n2128 );
buf ( n2130 , n2120 );
buf ( n2131 , n2130 );
buf ( n2132 , n2131 );
buf ( n2133 , n2132 );
not ( n2134 , n2133 );
buf ( n2135 , n2134 );
buf ( n2136 , n2135 );
buf ( n2137 , n559 );
nand ( n2138 , n2136 , n2137 );
buf ( n2139 , n2138 );
buf ( n2140 , n2139 );
buf ( n2141 , n2109 );
and ( n2142 , n2140 , n2141 );
nor ( n2143 , n2129 , n2142 );
buf ( n2144 , n2143 );
buf ( n2145 , n2144 );
buf ( n2146 , n1155 );
not ( n2147 , n2146 );
buf ( n2148 , n1060 );
not ( n2149 , n2148 );
or ( n2150 , n2147 , n2149 );
buf ( n2151 , n1074 );
buf ( n2152 , n555 );
buf ( n2153 , n588 );
xor ( n2154 , n2152 , n2153 );
buf ( n2155 , n2154 );
buf ( n2156 , n2155 );
nand ( n2157 , n2151 , n2156 );
buf ( n2158 , n2157 );
buf ( n2159 , n2158 );
nand ( n2160 , n2150 , n2159 );
buf ( n2161 , n2160 );
buf ( n2162 , n2161 );
xor ( n2163 , n2145 , n2162 );
buf ( n2164 , n2163 );
buf ( n2165 , n2164 );
not ( n2166 , n2165 );
buf ( n2167 , n2166 );
not ( n2168 , n2167 );
or ( n2169 , n2093 , n2168 );
buf ( n2170 , n2164 );
buf ( n2171 , n2089 );
nand ( n2172 , n2170 , n2171 );
buf ( n2173 , n2172 );
nand ( n2174 , n2169 , n2173 );
xnor ( n2175 , n2064 , n2174 );
not ( n2176 , n2175 );
and ( n2177 , n2043 , n2176 );
not ( n2178 , n2043 );
and ( n2179 , n2178 , n2175 );
nor ( n2180 , n2177 , n2179 );
buf ( n2181 , n2180 );
xor ( n2182 , n935 , n1092 );
and ( n2183 , n2182 , n1228 );
and ( n2184 , n935 , n1092 );
or ( n2185 , n2183 , n2184 );
buf ( n2186 , n2185 );
buf ( n2187 , n2186 );
nand ( n2188 , n2181 , n2187 );
buf ( n2189 , n2188 );
buf ( n2190 , n2189 );
buf ( n2191 , n2190 );
buf ( n2192 , n2191 );
not ( n2193 , n2180 );
buf ( n2194 , n2186 );
not ( n2195 , n2194 );
buf ( n2196 , n2195 );
nand ( n2197 , n2193 , n2196 );
nand ( n2198 , n2192 , n2197 );
not ( n2199 , n2198 );
buf ( n2200 , n1230 );
buf ( n2201 , n1292 );
nor ( n2202 , n2200 , n2201 );
buf ( n2203 , n2202 );
or ( n2204 , n2203 , n1589 );
nand ( n2205 , n2204 , n1303 );
not ( n2206 , n2205 );
buf ( n2207 , n1925 );
not ( n2208 , n2207 );
buf ( n2209 , n1298 );
buf ( n2210 , n1582 );
nand ( n2211 , n2208 , n2209 , n2210 );
buf ( n2212 , n2211 );
nand ( n2213 , n2206 , n2212 );
not ( n2214 , n2213 );
or ( n2215 , n2199 , n2214 );
nand ( n2216 , n2206 , n2212 , n2192 , n2197 );
nand ( n2217 , n2215 , n2216 );
not ( n2218 , n1596 );
not ( n2219 , n556 );
not ( n2220 , n1732 );
not ( n2221 , n2220 );
or ( n2222 , n2219 , n2221 );
nand ( n2223 , n1732 , n1625 );
nand ( n2224 , n2222 , n2223 );
not ( n2225 , n2224 );
or ( n2226 , n2218 , n2225 );
nand ( n2227 , n1627 , n1659 );
nand ( n2228 , n2226 , n2227 );
not ( n2229 , n558 );
or ( n2230 , n571 , n587 );
or ( n2231 , n570 , n586 );
nand ( n2232 , n2230 , n2231 );
not ( n2233 , n2232 );
not ( n2234 , n2233 );
not ( n2235 , n1754 );
or ( n2236 , n2234 , n2235 );
nand ( n2237 , n571 , n587 );
or ( n2238 , n1760 , n2237 );
nand ( n2239 , n2238 , n1758 );
not ( n2240 , n2239 );
nand ( n2241 , n2236 , n2240 );
nor ( n2242 , n569 , n585 );
not ( n2243 , n2242 );
nand ( n2244 , n569 , n585 );
nand ( n2245 , n2243 , n2244 );
not ( n2246 , n2245 );
and ( n2247 , n2241 , n2246 );
not ( n2248 , n2241 );
and ( n2249 , n2248 , n2245 );
nor ( n2250 , n2247 , n2249 );
buf ( n2251 , n2250 );
not ( n2252 , n2251 );
not ( n2253 , n2252 );
or ( n2254 , n2229 , n2253 );
not ( n2255 , n558 );
nand ( n2256 , n2255 , n2251 );
nand ( n2257 , n2254 , n2256 );
not ( n2258 , n2257 );
not ( n2259 , n559 );
or ( n2260 , n2258 , n2259 );
not ( n2261 , n1772 );
nand ( n2262 , n2261 , n1740 );
nand ( n2263 , n2260 , n2262 );
xor ( n2264 , n2228 , n2263 );
xor ( n2265 , n553 , n554 );
and ( n2266 , n1664 , n2265 );
not ( n2267 , n1668 );
not ( n2268 , n1651 );
not ( n2269 , n1681 );
or ( n2270 , n2268 , n2269 );
nand ( n2271 , n1838 , n554 );
nand ( n2272 , n2270 , n2271 );
not ( n2273 , n2272 );
or ( n2274 , n2267 , n2273 );
xnor ( n2275 , n555 , n556 );
and ( n2276 , n2275 , n1692 );
nand ( n2277 , n1683 , n2276 );
nand ( n2278 , n2274 , n2277 );
xor ( n2279 , n2266 , n2278 );
and ( n2280 , n1667 , n1696 );
xor ( n2281 , n2279 , n2280 );
xor ( n2282 , n2264 , n2281 );
not ( n2283 , n2282 );
not ( n2284 , n2283 );
xor ( n2285 , n1661 , n1697 );
and ( n2286 , n2285 , n1778 );
and ( n2287 , n1661 , n1697 );
or ( n2288 , n2286 , n2287 );
and ( n2289 , n2284 , n2288 );
not ( n2290 , n2284 );
not ( n2291 , n2288 );
and ( n2292 , n2290 , n2291 );
nor ( n2293 , n2289 , n2292 );
not ( n2294 , n1887 );
not ( n2295 , n1779 );
nand ( n2296 , n2295 , n1817 );
not ( n2297 , n2296 );
or ( n2298 , n2294 , n2297 );
nand ( n2299 , n1779 , n1816 );
nand ( n2300 , n2298 , n2299 );
buf ( n2301 , n2300 );
xor ( n2302 , n2293 , n2301 );
not ( n2303 , n2302 );
nor ( n2304 , n2217 , n2303 );
not ( n2305 , n2304 );
not ( n2306 , n2302 );
nand ( n2307 , n2306 , n2217 );
nand ( n2308 , n2305 , n2307 );
not ( n2309 , n2308 );
not ( n2310 , n2309 );
or ( n2311 , n1963 , n2310 );
not ( n2312 , n1962 );
nand ( n2313 , n2312 , n2308 );
nand ( n2314 , n2311 , n2313 );
nand ( n2315 , n2314 , n585 );
not ( n2316 , n2314 );
not ( n2317 , n585 );
nand ( n2318 , n2316 , n2317 );
nand ( n2319 , n2315 , n2318 );
nand ( n2320 , C1 , n1917 );
not ( n2321 , n2320 );
and ( n2322 , n2321 , C1 );
nor ( n2323 , C0 , n2322 );
not ( n2324 , n2323 );
not ( n2325 , n588 );
nand ( n2326 , n2324 , n2325 );
nand ( n2327 , n1960 , n1894 );
not ( n2328 , n2327 );
not ( n2329 , n2328 );
not ( n2330 , n1950 );
or ( n2331 , C0 , n2330 );
nand ( n2332 , n2331 , n1953 );
not ( n2333 , n2332 );
not ( n2334 , n2333 );
or ( n2335 , n2329 , n2334 );
nand ( n2336 , n2332 , n2327 );
nand ( n2337 , n2335 , n2336 );
not ( n2338 , n2337 );
nand ( n2339 , n2338 , n1766 );
nand ( n2340 , n1950 , n1953 );
not ( n2341 , n2340 );
and ( n2342 , n2341 , C1 );
nor ( n2343 , C0 , n2342 );
not ( n2344 , n2343 );
nand ( n2345 , n2344 , n1722 );
nor ( n2346 , n2337 , n586 );
buf ( n2347 , n2343 );
nand ( n2348 , n2347 , n587 );
or ( n2349 , n2346 , n2348 );
nand ( n2350 , n2337 , n586 );
nand ( n2351 , n2349 , n2350 );
not ( n2352 , n2351 );
nand ( n2353 , C1 , n2352 );
not ( n2354 , n2353 );
and ( n2355 , n2319 , n2354 );
not ( n2356 , n2319 );
and ( n2357 , n2356 , n2353 );
nor ( n2358 , n2355 , n2357 );
buf ( n2359 , n2358 );
buf ( n2360 , n2359 );
buf ( n2361 , n2360 );
buf ( n2362 , n2361 );
not ( n2363 , n2362 );
buf ( n2364 , n2363 );
buf ( n2365 , n2364 );
not ( n2366 , n2365 );
or ( n2367 , n829 , n2366 );
buf ( n2368 , n2361 );
buf ( n2369 , n596 );
not ( n2370 , n2369 );
buf ( n2371 , n2370 );
buf ( n2372 , n2371 );
nand ( n2373 , n2368 , n2372 );
buf ( n2374 , n2373 );
buf ( n2375 , n2374 );
nand ( n2376 , n2367 , n2375 );
buf ( n2377 , n2376 );
buf ( n2378 , n2377 );
not ( n2379 , n2378 );
or ( n2380 , n827 , n2379 );
nand ( n2381 , C1 , n2348 );
not ( n2382 , n2381 );
not ( n2383 , n2382 );
nand ( n2384 , n2339 , n2350 );
not ( n2385 , n2384 );
not ( n2386 , n2385 );
or ( n2387 , n2383 , n2386 );
nand ( n2388 , n2384 , n2381 );
nand ( n2389 , n2387 , n2388 );
buf ( n2390 , n2389 );
and ( n2391 , n2390 , n2371 );
not ( n2392 , n2390 );
and ( n2393 , n2392 , n596 );
or ( n2394 , n2391 , n2393 );
buf ( n2395 , n2394 );
buf ( n2396 , n2371 );
buf ( n2397 , n822 );
and ( n2398 , n2396 , n2397 );
buf ( n2399 , n596 );
buf ( n2400 , n597 );
and ( n2401 , n2399 , n2400 );
buf ( n2402 , n824 );
nor ( n2403 , n2398 , n2401 , n2402 );
buf ( n2404 , n2403 );
buf ( n2405 , n2404 );
nand ( n2406 , n2395 , n2405 );
buf ( n2407 , n2406 );
buf ( n2408 , n2407 );
nand ( n2409 , n2380 , n2408 );
buf ( n2410 , n2409 );
buf ( n2411 , n2410 );
xnor ( n2412 , C0 , n591 );
buf ( n2413 , n2412 );
buf ( n2414 , n592 );
not ( n2415 , n2414 );
buf ( n2416 , n2415 );
buf ( n2417 , n2416 );
nor ( n2418 , n2413 , n2417 );
buf ( n2419 , n2418 );
buf ( n2420 , n2419 );
buf ( n2421 , n592 );
not ( n2422 , n2421 );
xor ( n2423 , n590 , C0 );
xnor ( n2424 , n2423 , C0 );
not ( n2425 , n2424 );
buf ( n2426 , n2425 );
buf ( n2427 , n2426 );
buf ( n2428 , n2427 );
buf ( n2429 , n2428 );
not ( n2430 , n2429 );
buf ( n2431 , n2430 );
buf ( n2432 , n2431 );
not ( n2433 , n2432 );
or ( n2434 , n2422 , n2433 );
buf ( n2435 , n2425 );
not ( n2436 , n2435 );
buf ( n2437 , n2436 );
buf ( n2438 , n2437 );
not ( n2439 , n2438 );
buf ( n2440 , n2439 );
buf ( n2441 , n2440 );
buf ( n2442 , n2416 );
nand ( n2443 , n2441 , n2442 );
buf ( n2444 , n2443 );
buf ( n2445 , n2444 );
nand ( n2446 , n2434 , n2445 );
buf ( n2447 , n2446 );
buf ( n2448 , n2447 );
buf ( n2449 , n593 );
buf ( n2450 , n594 );
xor ( n2451 , n2449 , n2450 );
buf ( n2452 , n2451 );
buf ( n2453 , n2452 );
and ( n2454 , n2448 , n2453 );
buf ( n2455 , n593 );
not ( n2456 , n2455 );
buf ( n2457 , n2456 );
and ( n2458 , n2416 , n2457 );
and ( n2459 , n592 , n593 );
nor ( n2460 , n2458 , n2459 , n2452 );
buf ( n2461 , n2460 );
not ( n2462 , n2461 );
buf ( n2463 , n2412 );
buf ( n2464 , n592 );
and ( n2465 , n2463 , n2464 );
not ( n2466 , n2412 );
buf ( n2467 , n2466 );
buf ( n2468 , n2416 );
and ( n2469 , n2467 , n2468 );
nor ( n2470 , n2465 , n2469 );
buf ( n2471 , n2470 );
buf ( n2472 , n2471 );
nor ( n2473 , n2462 , n2472 );
buf ( n2474 , n2473 );
buf ( n2475 , n2474 );
nor ( n2476 , n2454 , n2475 );
buf ( n2477 , n2476 );
buf ( n2478 , n2477 );
buf ( n2479 , n594 );
not ( n2480 , n2479 );
buf ( n2481 , n2480 );
buf ( n2482 , n2481 );
buf ( n2483 , n2457 );
or ( n2484 , n2482 , n2483 );
buf ( n2485 , n593 );
buf ( n2486 , n594 );
or ( n2487 , n2485 , n2486 );
buf ( n2488 , n2466 );
nand ( n2489 , n2487 , n2488 );
buf ( n2490 , n2489 );
buf ( n2491 , n2490 );
buf ( n2492 , n592 );
nand ( n2493 , n2484 , n2491 , n2492 );
buf ( n2494 , n2493 );
buf ( n2495 , n2494 );
nor ( n2496 , n2478 , n2495 );
buf ( n2497 , n2496 );
buf ( n2498 , n2497 );
xor ( n2499 , n2420 , n2498 );
buf ( n2500 , n2416 );
not ( n2501 , n2500 );
buf ( n2502 , C0 );
and ( n2503 , C1 , n589 );
nor ( n2504 , C0 , n2503 );
or ( n2505 , n2502 , n2504 );
nand ( n2506 , C1 , n2505 );
buf ( n2507 , n2506 );
not ( n2508 , n2507 );
and ( n2509 , n2501 , n2508 );
buf ( n2510 , n2506 );
buf ( n2511 , n2510 );
buf ( n2512 , n2416 );
and ( n2513 , n2511 , n2512 );
nor ( n2514 , n2509 , n2513 );
buf ( n2515 , n2514 );
buf ( n2516 , n2515 );
buf ( n2517 , n2452 );
not ( n2518 , n2517 );
buf ( n2519 , n2518 );
buf ( n2520 , n2519 );
or ( n2521 , n2516 , n2520 );
buf ( n2522 , n2447 );
buf ( n2523 , n2460 );
nand ( n2524 , n2522 , n2523 );
buf ( n2525 , n2524 );
buf ( n2526 , n2525 );
nand ( n2527 , n2521 , n2526 );
buf ( n2528 , n2527 );
buf ( n2529 , n2528 );
xor ( n2530 , n2499 , n2529 );
buf ( n2531 , n2530 );
buf ( n2532 , n2531 );
not ( n2533 , n596 );
buf ( n2534 , n595 );
not ( n2535 , n2534 );
buf ( n2536 , n2535 );
not ( n2537 , n2536 );
and ( n2538 , n2533 , n2537 );
nor ( n2539 , n2371 , n595 );
nor ( n2540 , n2538 , n2539 );
not ( n2541 , n2540 );
buf ( n2542 , n2541 );
not ( n2543 , n2542 );
nand ( n2544 , n2343 , n587 );
nand ( n2545 , n2345 , n2544 );
not ( n2546 , n2545 );
not ( n2547 , n2546 );
or ( n2548 , C0 , n2547 );
nand ( n2549 , n2548 , C1 );
buf ( n2550 , n2549 );
buf ( n2551 , n2550 );
buf ( n2552 , n2551 );
buf ( n2553 , n2552 );
not ( n2554 , n2553 );
buf ( n2555 , n2554 );
buf ( n2556 , n2555 );
buf ( n2557 , n2556 );
buf ( n2558 , n2557 );
and ( n2559 , n2558 , n594 );
not ( n2560 , n2558 );
and ( n2561 , n2560 , n2481 );
or ( n2562 , n2559 , n2561 );
buf ( n2563 , n2562 );
not ( n2564 , n2563 );
or ( n2565 , n2543 , n2564 );
buf ( n2566 , n594 );
not ( n2567 , n2566 );
nand ( n2568 , n2326 , C1 );
and ( n2569 , n2568 , C1 );
nor ( n2570 , n2569 , C0 );
buf ( n2571 , n2570 );
buf ( n2572 , n2571 );
buf ( n2573 , n2572 );
buf ( n2574 , n2573 );
not ( n2575 , n2574 );
buf ( n2576 , n2575 );
buf ( n2577 , n2576 );
not ( n2578 , n2577 );
or ( n2579 , n2567 , n2578 );
buf ( n2580 , n2573 );
buf ( n2581 , n2481 );
nand ( n2582 , n2580 , n2581 );
buf ( n2583 , n2582 );
buf ( n2584 , n2583 );
nand ( n2585 , n2579 , n2584 );
buf ( n2586 , n2585 );
buf ( n2587 , n2586 );
and ( n2588 , n2536 , n2481 );
and ( n2589 , n595 , n594 );
nor ( n2590 , n2588 , n2589 );
nand ( n2591 , n2540 , n2590 );
not ( n2592 , n2591 );
buf ( n2593 , n2592 );
nand ( n2594 , n2587 , n2593 );
buf ( n2595 , n2594 );
buf ( n2596 , n2595 );
nand ( n2597 , n2565 , n2596 );
buf ( n2598 , n2597 );
buf ( n2599 , n2598 );
xor ( n2600 , n2532 , n2599 );
xor ( n2601 , n2494 , n2477 );
buf ( n2602 , n2601 );
buf ( n2603 , n2541 );
not ( n2604 , n2603 );
buf ( n2605 , n2586 );
not ( n2606 , n2605 );
or ( n2607 , n2604 , n2606 );
buf ( n2608 , n594 );
not ( n2609 , n2608 );
buf ( n2610 , n2506 );
not ( n2611 , n2610 );
buf ( n2612 , n2611 );
buf ( n2613 , n2612 );
not ( n2614 , n2613 );
or ( n2615 , n2609 , n2614 );
buf ( n2616 , n2510 );
buf ( n2617 , n2481 );
nand ( n2618 , n2616 , n2617 );
buf ( n2619 , n2618 );
buf ( n2620 , n2619 );
nand ( n2621 , n2615 , n2620 );
buf ( n2622 , n2621 );
buf ( n2623 , n2622 );
buf ( n2624 , n2592 );
nand ( n2625 , n2623 , n2624 );
buf ( n2626 , n2625 );
buf ( n2627 , n2626 );
nand ( n2628 , n2607 , n2627 );
buf ( n2629 , n2628 );
buf ( n2630 , n2629 );
xor ( n2631 , n2602 , n2630 );
buf ( n2632 , n2412 );
buf ( n2633 , n2519 );
nor ( n2634 , n2632 , n2633 );
buf ( n2635 , n2634 );
buf ( n2636 , n2635 );
buf ( n2637 , n2541 );
not ( n2638 , n2637 );
buf ( n2639 , n594 );
not ( n2640 , n2639 );
buf ( n2641 , n2437 );
not ( n2642 , n2641 );
or ( n2643 , n2640 , n2642 );
buf ( n2644 , n2428 );
buf ( n2645 , n2481 );
nand ( n2646 , n2644 , n2645 );
buf ( n2647 , n2646 );
buf ( n2648 , n2647 );
nand ( n2649 , n2643 , n2648 );
buf ( n2650 , n2649 );
buf ( n2651 , n2650 );
not ( n2652 , n2651 );
or ( n2653 , n2638 , n2652 );
buf ( n2654 , n2466 );
buf ( n2655 , n2592 );
buf ( n2656 , n594 );
not ( n2657 , n2656 );
and ( n2658 , n2655 , n2657 );
buf ( n2659 , n2658 );
buf ( n2660 , n2659 );
and ( n2661 , n2654 , n2660 );
buf ( n2662 , n2412 );
buf ( n2663 , n2592 );
buf ( n2664 , n594 );
nand ( n2665 , n2663 , n2664 );
buf ( n2666 , n2665 );
buf ( n2667 , n2666 );
not ( n2668 , n2667 );
buf ( n2669 , n2668 );
buf ( n2670 , n2669 );
and ( n2671 , n2662 , n2670 );
nor ( n2672 , n2661 , n2671 );
buf ( n2673 , n2672 );
buf ( n2674 , n2673 );
nand ( n2675 , n2653 , n2674 );
buf ( n2676 , n2675 );
buf ( n2677 , n2676 );
not ( n2678 , n2677 );
buf ( n2679 , n2371 );
buf ( n2680 , n2536 );
or ( n2681 , n2679 , n2680 );
buf ( n2682 , n595 );
buf ( n2683 , n596 );
or ( n2684 , n2682 , n2683 );
buf ( n2685 , n2466 );
nand ( n2686 , n2684 , n2685 );
buf ( n2687 , n2686 );
buf ( n2688 , n2687 );
buf ( n2689 , n594 );
nand ( n2690 , n2681 , n2688 , n2689 );
buf ( n2691 , n2690 );
buf ( n2692 , n2691 );
nor ( n2693 , n2678 , n2692 );
buf ( n2694 , n2693 );
buf ( n2695 , n2694 );
xor ( n2696 , n2636 , n2695 );
buf ( n2697 , n2541 );
not ( n2698 , n2697 );
buf ( n2699 , n2622 );
not ( n2700 , n2699 );
or ( n2701 , n2698 , n2700 );
buf ( n2702 , n2650 );
buf ( n2703 , n2592 );
nand ( n2704 , n2702 , n2703 );
buf ( n2705 , n2704 );
buf ( n2706 , n2705 );
nand ( n2707 , n2701 , n2706 );
buf ( n2708 , n2707 );
buf ( n2709 , n2708 );
and ( n2710 , n2696 , n2709 );
or ( n2711 , n2710 , C0 );
buf ( n2712 , n2711 );
buf ( n2713 , n2712 );
and ( n2714 , n2631 , n2713 );
and ( n2715 , n2602 , n2630 );
or ( n2716 , n2714 , n2715 );
buf ( n2717 , n2716 );
buf ( n2718 , n2717 );
xor ( n2719 , n2600 , n2718 );
buf ( n2720 , n2719 );
buf ( n2721 , n2720 );
xor ( n2722 , n2411 , n2721 );
buf ( n2723 , n825 );
not ( n2724 , n2723 );
buf ( n2725 , n2394 );
not ( n2726 , n2725 );
or ( n2727 , n2724 , n2726 );
buf ( n2728 , n596 );
not ( n2729 , n2728 );
buf ( n2730 , n2558 );
not ( n2731 , n2730 );
or ( n2732 , n2729 , n2731 );
buf ( n2733 , n2549 );
not ( n2734 , n2733 );
buf ( n2735 , n2734 );
buf ( n2736 , n2735 );
buf ( n2737 , n2736 );
buf ( n2738 , n2737 );
buf ( n2739 , n2738 );
not ( n2740 , n2739 );
buf ( n2741 , n2371 );
nand ( n2742 , n2740 , n2741 );
buf ( n2743 , n2742 );
buf ( n2744 , n2743 );
nand ( n2745 , n2732 , n2744 );
buf ( n2746 , n2745 );
buf ( n2747 , n2746 );
buf ( n2748 , n2404 );
nand ( n2749 , n2747 , n2748 );
buf ( n2750 , n2749 );
buf ( n2751 , n2750 );
nand ( n2752 , n2727 , n2751 );
buf ( n2753 , n2752 );
buf ( n2754 , n2753 );
xor ( n2755 , n2602 , n2630 );
xor ( n2756 , n2755 , n2713 );
buf ( n2757 , n2756 );
buf ( n2758 , n2757 );
xor ( n2759 , n2754 , n2758 );
xor ( n2760 , n2636 , n2695 );
xor ( n2761 , n2760 , n2709 );
buf ( n2762 , n2761 );
buf ( n2763 , n2762 );
buf ( n2764 , n825 );
not ( n2765 , n2764 );
buf ( n2766 , n2746 );
not ( n2767 , n2766 );
or ( n2768 , n2765 , n2767 );
buf ( n2769 , n596 );
not ( n2770 , n2769 );
buf ( n2771 , n2576 );
not ( n2772 , n2771 );
or ( n2773 , n2770 , n2772 );
buf ( n2774 , n2573 );
buf ( n2775 , n2371 );
nand ( n2776 , n2774 , n2775 );
buf ( n2777 , n2776 );
buf ( n2778 , n2777 );
nand ( n2779 , n2773 , n2778 );
buf ( n2780 , n2779 );
buf ( n2781 , n2780 );
buf ( n2782 , n2404 );
nand ( n2783 , n2781 , n2782 );
buf ( n2784 , n2783 );
buf ( n2785 , n2784 );
nand ( n2786 , n2768 , n2785 );
buf ( n2787 , n2786 );
buf ( n2788 , n2787 );
xor ( n2789 , n2763 , n2788 );
buf ( n2790 , n2691 );
not ( n2791 , n2790 );
buf ( n2792 , n2676 );
not ( n2793 , n2792 );
or ( n2794 , n2791 , n2793 );
buf ( n2795 , n2676 );
buf ( n2796 , n2691 );
or ( n2797 , n2795 , n2796 );
nand ( n2798 , n2794 , n2797 );
buf ( n2799 , n2798 );
buf ( n2800 , n2799 );
buf ( n2801 , n825 );
not ( n2802 , n2801 );
buf ( n2803 , n2780 );
not ( n2804 , n2803 );
or ( n2805 , n2802 , n2804 );
buf ( n2806 , n596 );
not ( n2807 , n2806 );
buf ( n2808 , n2612 );
not ( n2809 , n2808 );
or ( n2810 , n2807 , n2809 );
buf ( n2811 , n2510 );
buf ( n2812 , n2371 );
nand ( n2813 , n2811 , n2812 );
buf ( n2814 , n2813 );
buf ( n2815 , n2814 );
nand ( n2816 , n2810 , n2815 );
buf ( n2817 , n2816 );
buf ( n2818 , n2817 );
buf ( n2819 , n2404 );
nand ( n2820 , n2818 , n2819 );
buf ( n2821 , n2820 );
buf ( n2822 , n2821 );
nand ( n2823 , n2805 , n2822 );
buf ( n2824 , n2823 );
buf ( n2825 , n2824 );
xor ( n2826 , n2800 , n2825 );
buf ( n2827 , n2540 );
buf ( n2828 , n2412 );
nor ( n2829 , n2827 , n2828 );
buf ( n2830 , n2829 );
buf ( n2831 , n2830 );
not ( n2832 , n824 );
not ( n2833 , n596 );
not ( n2834 , n2431 );
or ( n2835 , n2833 , n2834 );
buf ( n2836 , n2440 );
buf ( n2837 , n2371 );
nand ( n2838 , n2836 , n2837 );
buf ( n2839 , n2838 );
nand ( n2840 , n2835 , n2839 );
not ( n2841 , n2840 );
or ( n2842 , n2832 , n2841 );
and ( n2843 , n2404 , n596 );
and ( n2844 , n2843 , n2412 );
and ( n2845 , n2404 , n2371 );
and ( n2846 , n2845 , n2466 );
nor ( n2847 , n2844 , n2846 );
nand ( n2848 , n2842 , n2847 );
buf ( n2849 , n2848 );
not ( n2850 , n2849 );
buf ( n2851 , n597 );
buf ( n2852 , n598 );
or ( n2853 , n2851 , n2852 );
buf ( n2854 , n2466 );
nand ( n2855 , n2853 , n2854 );
buf ( n2856 , n2855 );
buf ( n2857 , n2856 );
buf ( n2858 , n597 );
buf ( n2859 , n598 );
nand ( n2860 , n2858 , n2859 );
buf ( n2861 , n2860 );
buf ( n2862 , n2861 );
buf ( n2863 , n596 );
nand ( n2864 , n2857 , n2862 , n2863 );
buf ( n2865 , n2864 );
buf ( n2866 , n2865 );
nor ( n2867 , n2850 , n2866 );
buf ( n2868 , n2867 );
buf ( n2869 , n2868 );
xor ( n2870 , n2831 , n2869 );
buf ( n2871 , n825 );
not ( n2872 , n2871 );
buf ( n2873 , n2817 );
not ( n2874 , n2873 );
or ( n2875 , n2872 , n2874 );
buf ( n2876 , n2840 );
buf ( n2877 , n2404 );
nand ( n2878 , n2876 , n2877 );
buf ( n2879 , n2878 );
buf ( n2880 , n2879 );
nand ( n2881 , n2875 , n2880 );
buf ( n2882 , n2881 );
buf ( n2883 , n2882 );
and ( n2884 , n2870 , n2883 );
or ( n2885 , n2884 , C0 );
buf ( n2886 , n2885 );
buf ( n2887 , n2886 );
and ( n2888 , n2826 , n2887 );
and ( n2889 , n2800 , n2825 );
or ( n2890 , n2888 , n2889 );
buf ( n2891 , n2890 );
buf ( n2892 , n2891 );
and ( n2893 , n2789 , n2892 );
and ( n2894 , n2763 , n2788 );
or ( n2895 , n2893 , n2894 );
buf ( n2896 , n2895 );
buf ( n2897 , n2896 );
and ( n2898 , n2759 , n2897 );
and ( n2899 , n2754 , n2758 );
or ( n2900 , n2898 , n2899 );
buf ( n2901 , n2900 );
buf ( n2902 , n2901 );
and ( n2903 , n2722 , n2902 );
and ( n2904 , n2411 , n2721 );
or ( n2905 , n2903 , n2904 );
buf ( n2906 , n2905 );
buf ( n2907 , n2906 );
and ( n2908 , n601 , n602 );
not ( n2909 , n601 );
buf ( n2910 , n602 );
not ( n2911 , n2910 );
buf ( n2912 , n2911 );
and ( n2913 , n2909 , n2912 );
nor ( n2914 , n2908 , n2913 );
buf ( n2915 , n2914 );
buf ( n2916 , n2915 );
not ( n2917 , n2916 );
buf ( n2918 , n600 );
not ( n2919 , n2918 );
or ( n2920 , n553 , n554 );
nand ( n2921 , n2920 , n1798 );
nand ( n2922 , n553 , n554 );
and ( n2923 , n2921 , n2922 , n552 );
not ( n2924 , n2265 );
not ( n2925 , n552 );
not ( n2926 , n1855 );
or ( n2927 , n2925 , n2926 );
not ( n2928 , n552 );
nand ( n2929 , n2928 , n1791 );
nand ( n2930 , n2927 , n2929 );
not ( n2931 , n2930 );
or ( n2932 , n2924 , n2931 );
and ( n2933 , n552 , n1687 );
not ( n2934 , n552 );
and ( n2935 , n2934 , n1664 );
or ( n2936 , n2933 , n2935 );
xnor ( n2937 , n552 , n553 );
nor ( n2938 , n2265 , n2937 );
nand ( n2939 , n2936 , n2938 );
nand ( n2940 , n2932 , n2939 );
and ( n2941 , n2923 , n2940 );
not ( n2942 , n1659 );
not ( n2943 , n556 );
not ( n2944 , n1772 );
not ( n2945 , n2944 );
or ( n2946 , n2943 , n2945 );
nand ( n2947 , n1772 , n1625 );
nand ( n2948 , n2946 , n2947 );
not ( n2949 , n2948 );
or ( n2950 , n2942 , n2949 );
not ( n2951 , n1594 );
nor ( n2952 , n2951 , n1625 );
nand ( n2953 , n2952 , n2252 );
not ( n2954 , n2953 );
not ( n2955 , n1594 );
nor ( n2956 , n2955 , n556 );
and ( n2957 , n2251 , n2956 );
nor ( n2958 , n2954 , n2957 );
nand ( n2959 , n2950 , n2958 );
xor ( n2960 , n2941 , n2959 );
not ( n2961 , n1739 );
and ( n2962 , n568 , n584 );
not ( n2963 , n568 );
not ( n2964 , n584 );
and ( n2965 , n2963 , n2964 );
nor ( n2966 , n2962 , n2965 );
or ( n2967 , n571 , n587 );
or ( n2968 , n570 , n586 );
nand ( n2969 , n2967 , n2968 );
nor ( n2970 , n2969 , n2242 );
not ( n2971 , n2970 );
not ( n2972 , n1720 );
or ( n2973 , n2971 , n2972 );
not ( n2974 , n569 );
nand ( n2975 , n2974 , n2317 );
and ( n2976 , n2239 , n2975 );
not ( n2977 , n2244 );
nor ( n2978 , n2976 , n2977 );
nand ( n2979 , n2973 , n2978 );
xor ( n2980 , n2966 , n2979 );
buf ( n2981 , n2980 );
not ( n2982 , n2981 );
and ( n2983 , n558 , n2982 );
not ( n2984 , n558 );
and ( n2985 , n2984 , n2981 );
or ( n2986 , n2983 , n2985 );
not ( n2987 , n2986 );
or ( n2988 , n2961 , n2987 );
not ( n2989 , n558 );
nand ( n2990 , n567 , n583 );
not ( n2991 , n2990 );
nor ( n2992 , n567 , n583 );
nor ( n2993 , n2991 , n2992 );
not ( n2994 , n585 );
not ( n2995 , n569 );
nand ( n2996 , n2994 , n2995 );
not ( n2997 , n568 );
nand ( n2998 , n2964 , n2997 );
nand ( n2999 , n1617 , n2996 , n2998 );
nor ( n3000 , n2999 , n2232 );
not ( n3001 , n3000 );
not ( n3002 , n1607 );
not ( n3003 , n1604 );
or ( n3004 , n3002 , n3003 );
nand ( n3005 , n573 , n589 );
nand ( n3006 , n572 , n588 );
and ( n3007 , n3005 , n3006 );
nand ( n3008 , n3004 , n3007 );
not ( n3009 , n3008 );
or ( n3010 , n3001 , n3009 );
nand ( n3011 , n568 , n584 );
not ( n3012 , n3011 );
not ( n3013 , n584 );
not ( n3014 , n3013 );
not ( n3015 , n568 );
not ( n3016 , n3015 );
or ( n3017 , n3014 , n3016 );
nand ( n3018 , n3017 , n2975 );
not ( n3019 , n3018 );
or ( n3020 , n3012 , n3019 );
nand ( n3021 , n570 , n586 );
nand ( n3022 , n568 , n584 );
nand ( n3023 , n569 , n585 );
nand ( n3024 , n3021 , n3022 , n3023 );
not ( n3025 , n3024 );
not ( n3026 , n1766 );
not ( n3027 , n1764 );
or ( n3028 , n3026 , n3027 );
and ( n3029 , n571 , n587 );
nand ( n3030 , n3028 , n3029 );
nand ( n3031 , n3025 , n3030 );
nand ( n3032 , n3020 , n3031 );
nand ( n3033 , n3010 , n3032 );
buf ( n3034 , n3033 );
xor ( n3035 , n2993 , n3034 );
buf ( n3036 , n3035 );
not ( n3037 , n3036 );
not ( n3038 , n3037 );
or ( n3039 , n2989 , n3038 );
nand ( n3040 , n3036 , n1736 );
nand ( n3041 , n3039 , n3040 );
nand ( n3042 , n3041 , n559 );
nand ( n3043 , n2988 , n3042 );
and ( n3044 , n2960 , n3043 );
and ( n3045 , n2941 , n2959 );
or ( n3046 , n3044 , n3045 );
not ( n3047 , n2265 );
not ( n3048 , n552 );
not ( n3049 , n1624 );
not ( n3050 , n3049 );
or ( n3051 , n3048 , n3050 );
not ( n3052 , n552 );
nand ( n3053 , n3052 , n1624 );
nand ( n3054 , n3051 , n3053 );
not ( n3055 , n3054 );
or ( n3056 , n3047 , n3055 );
not ( n3057 , n552 );
not ( n3058 , n1652 );
or ( n3059 , n3057 , n3058 );
not ( n3060 , n552 );
nand ( n3061 , n3060 , n1651 );
nand ( n3062 , n3059 , n3061 );
nor ( n3063 , n2937 , n2265 );
buf ( n3064 , n3063 );
nand ( n3065 , n3062 , n3064 );
nand ( n3066 , n3056 , n3065 );
xor ( n3067 , n551 , n552 );
buf ( n3068 , n3067 );
not ( n3069 , n3068 );
not ( n3070 , n550 );
not ( n3071 , n1677 );
or ( n3072 , n3070 , n3071 );
not ( n3073 , n550 );
nand ( n3074 , n1680 , n3073 );
nand ( n3075 , n3072 , n3074 );
not ( n3076 , n3075 );
or ( n3077 , n3069 , n3076 );
not ( n3078 , n550 );
not ( n3079 , n1687 );
or ( n3080 , n3078 , n3079 );
nand ( n3081 , n1664 , n3073 );
nand ( n3082 , n3080 , n3081 );
xnor ( n3083 , n550 , n551 );
nor ( n3084 , n3067 , n3083 );
nand ( n3085 , n3082 , n3084 );
nand ( n3086 , n3077 , n3085 );
or ( n3087 , n551 , n552 );
not ( n3088 , n3087 );
not ( n3089 , n1664 );
or ( n3090 , n3088 , n3089 );
nand ( n3091 , n551 , n552 );
and ( n3092 , n3091 , n550 );
nand ( n3093 , n3090 , n3092 );
and ( n3094 , n3086 , n3093 );
not ( n3095 , n3086 );
not ( n3096 , n3093 );
and ( n3097 , n3095 , n3096 );
or ( n3098 , n3094 , n3097 );
xor ( n3099 , n3066 , n3098 );
not ( n3100 , n1596 );
not ( n3101 , n556 );
not ( n3102 , n2982 );
or ( n3103 , n3101 , n3102 );
not ( n3104 , n2982 );
nand ( n3105 , n3104 , n1625 );
nand ( n3106 , n3103 , n3105 );
not ( n3107 , n3106 );
or ( n3108 , n3100 , n3107 );
and ( n3109 , n1810 , n556 );
and ( n3110 , n2252 , n3109 );
not ( n3111 , n2252 );
and ( n3112 , n1659 , n1625 );
and ( n3113 , n3111 , n3112 );
nor ( n3114 , n3110 , n3113 );
nand ( n3115 , n3108 , n3114 );
xor ( n3116 , n3099 , n3115 );
xor ( n3117 , n3046 , n3116 );
buf ( n3118 , n1668 );
not ( n3119 , n3118 );
not ( n3120 , n554 );
not ( n3121 , n2944 );
or ( n3122 , n3120 , n3121 );
nand ( n3123 , n1772 , n1681 );
nand ( n3124 , n3122 , n3123 );
not ( n3125 , n3124 );
or ( n3126 , n3119 , n3125 );
not ( n3127 , n554 );
not ( n3128 , n1733 );
or ( n3129 , n3127 , n3128 );
nand ( n3130 , n1732 , n1681 );
nand ( n3131 , n3129 , n3130 );
nand ( n3132 , n3131 , n2276 );
nand ( n3133 , n3126 , n3132 );
and ( n3134 , n1664 , n3067 );
not ( n3135 , n2265 );
not ( n3136 , n3062 );
or ( n3137 , n3135 , n3136 );
nand ( n3138 , n2930 , n3063 );
nand ( n3139 , n3137 , n3138 );
xor ( n3140 , n3134 , n3139 );
not ( n3141 , n1668 );
not ( n3142 , n3131 );
or ( n3143 , n3141 , n3142 );
and ( n3144 , n1621 , n554 );
not ( n3145 , n1621 );
and ( n3146 , n3145 , n1681 );
or ( n3147 , n3144 , n3146 );
nand ( n3148 , n3147 , n2276 );
nand ( n3149 , n3143 , n3148 );
and ( n3150 , n3140 , n3149 );
and ( n3151 , n3134 , n3139 );
or ( n3152 , n3150 , n3151 );
xor ( n3153 , n3133 , n3152 );
not ( n3154 , n559 );
not ( n3155 , n558 );
not ( n3156 , n2992 );
not ( n3157 , n3156 );
not ( n3158 , n3033 );
or ( n3159 , n3157 , n3158 );
nand ( n3160 , n3159 , n2990 );
xnor ( n3161 , n566 , n582 );
not ( n3162 , n3161 );
and ( n3163 , n3160 , n3162 );
not ( n3164 , n3160 );
and ( n3165 , n3164 , n3161 );
nor ( n3166 , n3163 , n3165 );
buf ( n3167 , n3166 );
not ( n3168 , n3167 );
not ( n3169 , n3168 );
or ( n3170 , n3155 , n3169 );
not ( n3171 , n558 );
nand ( n3172 , n3171 , n3167 );
nand ( n3173 , n3170 , n3172 );
not ( n3174 , n3173 );
or ( n3175 , n3154 , n3174 );
nand ( n3176 , n3041 , n1739 );
nand ( n3177 , n3175 , n3176 );
xor ( n3178 , n3153 , n3177 );
and ( n3179 , n3117 , n3178 );
and ( n3180 , n3046 , n3116 );
or ( n3181 , n3179 , n3180 );
and ( n3182 , n3086 , n3096 );
not ( n3183 , n1659 );
not ( n3184 , n3106 );
or ( n3185 , n3183 , n3184 );
and ( n3186 , n3036 , n1625 );
not ( n3187 , n3036 );
and ( n3188 , n3187 , n556 );
or ( n3189 , n3186 , n3188 );
nand ( n3190 , n3189 , n1594 );
nand ( n3191 , n3185 , n3190 );
xor ( n3192 , n3182 , n3191 );
not ( n3193 , n3118 );
not ( n3194 , n554 );
not ( n3195 , n2251 );
not ( n3196 , n3195 );
or ( n3197 , n3194 , n3196 );
not ( n3198 , n3195 );
nand ( n3199 , n3198 , n1681 );
nand ( n3200 , n3197 , n3199 );
not ( n3201 , n3200 );
or ( n3202 , n3193 , n3201 );
nand ( n3203 , n3124 , n2276 );
nand ( n3204 , n3202 , n3203 );
xor ( n3205 , n3192 , n3204 );
xor ( n3206 , n3133 , n3152 );
and ( n3207 , n3206 , n3177 );
and ( n3208 , n3133 , n3152 );
or ( n3209 , n3207 , n3208 );
xor ( n3210 , n3205 , n3209 );
not ( n3211 , n1664 );
xor ( n3212 , n549 , n550 );
not ( n3213 , n3212 );
nor ( n3214 , n3211 , n3213 );
not ( n3215 , n3068 );
not ( n3216 , n550 );
not ( n3217 , n1652 );
or ( n3218 , n3216 , n3217 );
nand ( n3219 , n1651 , n3073 );
nand ( n3220 , n3218 , n3219 );
not ( n3221 , n3220 );
or ( n3222 , n3215 , n3221 );
nand ( n3223 , n3075 , n3084 );
nand ( n3224 , n3222 , n3223 );
xor ( n3225 , n3214 , n3224 );
not ( n3226 , n2265 );
not ( n3227 , n552 );
not ( n3228 , n1733 );
or ( n3229 , n3227 , n3228 );
not ( n3230 , n552 );
nand ( n3231 , n3230 , n1732 );
nand ( n3232 , n3229 , n3231 );
not ( n3233 , n3232 );
or ( n3234 , n3226 , n3233 );
nand ( n3235 , n3054 , n3064 );
nand ( n3236 , n3234 , n3235 );
xor ( n3237 , n3225 , n3236 );
not ( n3238 , n559 );
not ( n3239 , n566 );
not ( n3240 , n582 );
and ( n3241 , n3239 , n3240 );
nor ( n3242 , n3241 , n2992 );
not ( n3243 , n3242 );
not ( n3244 , n3033 );
or ( n3245 , n3243 , n3244 );
not ( n3246 , n566 );
not ( n3247 , n582 );
or ( n3248 , n3246 , n3247 );
nor ( n3249 , n566 , n582 );
nand ( n3250 , n567 , n583 );
or ( n3251 , n3249 , n3250 );
nand ( n3252 , n3248 , n3251 );
buf ( n3253 , n3252 );
not ( n3254 , n3253 );
nand ( n3255 , n3245 , n3254 );
or ( n3256 , n565 , n581 );
nand ( n3257 , n565 , n581 );
nand ( n3258 , n3256 , n3257 );
not ( n3259 , n3258 );
and ( n3260 , n3255 , n3259 );
not ( n3261 , n3255 );
and ( n3262 , n3261 , n3258 );
nor ( n3263 , n3260 , n3262 );
buf ( n3264 , n3263 );
not ( n3265 , n3264 );
and ( n3266 , n3265 , n558 );
not ( n3267 , n3265 );
and ( n3268 , n3267 , n1736 );
or ( n3269 , n3266 , n3268 );
not ( n3270 , n3269 );
or ( n3271 , n3238 , n3270 );
nand ( n3272 , n3173 , n1739 );
nand ( n3273 , n3271 , n3272 );
xor ( n3274 , n3237 , n3273 );
xor ( n3275 , n3066 , n3098 );
and ( n3276 , n3275 , n3115 );
and ( n3277 , n3066 , n3098 );
or ( n3278 , n3276 , n3277 );
xor ( n3279 , n3274 , n3278 );
xor ( n3280 , n3210 , n3279 );
buf ( n3281 , n3280 );
not ( n3282 , n3281 );
xor ( n3283 , n3181 , n3282 );
xor ( n3284 , n3134 , n3139 );
xor ( n3285 , n3284 , n3149 );
not ( n3286 , n1668 );
not ( n3287 , n3147 );
or ( n3288 , n3286 , n3287 );
nand ( n3289 , n2272 , n2276 );
nand ( n3290 , n3288 , n3289 );
xor ( n3291 , n2923 , n2940 );
xor ( n3292 , n3290 , n3291 );
not ( n3293 , n1596 );
not ( n3294 , n2948 );
or ( n3295 , n3293 , n3294 );
nand ( n3296 , n2224 , n1659 );
nand ( n3297 , n3295 , n3296 );
and ( n3298 , n3292 , n3297 );
and ( n3299 , n3290 , n3291 );
or ( n3300 , n3298 , n3299 );
xor ( n3301 , n3285 , n3300 );
xor ( n3302 , n2941 , n2959 );
xor ( n3303 , n3302 , n3043 );
and ( n3304 , n3301 , n3303 );
and ( n3305 , n3285 , n3300 );
or ( n3306 , n3304 , n3305 );
not ( n3307 , n3306 );
xor ( n3308 , n3046 , n3116 );
xor ( n3309 , n3308 , n3178 );
not ( n3310 , n3309 );
or ( n3311 , n3307 , n3310 );
xor ( n3312 , n3285 , n3300 );
xor ( n3313 , n3312 , n3303 );
not ( n3314 , n559 );
not ( n3315 , n2986 );
or ( n3316 , n3314 , n3315 );
nand ( n3317 , n2257 , n1739 );
nand ( n3318 , n3316 , n3317 );
xor ( n3319 , n2266 , n2278 );
and ( n3320 , n3319 , n2280 );
and ( n3321 , n2266 , n2278 );
or ( n3322 , n3320 , n3321 );
xor ( n3323 , n3318 , n3322 );
xor ( n3324 , n3290 , n3291 );
xor ( n3325 , n3324 , n3297 );
and ( n3326 , n3323 , n3325 );
and ( n3327 , n3318 , n3322 );
or ( n3328 , n3326 , n3327 );
nand ( n3329 , n3313 , n3328 );
nand ( n3330 , n3311 , n3329 );
not ( n3331 , n3330 );
not ( n3332 , n3309 );
not ( n3333 , n3306 );
nand ( n3334 , n3332 , n3333 );
not ( n3335 , n3334 );
or ( n3336 , n3331 , n3335 );
not ( n3337 , n3309 );
nand ( n3338 , n3337 , n3333 );
xor ( n3339 , n3318 , n3322 );
xor ( n3340 , n3339 , n3325 );
not ( n3341 , n3340 );
xor ( n3342 , n2228 , n2263 );
and ( n3343 , n3342 , n2281 );
and ( n3344 , n2228 , n2263 );
or ( n3345 , n3343 , n3344 );
not ( n3346 , n3345 );
nand ( n3347 , n3341 , n3346 );
not ( n3348 , n3347 );
not ( n3349 , n2284 );
not ( n3350 , n2288 );
or ( n3351 , n3349 , n3350 );
not ( n3352 , n2283 );
not ( n3353 , n2291 );
or ( n3354 , n3352 , n3353 );
nand ( n3355 , n3354 , n2300 );
nand ( n3356 , n3351 , n3355 );
not ( n3357 , n3356 );
or ( n3358 , n3348 , n3357 );
buf ( n3359 , n3340 );
nand ( n3360 , n3359 , n3345 );
nand ( n3361 , n3358 , n3360 );
not ( n3362 , n3313 );
not ( n3363 , n3328 );
nand ( n3364 , n3362 , n3363 );
nand ( n3365 , n3338 , n3361 , n3364 );
nand ( n3366 , n3336 , n3365 );
buf ( n3367 , n3366 );
xnor ( n3368 , n3283 , n3367 );
not ( n3369 , n3368 );
xor ( n3370 , n2005 , n2017 );
and ( n3371 , n3370 , n2034 );
and ( n3372 , n2005 , n2017 );
or ( n3373 , n3371 , n3372 );
buf ( n3374 , n2012 );
not ( n3375 , n3374 );
buf ( n3376 , n1110 );
not ( n3377 , n3376 );
or ( n3378 , n3375 , n3377 );
buf ( n3379 , n552 );
buf ( n3380 , n574 );
xor ( n3381 , n3379 , n3380 );
buf ( n3382 , n3381 );
buf ( n3383 , n3382 );
buf ( n3384 , n575 );
nand ( n3385 , n3383 , n3384 );
buf ( n3386 , n3385 );
buf ( n3387 , n3386 );
nand ( n3388 , n3378 , n3387 );
buf ( n3389 , n3388 );
buf ( n3390 , n3389 );
buf ( n3391 , n559 );
buf ( n3392 , n569 );
or ( n3393 , n3391 , n3392 );
buf ( n3394 , n570 );
nand ( n3395 , n3393 , n3394 );
buf ( n3396 , n3395 );
buf ( n3397 , n3396 );
buf ( n3398 , n559 );
buf ( n3399 , n569 );
nand ( n3400 , n3398 , n3399 );
buf ( n3401 , n3400 );
buf ( n3402 , n3401 );
buf ( n3403 , n568 );
nand ( n3404 , n3397 , n3402 , n3403 );
buf ( n3405 , n3404 );
buf ( n3406 , n3405 );
and ( n3407 , n3390 , n3406 );
not ( n3408 , n3390 );
buf ( n3409 , n3405 );
not ( n3410 , n3409 );
buf ( n3411 , n3410 );
buf ( n3412 , n3411 );
and ( n3413 , n3408 , n3412 );
nor ( n3414 , n3407 , n3413 );
buf ( n3415 , n3414 );
xor ( n3416 , n3373 , n3415 );
buf ( n3417 , n559 );
buf ( n3418 , n568 );
xor ( n3419 , n3417 , n3418 );
buf ( n3420 , n3419 );
buf ( n3421 , n3420 );
not ( n3422 , n3421 );
not ( n3423 , n2001 );
not ( n3424 , n568 );
nand ( n3425 , n3424 , n569 );
not ( n3426 , n569 );
nand ( n3427 , n3426 , n568 );
nand ( n3428 , n3425 , n3427 );
and ( n3429 , n3423 , n3428 );
buf ( n3430 , n3429 );
not ( n3431 , n3430 );
or ( n3432 , n3422 , n3431 );
and ( n3433 , n569 , n570 );
not ( n3434 , n569 );
and ( n3435 , n3434 , n1764 );
nor ( n3436 , n3433 , n3435 );
buf ( n3437 , n3436 );
buf ( n3438 , n3437 );
buf ( n3439 , n3438 );
buf ( n3440 , n3439 );
buf ( n3441 , n558 );
buf ( n3442 , n568 );
xor ( n3443 , n3441 , n3442 );
buf ( n3444 , n3443 );
buf ( n3445 , n3444 );
nand ( n3446 , n3440 , n3445 );
buf ( n3447 , n3446 );
buf ( n3448 , n3447 );
nand ( n3449 , n3432 , n3448 );
buf ( n3450 , n3449 );
buf ( n3451 , n3450 );
not ( n3452 , n3451 );
buf ( n3453 , n2028 );
not ( n3454 , n3453 );
buf ( n3455 , n884 );
not ( n3456 , n3455 );
or ( n3457 , n3454 , n3456 );
buf ( n3458 , n888 );
buf ( n3459 , n554 );
buf ( n3460 , n572 );
xor ( n3461 , n3459 , n3460 );
buf ( n3462 , n3461 );
buf ( n3463 , n3462 );
nand ( n3464 , n3458 , n3463 );
buf ( n3465 , n3464 );
buf ( n3466 , n3465 );
nand ( n3467 , n3457 , n3466 );
buf ( n3468 , n3467 );
buf ( n3469 , n3468 );
not ( n3470 , n3469 );
buf ( n3471 , n3470 );
buf ( n3472 , n3471 );
not ( n3473 , n3472 );
or ( n3474 , n3452 , n3473 );
buf ( n3475 , n3468 );
buf ( n3476 , n3450 );
not ( n3477 , n3476 );
buf ( n3478 , n3477 );
buf ( n3479 , n3478 );
nand ( n3480 , n3475 , n3479 );
buf ( n3481 , n3480 );
buf ( n3482 , n3481 );
nand ( n3483 , n3474 , n3482 );
buf ( n3484 , n3483 );
buf ( n3485 , n3484 );
buf ( n3486 , n1987 );
not ( n3487 , n3486 );
buf ( n3488 , n850 );
not ( n3489 , n3488 );
or ( n3490 , n3487 , n3489 );
buf ( n3491 , n856 );
buf ( n3492 , n556 );
buf ( n3493 , n570 );
xor ( n3494 , n3492 , n3493 );
buf ( n3495 , n3494 );
buf ( n3496 , n3495 );
nand ( n3497 , n3491 , n3496 );
buf ( n3498 , n3497 );
buf ( n3499 , n3498 );
nand ( n3500 , n3490 , n3499 );
buf ( n3501 , n3500 );
buf ( n3502 , n3501 );
and ( n3503 , n3485 , n3502 );
not ( n3504 , n3485 );
buf ( n3505 , n3501 );
not ( n3506 , n3505 );
buf ( n3507 , n3506 );
buf ( n3508 , n3507 );
and ( n3509 , n3504 , n3508 );
nor ( n3510 , n3503 , n3509 );
buf ( n3511 , n3510 );
and ( n3512 , n3416 , n3511 );
not ( n3513 , n3416 );
not ( n3514 , n3511 );
and ( n3515 , n3513 , n3514 );
or ( n3516 , n3512 , n3515 );
buf ( n3517 , n3516 );
buf ( n3518 , n2057 );
not ( n3519 , n3518 );
not ( n3520 , n2062 );
or ( n3521 , n3519 , n3520 );
not ( n3522 , n3518 );
not ( n3523 , n3522 );
not ( n3524 , n2063 );
or ( n3525 , n3523 , n3524 );
nand ( n3526 , n3525 , n2174 );
nand ( n3527 , n3521 , n3526 );
buf ( n3528 , n3527 );
xor ( n3529 , n3517 , n3528 );
xor ( n3530 , n1994 , n1999 );
and ( n3531 , n3530 , n2036 );
and ( n3532 , n1994 , n1999 );
or ( n3533 , n3531 , n3532 );
buf ( n3534 , n3533 );
buf ( n3535 , n3534 );
not ( n3536 , n2087 );
and ( n3537 , n2083 , n3536 );
not ( n3538 , n3537 );
buf ( n3539 , n3538 );
not ( n3540 , n3539 );
buf ( n3541 , n2167 );
not ( n3542 , n3541 );
or ( n3543 , n3540 , n3542 );
buf ( n3544 , n2087 );
buf ( n3545 , n2080 );
nand ( n3546 , n3544 , n3545 );
buf ( n3547 , n3546 );
buf ( n3548 , n3547 );
nand ( n3549 , n3543 , n3548 );
buf ( n3550 , n3549 );
buf ( n3551 , n3550 );
xor ( n3552 , n3535 , n3551 );
buf ( n3553 , n559 );
buf ( n3554 , n585 );
or ( n3555 , n3553 , n3554 );
buf ( n3556 , n586 );
nand ( n3557 , n3555 , n3556 );
buf ( n3558 , n3557 );
buf ( n3559 , n3558 );
buf ( n3560 , n559 );
buf ( n3561 , n585 );
nand ( n3562 , n3560 , n3561 );
buf ( n3563 , n3562 );
buf ( n3564 , n3563 );
buf ( n3565 , n584 );
nand ( n3566 , n3559 , n3564 , n3565 );
buf ( n3567 , n3566 );
buf ( n3568 , n3567 );
not ( n3569 , n3568 );
buf ( n3570 , n2105 );
not ( n3571 , n3570 );
buf ( n3572 , n984 );
not ( n3573 , n3572 );
or ( n3574 , n3571 , n3573 );
buf ( n3575 , n552 );
buf ( n3576 , n590 );
xor ( n3577 , n3575 , n3576 );
buf ( n3578 , n3577 );
buf ( n3579 , n3578 );
buf ( n3580 , n591 );
nand ( n3581 , n3579 , n3580 );
buf ( n3582 , n3581 );
buf ( n3583 , n3582 );
nand ( n3584 , n3574 , n3583 );
buf ( n3585 , n3584 );
buf ( n3586 , n3585 );
not ( n3587 , n3586 );
or ( n3588 , n3569 , n3587 );
buf ( n3589 , n3585 );
buf ( n3590 , n3567 );
or ( n3591 , n3589 , n3590 );
nand ( n3592 , n3588 , n3591 );
buf ( n3593 , n3592 );
buf ( n3594 , n3593 );
buf ( n3595 , n2109 );
not ( n3596 , n3595 );
buf ( n3597 , n3596 );
nand ( n3598 , n3597 , n2139 );
not ( n3599 , n3598 );
not ( n3600 , n2161 );
or ( n3601 , n3599 , n3600 );
not ( n3602 , n2139 );
nand ( n3603 , n3602 , n2109 );
nand ( n3604 , n3601 , n3603 );
buf ( n3605 , n3604 );
xor ( n3606 , n3594 , n3605 );
buf ( n3607 , n2074 );
not ( n3608 , n3607 );
buf ( n3609 , n586 );
buf ( n3610 , n587 );
xnor ( n3611 , n3609 , n3610 );
buf ( n3612 , n3611 );
buf ( n3613 , n3612 );
buf ( n3614 , n1169 );
nor ( n3615 , n3613 , n3614 );
buf ( n3616 , n3615 );
buf ( n3617 , n3616 );
not ( n3618 , n3617 );
or ( n3619 , n3608 , n3618 );
buf ( n3620 , n1036 );
buf ( n3621 , n556 );
buf ( n3622 , n586 );
xor ( n3623 , n3621 , n3622 );
buf ( n3624 , n3623 );
buf ( n3625 , n3624 );
nand ( n3626 , n3620 , n3625 );
buf ( n3627 , n3626 );
buf ( n3628 , n3627 );
nand ( n3629 , n3619 , n3628 );
buf ( n3630 , n3629 );
buf ( n3631 , n3630 );
buf ( n3632 , n2155 );
not ( n3633 , n3632 );
buf ( n3634 , n1057 );
not ( n3635 , n3634 );
buf ( n3636 , n3635 );
buf ( n3637 , n3636 );
not ( n3638 , n3637 );
buf ( n3639 , n3638 );
buf ( n3640 , n3639 );
not ( n3641 , n3640 );
or ( n3642 , n3633 , n3641 );
buf ( n3643 , n1071 );
buf ( n3644 , n554 );
buf ( n3645 , n588 );
xor ( n3646 , n3644 , n3645 );
buf ( n3647 , n3646 );
buf ( n3648 , n3647 );
nand ( n3649 , n3643 , n3648 );
buf ( n3650 , n3649 );
buf ( n3651 , n3650 );
nand ( n3652 , n3642 , n3651 );
buf ( n3653 , n3652 );
buf ( n3654 , n3653 );
xor ( n3655 , n3631 , n3654 );
buf ( n3656 , n559 );
buf ( n3657 , n584 );
xor ( n3658 , n3656 , n3657 );
buf ( n3659 , n3658 );
buf ( n3660 , n3659 );
not ( n3661 , n3660 );
xor ( n3662 , n585 , n584 );
nand ( n3663 , n3662 , n2120 );
not ( n3664 , n3663 );
buf ( n3665 , n3664 );
not ( n3666 , n3665 );
or ( n3667 , n3661 , n3666 );
buf ( n3668 , n2123 );
buf ( n3669 , n558 );
buf ( n3670 , n584 );
xor ( n3671 , n3669 , n3670 );
buf ( n3672 , n3671 );
buf ( n3673 , n3672 );
nand ( n3674 , n3668 , n3673 );
buf ( n3675 , n3674 );
buf ( n3676 , n3675 );
nand ( n3677 , n3667 , n3676 );
buf ( n3678 , n3677 );
buf ( n3679 , n3678 );
xor ( n3680 , n3655 , n3679 );
buf ( n3681 , n3680 );
buf ( n3682 , n3681 );
xor ( n3683 , n3606 , n3682 );
buf ( n3684 , n3683 );
buf ( n3685 , n3684 );
xor ( n3686 , n3552 , n3685 );
buf ( n3687 , n3686 );
buf ( n3688 , n3687 );
xor ( n3689 , n3529 , n3688 );
buf ( n3690 , n3689 );
buf ( n3691 , n3690 );
not ( n3692 , n3691 );
not ( n3693 , n2175 );
not ( n3694 , n1968 );
nand ( n3695 , n3694 , n2039 );
not ( n3696 , n3695 );
or ( n3697 , n3693 , n3696 );
nand ( n3698 , n1968 , n2038 );
nand ( n3699 , n3697 , n3698 );
buf ( n3700 , n3699 );
not ( n3701 , n3700 );
buf ( n3702 , n3701 );
buf ( n3703 , n3702 );
nand ( n3704 , n3692 , n3703 );
buf ( n3705 , n3704 );
buf ( n3706 , n3705 );
buf ( n3707 , n1298 );
buf ( n3708 , n1582 );
buf ( n3709 , n1928 );
and ( n3710 , n3707 , n3708 , n3709 );
buf ( n3711 , n3710 );
buf ( n3712 , n3711 );
buf ( n3713 , n2197 );
nand ( n3714 , n3706 , n3712 , n3713 );
buf ( n3715 , n3714 );
buf ( n3716 , n3690 );
not ( n3717 , n3716 );
buf ( n3718 , n3717 );
buf ( n3719 , n3718 );
buf ( n3720 , n3702 );
nand ( n3721 , n3719 , n3720 );
buf ( n3722 , n3721 );
nand ( n3723 , n3722 , n2197 , n2205 );
buf ( n3724 , n3722 );
buf ( n3725 , n2189 );
not ( n3726 , n3725 );
buf ( n3727 , n3726 );
buf ( n3728 , n3727 );
and ( n3729 , n3724 , n3728 );
buf ( n3730 , n3690 );
buf ( n3731 , n3699 );
nand ( n3732 , n3730 , n3731 );
buf ( n3733 , n3732 );
buf ( n3734 , n3733 );
not ( n3735 , n3734 );
buf ( n3736 , n3735 );
buf ( n3737 , n3736 );
nor ( n3738 , n3729 , n3737 );
buf ( n3739 , n3738 );
nand ( n3740 , n3715 , n3723 , n3739 );
buf ( n3741 , n3740 );
not ( n3742 , n3741 );
xor ( n3743 , n567 , n568 );
buf ( n3744 , n3743 );
buf ( n3745 , n559 );
and ( n3746 , n3744 , n3745 );
buf ( n3747 , n3746 );
buf ( n3748 , n3747 );
buf ( n3749 , n3382 );
not ( n3750 , n3749 );
buf ( n3751 , n1110 );
not ( n3752 , n3751 );
or ( n3753 , n3750 , n3752 );
buf ( n3754 , n551 );
buf ( n3755 , n574 );
xor ( n3756 , n3754 , n3755 );
buf ( n3757 , n3756 );
buf ( n3758 , n3757 );
buf ( n3759 , n575 );
nand ( n3760 , n3758 , n3759 );
buf ( n3761 , n3760 );
buf ( n3762 , n3761 );
nand ( n3763 , n3753 , n3762 );
buf ( n3764 , n3763 );
buf ( n3765 , n3764 );
xor ( n3766 , n3748 , n3765 );
buf ( n3767 , n3444 );
not ( n3768 , n3767 );
buf ( n3769 , n3429 );
not ( n3770 , n3769 );
or ( n3771 , n3768 , n3770 );
xor ( n3772 , n570 , n569 );
buf ( n3773 , n3772 );
buf ( n3774 , n557 );
buf ( n3775 , n568 );
xor ( n3776 , n3774 , n3775 );
buf ( n3777 , n3776 );
buf ( n3778 , n3777 );
nand ( n3779 , n3773 , n3778 );
buf ( n3780 , n3779 );
buf ( n3781 , n3780 );
nand ( n3782 , n3771 , n3781 );
buf ( n3783 , n3782 );
buf ( n3784 , n3783 );
xor ( n3785 , n3766 , n3784 );
buf ( n3786 , n3785 );
buf ( n3787 , n3786 );
not ( n3788 , n3468 );
not ( n3789 , n3450 );
or ( n3790 , n3788 , n3789 );
not ( n3791 , n3478 );
not ( n3792 , n3471 );
or ( n3793 , n3791 , n3792 );
nand ( n3794 , n3793 , n3501 );
nand ( n3795 , n3790 , n3794 );
buf ( n3796 , n3795 );
xor ( n3797 , n3787 , n3796 );
buf ( n3798 , n3462 );
not ( n3799 , n3798 );
buf ( n3800 , n1243 );
not ( n3801 , n3800 );
or ( n3802 , n3799 , n3801 );
buf ( n3803 , n888 );
buf ( n3804 , n553 );
buf ( n3805 , n572 );
xor ( n3806 , n3804 , n3805 );
buf ( n3807 , n3806 );
buf ( n3808 , n3807 );
nand ( n3809 , n3803 , n3808 );
buf ( n3810 , n3809 );
buf ( n3811 , n3810 );
nand ( n3812 , n3802 , n3811 );
buf ( n3813 , n3812 );
buf ( n3814 , n3813 );
buf ( n3815 , n3495 );
not ( n3816 , n3815 );
buf ( n3817 , n1973 );
not ( n3818 , n3817 );
or ( n3819 , n3816 , n3818 );
buf ( n3820 , n856 );
buf ( n3821 , n555 );
buf ( n3822 , n570 );
xor ( n3823 , n3821 , n3822 );
buf ( n3824 , n3823 );
buf ( n3825 , n3824 );
nand ( n3826 , n3820 , n3825 );
buf ( n3827 , n3826 );
buf ( n3828 , n3827 );
nand ( n3829 , n3819 , n3828 );
buf ( n3830 , n3829 );
buf ( n3831 , n3830 );
xor ( n3832 , n3814 , n3831 );
buf ( n3833 , n3389 );
buf ( n3834 , n3411 );
and ( n3835 , n3833 , n3834 );
buf ( n3836 , n3835 );
buf ( n3837 , n3836 );
xor ( n3838 , n3832 , n3837 );
buf ( n3839 , n3838 );
buf ( n3840 , n3839 );
xor ( n3841 , n3797 , n3840 );
buf ( n3842 , n3841 );
not ( n3843 , n3842 );
xor ( n3844 , n3535 , n3551 );
and ( n3845 , n3844 , n3685 );
and ( n3846 , n3535 , n3551 );
or ( n3847 , n3845 , n3846 );
buf ( n3848 , n3847 );
not ( n3849 , n3848 );
not ( n3850 , n3849 );
or ( n3851 , n3843 , n3850 );
not ( n3852 , n3842 );
nand ( n3853 , n3848 , n3852 );
nand ( n3854 , n3851 , n3853 );
not ( n3855 , n3373 );
nand ( n3856 , n3855 , n3415 );
not ( n3857 , n3856 );
not ( n3858 , n3511 );
or ( n3859 , n3857 , n3858 );
buf ( n3860 , n3415 );
not ( n3861 , n3860 );
buf ( n3862 , n3373 );
nand ( n3863 , n3861 , n3862 );
buf ( n3864 , n3863 );
nand ( n3865 , n3859 , n3864 );
buf ( n3866 , n3865 );
xor ( n3867 , n3594 , n3605 );
and ( n3868 , n3867 , n3682 );
and ( n3869 , n3594 , n3605 );
or ( n3870 , n3868 , n3869 );
buf ( n3871 , n3870 );
buf ( n3872 , n3871 );
xor ( n3873 , n3866 , n3872 );
buf ( n3874 , n583 );
buf ( n3875 , n584 );
xor ( n3876 , n3874 , n3875 );
buf ( n3877 , n3876 );
buf ( n3878 , n3877 );
not ( n3879 , n3878 );
buf ( n3880 , n3879 );
buf ( n3881 , n3880 );
not ( n3882 , n3881 );
buf ( n3883 , n3882 );
buf ( n3884 , n3883 );
buf ( n3885 , n559 );
and ( n3886 , n3884 , n3885 );
buf ( n3887 , n3886 );
buf ( n3888 , n3887 );
buf ( n3889 , n3578 );
not ( n3890 , n3889 );
buf ( n3891 , n984 );
not ( n3892 , n3891 );
or ( n3893 , n3890 , n3892 );
buf ( n3894 , n551 );
buf ( n3895 , n590 );
xor ( n3896 , n3894 , n3895 );
buf ( n3897 , n3896 );
buf ( n3898 , n3897 );
buf ( n3899 , n591 );
nand ( n3900 , n3898 , n3899 );
buf ( n3901 , n3900 );
buf ( n3902 , n3901 );
nand ( n3903 , n3893 , n3902 );
buf ( n3904 , n3903 );
buf ( n3905 , n3904 );
xor ( n3906 , n3888 , n3905 );
buf ( n3907 , n3672 );
not ( n3908 , n3907 );
buf ( n3909 , n3664 );
not ( n3910 , n3909 );
or ( n3911 , n3908 , n3910 );
buf ( n3912 , n2123 );
buf ( n3913 , n557 );
buf ( n3914 , n584 );
xor ( n3915 , n3913 , n3914 );
buf ( n3916 , n3915 );
buf ( n3917 , n3916 );
nand ( n3918 , n3912 , n3917 );
buf ( n3919 , n3918 );
buf ( n3920 , n3919 );
nand ( n3921 , n3911 , n3920 );
buf ( n3922 , n3921 );
buf ( n3923 , n3922 );
xor ( n3924 , n3906 , n3923 );
buf ( n3925 , n3924 );
buf ( n3926 , n3925 );
xor ( n3927 , n3631 , n3654 );
and ( n3928 , n3927 , n3679 );
and ( n3929 , n3631 , n3654 );
or ( n3930 , n3928 , n3929 );
buf ( n3931 , n3930 );
buf ( n3932 , n3931 );
xor ( n3933 , n3926 , n3932 );
buf ( n3934 , n3624 );
not ( n3935 , n3934 );
buf ( n3936 , n1177 );
not ( n3937 , n3936 );
or ( n3938 , n3935 , n3937 );
buf ( n3939 , n1036 );
buf ( n3940 , n555 );
buf ( n3941 , n586 );
xor ( n3942 , n3940 , n3941 );
buf ( n3943 , n3942 );
buf ( n3944 , n3943 );
nand ( n3945 , n3939 , n3944 );
buf ( n3946 , n3945 );
buf ( n3947 , n3946 );
nand ( n3948 , n3938 , n3947 );
buf ( n3949 , n3948 );
buf ( n3950 , n3949 );
not ( n3951 , n3950 );
buf ( n3952 , n3951 );
buf ( n3953 , n3952 );
not ( n3954 , n3953 );
buf ( n3955 , n3647 );
not ( n3956 , n3955 );
buf ( n3957 , n1263 );
not ( n3958 , n3957 );
or ( n3959 , n3956 , n3958 );
buf ( n3960 , n1074 );
buf ( n3961 , n553 );
buf ( n3962 , n588 );
xor ( n3963 , n3961 , n3962 );
buf ( n3964 , n3963 );
buf ( n3965 , n3964 );
nand ( n3966 , n3960 , n3965 );
buf ( n3967 , n3966 );
buf ( n3968 , n3967 );
nand ( n3969 , n3959 , n3968 );
buf ( n3970 , n3969 );
buf ( n3971 , n3970 );
not ( n3972 , n3971 );
or ( n3973 , n3954 , n3972 );
buf ( n3974 , n3647 );
not ( n3975 , n3974 );
buf ( n3976 , n1263 );
not ( n3977 , n3976 );
or ( n3978 , n3975 , n3977 );
buf ( n3979 , n3967 );
nand ( n3980 , n3978 , n3979 );
buf ( n3981 , n3980 );
buf ( n3982 , n3981 );
buf ( n3983 , n3952 );
or ( n3984 , n3982 , n3983 );
nand ( n3985 , n3973 , n3984 );
buf ( n3986 , n3985 );
buf ( n3987 , n3986 );
buf ( n3988 , n3567 );
not ( n3989 , n3988 );
buf ( n3990 , n3585 );
nand ( n3991 , n3989 , n3990 );
buf ( n3992 , n3991 );
buf ( n3993 , n3992 );
not ( n3994 , n3993 );
buf ( n3995 , n3994 );
buf ( n3996 , n3995 );
xor ( n3997 , n3987 , n3996 );
buf ( n3998 , n3997 );
buf ( n3999 , n3998 );
xor ( n4000 , n3933 , n3999 );
buf ( n4001 , n4000 );
buf ( n4002 , n4001 );
xor ( n4003 , n3873 , n4002 );
buf ( n4004 , n4003 );
and ( n4005 , n3854 , n4004 );
not ( n4006 , n3854 );
not ( n4007 , n4004 );
and ( n4008 , n4006 , n4007 );
nor ( n4009 , n4005 , n4008 );
not ( n4010 , n4009 );
xor ( n4011 , n3517 , n3528 );
and ( n4012 , n4011 , n3688 );
and ( n4013 , n3517 , n3528 );
or ( n4014 , n4012 , n4013 );
buf ( n4015 , n4014 );
not ( n4016 , n4015 );
and ( n4017 , n4010 , n4016 );
buf ( n4018 , n3777 );
not ( n4019 , n4018 );
nand ( n4020 , n3423 , n3428 );
not ( n4021 , n4020 );
buf ( n4022 , n4021 );
not ( n4023 , n4022 );
or ( n4024 , n4019 , n4023 );
buf ( n4025 , n3772 );
and ( n4026 , n556 , n568 );
not ( n4027 , n556 );
and ( n4028 , n4027 , n3015 );
nor ( n4029 , n4026 , n4028 );
buf ( n4030 , n4029 );
nand ( n4031 , n4025 , n4030 );
buf ( n4032 , n4031 );
buf ( n4033 , n4032 );
nand ( n4034 , n4024 , n4033 );
buf ( n4035 , n4034 );
buf ( n4036 , n559 );
buf ( n4037 , n566 );
xor ( n4038 , n4036 , n4037 );
buf ( n4039 , n4038 );
buf ( n4040 , n4039 );
not ( n4041 , n4040 );
xor ( n4042 , n567 , n566 );
xnor ( n4043 , n567 , n568 );
and ( n4044 , n4042 , n4043 );
buf ( n4045 , n4044 );
not ( n4046 , n4045 );
or ( n4047 , n4041 , n4046 );
buf ( n4048 , n3743 );
buf ( n4049 , n558 );
buf ( n4050 , n566 );
xor ( n4051 , n4049 , n4050 );
buf ( n4052 , n4051 );
buf ( n4053 , n4052 );
nand ( n4054 , n4048 , n4053 );
buf ( n4055 , n4054 );
buf ( n4056 , n4055 );
nand ( n4057 , n4047 , n4056 );
buf ( n4058 , n4057 );
xor ( n4059 , n4035 , n4058 );
buf ( n4060 , n3757 );
not ( n4061 , n4060 );
buf ( n4062 , n1110 );
not ( n4063 , n4062 );
or ( n4064 , n4061 , n4063 );
buf ( n4065 , n550 );
buf ( n4066 , n574 );
xor ( n4067 , n4065 , n4066 );
buf ( n4068 , n4067 );
buf ( n4069 , n4068 );
buf ( n4070 , n575 );
nand ( n4071 , n4069 , n4070 );
buf ( n4072 , n4071 );
buf ( n4073 , n4072 );
nand ( n4074 , n4064 , n4073 );
buf ( n4075 , n4074 );
xor ( n4076 , n4059 , n4075 );
buf ( n4077 , n4076 );
xor ( n4078 , n3814 , n3831 );
and ( n4079 , n4078 , n3837 );
and ( n4080 , n3814 , n3831 );
or ( n4081 , n4079 , n4080 );
buf ( n4082 , n4081 );
buf ( n4083 , n4082 );
xor ( n4084 , n4077 , n4083 );
buf ( n4085 , n3824 );
not ( n4086 , n4085 );
buf ( n4087 , n1973 );
not ( n4088 , n4087 );
or ( n4089 , n4086 , n4088 );
buf ( n4090 , n1982 );
buf ( n4091 , n554 );
buf ( n4092 , n570 );
xor ( n4093 , n4091 , n4092 );
buf ( n4094 , n4093 );
buf ( n4095 , n4094 );
nand ( n4096 , n4090 , n4095 );
buf ( n4097 , n4096 );
buf ( n4098 , n4097 );
nand ( n4099 , n4089 , n4098 );
buf ( n4100 , n4099 );
buf ( n4101 , n4100 );
not ( n4102 , n3807 );
not ( n4103 , n1243 );
or ( n4104 , n4102 , n4103 );
buf ( n4105 , n888 );
buf ( n4106 , n552 );
buf ( n4107 , n572 );
xor ( n4108 , n4106 , n4107 );
buf ( n4109 , n4108 );
buf ( n4110 , n4109 );
nand ( n4111 , n4105 , n4110 );
buf ( n4112 , n4111 );
nand ( n4113 , n4104 , n4112 );
buf ( n4114 , n559 );
buf ( n4115 , n567 );
nand ( n4116 , n4114 , n4115 );
buf ( n4117 , n4116 );
or ( n4118 , n559 , n567 );
nand ( n4119 , n4118 , n568 );
nand ( n4120 , n4117 , n4119 , n566 );
and ( n4121 , n4113 , n4120 );
not ( n4122 , n4113 );
not ( n4123 , n4120 );
and ( n4124 , n4122 , n4123 );
or ( n4125 , n4121 , n4124 );
buf ( n4126 , n4125 );
xor ( n4127 , n4101 , n4126 );
xor ( n4128 , n3748 , n3765 );
and ( n4129 , n4128 , n3784 );
and ( n4130 , n3748 , n3765 );
or ( n4131 , n4129 , n4130 );
buf ( n4132 , n4131 );
buf ( n4133 , n4132 );
xor ( n4134 , n4127 , n4133 );
buf ( n4135 , n4134 );
buf ( n4136 , n4135 );
xor ( n4137 , n4084 , n4136 );
buf ( n4138 , n4137 );
buf ( n4139 , n4138 );
xor ( n4140 , n3866 , n3872 );
and ( n4141 , n4140 , n4002 );
and ( n4142 , n3866 , n3872 );
or ( n4143 , n4141 , n4142 );
buf ( n4144 , n4143 );
buf ( n4145 , n4144 );
xor ( n4146 , n4139 , n4145 );
xor ( n4147 , n3787 , n3796 );
and ( n4148 , n4147 , n3840 );
and ( n4149 , n3787 , n3796 );
or ( n4150 , n4148 , n4149 );
buf ( n4151 , n4150 );
buf ( n4152 , n4151 );
xor ( n4153 , n3926 , n3932 );
and ( n4154 , n4153 , n3999 );
and ( n4155 , n3926 , n3932 );
or ( n4156 , n4154 , n4155 );
buf ( n4157 , n4156 );
buf ( n4158 , n4157 );
xor ( n4159 , n4152 , n4158 );
buf ( n4160 , n3952 );
not ( n4161 , n4160 );
buf ( n4162 , n3992 );
not ( n4163 , n4162 );
or ( n4164 , n4161 , n4163 );
buf ( n4165 , n3981 );
nand ( n4166 , n4164 , n4165 );
buf ( n4167 , n4166 );
buf ( n4168 , n4167 );
buf ( n4169 , n3995 );
buf ( n4170 , n3949 );
nand ( n4171 , n4169 , n4170 );
buf ( n4172 , n4171 );
buf ( n4173 , n4172 );
nand ( n4174 , n4168 , n4173 );
buf ( n4175 , n4174 );
buf ( n4176 , n4175 );
buf ( n4177 , n3897 );
not ( n4178 , n4177 );
buf ( n4179 , n984 );
not ( n4180 , n4179 );
or ( n4181 , n4178 , n4180 );
buf ( n4182 , n550 );
buf ( n4183 , n590 );
xor ( n4184 , n4182 , n4183 );
buf ( n4185 , n4184 );
buf ( n4186 , n4185 );
buf ( n4187 , n591 );
nand ( n4188 , n4186 , n4187 );
buf ( n4189 , n4188 );
buf ( n4190 , n4189 );
nand ( n4191 , n4181 , n4190 );
buf ( n4192 , n4191 );
buf ( n4193 , n4192 );
buf ( n4194 , n559 );
buf ( n4195 , n582 );
xor ( n4196 , n4194 , n4195 );
buf ( n4197 , n4196 );
buf ( n4198 , n4197 );
not ( n4199 , n4198 );
xnor ( n4200 , n583 , n584 );
xor ( n4201 , n583 , n582 );
nand ( n4202 , n4200 , n4201 );
buf ( n4203 , n4202 );
not ( n4204 , n4203 );
buf ( n4205 , n4204 );
buf ( n4206 , n4205 );
not ( n4207 , n4206 );
or ( n4208 , n4199 , n4207 );
buf ( n4209 , n3877 );
buf ( n4210 , n4209 );
buf ( n4211 , n4210 );
buf ( n4212 , n4211 );
buf ( n4213 , n558 );
buf ( n4214 , n582 );
xor ( n4215 , n4213 , n4214 );
buf ( n4216 , n4215 );
buf ( n4217 , n4216 );
nand ( n4218 , n4212 , n4217 );
buf ( n4219 , n4218 );
buf ( n4220 , n4219 );
nand ( n4221 , n4208 , n4220 );
buf ( n4222 , n4221 );
buf ( n4223 , n4222 );
xor ( n4224 , n4193 , n4223 );
buf ( n4225 , n3916 );
not ( n4226 , n4225 );
buf ( n4227 , n3664 );
not ( n4228 , n4227 );
or ( n4229 , n4226 , n4228 );
buf ( n4230 , n2132 );
not ( n4231 , n4230 );
buf ( n4232 , n4231 );
buf ( n4233 , n4232 );
buf ( n4234 , n556 );
buf ( n4235 , n584 );
xor ( n4236 , n4234 , n4235 );
buf ( n4237 , n4236 );
buf ( n4238 , n4237 );
nand ( n4239 , n4233 , n4238 );
buf ( n4240 , n4239 );
buf ( n4241 , n4240 );
nand ( n4242 , n4229 , n4241 );
buf ( n4243 , n4242 );
buf ( n4244 , n4243 );
xor ( n4245 , n4224 , n4244 );
buf ( n4246 , n4245 );
buf ( n4247 , n4246 );
xor ( n4248 , n4176 , n4247 );
buf ( n4249 , n3943 );
not ( n4250 , n4249 );
buf ( n4251 , n1177 );
not ( n4252 , n4251 );
or ( n4253 , n4250 , n4252 );
buf ( n4254 , n1036 );
and ( n4255 , n586 , n554 );
not ( n4256 , n586 );
not ( n4257 , n554 );
and ( n4258 , n4256 , n4257 );
nor ( n4259 , n4255 , n4258 );
buf ( n4260 , n4259 );
nand ( n4261 , n4254 , n4260 );
buf ( n4262 , n4261 );
buf ( n4263 , n4262 );
nand ( n4264 , n4253 , n4263 );
buf ( n4265 , n4264 );
buf ( n4266 , n4265 );
buf ( n4267 , n559 );
buf ( n4268 , n583 );
or ( n4269 , n4267 , n4268 );
buf ( n4270 , n584 );
nand ( n4271 , n4269 , n4270 );
buf ( n4272 , n4271 );
buf ( n4273 , n4272 );
buf ( n4274 , n559 );
buf ( n4275 , n583 );
nand ( n4276 , n4274 , n4275 );
buf ( n4277 , n4276 );
buf ( n4278 , n4277 );
buf ( n4279 , n582 );
and ( n4280 , n4273 , n4278 , n4279 );
buf ( n4281 , n4280 );
buf ( n4282 , n3964 );
not ( n4283 , n4282 );
not ( n4284 , n590 );
nand ( n4285 , n4284 , n589 );
and ( n4286 , n1049 , n1054 , n4285 );
buf ( n4287 , n4286 );
not ( n4288 , n4287 );
or ( n4289 , n4283 , n4288 );
buf ( n4290 , n1071 );
buf ( n4291 , n552 );
buf ( n4292 , n588 );
xor ( n4293 , n4291 , n4292 );
buf ( n4294 , n4293 );
buf ( n4295 , n4294 );
nand ( n4296 , n4290 , n4295 );
buf ( n4297 , n4296 );
buf ( n4298 , n4297 );
nand ( n4299 , n4289 , n4298 );
buf ( n4300 , n4299 );
xor ( n4301 , n4281 , n4300 );
buf ( n4302 , n4301 );
xor ( n4303 , n4266 , n4302 );
xor ( n4304 , n3888 , n3905 );
and ( n4305 , n4304 , n3923 );
and ( n4306 , n3888 , n3905 );
or ( n4307 , n4305 , n4306 );
buf ( n4308 , n4307 );
buf ( n4309 , n4308 );
xor ( n4310 , n4303 , n4309 );
buf ( n4311 , n4310 );
buf ( n4312 , n4311 );
xor ( n4313 , n4248 , n4312 );
buf ( n4314 , n4313 );
buf ( n4315 , n4314 );
xor ( n4316 , n4159 , n4315 );
buf ( n4317 , n4316 );
buf ( n4318 , n4317 );
xor ( n4319 , n4146 , n4318 );
buf ( n4320 , n4319 );
buf ( n4321 , n4320 );
nand ( n4322 , n3852 , n3849 );
not ( n4323 , n4322 );
not ( n4324 , n4004 );
or ( n4325 , n4323 , n4324 );
nand ( n4326 , n3842 , n3848 );
nand ( n4327 , n4325 , n4326 );
buf ( n4328 , n4327 );
nor ( n4329 , n4321 , n4328 );
buf ( n4330 , n4329 );
nor ( n4331 , n4017 , n4330 );
not ( n4332 , n4331 );
or ( n4333 , n3742 , n4332 );
buf ( n4334 , n4009 );
buf ( n4335 , n4015 );
nand ( n4336 , n4334 , n4335 );
buf ( n4337 , n4336 );
buf ( n4338 , n4337 );
buf ( n4339 , n4330 );
or ( n4340 , n4338 , n4339 );
buf ( n4341 , n4320 );
buf ( n4342 , n4327 );
nand ( n4343 , n4341 , n4342 );
buf ( n4344 , n4343 );
buf ( n4345 , n4344 );
nand ( n4346 , n4340 , n4345 );
buf ( n4347 , n4346 );
buf ( n4348 , n4347 );
not ( n4349 , n4348 );
buf ( n4350 , n4349 );
nand ( n4351 , n4333 , n4350 );
xor ( n4352 , n4139 , n4145 );
and ( n4353 , n4352 , n4318 );
and ( n4354 , n4139 , n4145 );
or ( n4355 , n4353 , n4354 );
buf ( n4356 , n4355 );
not ( n4357 , n4356 );
buf ( n4358 , n4068 );
not ( n4359 , n4358 );
buf ( n4360 , n1110 );
not ( n4361 , n4360 );
or ( n4362 , n4359 , n4361 );
and ( n4363 , n574 , n549 );
not ( n4364 , n574 );
not ( n4365 , n549 );
and ( n4366 , n4364 , n4365 );
nor ( n4367 , n4363 , n4366 );
buf ( n4368 , n4367 );
buf ( n4369 , n575 );
nand ( n4370 , n4368 , n4369 );
buf ( n4371 , n4370 );
buf ( n4372 , n4371 );
nand ( n4373 , n4362 , n4372 );
buf ( n4374 , n4373 );
buf ( n4375 , n4052 );
not ( n4376 , n4375 );
nand ( n4377 , n4043 , n4042 );
buf ( n4378 , n4377 );
not ( n4379 , n4378 );
buf ( n4380 , n4379 );
buf ( n4381 , n4380 );
not ( n4382 , n4381 );
or ( n4383 , n4376 , n4382 );
not ( n4384 , n4043 );
xor ( n4385 , n566 , n557 );
nand ( n4386 , n4384 , n4385 );
buf ( n4387 , n4386 );
nand ( n4388 , n4383 , n4387 );
buf ( n4389 , n4388 );
xor ( n4390 , n4374 , n4389 );
buf ( n4391 , n4094 );
not ( n4392 , n4391 );
buf ( n4393 , n850 );
not ( n4394 , n4393 );
or ( n4395 , n4392 , n4394 );
buf ( n4396 , n856 );
buf ( n4397 , n553 );
buf ( n4398 , n570 );
xor ( n4399 , n4397 , n4398 );
buf ( n4400 , n4399 );
buf ( n4401 , n4400 );
nand ( n4402 , n4396 , n4401 );
buf ( n4403 , n4402 );
buf ( n4404 , n4403 );
nand ( n4405 , n4395 , n4404 );
buf ( n4406 , n4405 );
xor ( n4407 , n4390 , n4406 );
buf ( n4408 , n4407 );
xor ( n4409 , n4101 , n4126 );
and ( n4410 , n4409 , n4133 );
and ( n4411 , n4101 , n4126 );
or ( n4412 , n4410 , n4411 );
buf ( n4413 , n4412 );
buf ( n4414 , n4413 );
xor ( n4415 , n4408 , n4414 );
nand ( n4416 , n4113 , n4123 );
not ( n4417 , n4075 );
not ( n4418 , n4035 );
or ( n4419 , n4417 , n4418 );
buf ( n4420 , n4075 );
buf ( n4421 , n4035 );
or ( n4422 , n4420 , n4421 );
buf ( n4423 , n4058 );
nand ( n4424 , n4422 , n4423 );
buf ( n4425 , n4424 );
nand ( n4426 , n4419 , n4425 );
xor ( n4427 , n4416 , n4426 );
xor ( n4428 , n565 , n566 );
buf ( n4429 , n4428 );
buf ( n4430 , n559 );
and ( n4431 , n4429 , n4430 );
buf ( n4432 , n4431 );
not ( n4433 , n4109 );
nand ( n4434 , n875 , n878 );
and ( n4435 , n882 , n4434 );
not ( n4436 , n4435 );
or ( n4437 , n4433 , n4436 );
buf ( n4438 , n551 );
buf ( n4439 , n572 );
xor ( n4440 , n4438 , n4439 );
buf ( n4441 , n4440 );
nand ( n4442 , n888 , n4441 );
nand ( n4443 , n4437 , n4442 );
xor ( n4444 , n4432 , n4443 );
not ( n4445 , n4029 );
not ( n4446 , n3429 );
or ( n4447 , n4445 , n4446 );
buf ( n4448 , n3772 );
buf ( n4449 , n555 );
buf ( n4450 , n568 );
xor ( n4451 , n4449 , n4450 );
buf ( n4452 , n4451 );
buf ( n4453 , n4452 );
nand ( n4454 , n4448 , n4453 );
buf ( n4455 , n4454 );
nand ( n4456 , n4447 , n4455 );
xnor ( n4457 , n4444 , n4456 );
buf ( n4458 , n4457 );
not ( n4459 , n4458 );
buf ( n4460 , n4459 );
xnor ( n4461 , n4427 , n4460 );
buf ( n4462 , n4461 );
xor ( n4463 , n4415 , n4462 );
buf ( n4464 , n4463 );
buf ( n4465 , n4464 );
xor ( n4466 , n4152 , n4158 );
and ( n4467 , n4466 , n4315 );
and ( n4468 , n4152 , n4158 );
or ( n4469 , n4467 , n4468 );
buf ( n4470 , n4469 );
buf ( n4471 , n4470 );
xor ( n4472 , n4465 , n4471 );
xor ( n4473 , n4077 , n4083 );
and ( n4474 , n4473 , n4136 );
and ( n4475 , n4077 , n4083 );
or ( n4476 , n4474 , n4475 );
buf ( n4477 , n4476 );
buf ( n4478 , n4477 );
xor ( n4479 , n4176 , n4247 );
and ( n4480 , n4479 , n4312 );
and ( n4481 , n4176 , n4247 );
or ( n4482 , n4480 , n4481 );
buf ( n4483 , n4482 );
buf ( n4484 , n4483 );
xor ( n4485 , n4478 , n4484 );
xor ( n4486 , n586 , n553 );
not ( n4487 , n4486 );
not ( n4488 , n1036 );
or ( n4489 , n4487 , n4488 );
nand ( n4490 , n1170 , n1175 , n4259 );
nand ( n4491 , n4489 , n4490 );
not ( n4492 , n984 );
not ( n4493 , n4185 );
or ( n4494 , n4492 , n4493 );
and ( n4495 , n590 , n549 );
not ( n4496 , n590 );
and ( n4497 , n4496 , n4365 );
nor ( n4498 , n4495 , n4497 );
buf ( n4499 , n4498 );
buf ( n4500 , n591 );
nand ( n4501 , n4499 , n4500 );
buf ( n4502 , n4501 );
nand ( n4503 , n4494 , n4502 );
nor ( n4504 , n4491 , n4503 );
nand ( n4505 , n4201 , n3880 );
not ( n4506 , n4505 );
nand ( n4507 , n4216 , n4506 );
buf ( n4508 , n4211 );
buf ( n4509 , n557 );
buf ( n4510 , n582 );
xor ( n4511 , n4509 , n4510 );
buf ( n4512 , n4511 );
buf ( n4513 , n4512 );
nand ( n4514 , n4508 , n4513 );
buf ( n4515 , n4514 );
and ( n4516 , n4507 , n4515 );
not ( n4517 , n4516 );
nand ( n4518 , n4504 , n4517 );
nand ( n4519 , n4517 , n4491 , n4503 );
not ( n4520 , n4503 );
nand ( n4521 , n4516 , n4491 , n4520 );
not ( n4522 , n4491 );
nand ( n4523 , n4516 , n4522 , n4503 );
nand ( n4524 , n4518 , n4519 , n4521 , n4523 );
buf ( n4525 , n4524 );
xor ( n4526 , n4266 , n4302 );
and ( n4527 , n4526 , n4309 );
and ( n4528 , n4266 , n4302 );
or ( n4529 , n4527 , n4528 );
buf ( n4530 , n4529 );
buf ( n4531 , n4530 );
xor ( n4532 , n4525 , n4531 );
buf ( n4533 , n4300 );
buf ( n4534 , n4281 );
and ( n4535 , n4533 , n4534 );
buf ( n4536 , n4535 );
buf ( n4537 , n4536 );
xor ( n4538 , n581 , n582 );
buf ( n4539 , n4538 );
not ( n4540 , n4539 );
buf ( n4541 , n4540 );
buf ( n4542 , n4541 );
not ( n4543 , n4542 );
buf ( n4544 , n4543 );
buf ( n4545 , n4544 );
buf ( n4546 , n559 );
and ( n4547 , n4545 , n4546 );
buf ( n4548 , n4547 );
buf ( n4549 , n4294 );
not ( n4550 , n4549 );
buf ( n4551 , n4286 );
not ( n4552 , n4551 );
or ( n4553 , n4550 , n4552 );
nand ( n4554 , n1643 , n590 );
nand ( n4555 , n4284 , n589 );
nand ( n4556 , n4554 , n4555 );
buf ( n4557 , n551 );
buf ( n4558 , n588 );
xor ( n4559 , n4557 , n4558 );
buf ( n4560 , n4559 );
nand ( n4561 , n4556 , n4560 );
buf ( n4562 , n4561 );
nand ( n4563 , n4553 , n4562 );
buf ( n4564 , n4563 );
xor ( n4565 , n4548 , n4564 );
buf ( n4566 , n4237 );
not ( n4567 , n4566 );
buf ( n4568 , n3664 );
not ( n4569 , n4568 );
or ( n4570 , n4567 , n4569 );
buf ( n4571 , n4232 );
buf ( n4572 , n555 );
buf ( n4573 , n584 );
xor ( n4574 , n4572 , n4573 );
buf ( n4575 , n4574 );
buf ( n4576 , n4575 );
nand ( n4577 , n4571 , n4576 );
buf ( n4578 , n4577 );
buf ( n4579 , n4578 );
nand ( n4580 , n4570 , n4579 );
buf ( n4581 , n4580 );
xor ( n4582 , n4565 , n4581 );
buf ( n4583 , n4582 );
xor ( n4584 , n4537 , n4583 );
xor ( n4585 , n4193 , n4223 );
and ( n4586 , n4585 , n4244 );
and ( n4587 , n4193 , n4223 );
or ( n4588 , n4586 , n4587 );
buf ( n4589 , n4588 );
buf ( n4590 , n4589 );
xor ( n4591 , n4584 , n4590 );
buf ( n4592 , n4591 );
buf ( n4593 , n4592 );
xor ( n4594 , n4532 , n4593 );
buf ( n4595 , n4594 );
buf ( n4596 , n4595 );
xor ( n4597 , n4485 , n4596 );
buf ( n4598 , n4597 );
buf ( n4599 , n4598 );
xor ( n4600 , n4472 , n4599 );
buf ( n4601 , n4600 );
not ( n4602 , n4601 );
or ( n4603 , n4357 , n4602 );
buf ( n4604 , n4601 );
not ( n4605 , n4604 );
buf ( n4606 , n4605 );
buf ( n4607 , n4356 );
not ( n4608 , n4607 );
buf ( n4609 , n4608 );
nand ( n4610 , n4606 , n4609 );
nand ( n4611 , n4603 , n4610 );
and ( n4612 , n4351 , n4611 );
not ( n4613 , n4351 );
not ( n4614 , n4611 );
and ( n4615 , n4613 , n4614 );
nor ( n4616 , n4612 , n4615 );
not ( n4617 , n4616 );
nand ( n4618 , n3369 , n4617 );
nand ( n4619 , n3368 , n4616 );
nand ( n4620 , n4618 , n4619 );
or ( n4621 , n1951 , n1961 );
buf ( n4622 , n2180 );
not ( n4623 , n4622 );
buf ( n4624 , n2196 );
nand ( n4625 , n4623 , n4624 );
buf ( n4626 , n4625 );
nand ( n4627 , n4626 , n2205 );
buf ( n4628 , n2180 );
not ( n4629 , n4628 );
buf ( n4630 , n2196 );
nand ( n4631 , n4629 , n4630 );
buf ( n4632 , n4631 );
buf ( n4633 , n2203 );
buf ( n4634 , n1368 );
nor ( n4635 , n4633 , n4634 );
buf ( n4636 , n4635 );
nand ( n4637 , n4632 , n4636 , n1582 );
nand ( n4638 , n4627 , n4637 , n2192 );
not ( n4639 , n3736 );
nand ( n4640 , n4639 , n3705 );
not ( n4641 , n4640 );
and ( n4642 , n4638 , n4641 );
not ( n4643 , n4638 );
and ( n4644 , n4643 , n4640 );
nor ( n4645 , n4642 , n4644 );
not ( n4646 , n4645 );
not ( n4647 , n3359 );
nand ( n4648 , n4647 , n3346 );
nand ( n4649 , n4648 , n3360 );
buf ( n4650 , n3356 );
and ( n4651 , n4649 , n4650 );
not ( n4652 , n4649 );
not ( n4653 , n4650 );
and ( n4654 , n4652 , n4653 );
nor ( n4655 , n4651 , n4654 );
not ( n4656 , n4655 );
nand ( n4657 , n4646 , n4656 );
nand ( n4658 , n4621 , n4657 , n2305 );
nand ( n4659 , n4645 , n4655 );
not ( n4660 , n4659 );
not ( n4661 , n4645 );
and ( n4662 , n4661 , n4656 );
nor ( n4663 , n4662 , n2307 );
nor ( n4664 , n4660 , n4663 );
nand ( n4665 , n4658 , n4664 );
buf ( n4666 , n4665 );
not ( n4667 , n4666 );
and ( n4668 , n3332 , n3333 );
not ( n4669 , n3332 );
and ( n4670 , n4669 , n3306 );
or ( n4671 , n4668 , n4670 );
not ( n4672 , n4671 );
not ( n4673 , n3313 );
nand ( n4674 , n4673 , n3363 );
not ( n4675 , n4674 );
buf ( n4676 , n3361 );
not ( n4677 , n4676 );
or ( n4678 , n4675 , n4677 );
nand ( n4679 , n3313 , n3328 );
nand ( n4680 , n4678 , n4679 );
not ( n4681 , n4680 );
or ( n4682 , n4672 , n4681 );
or ( n4683 , n4671 , n4680 );
nand ( n4684 , n4682 , n4683 );
buf ( n4685 , n4320 );
not ( n4686 , n4685 );
buf ( n4687 , n4327 );
not ( n4688 , n4687 );
buf ( n4689 , n4688 );
buf ( n4690 , n4689 );
nand ( n4691 , n4686 , n4690 );
buf ( n4692 , n4691 );
nand ( n4693 , n4344 , n4692 );
not ( n4694 , n4693 );
not ( n4695 , n4015 );
not ( n4696 , n4009 );
nand ( n4697 , n4695 , n4696 );
not ( n4698 , n4697 );
not ( n4699 , n3740 );
or ( n4700 , n4698 , n4699 );
nand ( n4701 , n4700 , n4337 );
not ( n4702 , n4701 );
and ( n4703 , n4694 , n4702 );
and ( n4704 , n4693 , n4701 );
nor ( n4705 , n4703 , n4704 );
nand ( n4706 , n4684 , n4705 );
buf ( n4707 , n3741 );
buf ( n4708 , n4697 );
buf ( n4709 , n4337 );
and ( n4710 , n4708 , n4709 );
buf ( n4711 , n4710 );
buf ( n4712 , n4711 );
xor ( n4713 , n4707 , n4712 );
buf ( n4714 , n4713 );
not ( n4715 , n4714 );
nand ( n4716 , n4674 , n4679 );
not ( n4717 , n4716 );
not ( n4718 , n4676 );
or ( n4719 , n4717 , n4718 );
or ( n4720 , n4676 , n4716 );
nand ( n4721 , n4719 , n4720 );
nand ( n4722 , n4715 , n4721 );
and ( n4723 , n4706 , n4722 );
not ( n4724 , n4723 );
or ( n4725 , n4667 , n4724 );
not ( n4726 , n4721 );
nand ( n4727 , n4726 , n4714 );
not ( n4728 , n4727 );
not ( n4729 , n4728 );
not ( n4730 , n4706 );
or ( n4731 , n4729 , n4730 );
not ( n4732 , n4684 );
not ( n4733 , n4705 );
nand ( n4734 , n4732 , n4733 );
nand ( n4735 , n4731 , n4734 );
not ( n4736 , n4735 );
nand ( n4737 , n4725 , n4736 );
xor ( n4738 , n4620 , n4737 );
not ( n4739 , n581 );
nand ( n4740 , n4738 , n4739 );
nand ( n4741 , C1 , n2352 );
nand ( n4742 , n2305 , n1961 );
nand ( n4743 , n2305 , n1951 );
nand ( n4744 , n4742 , n4743 , n2307 );
and ( n4745 , n4657 , n4659 );
and ( n4746 , n4744 , n4745 );
not ( n4747 , n4744 );
not ( n4748 , n4745 );
and ( n4749 , n4747 , n4748 );
nor ( n4750 , n4746 , n4749 );
not ( n4751 , n4750 );
nand ( n4752 , n4751 , n3013 );
nand ( n4753 , n4741 , n4752 , n2318 );
not ( n4754 , n4751 );
nand ( n4755 , n4754 , n584 );
not ( n4756 , n2315 );
nand ( n4757 , n4756 , n4752 );
nand ( n4758 , n4753 , n4755 , n4757 );
and ( n4759 , n4722 , n4727 );
and ( n4760 , n4759 , n4666 );
not ( n4761 , n4759 );
not ( n4762 , n4666 );
and ( n4763 , n4761 , n4762 );
nor ( n4764 , n4760 , n4763 );
not ( n4765 , n4764 );
not ( n4766 , n583 );
and ( n4767 , n4765 , n4766 );
not ( n4768 , n4722 );
not ( n4769 , n4665 );
or ( n4770 , n4768 , n4769 );
nand ( n4771 , n4770 , n4727 );
not ( n4772 , n4771 );
nand ( n4773 , n4706 , n4734 );
not ( n4774 , n4773 );
nand ( n4775 , n4772 , n4774 );
nand ( n4776 , n4771 , n4773 );
not ( n4777 , n582 );
and ( n4778 , n4775 , n4776 , n4777 );
nor ( n4779 , n4767 , n4778 );
nand ( n4780 , n4740 , n4758 , n4779 );
buf ( n4781 , n583 );
not ( n4782 , n4781 );
buf ( n4783 , n4782 );
not ( n4784 , n4783 );
nand ( n4785 , n4784 , n4764 );
or ( n4786 , n4778 , n4785 );
not ( n4787 , n4776 );
not ( n4788 , n4775 );
or ( n4789 , n4787 , n4788 );
nand ( n4790 , n4789 , n582 );
nand ( n4791 , n4786 , n4790 );
nand ( n4792 , n4791 , n4740 );
not ( n4793 , n4738 );
nand ( n4794 , n4793 , n581 );
nand ( n4795 , n4780 , n4792 , n4794 );
nand ( n4796 , n4735 , n4619 );
nand ( n4797 , n4616 , n3368 );
nand ( n4798 , n4723 , n4797 , n4666 );
nand ( n4799 , n4796 , n4798 , n4618 );
not ( n4800 , n4799 );
buf ( n4801 , n4692 );
buf ( n4802 , n4697 );
nand ( n4803 , n4801 , n4802 );
buf ( n4804 , n4803 );
buf ( n4805 , n4804 );
buf ( n4806 , n4601 );
buf ( n4807 , n4356 );
nor ( n4808 , n4806 , n4807 );
buf ( n4809 , n4808 );
buf ( n4810 , n4809 );
nor ( n4811 , n4805 , n4810 );
buf ( n4812 , n4811 );
not ( n4813 , n4812 );
not ( n4814 , n3741 );
or ( n4815 , n4813 , n4814 );
and ( n4816 , n4347 , n4610 );
and ( n4817 , n4601 , n4356 );
nor ( n4818 , n4816 , n4817 );
nand ( n4819 , n4815 , n4818 );
buf ( n4820 , n559 );
buf ( n4821 , n564 );
xor ( n4822 , n4820 , n4821 );
buf ( n4823 , n4822 );
buf ( n4824 , n4823 );
not ( n4825 , n4824 );
buf ( n4826 , n4428 );
not ( n4827 , n4826 );
buf ( n4828 , n4827 );
buf ( n4829 , n4828 );
xor ( n4830 , n564 , n565 );
buf ( n4831 , n4830 );
nand ( n4832 , n4829 , n4831 );
buf ( n4833 , n4832 );
buf ( n4834 , n4833 );
not ( n4835 , n4834 );
buf ( n4836 , n4835 );
buf ( n4837 , n4836 );
not ( n4838 , n4837 );
or ( n4839 , n4825 , n4838 );
buf ( n4840 , n4428 );
buf ( n4841 , n4840 );
buf ( n4842 , n558 );
buf ( n4843 , n564 );
xor ( n4844 , n4842 , n4843 );
buf ( n4845 , n4844 );
buf ( n4846 , n4845 );
nand ( n4847 , n4841 , n4846 );
buf ( n4848 , n4847 );
buf ( n4849 , n4848 );
nand ( n4850 , n4839 , n4849 );
buf ( n4851 , n4850 );
buf ( n4852 , n4851 );
buf ( n4853 , n4400 );
not ( n4854 , n4853 );
buf ( n4855 , n1973 );
not ( n4856 , n4855 );
or ( n4857 , n4854 , n4856 );
buf ( n4858 , n1982 );
buf ( n4859 , n552 );
buf ( n4860 , n570 );
xor ( n4861 , n4859 , n4860 );
buf ( n4862 , n4861 );
buf ( n4863 , n4862 );
nand ( n4864 , n4858 , n4863 );
buf ( n4865 , n4864 );
buf ( n4866 , n4865 );
nand ( n4867 , n4857 , n4866 );
buf ( n4868 , n4867 );
buf ( n4869 , n4868 );
xor ( n4870 , n4852 , n4869 );
buf ( n4871 , n559 );
buf ( n4872 , n565 );
or ( n4873 , n4871 , n4872 );
buf ( n4874 , n566 );
nand ( n4875 , n4873 , n4874 );
buf ( n4876 , n4875 );
buf ( n4877 , n4876 );
buf ( n4878 , n559 );
buf ( n4879 , n565 );
nand ( n4880 , n4878 , n4879 );
buf ( n4881 , n4880 );
buf ( n4882 , n4881 );
buf ( n4883 , n564 );
and ( n4884 , n4877 , n4882 , n4883 );
buf ( n4885 , n4884 );
buf ( n4886 , n4885 );
buf ( n4887 , n4441 );
not ( n4888 , n4887 );
buf ( n4889 , n884 );
not ( n4890 , n4889 );
or ( n4891 , n4888 , n4890 );
buf ( n4892 , n888 );
xor ( n4893 , n572 , n550 );
buf ( n4894 , n4893 );
nand ( n4895 , n4892 , n4894 );
buf ( n4896 , n4895 );
buf ( n4897 , n4896 );
nand ( n4898 , n4891 , n4897 );
buf ( n4899 , n4898 );
buf ( n4900 , n4899 );
xor ( n4901 , n4886 , n4900 );
buf ( n4902 , n4901 );
buf ( n4903 , n4902 );
xor ( n4904 , n4870 , n4903 );
buf ( n4905 , n4904 );
buf ( n4906 , n4905 );
not ( n4907 , n4416 );
not ( n4908 , n4907 );
not ( n4909 , n4460 );
or ( n4910 , n4908 , n4909 );
not ( n4911 , n4416 );
not ( n4912 , n4457 );
or ( n4913 , n4911 , n4912 );
nand ( n4914 , n4913 , n4426 );
nand ( n4915 , n4910 , n4914 );
buf ( n4916 , n4915 );
xor ( n4917 , n4906 , n4916 );
buf ( n4918 , n4374 );
not ( n4919 , n4918 );
buf ( n4920 , n4389 );
not ( n4921 , n4920 );
or ( n4922 , n4919 , n4921 );
buf ( n4923 , n4389 );
buf ( n4924 , n4374 );
or ( n4925 , n4923 , n4924 );
buf ( n4926 , n4406 );
nand ( n4927 , n4925 , n4926 );
buf ( n4928 , n4927 );
buf ( n4929 , n4928 );
nand ( n4930 , n4922 , n4929 );
buf ( n4931 , n4930 );
buf ( n4932 , n4931 );
buf ( n4933 , n4432 );
not ( n4934 , n4933 );
buf ( n4935 , n4443 );
not ( n4936 , n4935 );
or ( n4937 , n4934 , n4936 );
or ( n4938 , n4443 , n4432 );
nand ( n4939 , n4938 , n4456 );
buf ( n4940 , n4939 );
nand ( n4941 , n4937 , n4940 );
buf ( n4942 , n4941 );
buf ( n4943 , n4942 );
xor ( n4944 , n4932 , n4943 );
not ( n4945 , n575 );
buf ( n4946 , n548 );
buf ( n4947 , n574 );
xor ( n4948 , n4946 , n4947 );
buf ( n4949 , n4948 );
not ( n4950 , n4949 );
or ( n4951 , n4945 , n4950 );
not ( n4952 , n574 );
nor ( n4953 , n4952 , n575 );
nand ( n4954 , n4953 , n4367 );
nand ( n4955 , n4951 , n4954 );
buf ( n4956 , n4955 );
not ( n4957 , n4452 );
not ( n4958 , n4020 );
not ( n4959 , n4958 );
or ( n4960 , n4957 , n4959 );
buf ( n4961 , n2001 );
buf ( n4962 , n554 );
buf ( n4963 , n568 );
xor ( n4964 , n4962 , n4963 );
buf ( n4965 , n4964 );
buf ( n4966 , n4965 );
nand ( n4967 , n4961 , n4966 );
buf ( n4968 , n4967 );
nand ( n4969 , n4960 , n4968 );
buf ( n4970 , n4969 );
xor ( n4971 , n4956 , n4970 );
buf ( n4972 , n4385 );
not ( n4973 , n4972 );
buf ( n4974 , n4380 );
not ( n4975 , n4974 );
or ( n4976 , n4973 , n4975 );
buf ( n4977 , n3743 );
xor ( n4978 , n566 , n556 );
buf ( n4979 , n4978 );
nand ( n4980 , n4977 , n4979 );
buf ( n4981 , n4980 );
buf ( n4982 , n4981 );
nand ( n4983 , n4976 , n4982 );
buf ( n4984 , n4983 );
buf ( n4985 , n4984 );
xor ( n4986 , n4971 , n4985 );
buf ( n4987 , n4986 );
buf ( n4988 , n4987 );
xor ( n4989 , n4944 , n4988 );
buf ( n4990 , n4989 );
buf ( n4991 , n4990 );
xor ( n4992 , n4917 , n4991 );
buf ( n4993 , n4992 );
buf ( n4994 , n4993 );
xor ( n4995 , n4478 , n4484 );
and ( n4996 , n4995 , n4596 );
and ( n4997 , n4478 , n4484 );
or ( n4998 , n4996 , n4997 );
buf ( n4999 , n4998 );
buf ( n5000 , n4999 );
xor ( n5001 , n4994 , n5000 );
xor ( n5002 , n4408 , n4414 );
and ( n5003 , n5002 , n4462 );
and ( n5004 , n4408 , n4414 );
or ( n5005 , n5003 , n5004 );
buf ( n5006 , n5005 );
buf ( n5007 , n5006 );
xor ( n5008 , n4525 , n4531 );
and ( n5009 , n5008 , n4593 );
and ( n5010 , n4525 , n4531 );
or ( n5011 , n5009 , n5010 );
buf ( n5012 , n5011 );
buf ( n5013 , n5012 );
xor ( n5014 , n5007 , n5013 );
buf ( n5015 , n559 );
buf ( n5016 , n581 );
or ( n5017 , n5015 , n5016 );
buf ( n5018 , n582 );
nand ( n5019 , n5017 , n5018 );
buf ( n5020 , n5019 );
buf ( n5021 , n5020 );
buf ( n5022 , n559 );
buf ( n5023 , n581 );
nand ( n5024 , n5022 , n5023 );
buf ( n5025 , n5024 );
buf ( n5026 , n5025 );
buf ( n5027 , n580 );
and ( n5028 , n5021 , n5026 , n5027 );
buf ( n5029 , n5028 );
buf ( n5030 , n4560 );
not ( n5031 , n5030 );
buf ( n5032 , n1060 );
not ( n5033 , n5032 );
or ( n5034 , n5031 , n5033 );
buf ( n5035 , n1071 );
buf ( n5036 , n550 );
buf ( n5037 , n588 );
xor ( n5038 , n5036 , n5037 );
buf ( n5039 , n5038 );
buf ( n5040 , n5039 );
nand ( n5041 , n5035 , n5040 );
buf ( n5042 , n5041 );
buf ( n5043 , n5042 );
nand ( n5044 , n5034 , n5043 );
buf ( n5045 , n5044 );
xor ( n5046 , n5029 , n5045 );
not ( n5047 , n5046 );
buf ( n5048 , n559 );
buf ( n5049 , n580 );
xor ( n5050 , n5048 , n5049 );
buf ( n5051 , n5050 );
not ( n5052 , n5051 );
not ( n5053 , n580 );
not ( n5054 , n4739 );
or ( n5055 , n5053 , n5054 );
not ( n5056 , n580 );
nand ( n5057 , n5056 , n581 );
nand ( n5058 , n5055 , n5057 );
nand ( n5059 , n5058 , n4541 );
not ( n5060 , n5059 );
not ( n5061 , n5060 );
or ( n5062 , n5052 , n5061 );
buf ( n5063 , n4544 );
buf ( n5064 , n5063 );
buf ( n5065 , n5064 );
buf ( n5066 , n5065 );
buf ( n5067 , n558 );
buf ( n5068 , n580 );
xor ( n5069 , n5067 , n5068 );
buf ( n5070 , n5069 );
buf ( n5071 , n5070 );
nand ( n5072 , n5066 , n5071 );
buf ( n5073 , n5072 );
nand ( n5074 , n5062 , n5073 );
not ( n5075 , n4486 );
not ( n5076 , n1177 );
or ( n5077 , n5075 , n5076 );
buf ( n5078 , n1036 );
buf ( n5079 , n552 );
buf ( n5080 , n586 );
xor ( n5081 , n5079 , n5080 );
buf ( n5082 , n5081 );
buf ( n5083 , n5082 );
nand ( n5084 , n5078 , n5083 );
buf ( n5085 , n5084 );
nand ( n5086 , n5077 , n5085 );
not ( n5087 , n5086 );
and ( n5088 , n5074 , n5087 );
not ( n5089 , n5074 );
and ( n5090 , n5089 , n5086 );
nor ( n5091 , n5088 , n5090 );
not ( n5092 , n5091 );
or ( n5093 , n5047 , n5092 );
or ( n5094 , n5046 , n5091 );
nand ( n5095 , n5093 , n5094 );
buf ( n5096 , n5095 );
xor ( n5097 , n4537 , n4583 );
and ( n5098 , n5097 , n4590 );
and ( n5099 , n4537 , n4583 );
or ( n5100 , n5098 , n5099 );
buf ( n5101 , n5100 );
buf ( n5102 , n5101 );
xor ( n5103 , n5096 , n5102 );
not ( n5104 , n4520 );
not ( n5105 , n4522 );
or ( n5106 , n5104 , n5105 );
nand ( n5107 , n5106 , n4517 );
nand ( n5108 , n4491 , n4503 );
nand ( n5109 , n5107 , n5108 );
xor ( n5110 , n4548 , n4564 );
and ( n5111 , n5110 , n4581 );
and ( n5112 , n4548 , n4564 );
or ( n5113 , n5111 , n5112 );
xor ( n5114 , n5109 , n5113 );
not ( n5115 , n4498 );
not ( n5116 , n984 );
or ( n5117 , n5115 , n5116 );
xor ( n5118 , n590 , n548 );
nand ( n5119 , n5118 , n591 );
nand ( n5120 , n5117 , n5119 );
not ( n5121 , n4575 );
not ( n5122 , n3664 );
or ( n5123 , n5121 , n5122 );
buf ( n5124 , n2123 );
buf ( n5125 , n554 );
buf ( n5126 , n584 );
xor ( n5127 , n5125 , n5126 );
buf ( n5128 , n5127 );
buf ( n5129 , n5128 );
nand ( n5130 , n5124 , n5129 );
buf ( n5131 , n5130 );
nand ( n5132 , n5123 , n5131 );
xor ( n5133 , n5120 , n5132 );
buf ( n5134 , n556 );
buf ( n5135 , n582 );
xor ( n5136 , n5134 , n5135 );
buf ( n5137 , n5136 );
and ( n5138 , n4211 , n5137 );
and ( n5139 , n4205 , n4512 );
nor ( n5140 , n5138 , n5139 );
not ( n5141 , n5140 );
xor ( n5142 , n5133 , n5141 );
xor ( n5143 , n5114 , n5142 );
buf ( n5144 , n5143 );
xor ( n5145 , n5103 , n5144 );
buf ( n5146 , n5145 );
buf ( n5147 , n5146 );
xor ( n5148 , n5014 , n5147 );
buf ( n5149 , n5148 );
buf ( n5150 , n5149 );
xor ( n5151 , n5001 , n5150 );
buf ( n5152 , n5151 );
buf ( n5153 , n5152 );
not ( n5154 , n5153 );
buf ( n5155 , n5154 );
xor ( n5156 , n4465 , n4471 );
and ( n5157 , n5156 , n4599 );
and ( n5158 , n4465 , n4471 );
or ( n5159 , n5157 , n5158 );
buf ( n5160 , n5159 );
buf ( n5161 , n5160 );
not ( n5162 , n5161 );
buf ( n5163 , n5162 );
nand ( n5164 , n5155 , n5163 );
not ( n5165 , n5164 );
nand ( n5166 , n5152 , n5160 );
not ( n5167 , n5166 );
nor ( n5168 , n5165 , n5167 );
buf ( n5169 , n5168 );
and ( n5170 , n4819 , n5169 );
not ( n5171 , n4819 );
buf ( n5172 , n5168 );
not ( n5173 , n5172 );
buf ( n5174 , n5173 );
and ( n5175 , n5171 , n5174 );
or ( n5176 , n5170 , n5175 );
xor ( n5177 , n3205 , n3209 );
and ( n5178 , n5177 , n3279 );
and ( n5179 , n3205 , n3209 );
or ( n5180 , n5178 , n5179 );
not ( n5181 , n5180 );
not ( n5182 , n2276 );
not ( n5183 , n3200 );
or ( n5184 , n5182 , n5183 );
not ( n5185 , n554 );
not ( n5186 , n2981 );
not ( n5187 , n5186 );
or ( n5188 , n5185 , n5187 );
not ( n5189 , n554 );
nand ( n5190 , n5189 , n2981 );
nand ( n5191 , n5188 , n5190 );
nand ( n5192 , n5191 , n3118 );
nand ( n5193 , n5184 , n5192 );
xor ( n5194 , n3214 , n3224 );
and ( n5195 , n5194 , n3236 );
and ( n5196 , n3214 , n3224 );
or ( n5197 , n5195 , n5196 );
xor ( n5198 , n5193 , n5197 );
not ( n5199 , n1596 );
not ( n5200 , n556 );
not ( n5201 , n3167 );
not ( n5202 , n5201 );
or ( n5203 , n5200 , n5202 );
nand ( n5204 , n3167 , n1625 );
nand ( n5205 , n5203 , n5204 );
not ( n5206 , n5205 );
or ( n5207 , n5199 , n5206 );
nand ( n5208 , n3189 , n1659 );
nand ( n5209 , n5207 , n5208 );
xor ( n5210 , n5198 , n5209 );
xor ( n5211 , n3237 , n3273 );
and ( n5212 , n5211 , n3278 );
and ( n5213 , n3237 , n3273 );
or ( n5214 , n5212 , n5213 );
xor ( n5215 , n5210 , n5214 );
not ( n5216 , n559 );
not ( n5217 , n558 );
nand ( n5218 , n564 , n580 );
not ( n5219 , n5218 );
nor ( n5220 , n564 , n580 );
nor ( n5221 , n5219 , n5220 );
not ( n5222 , n5221 );
and ( n5223 , n3242 , n3256 );
not ( n5224 , n5223 );
not ( n5225 , n3008 );
not ( n5226 , n3000 );
or ( n5227 , n5225 , n5226 );
not ( n5228 , n3025 );
not ( n5229 , n3030 );
or ( n5230 , n5228 , n5229 );
nand ( n5231 , n3018 , n3011 );
nand ( n5232 , n5230 , n5231 );
nand ( n5233 , n5227 , n5232 );
not ( n5234 , n5233 );
or ( n5235 , n5224 , n5234 );
and ( n5236 , n3256 , n3252 );
not ( n5237 , n3257 );
nor ( n5238 , n5236 , n5237 );
nand ( n5239 , n5235 , n5238 );
not ( n5240 , n5239 );
not ( n5241 , n5240 );
or ( n5242 , n5222 , n5241 );
not ( n5243 , n5218 );
or ( n5244 , n5243 , n5220 );
nand ( n5245 , n5244 , n5239 );
nand ( n5246 , n5242 , n5245 );
not ( n5247 , n5246 );
not ( n5248 , n5247 );
or ( n5249 , n5217 , n5248 );
not ( n5250 , n5247 );
nand ( n5251 , n5250 , n1736 );
nand ( n5252 , n5249 , n5251 );
not ( n5253 , n5252 );
or ( n5254 , n5216 , n5253 );
nand ( n5255 , n3269 , n1739 );
nand ( n5256 , n5254 , n5255 );
not ( n5257 , n3068 );
not ( n5258 , n550 );
not ( n5259 , n3049 );
or ( n5260 , n5258 , n5259 );
not ( n5261 , n1621 );
nand ( n5262 , n5261 , n3073 );
nand ( n5263 , n5260 , n5262 );
not ( n5264 , n5263 );
or ( n5265 , n5257 , n5264 );
not ( n5266 , n3083 );
not ( n5267 , n3067 );
and ( n5268 , n5266 , n5267 );
nand ( n5269 , n3220 , n5268 );
nand ( n5270 , n5265 , n5269 );
or ( n5271 , n549 , n550 );
nand ( n5272 , n5271 , n1664 );
nand ( n5273 , n549 , n550 );
and ( n5274 , n5272 , n5273 , n548 );
not ( n5275 , n3212 );
not ( n5276 , n548 );
not ( n5277 , n1677 );
or ( n5278 , n5276 , n5277 );
not ( n5279 , n548 );
nand ( n5280 , n1680 , n5279 );
nand ( n5281 , n5278 , n5280 );
not ( n5282 , n5281 );
or ( n5283 , n5275 , n5282 );
not ( n5284 , n548 );
not ( n5285 , n1687 );
or ( n5286 , n5284 , n5285 );
nand ( n5287 , n1664 , n5279 );
nand ( n5288 , n5286 , n5287 );
xnor ( n5289 , n548 , n549 );
and ( n5290 , n549 , n3073 );
not ( n5291 , n549 );
and ( n5292 , n5291 , n550 );
or ( n5293 , n5290 , n5292 );
nor ( n5294 , n5289 , n5293 );
nand ( n5295 , n5288 , n5294 );
nand ( n5296 , n5283 , n5295 );
xor ( n5297 , n5274 , n5296 );
xor ( n5298 , n5270 , n5297 );
buf ( n5299 , n2265 );
not ( n5300 , n5299 );
not ( n5301 , n552 );
not ( n5302 , n1776 );
or ( n5303 , n5301 , n5302 );
not ( n5304 , n1772 );
or ( n5305 , n5304 , n552 );
nand ( n5306 , n5303 , n5305 );
not ( n5307 , n5306 );
or ( n5308 , n5300 , n5307 );
nand ( n5309 , n3064 , n3232 );
nand ( n5310 , n5308 , n5309 );
xor ( n5311 , n5298 , n5310 );
xor ( n5312 , n5256 , n5311 );
xor ( n5313 , n3182 , n3191 );
and ( n5314 , n5313 , n3204 );
and ( n5315 , n3182 , n3191 );
or ( n5316 , n5314 , n5315 );
xor ( n5317 , n5312 , n5316 );
xor ( n5318 , n5215 , n5317 );
not ( n5319 , n5318 );
or ( n5320 , n5181 , n5319 );
nor ( n5321 , n5318 , n5180 );
not ( n5322 , n5321 );
nand ( n5323 , n5320 , n5322 );
not ( n5324 , n5323 );
not ( n5325 , n3280 );
not ( n5326 , n3181 );
nand ( n5327 , n5325 , n5326 );
nand ( n5328 , n3366 , n5327 );
not ( n5329 , n5328 );
not ( n5330 , n5329 );
nand ( n5331 , n3281 , n3181 );
nand ( n5332 , n5330 , n5331 );
not ( n5333 , n5332 );
or ( n5334 , n5324 , n5333 );
not ( n5335 , n5329 );
nand ( n5336 , n5335 , n5331 );
or ( n5337 , n5336 , n5323 );
nand ( n5338 , n5334 , n5337 );
nor ( n5339 , n5176 , n5338 );
not ( n5340 , n5339 );
and ( n5341 , n4819 , n5169 );
not ( n5342 , n4819 );
and ( n5343 , n5342 , n5174 );
nor ( n5344 , n5341 , n5343 );
not ( n5345 , n5344 );
not ( n5346 , n5323 );
not ( n5347 , n5332 );
or ( n5348 , n5346 , n5347 );
or ( n5349 , n5323 , n5336 );
nand ( n5350 , n5348 , n5349 );
nand ( n5351 , n5345 , n5350 );
nand ( n5352 , n5340 , n5351 );
and ( n5353 , n4800 , n5352 );
not ( n5354 , n4800 );
not ( n5355 , n5352 );
and ( n5356 , n5354 , n5355 );
nor ( n5357 , n5353 , n5356 );
nor ( n5358 , n580 , n5357 );
not ( n5359 , n5358 );
and ( n5360 , n4800 , n5352 );
not ( n5361 , n4800 );
and ( n5362 , n5361 , n5355 );
nor ( n5363 , n5360 , n5362 );
nand ( n5364 , n5363 , n580 );
nand ( n5365 , n5359 , n5364 );
or ( n5366 , n4795 , n5365 );
nand ( n5367 , n4795 , n5365 );
nand ( n5368 , n5366 , n5367 );
not ( n5369 , n5368 );
buf ( n5370 , n5369 );
not ( n5371 , n5370 );
or ( n5372 , n2919 , n5371 );
buf ( n5373 , n5368 );
buf ( n5374 , n5373 );
not ( n5375 , n5374 );
buf ( n5376 , n5375 );
buf ( n5377 , n5376 );
not ( n5378 , n5377 );
buf ( n5379 , n5378 );
buf ( n5380 , n5379 );
not ( n5381 , n600 );
buf ( n5382 , n5381 );
buf ( n5383 , n5382 );
buf ( n5384 , n5383 );
nand ( n5385 , n5380 , n5384 );
buf ( n5386 , n5385 );
buf ( n5387 , n5386 );
nand ( n5388 , n5372 , n5387 );
buf ( n5389 , n5388 );
buf ( n5390 , n5389 );
not ( n5391 , n5390 );
or ( n5392 , n2917 , n5391 );
buf ( n5393 , n600 );
not ( n5394 , n5393 );
nand ( n5395 , n4738 , n4739 );
nand ( n5396 , n5395 , n4794 );
not ( n5397 , n5396 );
not ( n5398 , n4779 );
not ( n5399 , n4758 );
or ( n5400 , n5398 , n5399 );
not ( n5401 , n4791 );
nand ( n5402 , n5400 , n5401 );
not ( n5403 , n5402 );
or ( n5404 , n5397 , n5403 );
or ( n5405 , n5402 , n5396 );
nand ( n5406 , n5404 , n5405 );
not ( n5407 , n5406 );
buf ( n5408 , n5407 );
not ( n5409 , n5408 );
or ( n5410 , n5394 , n5409 );
buf ( n5411 , n5406 );
buf ( n5412 , n5411 );
buf ( n5413 , n5383 );
nand ( n5414 , n5412 , n5413 );
buf ( n5415 , n5414 );
buf ( n5416 , n5415 );
nand ( n5417 , n5410 , n5416 );
buf ( n5418 , n5417 );
buf ( n5419 , n5418 );
buf ( n5420 , n600 );
buf ( n5421 , n601 );
and ( n5422 , n5420 , n5421 );
buf ( n5423 , n2914 );
buf ( n5424 , n600 );
buf ( n5425 , n601 );
nor ( n5426 , n5424 , n5425 );
buf ( n5427 , n5426 );
buf ( n5428 , n5427 );
nor ( n5429 , n5422 , n5423 , n5428 );
buf ( n5430 , n5429 );
buf ( n5431 , n5430 );
nand ( n5432 , n5419 , n5431 );
buf ( n5433 , n5432 );
buf ( n5434 , n5433 );
nand ( n5435 , n5392 , n5434 );
buf ( n5436 , n5435 );
buf ( n5437 , n5436 );
xor ( n5438 , n2907 , n5437 );
buf ( n5439 , n825 );
not ( n5440 , n5439 );
buf ( n5441 , n596 );
not ( n5442 , n5441 );
not ( n5443 , n2352 );
or ( n5444 , n5443 , C0 );
or ( n5445 , n2314 , n585 );
nand ( n5446 , n5444 , n5445 );
nand ( n5447 , n5446 , n2315 );
not ( n5448 , n5447 );
not ( n5449 , n5448 );
nand ( n5450 , n4755 , n4752 );
not ( n5451 , n5450 );
not ( n5452 , n5451 );
or ( n5453 , n5449 , n5452 );
nand ( n5454 , n5450 , n5447 );
nand ( n5455 , n5453 , n5454 );
buf ( n5456 , n5455 );
not ( n5457 , n5456 );
buf ( n5458 , n5457 );
buf ( n5459 , n5458 );
not ( n5460 , n5459 );
or ( n5461 , n5442 , n5460 );
buf ( n5462 , n5455 );
buf ( n5463 , n5462 );
buf ( n5464 , n5463 );
buf ( n5465 , n5464 );
buf ( n5466 , n2371 );
nand ( n5467 , n5465 , n5466 );
buf ( n5468 , n5467 );
buf ( n5469 , n5468 );
nand ( n5470 , n5461 , n5469 );
buf ( n5471 , n5470 );
buf ( n5472 , n5471 );
not ( n5473 , n5472 );
or ( n5474 , n5440 , n5473 );
buf ( n5475 , n2377 );
buf ( n5476 , n2404 );
nand ( n5477 , n5475 , n5476 );
buf ( n5478 , n5477 );
buf ( n5479 , n5478 );
nand ( n5480 , n5474 , n5479 );
buf ( n5481 , n5480 );
buf ( n5482 , n5481 );
buf ( n5483 , n2541 );
not ( n5484 , n5483 );
buf ( n5485 , n594 );
not ( n5486 , n5485 );
not ( n5487 , n2389 );
buf ( n5488 , n5487 );
not ( n5489 , n5488 );
or ( n5490 , n5486 , n5489 );
buf ( n5491 , n2390 );
buf ( n5492 , n2481 );
nand ( n5493 , n5491 , n5492 );
buf ( n5494 , n5493 );
buf ( n5495 , n5494 );
nand ( n5496 , n5490 , n5495 );
buf ( n5497 , n5496 );
buf ( n5498 , n5497 );
not ( n5499 , n5498 );
or ( n5500 , n5484 , n5499 );
buf ( n5501 , n2562 );
buf ( n5502 , n2592 );
nand ( n5503 , n5501 , n5502 );
buf ( n5504 , n5503 );
buf ( n5505 , n5504 );
nand ( n5506 , n5500 , n5505 );
buf ( n5507 , n5506 );
buf ( n5508 , n5507 );
buf ( n5509 , n2440 );
buf ( n5510 , n592 );
and ( n5511 , n5509 , n5510 );
buf ( n5512 , n5511 );
buf ( n5513 , n5512 );
xor ( n5514 , n2420 , n2498 );
and ( n5515 , n5514 , n2529 );
or ( n5516 , n5515 , C0 );
buf ( n5517 , n5516 );
buf ( n5518 , n5517 );
xor ( n5519 , n5513 , n5518 );
and ( n5520 , n2573 , n2416 );
not ( n5521 , n2573 );
and ( n5522 , n5521 , n592 );
nor ( n5523 , n5520 , n5522 );
or ( n5524 , n5523 , n2519 );
buf ( n5525 , n2515 );
not ( n5526 , n5525 );
buf ( n5527 , n2460 );
nand ( n5528 , n5526 , n5527 );
buf ( n5529 , n5528 );
nand ( n5530 , n5524 , n5529 );
buf ( n5531 , n5530 );
xor ( n5532 , n5519 , n5531 );
buf ( n5533 , n5532 );
buf ( n5534 , n5533 );
xor ( n5535 , n5508 , n5534 );
xor ( n5536 , n2532 , n2599 );
and ( n5537 , n5536 , n2718 );
and ( n5538 , n2532 , n2599 );
or ( n5539 , n5537 , n5538 );
buf ( n5540 , n5539 );
buf ( n5541 , n5540 );
xor ( n5542 , n5535 , n5541 );
buf ( n5543 , n5542 );
buf ( n5544 , n5543 );
xor ( n5545 , n5482 , n5544 );
and ( n5546 , n599 , n600 );
not ( n5547 , n599 );
and ( n5548 , n5547 , n5381 );
nor ( n5549 , n5546 , n5548 );
buf ( n5550 , n5549 );
buf ( n5551 , n5550 );
not ( n5552 , n5551 );
buf ( n5553 , n598 );
not ( n5554 , n5553 );
and ( n5555 , n4759 , n4762 );
not ( n5556 , n4759 );
and ( n5557 , n5556 , n4666 );
nor ( n5558 , n5555 , n5557 );
nand ( n5559 , n4783 , n5558 );
not ( n5560 , n5559 );
not ( n5561 , n4758 );
or ( n5562 , n5560 , n5561 );
buf ( n5563 , n4785 );
nand ( n5564 , n5562 , n5563 );
not ( n5565 , n4778 );
nand ( n5566 , n5565 , n4790 );
not ( n5567 , n5566 );
and ( n5568 , n5564 , n5567 );
not ( n5569 , n5564 );
and ( n5570 , n5569 , n5566 );
nor ( n5571 , n5568 , n5570 );
not ( n5572 , n5571 );
buf ( n5573 , n5572 );
not ( n5574 , n5573 );
or ( n5575 , n5554 , n5574 );
buf ( n5576 , n5571 );
buf ( n5577 , n5576 );
buf ( n5578 , n818 );
nand ( n5579 , n5577 , n5578 );
buf ( n5580 , n5579 );
buf ( n5581 , n5580 );
nand ( n5582 , n5575 , n5581 );
buf ( n5583 , n5582 );
buf ( n5584 , n5583 );
not ( n5585 , n5584 );
or ( n5586 , n5552 , n5585 );
buf ( n5587 , n598 );
not ( n5588 , n5587 );
not ( n5589 , n583 );
not ( n5590 , n4764 );
or ( n5591 , n5589 , n5590 );
nand ( n5592 , n5591 , n5559 );
nand ( n5593 , n4753 , n4755 , n4757 );
and ( n5594 , n5592 , n5593 );
not ( n5595 , n5592 );
not ( n5596 , n5593 );
and ( n5597 , n5595 , n5596 );
nor ( n5598 , n5594 , n5597 );
buf ( n5599 , n5598 );
buf ( n5600 , n5599 );
buf ( n5601 , n5600 );
buf ( n5602 , n5601 );
not ( n5603 , n5602 );
or ( n5604 , n5588 , n5603 );
buf ( n5605 , n5601 );
not ( n5606 , n5605 );
buf ( n5607 , n5606 );
buf ( n5608 , n5607 );
buf ( n5609 , n818 );
nand ( n5610 , n5608 , n5609 );
buf ( n5611 , n5610 );
buf ( n5612 , n5611 );
nand ( n5613 , n5604 , n5612 );
buf ( n5614 , n5613 );
buf ( n5615 , n5614 );
buf ( n5616 , n5549 );
not ( n5617 , n5616 );
buf ( n5618 , n5617 );
buf ( n5619 , n5618 );
buf ( n5620 , n599 );
buf ( n5621 , n598 );
and ( n5622 , n5620 , n5621 );
not ( n5623 , n5620 );
buf ( n5624 , n818 );
and ( n5625 , n5623 , n5624 );
nor ( n5626 , n5622 , n5625 );
buf ( n5627 , n5626 );
buf ( n5628 , n5627 );
and ( n5629 , n5619 , n5628 );
buf ( n5630 , n5629 );
buf ( n5631 , n5630 );
buf ( n5632 , n5631 );
nand ( n5633 , n5615 , n5632 );
buf ( n5634 , n5633 );
buf ( n5635 , n5634 );
nand ( n5636 , n5586 , n5635 );
buf ( n5637 , n5636 );
buf ( n5638 , n5637 );
xor ( n5639 , n5545 , n5638 );
buf ( n5640 , n5639 );
buf ( n5641 , n5640 );
and ( n5642 , n5438 , n5641 );
and ( n5643 , n2907 , n5437 );
or ( n5644 , n5642 , n5643 );
buf ( n5645 , n5644 );
buf ( n5646 , n5645 );
or ( n5647 , n603 , n604 );
buf ( n5648 , n603 );
buf ( n5649 , n604 );
nand ( n5650 , n5648 , n5649 );
buf ( n5651 , n5650 );
nand ( n5652 , n5647 , n5651 );
buf ( n5653 , n5652 );
not ( n5654 , n5653 );
buf ( n5655 , n5654 );
buf ( n5656 , n5655 );
not ( n5657 , n5656 );
buf ( n5658 , n602 );
not ( n5659 , n5658 );
xor ( n5660 , n4852 , n4869 );
and ( n5661 , n5660 , n4903 );
and ( n5662 , n4852 , n4869 );
or ( n5663 , n5661 , n5662 );
buf ( n5664 , n5663 );
not ( n5665 , n5664 );
buf ( n5666 , n547 );
buf ( n5667 , n574 );
xor ( n5668 , n5666 , n5667 );
buf ( n5669 , n5668 );
not ( n5670 , n5669 );
not ( n5671 , n575 );
or ( n5672 , n5670 , n5671 );
nand ( n5673 , n4949 , n4953 );
nand ( n5674 , n5672 , n5673 );
not ( n5675 , n4845 );
not ( n5676 , n4830 );
xor ( n5677 , n565 , n566 );
nor ( n5678 , n5676 , n5677 );
not ( n5679 , n5678 );
or ( n5680 , n5675 , n5679 );
buf ( n5681 , n4840 );
buf ( n5682 , n557 );
buf ( n5683 , n564 );
xor ( n5684 , n5682 , n5683 );
buf ( n5685 , n5684 );
buf ( n5686 , n5685 );
nand ( n5687 , n5681 , n5686 );
buf ( n5688 , n5687 );
nand ( n5689 , n5680 , n5688 );
xor ( n5690 , n5674 , n5689 );
not ( n5691 , n4978 );
not ( n5692 , n4380 );
or ( n5693 , n5691 , n5692 );
buf ( n5694 , n3743 );
buf ( n5695 , n555 );
buf ( n5696 , n566 );
xor ( n5697 , n5695 , n5696 );
buf ( n5698 , n5697 );
buf ( n5699 , n5698 );
nand ( n5700 , n5694 , n5699 );
buf ( n5701 , n5700 );
nand ( n5702 , n5693 , n5701 );
xor ( n5703 , n5690 , n5702 );
not ( n5704 , n5703 );
buf ( n5705 , n563 );
buf ( n5706 , n564 );
xor ( n5707 , n5705 , n5706 );
buf ( n5708 , n5707 );
buf ( n5709 , n5708 );
not ( n5710 , n5709 );
buf ( n5711 , n1490 );
nor ( n5712 , n5710 , n5711 );
buf ( n5713 , n5712 );
buf ( n5714 , n5713 );
buf ( n5715 , n4893 );
not ( n5716 , n5715 );
buf ( n5717 , n4435 );
not ( n5718 , n5717 );
or ( n5719 , n5716 , n5718 );
buf ( n5720 , n888 );
xor ( n5721 , n572 , n549 );
buf ( n5722 , n5721 );
nand ( n5723 , n5720 , n5722 );
buf ( n5724 , n5723 );
buf ( n5725 , n5724 );
nand ( n5726 , n5719 , n5725 );
buf ( n5727 , n5726 );
buf ( n5728 , n5727 );
xor ( n5729 , n5714 , n5728 );
buf ( n5730 , n4965 );
not ( n5731 , n5730 );
buf ( n5732 , n4021 );
not ( n5733 , n5732 );
or ( n5734 , n5731 , n5733 );
buf ( n5735 , n3436 );
xor ( n5736 , n568 , n553 );
buf ( n5737 , n5736 );
nand ( n5738 , n5735 , n5737 );
buf ( n5739 , n5738 );
buf ( n5740 , n5739 );
nand ( n5741 , n5734 , n5740 );
buf ( n5742 , n5741 );
buf ( n5743 , n5742 );
xor ( n5744 , n5729 , n5743 );
buf ( n5745 , n5744 );
not ( n5746 , n5745 );
nand ( n5747 , n5704 , n5746 );
not ( n5748 , n5747 );
or ( n5749 , n5665 , n5748 );
nand ( n5750 , n5703 , n5745 );
nand ( n5751 , n5749 , n5750 );
buf ( n5752 , n5751 );
xor ( n5753 , n5714 , n5728 );
and ( n5754 , n5753 , n5743 );
and ( n5755 , n5714 , n5728 );
or ( n5756 , n5754 , n5755 );
buf ( n5757 , n5756 );
buf ( n5758 , n5669 );
not ( n5759 , n5758 );
buf ( n5760 , n1110 );
not ( n5761 , n5760 );
or ( n5762 , n5759 , n5761 );
xor ( n5763 , n546 , n574 );
nand ( n5764 , n5763 , n575 );
buf ( n5765 , n5764 );
nand ( n5766 , n5762 , n5765 );
buf ( n5767 , n5766 );
buf ( n5768 , n5767 );
buf ( n5769 , n559 );
buf ( n5770 , n563 );
nand ( n5771 , n5769 , n5770 );
buf ( n5772 , n5771 );
or ( n5773 , n559 , n563 );
nand ( n5774 , n5773 , n564 );
nand ( n5775 , n5772 , n5774 , n562 );
not ( n5776 , n5775 );
buf ( n5777 , n5776 );
and ( n5778 , n5768 , n5777 );
not ( n5779 , n5768 );
buf ( n5780 , n5775 );
and ( n5781 , n5779 , n5780 );
nor ( n5782 , n5778 , n5781 );
buf ( n5783 , n5782 );
not ( n5784 , n5783 );
and ( n5785 , n5757 , n5784 );
not ( n5786 , n5757 );
and ( n5787 , n5786 , n5783 );
nor ( n5788 , n5785 , n5787 );
xor ( n5789 , n5674 , n5689 );
and ( n5790 , n5789 , n5702 );
and ( n5791 , n5674 , n5689 );
or ( n5792 , n5790 , n5791 );
xor ( n5793 , n5788 , n5792 );
not ( n5794 , n5793 );
and ( n5795 , n5752 , n5794 );
not ( n5796 , n5752 );
and ( n5797 , n5796 , n5793 );
nor ( n5798 , n5795 , n5797 );
buf ( n5799 , n5708 );
buf ( n5800 , n5799 );
buf ( n5801 , n5800 );
not ( n5802 , n5801 );
buf ( n5803 , n558 );
buf ( n5804 , n562 );
xor ( n5805 , n5803 , n5804 );
buf ( n5806 , n5805 );
not ( n5807 , n5806 );
or ( n5808 , n5802 , n5807 );
not ( n5809 , n563 );
or ( n5810 , n5809 , n564 );
not ( n5811 , n564 );
or ( n5812 , n5811 , n563 );
nand ( n5813 , n5810 , n5812 );
not ( n5814 , n5813 );
buf ( n5815 , n562 );
buf ( n5816 , n563 );
xnor ( n5817 , n5815 , n5816 );
buf ( n5818 , n5817 );
not ( n5819 , n5818 );
xor ( n5820 , n559 , n562 );
nand ( n5821 , n5814 , n5819 , n5820 );
nand ( n5822 , n5808 , n5821 );
buf ( n5823 , n5822 );
buf ( n5824 , n551 );
buf ( n5825 , n570 );
xor ( n5826 , n5824 , n5825 );
buf ( n5827 , n5826 );
buf ( n5828 , n5827 );
not ( n5829 , n5828 );
buf ( n5830 , n850 );
not ( n5831 , n5830 );
or ( n5832 , n5829 , n5831 );
buf ( n5833 , n1979 );
buf ( n5834 , n550 );
buf ( n5835 , n570 );
xor ( n5836 , n5834 , n5835 );
buf ( n5837 , n5836 );
buf ( n5838 , n5837 );
nand ( n5839 , n5833 , n5838 );
buf ( n5840 , n5839 );
buf ( n5841 , n5840 );
nand ( n5842 , n5832 , n5841 );
buf ( n5843 , n5842 );
buf ( n5844 , n5843 );
xor ( n5845 , n5823 , n5844 );
buf ( n5846 , n5685 );
not ( n5847 , n5846 );
buf ( n5848 , n4836 );
not ( n5849 , n5848 );
or ( n5850 , n5847 , n5849 );
buf ( n5851 , n4840 );
buf ( n5852 , n556 );
buf ( n5853 , n564 );
xor ( n5854 , n5852 , n5853 );
buf ( n5855 , n5854 );
buf ( n5856 , n5855 );
nand ( n5857 , n5851 , n5856 );
buf ( n5858 , n5857 );
buf ( n5859 , n5858 );
nand ( n5860 , n5850 , n5859 );
buf ( n5861 , n5860 );
buf ( n5862 , n5861 );
xor ( n5863 , n5845 , n5862 );
buf ( n5864 , n5863 );
buf ( n5865 , n5864 );
not ( n5866 , n3772 );
xor ( n5867 , n552 , n568 );
not ( n5868 , n5867 );
or ( n5869 , n5866 , n5868 );
nand ( n5870 , n4958 , n5736 );
nand ( n5871 , n5869 , n5870 );
buf ( n5872 , n5871 );
not ( n5873 , n5721 );
not ( n5874 , n884 );
or ( n5875 , n5873 , n5874 );
buf ( n5876 , n548 );
buf ( n5877 , n572 );
xor ( n5878 , n5876 , n5877 );
buf ( n5879 , n5878 );
nand ( n5880 , n5879 , n888 );
nand ( n5881 , n5875 , n5880 );
buf ( n5882 , n5881 );
xor ( n5883 , n5872 , n5882 );
buf ( n5884 , n5698 );
not ( n5885 , n5884 );
buf ( n5886 , n4380 );
not ( n5887 , n5886 );
or ( n5888 , n5885 , n5887 );
buf ( n5889 , n3743 );
buf ( n5890 , n554 );
buf ( n5891 , n566 );
xor ( n5892 , n5890 , n5891 );
buf ( n5893 , n5892 );
buf ( n5894 , n5893 );
nand ( n5895 , n5889 , n5894 );
buf ( n5896 , n5895 );
buf ( n5897 , n5896 );
nand ( n5898 , n5888 , n5897 );
buf ( n5899 , n5898 );
buf ( n5900 , n5899 );
xor ( n5901 , n5883 , n5900 );
buf ( n5902 , n5901 );
buf ( n5903 , n5902 );
xor ( n5904 , n5865 , n5903 );
buf ( n5905 , n4862 );
not ( n5906 , n5905 );
buf ( n5907 , n850 );
not ( n5908 , n5907 );
or ( n5909 , n5906 , n5908 );
buf ( n5910 , n1982 );
buf ( n5911 , n5827 );
nand ( n5912 , n5910 , n5911 );
buf ( n5913 , n5912 );
buf ( n5914 , n5913 );
nand ( n5915 , n5909 , n5914 );
buf ( n5916 , n5915 );
buf ( n5917 , n5916 );
xor ( n5918 , n4956 , n4970 );
and ( n5919 , n5918 , n4985 );
and ( n5920 , n4956 , n4970 );
or ( n5921 , n5919 , n5920 );
buf ( n5922 , n5921 );
buf ( n5923 , n5922 );
xor ( n5924 , n5917 , n5923 );
and ( n5925 , n4886 , n4900 );
buf ( n5926 , n5925 );
buf ( n5927 , n5926 );
and ( n5928 , n5924 , n5927 );
and ( n5929 , n5917 , n5923 );
or ( n5930 , n5928 , n5929 );
buf ( n5931 , n5930 );
buf ( n5932 , n5931 );
xor ( n5933 , n5904 , n5932 );
buf ( n5934 , n5933 );
and ( n5935 , n5798 , n5934 );
not ( n5936 , n5798 );
not ( n5937 , n5934 );
and ( n5938 , n5936 , n5937 );
nor ( n5939 , n5935 , n5938 );
buf ( n5940 , n5939 );
xor ( n5941 , n4906 , n4916 );
and ( n5942 , n5941 , n4991 );
and ( n5943 , n4906 , n4916 );
or ( n5944 , n5942 , n5943 );
buf ( n5945 , n5944 );
buf ( n5946 , n5945 );
xor ( n5947 , n5096 , n5102 );
and ( n5948 , n5947 , n5144 );
and ( n5949 , n5096 , n5102 );
or ( n5950 , n5948 , n5949 );
buf ( n5951 , n5950 );
buf ( n5952 , n5951 );
xor ( n5953 , n5946 , n5952 );
buf ( n5954 , n5082 );
not ( n5955 , n5954 );
buf ( n5956 , n1177 );
not ( n5957 , n5956 );
or ( n5958 , n5955 , n5957 );
buf ( n5959 , n1036 );
buf ( n5960 , n551 );
buf ( n5961 , n586 );
xor ( n5962 , n5960 , n5961 );
buf ( n5963 , n5962 );
buf ( n5964 , n5963 );
nand ( n5965 , n5959 , n5964 );
buf ( n5966 , n5965 );
buf ( n5967 , n5966 );
nand ( n5968 , n5958 , n5967 );
buf ( n5969 , n5968 );
buf ( n5970 , n5969 );
buf ( n5971 , n5045 );
buf ( n5972 , n5029 );
nand ( n5973 , n5971 , n5972 );
buf ( n5974 , n5973 );
buf ( n5975 , n5974 );
xor ( n5976 , n5970 , n5975 );
not ( n5977 , n5120 );
not ( n5978 , n5977 );
not ( n5979 , n5140 );
or ( n5980 , n5978 , n5979 );
nand ( n5981 , n5980 , n5132 );
nand ( n5982 , n5141 , n5120 );
nand ( n5983 , n5981 , n5982 );
buf ( n5984 , n5983 );
xnor ( n5985 , n5976 , n5984 );
buf ( n5986 , n5985 );
buf ( n5987 , n5986 );
xor ( n5988 , n5109 , n5113 );
and ( n5989 , n5988 , n5142 );
and ( n5990 , n5109 , n5113 );
or ( n5991 , n5989 , n5990 );
buf ( n5992 , n5991 );
xor ( n5993 , n5987 , n5992 );
buf ( n5994 , n579 );
buf ( n5995 , n580 );
xor ( n5996 , n5994 , n5995 );
buf ( n5997 , n5996 );
buf ( n5998 , n5997 );
buf ( n5999 , n559 );
and ( n6000 , n5998 , n5999 );
buf ( n6001 , n6000 );
buf ( n6002 , n6001 );
not ( n6003 , n6002 );
buf ( n6004 , n5039 );
not ( n6005 , n6004 );
buf ( n6006 , n4286 );
not ( n6007 , n6006 );
or ( n6008 , n6005 , n6007 );
buf ( n6009 , n549 );
buf ( n6010 , n588 );
xor ( n6011 , n6009 , n6010 );
buf ( n6012 , n6011 );
nand ( n6013 , n6012 , n4556 );
buf ( n6014 , n6013 );
nand ( n6015 , n6008 , n6014 );
buf ( n6016 , n6015 );
buf ( n6017 , n6016 );
not ( n6018 , n6017 );
buf ( n6019 , n6018 );
buf ( n6020 , n6019 );
not ( n6021 , n6020 );
or ( n6022 , n6003 , n6021 );
buf ( n6023 , n6016 );
buf ( n6024 , n5997 );
buf ( n6025 , n559 );
nand ( n6026 , n6024 , n6025 );
buf ( n6027 , n6026 );
buf ( n6028 , n6027 );
nand ( n6029 , n6023 , n6028 );
buf ( n6030 , n6029 );
buf ( n6031 , n6030 );
nand ( n6032 , n6022 , n6031 );
buf ( n6033 , n6032 );
buf ( n6034 , n6033 );
buf ( n6035 , n5128 );
not ( n6036 , n6035 );
buf ( n6037 , n3664 );
not ( n6038 , n6037 );
or ( n6039 , n6036 , n6038 );
buf ( n6040 , n2135 );
and ( n6041 , n553 , n584 );
not ( n6042 , n553 );
and ( n6043 , n6042 , n2964 );
nor ( n6044 , n6041 , n6043 );
buf ( n6045 , n6044 );
nand ( n6046 , n6040 , n6045 );
buf ( n6047 , n6046 );
buf ( n6048 , n6047 );
nand ( n6049 , n6039 , n6048 );
buf ( n6050 , n6049 );
buf ( n6051 , n6050 );
not ( n6052 , n6051 );
buf ( n6053 , n6052 );
buf ( n6054 , n6053 );
and ( n6055 , n6034 , n6054 );
not ( n6056 , n6034 );
buf ( n6057 , n6050 );
and ( n6058 , n6056 , n6057 );
nor ( n6059 , n6055 , n6058 );
buf ( n6060 , n6059 );
not ( n6061 , n6060 );
not ( n6062 , n6061 );
buf ( n6063 , n5118 );
not ( n6064 , n6063 );
buf ( n6065 , n984 );
not ( n6066 , n6065 );
or ( n6067 , n6064 , n6066 );
buf ( n6068 , n547 );
buf ( n6069 , n590 );
xor ( n6070 , n6068 , n6069 );
buf ( n6071 , n6070 );
buf ( n6072 , n6071 );
buf ( n6073 , n591 );
nand ( n6074 , n6072 , n6073 );
buf ( n6075 , n6074 );
buf ( n6076 , n6075 );
nand ( n6077 , n6067 , n6076 );
buf ( n6078 , n6077 );
buf ( n6079 , n6078 );
buf ( n6080 , n5137 );
not ( n6081 , n6080 );
buf ( n6082 , n4506 );
not ( n6083 , n6082 );
or ( n6084 , n6081 , n6083 );
buf ( n6085 , n3883 );
buf ( n6086 , n555 );
buf ( n6087 , n582 );
xor ( n6088 , n6086 , n6087 );
buf ( n6089 , n6088 );
buf ( n6090 , n6089 );
nand ( n6091 , n6085 , n6090 );
buf ( n6092 , n6091 );
buf ( n6093 , n6092 );
nand ( n6094 , n6084 , n6093 );
buf ( n6095 , n6094 );
buf ( n6096 , n6095 );
xor ( n6097 , n6079 , n6096 );
buf ( n6098 , n5070 );
not ( n6099 , n6098 );
buf ( n6100 , n5060 );
not ( n6101 , n6100 );
or ( n6102 , n6099 , n6101 );
buf ( n6103 , n4544 );
buf ( n6104 , n557 );
buf ( n6105 , n580 );
xor ( n6106 , n6104 , n6105 );
buf ( n6107 , n6106 );
buf ( n6108 , n6107 );
nand ( n6109 , n6103 , n6108 );
buf ( n6110 , n6109 );
buf ( n6111 , n6110 );
nand ( n6112 , n6102 , n6111 );
buf ( n6113 , n6112 );
buf ( n6114 , n6113 );
xor ( n6115 , n6097 , n6114 );
buf ( n6116 , n6115 );
not ( n6117 , n6116 );
or ( n6118 , n6062 , n6117 );
not ( n6119 , n6116 );
nand ( n6120 , n6119 , n6060 );
nand ( n6121 , n6118 , n6120 );
buf ( n6122 , n5074 );
not ( n6123 , n6122 );
buf ( n6124 , n5087 );
nand ( n6125 , n6123 , n6124 );
buf ( n6126 , n6125 );
buf ( n6127 , n6126 );
not ( n6128 , n6127 );
buf ( n6129 , n5046 );
not ( n6130 , n6129 );
or ( n6131 , n6128 , n6130 );
buf ( n6132 , n5086 );
buf ( n6133 , n5074 );
nand ( n6134 , n6132 , n6133 );
buf ( n6135 , n6134 );
buf ( n6136 , n6135 );
nand ( n6137 , n6131 , n6136 );
buf ( n6138 , n6137 );
not ( n6139 , n6138 );
and ( n6140 , n6121 , n6139 );
not ( n6141 , n6121 );
and ( n6142 , n6141 , n6138 );
nor ( n6143 , n6140 , n6142 );
buf ( n6144 , n6143 );
xor ( n6145 , n5993 , n6144 );
buf ( n6146 , n6145 );
buf ( n6147 , n6146 );
and ( n6148 , n5953 , n6147 );
and ( n6149 , n5946 , n5952 );
or ( n6150 , n6148 , n6149 );
buf ( n6151 , n6150 );
buf ( n6152 , n6151 );
xor ( n6153 , n5940 , n6152 );
xor ( n6154 , n4932 , n4943 );
and ( n6155 , n6154 , n4988 );
and ( n6156 , n4932 , n4943 );
or ( n6157 , n6155 , n6156 );
buf ( n6158 , n6157 );
not ( n6159 , n6158 );
xor ( n6160 , n5917 , n5923 );
xor ( n6161 , n6160 , n5927 );
buf ( n6162 , n6161 );
not ( n6163 , n6162 );
nand ( n6164 , n6159 , n6163 );
not ( n6165 , n6164 );
buf ( n6166 , n5664 );
not ( n6167 , n6166 );
not ( n6168 , n5704 );
not ( n6169 , n5745 );
and ( n6170 , n6168 , n6169 );
and ( n6171 , n5704 , n5745 );
nor ( n6172 , n6170 , n6171 );
not ( n6173 , n6172 );
or ( n6174 , n6167 , n6173 );
or ( n6175 , n6172 , n6166 );
nand ( n6176 , n6174 , n6175 );
not ( n6177 , n6176 );
or ( n6178 , n6165 , n6177 );
nand ( n6179 , n6162 , n6158 );
nand ( n6180 , n6178 , n6179 );
buf ( n6181 , n6180 );
xor ( n6182 , n5987 , n5992 );
and ( n6183 , n6182 , n6144 );
and ( n6184 , n5987 , n5992 );
or ( n6185 , n6183 , n6184 );
buf ( n6186 , n6185 );
buf ( n6187 , n6186 );
xor ( n6188 , n6181 , n6187 );
buf ( n6189 , n6060 );
not ( n6190 , n6189 );
buf ( n6191 , n6119 );
not ( n6192 , n6191 );
or ( n6193 , n6190 , n6192 );
buf ( n6194 , n6138 );
nand ( n6195 , n6193 , n6194 );
buf ( n6196 , n6195 );
buf ( n6197 , n6196 );
buf ( n6198 , n6060 );
not ( n6199 , n6198 );
buf ( n6200 , n6116 );
nand ( n6201 , n6199 , n6200 );
buf ( n6202 , n6201 );
buf ( n6203 , n6202 );
nand ( n6204 , n6197 , n6203 );
buf ( n6205 , n6204 );
buf ( n6206 , n6205 );
buf ( n6207 , n6027 );
not ( n6208 , n6207 );
buf ( n6209 , n6019 );
not ( n6210 , n6209 );
or ( n6211 , n6208 , n6210 );
buf ( n6212 , n6050 );
nand ( n6213 , n6211 , n6212 );
buf ( n6214 , n6213 );
buf ( n6215 , n6214 );
buf ( n6216 , n6019 );
not ( n6217 , n6216 );
buf ( n6218 , n6001 );
nand ( n6219 , n6217 , n6218 );
buf ( n6220 , n6219 );
buf ( n6221 , n6220 );
nand ( n6222 , n6215 , n6221 );
buf ( n6223 , n6222 );
buf ( n6224 , n559 );
buf ( n6225 , n579 );
or ( n6226 , n6224 , n6225 );
buf ( n6227 , n580 );
nand ( n6228 , n6226 , n6227 );
buf ( n6229 , n6228 );
buf ( n6230 , n559 );
buf ( n6231 , n579 );
nand ( n6232 , n6230 , n6231 );
buf ( n6233 , n6232 );
and ( n6234 , n6229 , n6233 , n578 );
buf ( n6235 , n6071 );
not ( n6236 , n6235 );
buf ( n6237 , n984 );
not ( n6238 , n6237 );
or ( n6239 , n6236 , n6238 );
buf ( n6240 , n546 );
buf ( n6241 , n590 );
xor ( n6242 , n6240 , n6241 );
buf ( n6243 , n6242 );
buf ( n6244 , n6243 );
buf ( n6245 , n591 );
nand ( n6246 , n6244 , n6245 );
buf ( n6247 , n6246 );
buf ( n6248 , n6247 );
nand ( n6249 , n6239 , n6248 );
buf ( n6250 , n6249 );
xor ( n6251 , n6234 , n6250 );
buf ( n6252 , n6251 );
xor ( n6253 , n6079 , n6096 );
and ( n6254 , n6253 , n6114 );
and ( n6255 , n6079 , n6096 );
or ( n6256 , n6254 , n6255 );
buf ( n6257 , n6256 );
nand ( n6258 , n6223 , n6252 , n6257 );
buf ( n6259 , n6214 );
buf ( n6260 , n6220 );
nand ( n6261 , n6259 , n6260 );
buf ( n6262 , n6261 );
nor ( n6263 , n6262 , n6252 );
nand ( n6264 , n6263 , n6257 );
not ( n6265 , n6223 );
not ( n6266 , n6257 );
nand ( n6267 , n6265 , n6266 , n6252 );
not ( n6268 , n6252 );
nand ( n6269 , n6268 , n6266 , n6223 );
nand ( n6270 , n6258 , n6264 , n6267 , n6269 );
buf ( n6271 , n6270 );
xor ( n6272 , n6206 , n6271 );
not ( n6273 , n6012 );
not ( n6274 , n4286 );
or ( n6275 , n6273 , n6274 );
buf ( n6276 , n548 );
buf ( n6277 , n588 );
xor ( n6278 , n6276 , n6277 );
buf ( n6279 , n6278 );
nand ( n6280 , n4556 , n6279 );
nand ( n6281 , n6275 , n6280 );
not ( n6282 , n2117 );
buf ( n6283 , n552 );
buf ( n6284 , n584 );
xor ( n6285 , n6283 , n6284 );
buf ( n6286 , n6285 );
not ( n6287 , n6286 );
or ( n6288 , n6282 , n6287 );
nand ( n6289 , n3662 , n2120 , n6044 );
nand ( n6290 , n6288 , n6289 );
not ( n6291 , n6290 );
xor ( n6292 , n6281 , n6291 );
not ( n6293 , n6089 );
not ( n6294 , n4506 );
or ( n6295 , n6293 , n6294 );
buf ( n6296 , n4211 );
buf ( n6297 , n554 );
buf ( n6298 , n582 );
xor ( n6299 , n6297 , n6298 );
buf ( n6300 , n6299 );
buf ( n6301 , n6300 );
nand ( n6302 , n6296 , n6301 );
buf ( n6303 , n6302 );
nand ( n6304 , n6295 , n6303 );
xor ( n6305 , n6292 , n6304 );
not ( n6306 , n3616 );
not ( n6307 , n5963 );
or ( n6308 , n6306 , n6307 );
and ( n6309 , n586 , n550 );
not ( n6310 , n586 );
not ( n6311 , n550 );
and ( n6312 , n6310 , n6311 );
nor ( n6313 , n6309 , n6312 );
nand ( n6314 , n6313 , n1036 );
nand ( n6315 , n6308 , n6314 );
buf ( n6316 , n6315 );
buf ( n6317 , n6107 );
not ( n6318 , n6317 );
buf ( n6319 , n5060 );
not ( n6320 , n6319 );
or ( n6321 , n6318 , n6320 );
buf ( n6322 , n4544 );
buf ( n6323 , n556 );
buf ( n6324 , n580 );
xor ( n6325 , n6323 , n6324 );
buf ( n6326 , n6325 );
buf ( n6327 , n6326 );
nand ( n6328 , n6322 , n6327 );
buf ( n6329 , n6328 );
buf ( n6330 , n6329 );
nand ( n6331 , n6321 , n6330 );
buf ( n6332 , n6331 );
buf ( n6333 , n6332 );
xor ( n6334 , n6316 , n6333 );
buf ( n6335 , n559 );
buf ( n6336 , n578 );
xor ( n6337 , n6335 , n6336 );
buf ( n6338 , n6337 );
buf ( n6339 , n6338 );
not ( n6340 , n6339 );
and ( n6341 , n579 , n580 );
not ( n6342 , n579 );
and ( n6343 , n6342 , n5056 );
nor ( n6344 , n6341 , n6343 );
not ( n6345 , n578 );
and ( n6346 , n579 , n6345 );
not ( n6347 , n579 );
and ( n6348 , n6347 , n578 );
nor ( n6349 , n6346 , n6348 );
nor ( n6350 , n6344 , n6349 );
buf ( n6351 , n6350 );
not ( n6352 , n6351 );
or ( n6353 , n6340 , n6352 );
buf ( n6354 , n5997 );
buf ( n6355 , n558 );
buf ( n6356 , n578 );
xor ( n6357 , n6355 , n6356 );
buf ( n6358 , n6357 );
buf ( n6359 , n6358 );
nand ( n6360 , n6354 , n6359 );
buf ( n6361 , n6360 );
buf ( n6362 , n6361 );
nand ( n6363 , n6353 , n6362 );
buf ( n6364 , n6363 );
buf ( n6365 , n6364 );
xor ( n6366 , n6334 , n6365 );
buf ( n6367 , n6366 );
xnor ( n6368 , n6305 , n6367 );
buf ( n6369 , n5969 );
not ( n6370 , n6369 );
buf ( n6371 , n5974 );
not ( n6372 , n6371 );
buf ( n6373 , n6372 );
buf ( n6374 , n6373 );
not ( n6375 , n6374 );
or ( n6376 , n6370 , n6375 );
buf ( n6377 , n5969 );
not ( n6378 , n6377 );
buf ( n6379 , n6378 );
buf ( n6380 , n6379 );
not ( n6381 , n6380 );
buf ( n6382 , n5974 );
not ( n6383 , n6382 );
or ( n6384 , n6381 , n6383 );
buf ( n6385 , n5983 );
nand ( n6386 , n6384 , n6385 );
buf ( n6387 , n6386 );
buf ( n6388 , n6387 );
nand ( n6389 , n6376 , n6388 );
buf ( n6390 , n6389 );
xor ( n6391 , n6368 , n6390 );
buf ( n6392 , n6391 );
xor ( n6393 , n6272 , n6392 );
buf ( n6394 , n6393 );
buf ( n6395 , n6394 );
xor ( n6396 , n6188 , n6395 );
buf ( n6397 , n6396 );
buf ( n6398 , n6397 );
xor ( n6399 , n6153 , n6398 );
buf ( n6400 , n6399 );
not ( n6401 , n6176 );
nand ( n6402 , n6179 , n6164 );
not ( n6403 , n6402 );
or ( n6404 , n6401 , n6403 );
not ( n6405 , n6176 );
xor ( n6406 , n6158 , n6162 );
nand ( n6407 , n6405 , n6406 );
nand ( n6408 , n6404 , n6407 );
buf ( n6409 , n6408 );
xor ( n6410 , n5007 , n5013 );
and ( n6411 , n6410 , n5147 );
and ( n6412 , n5007 , n5013 );
or ( n6413 , n6411 , n6412 );
buf ( n6414 , n6413 );
buf ( n6415 , n6414 );
xor ( n6416 , n6409 , n6415 );
xor ( n6417 , n5946 , n5952 );
xor ( n6418 , n6417 , n6147 );
buf ( n6419 , n6418 );
buf ( n6420 , n6419 );
and ( n6421 , n6416 , n6420 );
and ( n6422 , n6409 , n6415 );
or ( n6423 , n6421 , n6422 );
buf ( n6424 , n6423 );
nor ( n6425 , n6400 , n6424 );
xor ( n6426 , n6409 , n6415 );
xor ( n6427 , n6426 , n6420 );
buf ( n6428 , n6427 );
xor ( n6429 , n4994 , n5000 );
and ( n6430 , n6429 , n5150 );
and ( n6431 , n4994 , n5000 );
or ( n6432 , n6430 , n6431 );
buf ( n6433 , n6432 );
nand ( n6434 , n6428 , n6433 );
or ( n6435 , n6425 , n6434 );
nand ( n6436 , n6400 , n6424 );
nand ( n6437 , n6435 , n6436 );
buf ( n6438 , n6437 );
not ( n6439 , n6438 );
nand ( n6440 , n4610 , n5164 , n4331 );
not ( n6441 , n6440 );
buf ( n6442 , n6441 );
not ( n6443 , n6400 );
not ( n6444 , n6424 );
and ( n6445 , n6443 , n6444 );
not ( n6446 , n6428 );
not ( n6447 , n6433 );
and ( n6448 , n6446 , n6447 );
nor ( n6449 , n6445 , n6448 );
buf ( n6450 , n6449 );
buf ( n6451 , n6450 );
buf ( n6452 , n6451 );
buf ( n6453 , n6452 );
buf ( n6454 , n3741 );
buf ( n6455 , n6454 );
nand ( n6456 , n6442 , n6453 , n6455 );
buf ( n6457 , n6456 );
buf ( n6458 , n6457 );
not ( n6459 , n4347 );
not ( n6460 , n5152 );
not ( n6461 , n5160 );
and ( n6462 , n6460 , n6461 );
nor ( n6463 , n6462 , n4809 );
not ( n6464 , n6463 );
or ( n6465 , n6459 , n6464 );
nor ( n6466 , n4606 , n4609 );
and ( n6467 , n6466 , n5164 );
nor ( n6468 , n6467 , n5167 );
nand ( n6469 , n6465 , n6468 );
not ( n6470 , n6469 );
not ( n6471 , n6470 );
nand ( n6472 , n6452 , n6471 );
buf ( n6473 , n6472 );
nand ( n6474 , n6439 , n6458 , n6473 );
buf ( n6475 , n6474 );
buf ( n6476 , n6475 );
buf ( n6477 , n5806 );
not ( n6478 , n6477 );
nor ( n6479 , n5818 , n5813 );
buf ( n6480 , n6479 );
not ( n6481 , n6480 );
or ( n6482 , n6478 , n6481 );
buf ( n6483 , n5801 );
buf ( n6484 , n557 );
buf ( n6485 , n562 );
xor ( n6486 , n6484 , n6485 );
buf ( n6487 , n6486 );
buf ( n6488 , n6487 );
nand ( n6489 , n6483 , n6488 );
buf ( n6490 , n6489 );
buf ( n6491 , n6490 );
nand ( n6492 , n6482 , n6491 );
buf ( n6493 , n6492 );
buf ( n6494 , n6493 );
buf ( n6495 , n5855 );
not ( n6496 , n6495 );
buf ( n6497 , n4836 );
not ( n6498 , n6497 );
or ( n6499 , n6496 , n6498 );
buf ( n6500 , n4840 );
buf ( n6501 , n555 );
buf ( n6502 , n564 );
xor ( n6503 , n6501 , n6502 );
buf ( n6504 , n6503 );
buf ( n6505 , n6504 );
nand ( n6506 , n6500 , n6505 );
buf ( n6507 , n6506 );
buf ( n6508 , n6507 );
nand ( n6509 , n6499 , n6508 );
buf ( n6510 , n6509 );
buf ( n6511 , n6510 );
xor ( n6512 , n6494 , n6511 );
buf ( n6513 , n5767 );
buf ( n6514 , n5776 );
and ( n6515 , n6513 , n6514 );
buf ( n6516 , n6515 );
buf ( n6517 , n6516 );
xor ( n6518 , n6512 , n6517 );
buf ( n6519 , n6518 );
not ( n6520 , n6519 );
xor ( n6521 , n568 , n551 );
not ( n6522 , n6521 );
not ( n6523 , n3772 );
or ( n6524 , n6522 , n6523 );
nand ( n6525 , n3425 , n3427 );
nand ( n6526 , n3423 , n5867 , n6525 );
nand ( n6527 , n6524 , n6526 );
not ( n6528 , n5837 );
not ( n6529 , n850 );
or ( n6530 , n6528 , n6529 );
buf ( n6531 , n856 );
buf ( n6532 , n549 );
buf ( n6533 , n570 );
xor ( n6534 , n6532 , n6533 );
buf ( n6535 , n6534 );
buf ( n6536 , n6535 );
nand ( n6537 , n6531 , n6536 );
buf ( n6538 , n6537 );
nand ( n6539 , n6530 , n6538 );
xor ( n6540 , n6527 , n6539 );
not ( n6541 , n5893 );
not ( n6542 , n4044 );
or ( n6543 , n6541 , n6542 );
buf ( n6544 , n3743 );
buf ( n6545 , n553 );
buf ( n6546 , n566 );
xor ( n6547 , n6545 , n6546 );
buf ( n6548 , n6547 );
buf ( n6549 , n6548 );
nand ( n6550 , n6544 , n6549 );
buf ( n6551 , n6550 );
nand ( n6552 , n6543 , n6551 );
xnor ( n6553 , n6540 , n6552 );
not ( n6554 , n6553 );
or ( n6555 , n6520 , n6554 );
not ( n6556 , n6519 );
not ( n6557 , n6553 );
nand ( n6558 , n6556 , n6557 );
nand ( n6559 , n6555 , n6558 );
not ( n6560 , n5757 );
not ( n6561 , n5783 );
or ( n6562 , n6560 , n6561 );
buf ( n6563 , n5757 );
buf ( n6564 , n5783 );
or ( n6565 , n6563 , n6564 );
buf ( n6566 , n5792 );
nand ( n6567 , n6565 , n6566 );
buf ( n6568 , n6567 );
nand ( n6569 , n6562 , n6568 );
and ( n6570 , n6559 , n6569 );
not ( n6571 , n6559 );
not ( n6572 , n6569 );
and ( n6573 , n6571 , n6572 );
nor ( n6574 , n6570 , n6573 );
buf ( n6575 , n6574 );
xor ( n6576 , n5872 , n5882 );
and ( n6577 , n6576 , n5900 );
and ( n6578 , n5872 , n5882 );
or ( n6579 , n6577 , n6578 );
buf ( n6580 , n6579 );
buf ( n6581 , n6580 );
not ( n6582 , n6581 );
buf ( n6583 , n6582 );
buf ( n6584 , n6583 );
not ( n6585 , n905 );
not ( n6586 , n5763 );
or ( n6587 , n6585 , n6586 );
and ( n6588 , n574 , n545 );
not ( n6589 , n574 );
not ( n6590 , n545 );
and ( n6591 , n6589 , n6590 );
nor ( n6592 , n6588 , n6591 );
nand ( n6593 , n6592 , n575 );
nand ( n6594 , n6587 , n6593 );
xor ( n6595 , n561 , n562 );
buf ( n6596 , n6595 );
buf ( n6597 , n559 );
nand ( n6598 , n6596 , n6597 );
buf ( n6599 , n6598 );
xor ( n6600 , n6594 , n6599 );
buf ( n6601 , n5879 );
not ( n6602 , n6601 );
buf ( n6603 , n884 );
not ( n6604 , n6603 );
or ( n6605 , n6602 , n6604 );
buf ( n6606 , n888 );
buf ( n6607 , n547 );
buf ( n6608 , n572 );
xor ( n6609 , n6607 , n6608 );
buf ( n6610 , n6609 );
buf ( n6611 , n6610 );
nand ( n6612 , n6606 , n6611 );
buf ( n6613 , n6612 );
buf ( n6614 , n6613 );
nand ( n6615 , n6605 , n6614 );
buf ( n6616 , n6615 );
xor ( n6617 , n6600 , n6616 );
buf ( n6618 , n6617 );
and ( n6619 , n6584 , n6618 );
not ( n6620 , n6584 );
buf ( n6621 , n6617 );
not ( n6622 , n6621 );
buf ( n6623 , n6622 );
buf ( n6624 , n6623 );
and ( n6625 , n6620 , n6624 );
nor ( n6626 , n6619 , n6625 );
buf ( n6627 , n6626 );
buf ( n6628 , n6627 );
xor ( n6629 , n5823 , n5844 );
and ( n6630 , n6629 , n5862 );
and ( n6631 , n5823 , n5844 );
or ( n6632 , n6630 , n6631 );
buf ( n6633 , n6632 );
buf ( n6634 , n6633 );
and ( n6635 , n6628 , n6634 );
not ( n6636 , n6628 );
buf ( n6637 , n6633 );
not ( n6638 , n6637 );
buf ( n6639 , n6638 );
buf ( n6640 , n6639 );
and ( n6641 , n6636 , n6640 );
nor ( n6642 , n6635 , n6641 );
buf ( n6643 , n6642 );
buf ( n6644 , n6643 );
and ( n6645 , n6575 , n6644 );
not ( n6646 , n6575 );
buf ( n6647 , n6643 );
not ( n6648 , n6647 );
buf ( n6649 , n6648 );
buf ( n6650 , n6649 );
and ( n6651 , n6646 , n6650 );
nor ( n6652 , n6645 , n6651 );
buf ( n6653 , n6652 );
xor ( n6654 , n5865 , n5903 );
and ( n6655 , n6654 , n5932 );
and ( n6656 , n5865 , n5903 );
or ( n6657 , n6655 , n6656 );
buf ( n6658 , n6657 );
xor ( n6659 , n6653 , n6658 );
buf ( n6660 , n6659 );
xor ( n6661 , n6181 , n6187 );
and ( n6662 , n6661 , n6395 );
and ( n6663 , n6181 , n6187 );
or ( n6664 , n6662 , n6663 );
buf ( n6665 , n6664 );
buf ( n6666 , n6665 );
xor ( n6667 , n6660 , n6666 );
not ( n6668 , n5751 );
nand ( n6669 , n6668 , n5793 );
not ( n6670 , n6669 );
not ( n6671 , n5934 );
or ( n6672 , n6670 , n6671 );
nand ( n6673 , n5752 , n5794 );
nand ( n6674 , n6672 , n6673 );
xor ( n6675 , n6206 , n6271 );
and ( n6676 , n6675 , n6392 );
and ( n6677 , n6206 , n6271 );
or ( n6678 , n6676 , n6677 );
buf ( n6679 , n6678 );
xor ( n6680 , n6674 , n6679 );
buf ( n6681 , n6367 );
not ( n6682 , n6681 );
buf ( n6683 , n6682 );
nand ( n6684 , n6683 , n6305 );
nand ( n6685 , n6684 , n6390 );
buf ( n6686 , n6685 );
buf ( n6687 , n6305 );
not ( n6688 , n6687 );
buf ( n6689 , n6367 );
nand ( n6690 , n6688 , n6689 );
buf ( n6691 , n6690 );
buf ( n6692 , n6691 );
nand ( n6693 , n6686 , n6692 );
buf ( n6694 , n6693 );
buf ( n6695 , n6694 );
buf ( n6696 , n577 );
buf ( n6697 , n578 );
xor ( n6698 , n6696 , n6697 );
buf ( n6699 , n6698 );
buf ( n6700 , n6699 );
buf ( n6701 , n559 );
and ( n6702 , n6700 , n6701 );
buf ( n6703 , n6702 );
buf ( n6704 , n6703 );
not ( n6705 , n591 );
buf ( n6706 , n545 );
buf ( n6707 , n590 );
xor ( n6708 , n6706 , n6707 );
buf ( n6709 , n6708 );
not ( n6710 , n6709 );
or ( n6711 , n6705 , n6710 );
nand ( n6712 , n6243 , n984 );
nand ( n6713 , n6711 , n6712 );
buf ( n6714 , n6713 );
xor ( n6715 , n6704 , n6714 );
buf ( n6716 , n6279 );
not ( n6717 , n6716 );
buf ( n6718 , n4286 );
not ( n6719 , n6718 );
or ( n6720 , n6717 , n6719 );
buf ( n6721 , n547 );
buf ( n6722 , n588 );
xor ( n6723 , n6721 , n6722 );
buf ( n6724 , n6723 );
nand ( n6725 , n6724 , n4556 );
buf ( n6726 , n6725 );
nand ( n6727 , n6720 , n6726 );
buf ( n6728 , n6727 );
buf ( n6729 , n6728 );
xor ( n6730 , n6715 , n6729 );
buf ( n6731 , n6730 );
buf ( n6732 , n6731 );
nor ( n6733 , n6304 , n6281 );
or ( n6734 , n6733 , n6291 );
nand ( n6735 , n6304 , n6281 );
nand ( n6736 , n6734 , n6735 );
buf ( n6737 , n6736 );
xor ( n6738 , n6732 , n6737 );
xor ( n6739 , n6316 , n6333 );
and ( n6740 , n6739 , n6365 );
and ( n6741 , n6316 , n6333 );
or ( n6742 , n6740 , n6741 );
buf ( n6743 , n6742 );
buf ( n6744 , n6743 );
xor ( n6745 , n6738 , n6744 );
buf ( n6746 , n6745 );
buf ( n6747 , n6746 );
xor ( n6748 , n6695 , n6747 );
not ( n6749 , n6257 );
not ( n6750 , n6263 );
not ( n6751 , n6750 );
or ( n6752 , n6749 , n6751 );
nand ( n6753 , n6262 , n6252 );
nand ( n6754 , n6752 , n6753 );
not ( n6755 , n6754 );
buf ( n6756 , n6286 );
not ( n6757 , n6756 );
and ( n6758 , n3662 , n2120 );
buf ( n6759 , n6758 );
not ( n6760 , n6759 );
or ( n6761 , n6757 , n6760 );
buf ( n6762 , n2123 );
buf ( n6763 , n551 );
buf ( n6764 , n584 );
xor ( n6765 , n6763 , n6764 );
buf ( n6766 , n6765 );
buf ( n6767 , n6766 );
nand ( n6768 , n6762 , n6767 );
buf ( n6769 , n6768 );
buf ( n6770 , n6769 );
nand ( n6771 , n6761 , n6770 );
buf ( n6772 , n6771 );
buf ( n6773 , n6300 );
not ( n6774 , n6773 );
buf ( n6775 , n4506 );
not ( n6776 , n6775 );
or ( n6777 , n6774 , n6776 );
buf ( n6778 , n4211 );
buf ( n6779 , n553 );
buf ( n6780 , n582 );
xor ( n6781 , n6779 , n6780 );
buf ( n6782 , n6781 );
buf ( n6783 , n6782 );
nand ( n6784 , n6778 , n6783 );
buf ( n6785 , n6784 );
buf ( n6786 , n6785 );
nand ( n6787 , n6777 , n6786 );
buf ( n6788 , n6787 );
buf ( n6789 , n6788 );
not ( n6790 , n6789 );
buf ( n6791 , n6790 );
and ( n6792 , n6772 , n6791 );
not ( n6793 , n6772 );
and ( n6794 , n6793 , n6788 );
or ( n6795 , n6792 , n6794 );
not ( n6796 , n1036 );
buf ( n6797 , n549 );
buf ( n6798 , n586 );
xor ( n6799 , n6797 , n6798 );
buf ( n6800 , n6799 );
not ( n6801 , n6800 );
or ( n6802 , n6796 , n6801 );
nand ( n6803 , n1175 , n1170 , n6313 );
nand ( n6804 , n6802 , n6803 );
not ( n6805 , n6804 );
and ( n6806 , n6795 , n6805 );
not ( n6807 , n6795 );
and ( n6808 , n6807 , n6804 );
or ( n6809 , n6806 , n6808 );
buf ( n6810 , n6358 );
not ( n6811 , n6810 );
buf ( n6812 , n6350 );
not ( n6813 , n6812 );
or ( n6814 , n6811 , n6813 );
buf ( n6815 , n5997 );
buf ( n6816 , n557 );
buf ( n6817 , n578 );
xor ( n6818 , n6816 , n6817 );
buf ( n6819 , n6818 );
buf ( n6820 , n6819 );
nand ( n6821 , n6815 , n6820 );
buf ( n6822 , n6821 );
buf ( n6823 , n6822 );
nand ( n6824 , n6814 , n6823 );
buf ( n6825 , n6824 );
buf ( n6826 , n6250 );
buf ( n6827 , n6234 );
and ( n6828 , n6826 , n6827 );
buf ( n6829 , n6828 );
and ( n6830 , n6825 , n6829 );
not ( n6831 , n6825 );
not ( n6832 , n6829 );
and ( n6833 , n6831 , n6832 );
or ( n6834 , n6830 , n6833 );
buf ( n6835 , n6326 );
not ( n6836 , n6835 );
buf ( n6837 , n5060 );
not ( n6838 , n6837 );
or ( n6839 , n6836 , n6838 );
not ( n6840 , n580 );
not ( n6841 , n1031 );
or ( n6842 , n6840 , n6841 );
not ( n6843 , n580 );
nand ( n6844 , n6843 , n555 );
nand ( n6845 , n6842 , n6844 );
nand ( n6846 , n6845 , n5065 );
buf ( n6847 , n6846 );
nand ( n6848 , n6839 , n6847 );
buf ( n6849 , n6848 );
not ( n6850 , n6849 );
and ( n6851 , n6834 , n6850 );
not ( n6852 , n6834 );
and ( n6853 , n6852 , n6849 );
nor ( n6854 , n6851 , n6853 );
not ( n6855 , n6854 );
and ( n6856 , n6809 , n6855 );
not ( n6857 , n6809 );
and ( n6858 , n6857 , n6854 );
nor ( n6859 , n6856 , n6858 );
not ( n6860 , n6859 );
or ( n6861 , n6755 , n6860 );
or ( n6862 , n6754 , n6859 );
nand ( n6863 , n6861 , n6862 );
buf ( n6864 , n6863 );
xor ( n6865 , n6748 , n6864 );
buf ( n6866 , n6865 );
xor ( n6867 , n6680 , n6866 );
buf ( n6868 , n6867 );
xor ( n6869 , n6667 , n6868 );
buf ( n6870 , n6869 );
buf ( n6871 , n6870 );
xor ( n6872 , n5940 , n6152 );
and ( n6873 , n6872 , n6398 );
and ( n6874 , n5940 , n6152 );
or ( n6875 , n6873 , n6874 );
buf ( n6876 , n6875 );
buf ( n6877 , n6876 );
nor ( n6878 , n6871 , n6877 );
buf ( n6879 , n6878 );
buf ( n6880 , n6879 );
not ( n6881 , n6880 );
buf ( n6882 , n6881 );
buf ( n6883 , n6882 );
buf ( n6884 , n6870 );
buf ( n6885 , n6876 );
nand ( n6886 , n6884 , n6885 );
buf ( n6887 , n6886 );
buf ( n6888 , n6887 );
buf ( n6889 , n6888 );
buf ( n6890 , n6889 );
buf ( n6891 , n6890 );
nand ( n6892 , n6883 , n6891 );
buf ( n6893 , n6892 );
buf ( n6894 , n6893 );
not ( n6895 , n6894 );
buf ( n6896 , n6895 );
buf ( n6897 , n6896 );
and ( n6898 , n6476 , n6897 );
not ( n6899 , n6476 );
buf ( n6900 , n6893 );
and ( n6901 , n6899 , n6900 );
nor ( n6902 , n6898 , n6901 );
buf ( n6903 , n6902 );
not ( n6904 , n6903 );
not ( n6905 , n2276 );
not ( n6906 , n6905 );
not ( n6907 , n6906 );
buf ( n6908 , n3167 );
and ( n6909 , n6908 , n1681 );
not ( n6910 , n6908 );
and ( n6911 , n6910 , n554 );
or ( n6912 , n6909 , n6911 );
not ( n6913 , n6912 );
or ( n6914 , n6907 , n6913 );
not ( n6915 , n554 );
not ( n6916 , n3265 );
or ( n6917 , n6915 , n6916 );
not ( n6918 , n3265 );
nand ( n6919 , n6918 , n1681 );
nand ( n6920 , n6917 , n6919 );
nand ( n6921 , n6920 , n3118 );
nand ( n6922 , n6914 , n6921 );
not ( n6923 , n3213 );
not ( n6924 , n6923 );
not ( n6925 , n548 );
not ( n6926 , n1621 );
or ( n6927 , n6925 , n6926 );
nand ( n6928 , n1624 , n5279 );
nand ( n6929 , n6927 , n6928 );
not ( n6930 , n6929 );
or ( n6931 , n6924 , n6930 );
not ( n6932 , n1838 );
not ( n6933 , n6932 );
not ( n6934 , n5279 );
or ( n6935 , n6933 , n6934 );
nand ( n6936 , n548 , n1652 );
nand ( n6937 , n6935 , n6936 );
nor ( n6938 , n5289 , n5293 );
buf ( n6939 , n6938 );
nand ( n6940 , n6937 , n6939 );
nand ( n6941 , n6931 , n6940 );
buf ( n6942 , n1854 );
not ( n6943 , n6942 );
not ( n6944 , n6943 );
xor ( n6945 , n547 , n548 );
and ( n6946 , n6945 , n546 );
not ( n6947 , n6946 );
or ( n6948 , n6944 , n6947 );
not ( n6949 , n546 );
nand ( n6950 , n1791 , n6945 , n6949 );
not ( n6951 , n546 );
nand ( n6952 , n6951 , n548 , n547 );
not ( n6953 , n6952 );
and ( n6954 , n1664 , n6953 );
not ( n6955 , n1664 );
not ( n6956 , n546 );
nor ( n6957 , n6956 , n548 , n547 );
and ( n6958 , n6955 , n6957 );
nor ( n6959 , n6954 , n6958 );
and ( n6960 , n6950 , n6959 );
nand ( n6961 , n6948 , n6960 );
or ( n6962 , n547 , n548 );
not ( n6963 , n6962 );
not ( n6964 , n1664 );
or ( n6965 , n6963 , n6964 );
nand ( n6966 , n547 , n548 );
and ( n6967 , n6966 , n546 );
nand ( n6968 , n6965 , n6967 );
not ( n6969 , n6968 );
and ( n6970 , n6961 , n6969 );
not ( n6971 , n6961 );
and ( n6972 , n6971 , n6968 );
nor ( n6973 , n6970 , n6972 );
xor ( n6974 , n6941 , n6973 );
not ( n6975 , n3068 );
not ( n6976 , n550 );
not ( n6977 , n2944 );
or ( n6978 , n6976 , n6977 );
nand ( n6979 , n1772 , n3073 );
nand ( n6980 , n6978 , n6979 );
not ( n6981 , n6980 );
or ( n6982 , n6975 , n6981 );
not ( n6983 , n550 );
not ( n6984 , n2220 );
or ( n6985 , n6983 , n6984 );
nand ( n6986 , n1732 , n3073 );
nand ( n6987 , n6985 , n6986 );
nand ( n6988 , n6987 , n5268 );
nand ( n6989 , n6982 , n6988 );
and ( n6990 , n6974 , n6989 );
and ( n6991 , n6941 , n6973 );
or ( n6992 , n6990 , n6991 );
xor ( n6993 , n6922 , n6992 );
not ( n6994 , n6923 );
and ( n6995 , n1732 , n5279 );
not ( n6996 , n1732 );
and ( n6997 , n6996 , n548 );
or ( n6998 , n6995 , n6997 );
not ( n6999 , n6998 );
or ( n7000 , n6994 , n6999 );
nand ( n7001 , n6929 , n6939 );
nand ( n7002 , n7000 , n7001 );
not ( n7003 , n5268 );
not ( n7004 , n6980 );
or ( n7005 , n7003 , n7004 );
and ( n7006 , n2251 , n550 );
not ( n7007 , n2251 );
and ( n7008 , n7007 , n3073 );
nor ( n7009 , n7006 , n7008 );
nand ( n7010 , n7009 , n3068 );
nand ( n7011 , n7005 , n7010 );
xor ( n7012 , n7002 , n7011 );
not ( n7013 , n2265 );
not ( n7014 , n552 );
not ( n7015 , n3036 );
not ( n7016 , n7015 );
or ( n7017 , n7014 , n7016 );
not ( n7018 , n552 );
nand ( n7019 , n7018 , n3036 );
nand ( n7020 , n7017 , n7019 );
not ( n7021 , n7020 );
or ( n7022 , n7013 , n7021 );
and ( n7023 , n552 , n2982 );
not ( n7024 , n552 );
and ( n7025 , n7024 , n2981 );
or ( n7026 , n7023 , n7025 );
not ( n7027 , n7026 );
not ( n7028 , n3064 );
or ( n7029 , n7027 , n7028 );
nand ( n7030 , n7022 , n7029 );
xor ( n7031 , n7012 , n7030 );
xor ( n7032 , n6993 , n7031 );
not ( n7033 , n3068 );
not ( n7034 , n6987 );
or ( n7035 , n7033 , n7034 );
nand ( n7036 , n5263 , n5268 );
nand ( n7037 , n7035 , n7036 );
not ( n7038 , n2276 );
not ( n7039 , n5191 );
or ( n7040 , n7038 , n7039 );
not ( n7041 , n554 );
not ( n7042 , n7015 );
or ( n7043 , n7041 , n7042 );
nand ( n7044 , n3036 , n1681 );
nand ( n7045 , n7043 , n7044 );
nand ( n7046 , n7045 , n3118 );
nand ( n7047 , n7040 , n7046 );
xor ( n7048 , n7037 , n7047 );
not ( n7049 , n3064 );
not ( n7050 , n5306 );
or ( n7051 , n7049 , n7050 );
not ( n7052 , n552 );
not ( n7053 , n2252 );
or ( n7054 , n7052 , n7053 );
not ( n7055 , n552 );
nand ( n7056 , n7055 , n3198 );
nand ( n7057 , n7054 , n7056 );
nand ( n7058 , n7057 , n2265 );
nand ( n7059 , n7051 , n7058 );
and ( n7060 , n7048 , n7059 );
and ( n7061 , n7037 , n7047 );
or ( n7062 , n7060 , n7061 );
not ( n7063 , n1659 );
not ( n7064 , n5205 );
or ( n7065 , n7063 , n7064 );
or ( n7066 , n1625 , n3264 );
nand ( n7067 , n3264 , n1625 );
nand ( n7068 , n7066 , n7067 );
buf ( n7069 , n1594 );
nand ( n7070 , n7068 , n7069 );
nand ( n7071 , n7065 , n7070 );
not ( n7072 , n6945 );
nor ( n7073 , n7072 , n1687 );
not ( n7074 , n5293 );
not ( n7075 , n6937 );
or ( n7076 , n7074 , n7075 );
nand ( n7077 , n5281 , n6938 );
nand ( n7078 , n7076 , n7077 );
xor ( n7079 , n7073 , n7078 );
and ( n7080 , n5296 , n5274 );
xor ( n7081 , n7079 , n7080 );
xor ( n7082 , n7071 , n7081 );
not ( n7083 , n1739 );
not ( n7084 , n5252 );
or ( n7085 , n7083 , n7084 );
not ( n7086 , n558 );
or ( n7087 , n566 , n582 );
or ( n7088 , n567 , n583 );
nand ( n7089 , n7087 , n7088 );
not ( n7090 , n7089 );
not ( n7091 , n565 );
not ( n7092 , n581 );
and ( n7093 , n7091 , n7092 );
nor ( n7094 , n7093 , n5220 );
nand ( n7095 , n7090 , n7094 );
not ( n7096 , n7095 );
not ( n7097 , n7096 );
not ( n7098 , n5233 );
or ( n7099 , n7097 , n7098 );
not ( n7100 , n565 );
not ( n7101 , n581 );
and ( n7102 , n7100 , n7101 );
nor ( n7103 , n564 , n580 );
nor ( n7104 , n7102 , n7103 );
not ( n7105 , n7104 );
not ( n7106 , n3252 );
or ( n7107 , n7105 , n7106 );
not ( n7108 , n7103 );
not ( n7109 , n3257 );
and ( n7110 , n7108 , n7109 );
nor ( n7111 , n7110 , n5243 );
nand ( n7112 , n7107 , n7111 );
not ( n7113 , n7112 );
nand ( n7114 , n7099 , n7113 );
not ( n7115 , n7114 );
and ( n7116 , n563 , n579 );
nor ( n7117 , n563 , n579 );
nor ( n7118 , n7116 , n7117 );
buf ( n7119 , n7118 );
nand ( n7120 , n7115 , n7119 );
not ( n7121 , n7119 );
nand ( n7122 , n7114 , n7121 );
nand ( n7123 , n7120 , n7122 );
buf ( n7124 , n7123 );
not ( n7125 , n7124 );
not ( n7126 , n7125 );
or ( n7127 , n7086 , n7126 );
not ( n7128 , n7122 );
not ( n7129 , n7120 );
or ( n7130 , n7128 , n7129 );
nand ( n7131 , n7130 , n1736 );
nand ( n7132 , n7127 , n7131 );
nand ( n7133 , n7132 , n559 );
nand ( n7134 , n7085 , n7133 );
and ( n7135 , n7082 , n7134 );
and ( n7136 , n7071 , n7081 );
or ( n7137 , n7135 , n7136 );
xor ( n7138 , n7062 , n7137 );
not ( n7139 , n5299 );
not ( n7140 , n7026 );
or ( n7141 , n7139 , n7140 );
nand ( n7142 , n7057 , n3064 );
nand ( n7143 , n7141 , n7142 );
not ( n7144 , n1659 );
not ( n7145 , n7068 );
or ( n7146 , n7144 , n7145 );
buf ( n7147 , n5246 );
nand ( n7148 , n7147 , n1625 );
not ( n7149 , n7148 );
not ( n7150 , n7147 );
nand ( n7151 , n7150 , n556 );
not ( n7152 , n7151 );
or ( n7153 , n7149 , n7152 );
nand ( n7154 , n7153 , n7069 );
nand ( n7155 , n7146 , n7154 );
xor ( n7156 , n7143 , n7155 );
xor ( n7157 , n7073 , n7078 );
and ( n7158 , n7157 , n7080 );
and ( n7159 , n7073 , n7078 );
or ( n7160 , n7158 , n7159 );
xor ( n7161 , n7156 , n7160 );
and ( n7162 , n7138 , n7161 );
and ( n7163 , n7062 , n7137 );
or ( n7164 , n7162 , n7163 );
xor ( n7165 , n7032 , n7164 );
xor ( n7166 , n7143 , n7155 );
and ( n7167 , n7166 , n7160 );
and ( n7168 , n7143 , n7155 );
or ( n7169 , n7167 , n7168 );
xor ( n7170 , n545 , n546 );
and ( n7171 , n1664 , n7170 );
not ( n7172 , n546 );
not ( n7173 , n1838 );
or ( n7174 , n7172 , n7173 );
nand ( n7175 , n1837 , n6949 );
nand ( n7176 , n7174 , n7175 );
not ( n7177 , n7176 );
not ( n7178 , n6945 );
not ( n7179 , n7178 );
not ( n7180 , n7179 );
or ( n7181 , n7177 , n7180 );
and ( n7182 , n1791 , n6953 );
not ( n7183 , n1791 );
not ( n7184 , n546 );
nor ( n7185 , n7184 , n547 , n548 );
and ( n7186 , n7183 , n7185 );
nor ( n7187 , n7182 , n7186 );
nand ( n7188 , n7181 , n7187 );
xor ( n7189 , n7171 , n7188 );
and ( n7190 , n6943 , n6946 );
not ( n7191 , n6950 );
not ( n7192 , n6959 );
nor ( n7193 , n7190 , n7191 , n7192 );
nor ( n7194 , n7193 , n6968 );
xor ( n7195 , n7189 , n7194 );
not ( n7196 , n7147 );
nand ( n7197 , n7196 , n3109 );
not ( n7198 , n1625 );
nand ( n7199 , n7198 , n1596 );
not ( n7200 , n7199 );
not ( n7201 , n7124 );
nand ( n7202 , n7200 , n7201 );
nand ( n7203 , n7147 , n3112 );
nand ( n7204 , n7124 , n2956 );
nand ( n7205 , n7197 , n7202 , n7203 , n7204 );
xor ( n7206 , n7195 , n7205 );
not ( n7207 , n1739 );
not ( n7208 , n558 );
xor ( n7209 , n562 , n578 );
nor ( n7210 , n7095 , n7117 );
not ( n7211 , n7210 );
not ( n7212 , n3034 );
or ( n7213 , n7211 , n7212 );
not ( n7214 , n7117 );
not ( n7215 , n7214 );
not ( n7216 , n7112 );
or ( n7217 , n7215 , n7216 );
nand ( n7218 , n563 , n579 );
nand ( n7219 , n7217 , n7218 );
not ( n7220 , n7219 );
nand ( n7221 , n7213 , n7220 );
xor ( n7222 , n7209 , n7221 );
not ( n7223 , n7222 );
not ( n7224 , n7223 );
or ( n7225 , n7208 , n7224 );
nand ( n7226 , n7222 , n1736 );
nand ( n7227 , n7225 , n7226 );
not ( n7228 , n7227 );
or ( n7229 , n7207 , n7228 );
not ( n7230 , n558 );
or ( n7231 , n577 , n561 );
nand ( n7232 , n577 , n561 );
nand ( n7233 , n7231 , n7232 );
not ( n7234 , n7233 );
not ( n7235 , n7234 );
not ( n7236 , n562 );
not ( n7237 , n578 );
and ( n7238 , n7236 , n7237 );
nor ( n7239 , n7238 , n7117 );
not ( n7240 , n580 );
nand ( n7241 , n5811 , n7240 );
and ( n7242 , n7239 , n3242 , n3256 , n7241 );
not ( n7243 , n7242 );
not ( n7244 , n5233 );
or ( n7245 , n7243 , n7244 );
not ( n7246 , n3252 );
not ( n7247 , n7104 );
or ( n7248 , n7246 , n7247 );
nand ( n7249 , n7248 , n7111 );
not ( n7250 , n562 );
not ( n7251 , n578 );
and ( n7252 , n7250 , n7251 );
nor ( n7253 , n7252 , n7117 );
and ( n7254 , n7249 , n7253 );
nor ( n7255 , n562 , n578 );
or ( n7256 , n7255 , n7218 );
nand ( n7257 , n562 , n578 );
nand ( n7258 , n7256 , n7257 );
nor ( n7259 , n7254 , n7258 );
nand ( n7260 , n7245 , n7259 );
not ( n7261 , n7260 );
not ( n7262 , n7261 );
or ( n7263 , n7235 , n7262 );
not ( n7264 , n7232 );
nor ( n7265 , n561 , n577 );
nor ( n7266 , n7264 , n7265 );
not ( n7267 , n7266 );
nand ( n7268 , n7267 , n7260 );
nand ( n7269 , n7263 , n7268 );
not ( n7270 , n7269 );
not ( n7271 , n7270 );
or ( n7272 , n7230 , n7271 );
and ( n7273 , n7260 , n7266 );
not ( n7274 , n7260 );
and ( n7275 , n7274 , n7233 );
nor ( n7276 , n7273 , n7275 );
nand ( n7277 , n7276 , n1736 );
nand ( n7278 , n7272 , n7277 );
nand ( n7279 , n7278 , n559 );
nand ( n7280 , n7229 , n7279 );
xor ( n7281 , n7206 , n7280 );
xor ( n7282 , n7169 , n7281 );
not ( n7283 , n559 );
not ( n7284 , n7227 );
or ( n7285 , n7283 , n7284 );
nand ( n7286 , n7132 , n1739 );
nand ( n7287 , n7285 , n7286 );
not ( n7288 , n3118 );
not ( n7289 , n6912 );
or ( n7290 , n7288 , n7289 );
nand ( n7291 , n7045 , n6906 );
nand ( n7292 , n7290 , n7291 );
xor ( n7293 , n7287 , n7292 );
xor ( n7294 , n6941 , n6973 );
xor ( n7295 , n7294 , n6989 );
and ( n7296 , n7293 , n7295 );
and ( n7297 , n7287 , n7292 );
or ( n7298 , n7296 , n7297 );
xor ( n7299 , n7282 , n7298 );
xor ( n7300 , n7165 , n7299 );
buf ( n7301 , n7300 );
xor ( n7302 , n7287 , n7292 );
xor ( n7303 , n7302 , n7295 );
xor ( n7304 , n5270 , n5297 );
and ( n7305 , n7304 , n5310 );
and ( n7306 , n5270 , n5297 );
or ( n7307 , n7305 , n7306 );
xor ( n7308 , n7037 , n7047 );
xor ( n7309 , n7308 , n7059 );
xor ( n7310 , n7307 , n7309 );
xor ( n7311 , n5193 , n5197 );
and ( n7312 , n7311 , n5209 );
and ( n7313 , n5193 , n5197 );
or ( n7314 , n7312 , n7313 );
and ( n7315 , n7310 , n7314 );
and ( n7316 , n7307 , n7309 );
or ( n7317 , n7315 , n7316 );
xor ( n7318 , n7303 , n7317 );
xor ( n7319 , n7062 , n7137 );
xor ( n7320 , n7319 , n7161 );
and ( n7321 , n7318 , n7320 );
and ( n7322 , n7303 , n7317 );
or ( n7323 , n7321 , n7322 );
nand ( n7324 , n7301 , n7323 );
not ( n7325 , n7324 );
nor ( n7326 , n7301 , n7323 );
nor ( n7327 , n7325 , n7326 );
not ( n7328 , n5180 );
not ( n7329 , n5318 );
or ( n7330 , n7328 , n7329 );
nand ( n7331 , n3181 , n3280 );
nand ( n7332 , n7330 , n7331 );
or ( n7333 , n5329 , n7332 );
xor ( n7334 , n7071 , n7081 );
xor ( n7335 , n7334 , n7134 );
xor ( n7336 , n5256 , n5311 );
and ( n7337 , n7336 , n5316 );
and ( n7338 , n5256 , n5311 );
or ( n7339 , n7337 , n7338 );
xor ( n7340 , n7335 , n7339 );
xor ( n7341 , n7307 , n7309 );
xor ( n7342 , n7341 , n7314 );
xor ( n7343 , n7340 , n7342 );
xor ( n7344 , n5210 , n5214 );
and ( n7345 , n7344 , n5317 );
and ( n7346 , n5210 , n5214 );
or ( n7347 , n7345 , n7346 );
nor ( n7348 , n7343 , n7347 );
nor ( n7349 , n7348 , n5321 );
nand ( n7350 , n7333 , n7349 );
xor ( n7351 , n7303 , n7317 );
xor ( n7352 , n7351 , n7320 );
xor ( n7353 , n7335 , n7339 );
and ( n7354 , n7353 , n7342 );
and ( n7355 , n7335 , n7339 );
or ( n7356 , n7354 , n7355 );
nand ( n7357 , n7352 , n7356 );
buf ( n7358 , n7343 );
nand ( n7359 , n7358 , n7347 );
nand ( n7360 , n7350 , n7357 , n7359 );
or ( n7361 , n7352 , n7356 );
nand ( n7362 , n7360 , n7361 );
and ( n7363 , n7327 , n7362 );
not ( n7364 , n7327 );
not ( n7365 , n7362 );
and ( n7366 , n7364 , n7365 );
nor ( n7367 , n7363 , n7366 );
not ( n7368 , n7367 );
nand ( n7369 , n6904 , n7368 );
not ( n7370 , n7369 );
nand ( n7371 , n6903 , n7367 );
not ( n7372 , n7371 );
nor ( n7373 , n7370 , n7372 );
not ( n7374 , n7373 );
not ( n7375 , n7374 );
not ( n7376 , n7375 );
not ( n7377 , n5350 );
not ( n7378 , n5345 );
or ( n7379 , n7377 , n7378 );
nand ( n7380 , n7379 , n4797 );
not ( n7381 , n7380 );
and ( n7382 , n7381 , n4723 );
not ( n7383 , n7382 );
not ( n7384 , n7383 );
not ( n7385 , n5322 );
not ( n7386 , n7332 );
or ( n7387 , n7385 , n7386 );
nand ( n7388 , n3282 , n5326 );
nand ( n7389 , n3367 , n7388 , n5322 );
nand ( n7390 , n7387 , n7389 );
not ( n7391 , n7348 );
nand ( n7392 , n7391 , n7359 );
xnor ( n7393 , n7390 , n7392 );
not ( n7394 , n7393 );
not ( n7395 , n6454 );
not ( n7396 , n6441 );
or ( n7397 , n7395 , n7396 );
nand ( n7398 , n7397 , n6470 );
or ( n7399 , n6433 , n6428 );
not ( n7400 , n7399 );
not ( n7401 , n6434 );
nor ( n7402 , n7400 , n7401 );
and ( n7403 , n7398 , n7402 );
not ( n7404 , n7398 );
not ( n7405 , n7401 );
nand ( n7406 , n7399 , n7405 );
and ( n7407 , n7404 , n7406 );
nor ( n7408 , n7403 , n7407 );
nor ( n7409 , n7394 , n7408 );
not ( n7410 , n7409 );
nor ( n7411 , n6400 , n6424 );
buf ( n7412 , n7411 );
not ( n7413 , n7412 );
buf ( n7414 , n6436 );
nand ( n7415 , n7413 , n7414 );
buf ( n7416 , n7415 );
not ( n7417 , n7416 );
not ( n7418 , n7417 );
nand ( n7419 , n6471 , n7399 );
nand ( n7420 , n6454 , n7399 );
not ( n7421 , n7420 );
nand ( n7422 , n7421 , n6441 );
nand ( n7423 , n7419 , n7422 , n7405 );
not ( n7424 , n7423 );
or ( n7425 , n7418 , n7424 );
nand ( n7426 , n7419 , n7416 , n7422 , n7405 );
nand ( n7427 , n7425 , n7426 );
not ( n7428 , n7391 );
not ( n7429 , n7390 );
or ( n7430 , n7428 , n7429 );
buf ( n7431 , n7359 );
nand ( n7432 , n7430 , n7431 );
nand ( n7433 , n7361 , n7357 );
not ( n7434 , n7433 );
and ( n7435 , n7432 , n7434 );
not ( n7436 , n7432 );
and ( n7437 , n7436 , n7433 );
nor ( n7438 , n7435 , n7437 );
nand ( n7439 , n7427 , n7438 );
and ( n7440 , n7410 , n7439 );
buf ( n7441 , n4666 );
nand ( n7442 , n7384 , n7440 , n7441 );
not ( n7443 , n7439 );
nand ( n7444 , n7408 , n7394 );
not ( n7445 , n7444 );
not ( n7446 , n7445 );
or ( n7447 , n7443 , n7446 );
not ( n7448 , n7438 );
not ( n7449 , n7427 );
nand ( n7450 , n7448 , n7449 );
nand ( n7451 , n7447 , n7450 );
not ( n7452 , n7451 );
not ( n7453 , n4735 );
not ( n7454 , n7381 );
or ( n7455 , n7453 , n7454 );
nor ( n7456 , n3368 , n4616 );
nand ( n7457 , n5345 , n5350 );
and ( n7458 , n7456 , n7457 );
nor ( n7459 , n7458 , n5339 );
nand ( n7460 , n7455 , n7459 );
buf ( n7461 , n7460 );
not ( n7462 , n7439 );
nor ( n7463 , n7394 , n7408 );
nor ( n7464 , n7462 , n7463 );
nand ( n7465 , n7461 , n7464 );
nand ( n7466 , n7442 , n7452 , n7465 );
not ( n7467 , n7466 );
not ( n7468 , n7467 );
or ( n7469 , n7376 , n7468 );
not ( n7470 , n7373 );
nand ( n7471 , n7470 , n7466 );
nand ( n7472 , n7469 , n7471 );
not ( n7473 , n7472 );
not ( n7474 , n577 );
and ( n7475 , n7473 , n7474 );
and ( n7476 , n7472 , n577 );
nor ( n7477 , n7475 , n7476 );
not ( n7478 , n7463 );
not ( n7479 , n7445 );
nand ( n7480 , n7478 , n7479 );
and ( n7481 , n4706 , n4771 );
not ( n7482 , n7481 );
not ( n7483 , n7381 );
or ( n7484 , n7482 , n7483 );
not ( n7485 , n4734 );
and ( n7486 , n7381 , n7485 );
not ( n7487 , n7456 );
not ( n7488 , n5351 );
or ( n7489 , n7487 , n7488 );
not ( n7490 , n5339 );
nand ( n7491 , n7489 , n7490 );
nor ( n7492 , n7486 , n7491 );
nand ( n7493 , n7484 , n7492 );
and ( n7494 , n7480 , n7493 );
not ( n7495 , n7480 );
not ( n7496 , n7493 );
and ( n7497 , n7495 , n7496 );
nor ( n7498 , n7494 , n7497 );
not ( n7499 , n7498 );
nor ( n7500 , n7499 , n579 );
not ( n7501 , n7462 );
nand ( n7502 , n7501 , n7450 );
and ( n7503 , n7502 , n6345 );
not ( n7504 , n7503 );
nand ( n7505 , n7382 , n7410 , n7441 );
nand ( n7506 , n7478 , n7460 );
nand ( n7507 , n7505 , n7506 , n7479 );
not ( n7508 , n7507 );
not ( n7509 , n7508 );
or ( n7510 , n7504 , n7509 );
nor ( n7511 , n7502 , n578 );
nand ( n7512 , n7507 , n7511 );
nand ( n7513 , n7510 , n7512 );
nor ( n7514 , n7500 , n7513 );
not ( n7515 , n7514 );
not ( n7516 , n5358 );
buf ( n7517 , n4779 );
buf ( n7518 , n4758 );
nand ( n7519 , n7516 , n7517 , n4740 , n7518 );
not ( n7520 , n7519 );
not ( n7521 , n7520 );
or ( n7522 , n7515 , n7521 );
not ( n7523 , n4791 );
not ( n7524 , n5357 );
not ( n7525 , n580 );
and ( n7526 , n7524 , n7525 );
not ( n7527 , n5395 );
nor ( n7528 , n7526 , n7527 );
not ( n7529 , n7528 );
or ( n7530 , n7523 , n7529 );
not ( n7531 , n5364 );
not ( n7532 , n5357 );
not ( n7533 , n580 );
and ( n7534 , n7532 , n7533 );
nor ( n7535 , n7534 , n4794 );
nor ( n7536 , n7531 , n7535 );
nand ( n7537 , n7530 , n7536 );
and ( n7538 , n7514 , n7537 );
not ( n7539 , n7513 );
not ( n7540 , n7539 );
not ( n7541 , n7498 );
nand ( n7542 , n7541 , n579 );
not ( n7543 , n7542 );
not ( n7544 , n7543 );
or ( n7545 , n7540 , n7544 );
nand ( n7546 , n7507 , n7502 );
not ( n7547 , n7546 );
not ( n7548 , n7502 );
nand ( n7549 , n7508 , n7548 );
not ( n7550 , n7549 );
or ( n7551 , n7547 , n7550 );
nand ( n7552 , n7551 , n578 );
nand ( n7553 , n7545 , n7552 );
nor ( n7554 , n7538 , n7553 );
nand ( n7555 , n7522 , n7554 );
xor ( n7556 , n7477 , n7555 );
buf ( n7557 , n7556 );
buf ( n7558 , n7557 );
buf ( n7559 , n7558 );
buf ( n7560 , n7559 );
not ( n7561 , n7560 );
buf ( n7562 , n7561 );
buf ( n7563 , n7562 );
not ( n7564 , n7563 );
or ( n7565 , n5659 , n7564 );
buf ( n7566 , n7559 );
buf ( n7567 , n2912 );
nand ( n7568 , n7566 , n7567 );
buf ( n7569 , n7568 );
buf ( n7570 , n7569 );
nand ( n7571 , n7565 , n7570 );
buf ( n7572 , n7571 );
buf ( n7573 , n7572 );
not ( n7574 , n7573 );
or ( n7575 , n5657 , n7574 );
buf ( n7576 , n602 );
not ( n7577 , n7576 );
not ( n7578 , n579 );
not ( n7579 , n7499 );
nand ( n7580 , n7578 , n7579 );
nand ( n7581 , n7537 , n7580 );
not ( n7582 , n7500 );
nand ( n7583 , n7582 , n7528 , n7517 , n7518 );
nand ( n7584 , n7499 , n579 );
nand ( n7585 , n7581 , n7583 , n7584 );
not ( n7586 , n7585 );
not ( n7587 , n7586 );
nand ( n7588 , n7552 , n7539 );
not ( n7589 , n7588 );
not ( n7590 , n7589 );
and ( n7591 , n7587 , n7590 );
and ( n7592 , n7586 , n7589 );
nor ( n7593 , n7591 , n7592 );
buf ( n7594 , n7593 );
not ( n7595 , n7594 );
or ( n7596 , n7577 , n7595 );
buf ( n7597 , n7593 );
not ( n7598 , n7597 );
buf ( n7599 , n7598 );
buf ( n7600 , n7599 );
buf ( n7601 , n2912 );
nand ( n7602 , n7600 , n7601 );
buf ( n7603 , n7602 );
buf ( n7604 , n7603 );
nand ( n7605 , n7596 , n7604 );
buf ( n7606 , n7605 );
buf ( n7607 , n7606 );
buf ( n7608 , n5652 );
buf ( n7609 , n603 );
buf ( n7610 , n602 );
and ( n7611 , n7609 , n7610 );
not ( n7612 , n7609 );
buf ( n7613 , n2912 );
and ( n7614 , n7612 , n7613 );
nor ( n7615 , n7611 , n7614 );
buf ( n7616 , n7615 );
buf ( n7617 , n7616 );
and ( n7618 , n7608 , n7617 );
buf ( n7619 , n7618 );
buf ( n7620 , n7619 );
nand ( n7621 , n7607 , n7620 );
buf ( n7622 , n7621 );
buf ( n7623 , n7622 );
nand ( n7624 , n7575 , n7623 );
buf ( n7625 , n7624 );
buf ( n7626 , n7625 );
xor ( n7627 , n5646 , n7626 );
xor ( n7628 , n5482 , n5544 );
and ( n7629 , n7628 , n5638 );
and ( n7630 , n5482 , n5544 );
or ( n7631 , n7629 , n7630 );
buf ( n7632 , n7631 );
buf ( n7633 , n7632 );
not ( n7634 , n5430 );
not ( n7635 , n5389 );
or ( n7636 , n7634 , n7635 );
not ( n7637 , n7537 );
nand ( n7638 , n7637 , n7519 );
not ( n7639 , n7578 );
not ( n7640 , n7579 );
or ( n7641 , n7639 , n7640 );
nand ( n7642 , n7641 , n7584 );
not ( n7643 , n7642 );
and ( n7644 , n7638 , n7643 );
not ( n7645 , n7638 );
and ( n7646 , n7645 , n7642 );
nor ( n7647 , n7644 , n7646 );
buf ( n7648 , n7647 );
or ( n7649 , n7648 , n5381 );
not ( n7650 , n600 );
nand ( n7651 , n7647 , n7650 );
nand ( n7652 , n7649 , n7651 );
nand ( n7653 , n7652 , n2915 );
nand ( n7654 , n7636 , n7653 );
buf ( n7655 , n7654 );
xor ( n7656 , n7633 , n7655 );
xor ( n7657 , n5508 , n5534 );
and ( n7658 , n7657 , n5541 );
and ( n7659 , n5508 , n5534 );
or ( n7660 , n7658 , n7659 );
buf ( n7661 , n7660 );
buf ( n7662 , n7661 );
buf ( n7663 , n5550 );
not ( n7664 , n7663 );
buf ( n7665 , n598 );
not ( n7666 , n7665 );
buf ( n7667 , n5407 );
not ( n7668 , n7667 );
or ( n7669 , n7666 , n7668 );
buf ( n7670 , n5411 );
buf ( n7671 , n818 );
nand ( n7672 , n7670 , n7671 );
buf ( n7673 , n7672 );
buf ( n7674 , n7673 );
nand ( n7675 , n7669 , n7674 );
buf ( n7676 , n7675 );
buf ( n7677 , n7676 );
not ( n7678 , n7677 );
or ( n7679 , n7664 , n7678 );
buf ( n7680 , n5631 );
buf ( n7681 , n5583 );
nand ( n7682 , n7680 , n7681 );
buf ( n7683 , n7682 );
buf ( n7684 , n7683 );
nand ( n7685 , n7679 , n7684 );
buf ( n7686 , n7685 );
buf ( n7687 , n7686 );
xor ( n7688 , n7662 , n7687 );
buf ( n7689 , n2541 );
not ( n7690 , n7689 );
and ( n7691 , n2361 , n2481 );
not ( n7692 , n2361 );
and ( n7693 , n7692 , n594 );
or ( n7694 , n7691 , n7693 );
buf ( n7695 , n7694 );
not ( n7696 , n7695 );
or ( n7697 , n7690 , n7696 );
buf ( n7698 , n5497 );
buf ( n7699 , n2592 );
nand ( n7700 , n7698 , n7699 );
buf ( n7701 , n7700 );
buf ( n7702 , n7701 );
nand ( n7703 , n7697 , n7702 );
buf ( n7704 , n7703 );
buf ( n7705 , n7704 );
buf ( n7706 , n2510 );
buf ( n7707 , n592 );
and ( n7708 , n7706 , n7707 );
buf ( n7709 , n7708 );
buf ( n7710 , n7709 );
not ( n7711 , n2452 );
buf ( n7712 , n592 );
not ( n7713 , n7712 );
buf ( n7714 , n2735 );
not ( n7715 , n7714 );
or ( n7716 , n7713 , n7715 );
buf ( n7717 , n2735 );
not ( n7718 , n7717 );
buf ( n7719 , n7718 );
buf ( n7720 , n7719 );
buf ( n7721 , n2416 );
nand ( n7722 , n7720 , n7721 );
buf ( n7723 , n7722 );
buf ( n7724 , n7723 );
nand ( n7725 , n7716 , n7724 );
buf ( n7726 , n7725 );
not ( n7727 , n7726 );
or ( n7728 , n7711 , n7727 );
not ( n7729 , n5523 );
nand ( n7730 , n7729 , n2460 );
nand ( n7731 , n7728 , n7730 );
buf ( n7732 , n7731 );
xor ( n7733 , n7710 , n7732 );
xor ( n7734 , n5513 , n5518 );
and ( n7735 , n7734 , n5531 );
and ( n7736 , n5513 , n5518 );
or ( n7737 , n7735 , n7736 );
buf ( n7738 , n7737 );
buf ( n7739 , n7738 );
xor ( n7740 , n7733 , n7739 );
buf ( n7741 , n7740 );
buf ( n7742 , n7741 );
xor ( n7743 , n7705 , n7742 );
buf ( n7744 , n825 );
not ( n7745 , n7744 );
buf ( n7746 , n596 );
not ( n7747 , n7746 );
buf ( n7748 , n5601 );
not ( n7749 , n7748 );
or ( n7750 , n7747 , n7749 );
not ( n7751 , n5598 );
buf ( n7752 , n7751 );
not ( n7753 , n7752 );
buf ( n7754 , n7753 );
buf ( n7755 , n7754 );
not ( n7756 , n7755 );
buf ( n7757 , n7756 );
buf ( n7758 , n7757 );
buf ( n7759 , n2371 );
nand ( n7760 , n7758 , n7759 );
buf ( n7761 , n7760 );
buf ( n7762 , n7761 );
nand ( n7763 , n7750 , n7762 );
buf ( n7764 , n7763 );
buf ( n7765 , n7764 );
not ( n7766 , n7765 );
or ( n7767 , n7745 , n7766 );
buf ( n7768 , n5471 );
buf ( n7769 , n2404 );
nand ( n7770 , n7768 , n7769 );
buf ( n7771 , n7770 );
buf ( n7772 , n7771 );
nand ( n7773 , n7767 , n7772 );
buf ( n7774 , n7773 );
buf ( n7775 , n7774 );
xor ( n7776 , n7743 , n7775 );
buf ( n7777 , n7776 );
buf ( n7778 , n7777 );
xor ( n7779 , n7688 , n7778 );
buf ( n7780 , n7779 );
buf ( n7781 , n7780 );
xor ( n7782 , n7656 , n7781 );
buf ( n7783 , n7782 );
buf ( n7784 , n7783 );
xor ( n7785 , n7627 , n7784 );
buf ( n7786 , n7785 );
buf ( n7787 , n7786 );
xor ( n7788 , n605 , n606 );
buf ( n7789 , n7788 );
buf ( n7790 , n7789 );
buf ( n7791 , n7790 );
not ( n7792 , n7791 );
nand ( n7793 , n7373 , n7467 );
not ( n7794 , n577 );
nand ( n7795 , n7793 , n7471 , n7794 );
not ( n7796 , n7795 );
not ( n7797 , n7553 );
or ( n7798 , n7796 , n7797 );
not ( n7799 , n7794 );
nand ( n7800 , n7799 , n7472 );
nand ( n7801 , n7798 , n7800 );
not ( n7802 , n7801 );
or ( n7803 , n7520 , n7537 );
and ( n7804 , n7795 , n7514 );
nand ( n7805 , n7803 , n7804 );
nand ( n7806 , n7802 , n7805 );
buf ( n7807 , n576 );
not ( n7808 , n7807 );
buf ( n7809 , n7808 );
not ( n7810 , n7809 );
buf ( n7811 , n6882 );
not ( n7812 , n7811 );
buf ( n7813 , n6437 );
not ( n7814 , n7813 );
or ( n7815 , n7812 , n7814 );
buf ( n7816 , n6890 );
nand ( n7817 , n7815 , n7816 );
buf ( n7818 , n7817 );
not ( n7819 , n7818 );
buf ( n7820 , n6441 );
buf ( n7821 , n6452 );
buf ( n7822 , n6882 );
buf ( n7823 , n6454 );
nand ( n7824 , n7820 , n7821 , n7822 , n7823 );
buf ( n7825 , n7824 );
nand ( n7826 , n6471 , n6452 , n6882 );
nand ( n7827 , n7819 , n7825 , n7826 );
not ( n7828 , n6569 );
not ( n7829 , n6557 );
nand ( n7830 , n7829 , n6556 );
not ( n7831 , n7830 );
or ( n7832 , n7828 , n7831 );
not ( n7833 , n6556 );
nand ( n7834 , n7833 , n6557 );
nand ( n7835 , n7832 , n7834 );
not ( n7836 , n6539 );
not ( n7837 , n6552 );
or ( n7838 , n7836 , n7837 );
or ( n7839 , n6552 , n6539 );
nand ( n7840 , n7839 , n6527 );
nand ( n7841 , n7838 , n7840 );
buf ( n7842 , n7841 );
not ( n7843 , n7842 );
buf ( n7844 , n7843 );
not ( n7845 , n7844 );
buf ( n7846 , n6548 );
not ( n7847 , n7846 );
buf ( n7848 , n4044 );
not ( n7849 , n7848 );
or ( n7850 , n7847 , n7849 );
buf ( n7851 , n3743 );
buf ( n7852 , n552 );
buf ( n7853 , n566 );
xor ( n7854 , n7852 , n7853 );
buf ( n7855 , n7854 );
buf ( n7856 , n7855 );
nand ( n7857 , n7851 , n7856 );
buf ( n7858 , n7857 );
buf ( n7859 , n7858 );
nand ( n7860 , n7850 , n7859 );
buf ( n7861 , n7860 );
buf ( n7862 , n7861 );
not ( n7863 , n7862 );
buf ( n7864 , n7863 );
buf ( n7865 , n7864 );
not ( n7866 , n7865 );
buf ( n7867 , n6535 );
not ( n7868 , n7867 );
buf ( n7869 , n842 );
buf ( n7870 , n844 );
and ( n7871 , n7869 , n7870 );
buf ( n7872 , n7871 );
buf ( n7873 , n7872 );
not ( n7874 , n7873 );
or ( n7875 , n7868 , n7874 );
buf ( n7876 , n1979 );
buf ( n7877 , n548 );
buf ( n7878 , n570 );
xor ( n7879 , n7877 , n7878 );
buf ( n7880 , n7879 );
buf ( n7881 , n7880 );
nand ( n7882 , n7876 , n7881 );
buf ( n7883 , n7882 );
buf ( n7884 , n7883 );
nand ( n7885 , n7875 , n7884 );
buf ( n7886 , n7885 );
buf ( n7887 , n7886 );
not ( n7888 , n7887 );
and ( n7889 , n7866 , n7888 );
buf ( n7890 , n7886 );
buf ( n7891 , n7864 );
and ( n7892 , n7890 , n7891 );
nor ( n7893 , n7889 , n7892 );
buf ( n7894 , n7893 );
buf ( n7895 , n6504 );
not ( n7896 , n7895 );
buf ( n7897 , n4836 );
not ( n7898 , n7897 );
or ( n7899 , n7896 , n7898 );
buf ( n7900 , n4840 );
xor ( n7901 , n564 , n554 );
buf ( n7902 , n7901 );
nand ( n7903 , n7900 , n7902 );
buf ( n7904 , n7903 );
buf ( n7905 , n7904 );
nand ( n7906 , n7899 , n7905 );
buf ( n7907 , n7906 );
and ( n7908 , n7894 , n7907 );
not ( n7909 , n7894 );
buf ( n7910 , n7907 );
not ( n7911 , n7910 );
buf ( n7912 , n7911 );
and ( n7913 , n7909 , n7912 );
nor ( n7914 , n7908 , n7913 );
not ( n7915 , n7914 );
not ( n7916 , n7915 );
or ( n7917 , n7845 , n7916 );
nand ( n7918 , n7841 , n7914 );
nand ( n7919 , n7917 , n7918 );
buf ( n7920 , n6610 );
not ( n7921 , n7920 );
buf ( n7922 , n4435 );
not ( n7923 , n7922 );
or ( n7924 , n7921 , n7923 );
buf ( n7925 , n888 );
xor ( n7926 , n572 , n546 );
buf ( n7927 , n7926 );
nand ( n7928 , n7925 , n7927 );
buf ( n7929 , n7928 );
buf ( n7930 , n7929 );
nand ( n7931 , n7924 , n7930 );
buf ( n7932 , n7931 );
buf ( n7933 , n6521 );
not ( n7934 , n7933 );
buf ( n7935 , n4021 );
not ( n7936 , n7935 );
or ( n7937 , n7934 , n7936 );
buf ( n7938 , n3436 );
buf ( n7939 , n550 );
buf ( n7940 , n568 );
xor ( n7941 , n7939 , n7940 );
buf ( n7942 , n7941 );
buf ( n7943 , n7942 );
nand ( n7944 , n7938 , n7943 );
buf ( n7945 , n7944 );
buf ( n7946 , n7945 );
nand ( n7947 , n7937 , n7946 );
buf ( n7948 , n7947 );
xor ( n7949 , n7932 , n7948 );
buf ( n7950 , n7949 );
not ( n7951 , n6595 );
buf ( n7952 , n558 );
buf ( n7953 , n560 );
xor ( n7954 , n7952 , n7953 );
buf ( n7955 , n7954 );
not ( n7956 , n7955 );
or ( n7957 , n7951 , n7956 );
not ( n7958 , n560 );
nor ( n7959 , n561 , n562 );
not ( n7960 , n7959 );
or ( n7961 , n7958 , n7960 );
not ( n7962 , n560 );
nand ( n7963 , n7962 , n561 , n562 );
nand ( n7964 , n7961 , n7963 );
xor ( n7965 , n560 , n559 );
nand ( n7966 , n7964 , n7965 );
nand ( n7967 , n7957 , n7966 );
buf ( n7968 , n7967 );
xor ( n7969 , n7950 , n7968 );
buf ( n7970 , n7969 );
xnor ( n7971 , n7919 , n7970 );
xor ( n7972 , n7835 , n7971 );
xor ( n7973 , n6494 , n6511 );
and ( n7974 , n7973 , n6517 );
and ( n7975 , n6494 , n6511 );
or ( n7976 , n7974 , n7975 );
buf ( n7977 , n7976 );
buf ( n7978 , n7977 );
buf ( n7979 , n6487 );
not ( n7980 , n7979 );
buf ( n7981 , n5818 );
buf ( n7982 , n5813 );
nor ( n7983 , n7981 , n7982 );
buf ( n7984 , n7983 );
buf ( n7985 , n7984 );
not ( n7986 , n7985 );
or ( n7987 , n7980 , n7986 );
buf ( n7988 , n5801 );
buf ( n7989 , n556 );
buf ( n7990 , n562 );
xor ( n7991 , n7989 , n7990 );
buf ( n7992 , n7991 );
buf ( n7993 , n7992 );
nand ( n7994 , n7988 , n7993 );
buf ( n7995 , n7994 );
buf ( n7996 , n7995 );
nand ( n7997 , n7987 , n7996 );
buf ( n7998 , n7997 );
buf ( n7999 , n7998 );
buf ( n8000 , n559 );
buf ( n8001 , n561 );
or ( n8002 , n8000 , n8001 );
buf ( n8003 , n562 );
nand ( n8004 , n8002 , n8003 );
buf ( n8005 , n8004 );
buf ( n8006 , n8005 );
buf ( n8007 , n559 );
buf ( n8008 , n561 );
nand ( n8009 , n8007 , n8008 );
buf ( n8010 , n8009 );
buf ( n8011 , n8010 );
buf ( n8012 , n560 );
nand ( n8013 , n8006 , n8011 , n8012 );
buf ( n8014 , n8013 );
buf ( n8015 , n8014 );
not ( n8016 , n8015 );
buf ( n8017 , n6592 );
not ( n8018 , n8017 );
buf ( n8019 , n4953 );
not ( n8020 , n8019 );
or ( n8021 , n8018 , n8020 );
buf ( n8022 , n544 );
buf ( n8023 , n574 );
xor ( n8024 , n8022 , n8023 );
buf ( n8025 , n8024 );
buf ( n8026 , n8025 );
buf ( n8027 , n575 );
nand ( n8028 , n8026 , n8027 );
buf ( n8029 , n8028 );
buf ( n8030 , n8029 );
nand ( n8031 , n8021 , n8030 );
buf ( n8032 , n8031 );
buf ( n8033 , n8032 );
not ( n8034 , n8033 );
or ( n8035 , n8016 , n8034 );
buf ( n8036 , n8032 );
buf ( n8037 , n8014 );
or ( n8038 , n8036 , n8037 );
nand ( n8039 , n8035 , n8038 );
buf ( n8040 , n8039 );
buf ( n8041 , n8040 );
xor ( n8042 , n7999 , n8041 );
buf ( n8043 , n6599 );
not ( n8044 , n8043 );
buf ( n8045 , n6594 );
not ( n8046 , n8045 );
buf ( n8047 , n8046 );
buf ( n8048 , n8047 );
not ( n8049 , n8048 );
or ( n8050 , n8044 , n8049 );
buf ( n8051 , n6616 );
nand ( n8052 , n8050 , n8051 );
buf ( n8053 , n8052 );
buf ( n8054 , n8053 );
buf ( n8055 , n6599 );
not ( n8056 , n8055 );
buf ( n8057 , n6594 );
nand ( n8058 , n8056 , n8057 );
buf ( n8059 , n8058 );
buf ( n8060 , n8059 );
nand ( n8061 , n8054 , n8060 );
buf ( n8062 , n8061 );
buf ( n8063 , n8062 );
xor ( n8064 , n8042 , n8063 );
buf ( n8065 , n8064 );
buf ( n8066 , n8065 );
xor ( n8067 , n7978 , n8066 );
buf ( n8068 , n6617 );
not ( n8069 , n8068 );
buf ( n8070 , n6583 );
not ( n8071 , n8070 );
or ( n8072 , n8069 , n8071 );
buf ( n8073 , n6633 );
nand ( n8074 , n8072 , n8073 );
buf ( n8075 , n8074 );
buf ( n8076 , n8075 );
buf ( n8077 , n6580 );
buf ( n8078 , n6623 );
nand ( n8079 , n8077 , n8078 );
buf ( n8080 , n8079 );
buf ( n8081 , n8080 );
nand ( n8082 , n8076 , n8081 );
buf ( n8083 , n8082 );
buf ( n8084 , n8083 );
xor ( n8085 , n8067 , n8084 );
buf ( n8086 , n8085 );
xnor ( n8087 , n7972 , n8086 );
buf ( n8088 , n8087 );
xor ( n8089 , n6674 , n6679 );
and ( n8090 , n8089 , n6866 );
and ( n8091 , n6674 , n6679 );
or ( n8092 , n8090 , n8091 );
buf ( n8093 , n8092 );
xor ( n8094 , n8088 , n8093 );
buf ( n8095 , n6658 );
not ( n8096 , n8095 );
buf ( n8097 , n6574 );
not ( n8098 , n8097 );
or ( n8099 , n8096 , n8098 );
buf ( n8100 , n6658 );
buf ( n8101 , n6574 );
or ( n8102 , n8100 , n8101 );
buf ( n8103 , n6643 );
nand ( n8104 , n8102 , n8103 );
buf ( n8105 , n8104 );
buf ( n8106 , n8105 );
nand ( n8107 , n8099 , n8106 );
buf ( n8108 , n8107 );
buf ( n8109 , n8108 );
xor ( n8110 , n6695 , n6747 );
and ( n8111 , n8110 , n6864 );
and ( n8112 , n6695 , n6747 );
or ( n8113 , n8111 , n8112 );
buf ( n8114 , n8113 );
buf ( n8115 , n8114 );
xor ( n8116 , n8109 , n8115 );
not ( n8117 , n4538 );
and ( n8118 , n580 , n4257 );
not ( n8119 , n580 );
and ( n8120 , n8119 , n554 );
or ( n8121 , n8118 , n8120 );
not ( n8122 , n8121 );
or ( n8123 , n8117 , n8122 );
nand ( n8124 , n5058 , n6845 , n4541 );
nand ( n8125 , n8123 , n8124 );
buf ( n8126 , n6800 );
not ( n8127 , n8126 );
buf ( n8128 , n3616 );
not ( n8129 , n8128 );
or ( n8130 , n8127 , n8129 );
and ( n8131 , n548 , n586 );
not ( n8132 , n548 );
and ( n8133 , n8132 , n1766 );
nor ( n8134 , n8131 , n8133 );
nand ( n8135 , n1169 , n8134 );
buf ( n8136 , n8135 );
nand ( n8137 , n8130 , n8136 );
buf ( n8138 , n8137 );
xor ( n8139 , n8125 , n8138 );
buf ( n8140 , n6782 );
not ( n8141 , n8140 );
buf ( n8142 , n4205 );
not ( n8143 , n8142 );
or ( n8144 , n8141 , n8143 );
buf ( n8145 , n4211 );
buf ( n8146 , n552 );
buf ( n8147 , n582 );
xor ( n8148 , n8146 , n8147 );
buf ( n8149 , n8148 );
buf ( n8150 , n8149 );
nand ( n8151 , n8145 , n8150 );
buf ( n8152 , n8151 );
buf ( n8153 , n8152 );
nand ( n8154 , n8144 , n8153 );
buf ( n8155 , n8154 );
xor ( n8156 , n8139 , n8155 );
not ( n8157 , n8156 );
not ( n8158 , n6804 );
not ( n8159 , n6788 );
or ( n8160 , n8158 , n8159 );
not ( n8161 , n6805 );
not ( n8162 , n6791 );
or ( n8163 , n8161 , n8162 );
nand ( n8164 , n8163 , n6772 );
nand ( n8165 , n8160 , n8164 );
not ( n8166 , n8165 );
not ( n8167 , n8166 );
or ( n8168 , n8157 , n8167 );
or ( n8169 , n8166 , n8156 );
nand ( n8170 , n8168 , n8169 );
buf ( n8171 , n8170 );
not ( n8172 , n6724 );
not ( n8173 , n4286 );
or ( n8174 , n8172 , n8173 );
not ( n8175 , n4555 );
not ( n8176 , n4554 );
or ( n8177 , n8175 , n8176 );
buf ( n8178 , n546 );
buf ( n8179 , n588 );
xor ( n8180 , n8178 , n8179 );
buf ( n8181 , n8180 );
nand ( n8182 , n8177 , n8181 );
nand ( n8183 , n8174 , n8182 );
buf ( n8184 , n559 );
buf ( n8185 , n576 );
xor ( n8186 , n8184 , n8185 );
buf ( n8187 , n8186 );
not ( n8188 , n8187 );
buf ( n8189 , n6699 );
buf ( n8190 , n576 );
buf ( n8191 , n577 );
xnor ( n8192 , n8190 , n8191 );
buf ( n8193 , n8192 );
buf ( n8194 , n8193 );
nor ( n8195 , n8189 , n8194 );
buf ( n8196 , n8195 );
not ( n8197 , n8196 );
or ( n8198 , n8188 , n8197 );
buf ( n8199 , n6699 );
buf ( n8200 , n558 );
buf ( n8201 , n576 );
xor ( n8202 , n8200 , n8201 );
buf ( n8203 , n8202 );
buf ( n8204 , n8203 );
nand ( n8205 , n8199 , n8204 );
buf ( n8206 , n8205 );
nand ( n8207 , n8198 , n8206 );
xor ( n8208 , n8183 , n8207 );
not ( n8209 , n6766 );
not ( n8210 , n3664 );
or ( n8211 , n8209 , n8210 );
buf ( n8212 , n2135 );
buf ( n8213 , n550 );
buf ( n8214 , n584 );
xor ( n8215 , n8213 , n8214 );
buf ( n8216 , n8215 );
buf ( n8217 , n8216 );
nand ( n8218 , n8212 , n8217 );
buf ( n8219 , n8218 );
nand ( n8220 , n8211 , n8219 );
xnor ( n8221 , n8208 , n8220 );
buf ( n8222 , n8221 );
buf ( n8223 , n8222 );
buf ( n8224 , n8223 );
buf ( n8225 , n8224 );
xnor ( n8226 , n8171 , n8225 );
buf ( n8227 , n8226 );
buf ( n8228 , n8227 );
not ( n8229 , n6257 );
not ( n8230 , n6750 );
or ( n8231 , n8229 , n8230 );
nand ( n8232 , n8231 , n6753 );
not ( n8233 , n8232 );
not ( n8234 , n6809 );
nand ( n8235 , n8234 , n6855 );
not ( n8236 , n8235 );
or ( n8237 , n8233 , n8236 );
nand ( n8238 , n6809 , n6854 );
nand ( n8239 , n8237 , n8238 );
buf ( n8240 , n8239 );
xor ( n8241 , n8228 , n8240 );
not ( n8242 , n6825 );
nand ( n8243 , n8242 , n6832 );
not ( n8244 , n8243 );
not ( n8245 , n6849 );
or ( n8246 , n8244 , n8245 );
not ( n8247 , n6832 );
nand ( n8248 , n8247 , n6825 );
nand ( n8249 , n8246 , n8248 );
buf ( n8250 , n8249 );
buf ( n8251 , n559 );
buf ( n8252 , n577 );
or ( n8253 , n8251 , n8252 );
buf ( n8254 , n578 );
nand ( n8255 , n8253 , n8254 );
buf ( n8256 , n8255 );
buf ( n8257 , n8256 );
buf ( n8258 , n559 );
buf ( n8259 , n577 );
nand ( n8260 , n8258 , n8259 );
buf ( n8261 , n8260 );
buf ( n8262 , n8261 );
buf ( n8263 , n576 );
and ( n8264 , n8257 , n8262 , n8263 );
buf ( n8265 , n8264 );
buf ( n8266 , n8265 );
buf ( n8267 , n6709 );
not ( n8268 , n8267 );
buf ( n8269 , n984 );
not ( n8270 , n8269 );
or ( n8271 , n8268 , n8270 );
buf ( n8272 , n544 );
buf ( n8273 , n590 );
xor ( n8274 , n8272 , n8273 );
buf ( n8275 , n8274 );
buf ( n8276 , n8275 );
buf ( n8277 , n591 );
nand ( n8278 , n8276 , n8277 );
buf ( n8279 , n8278 );
buf ( n8280 , n8279 );
nand ( n8281 , n8271 , n8280 );
buf ( n8282 , n8281 );
buf ( n8283 , n8282 );
xor ( n8284 , n8266 , n8283 );
buf ( n8285 , n8284 );
buf ( n8286 , n8285 );
buf ( n8287 , n6819 );
not ( n8288 , n8287 );
buf ( n8289 , n6350 );
not ( n8290 , n8289 );
or ( n8291 , n8288 , n8290 );
buf ( n8292 , n5997 );
buf ( n8293 , n8292 );
buf ( n8294 , n8293 );
buf ( n8295 , n8294 );
xor ( n8296 , n578 , n556 );
buf ( n8297 , n8296 );
nand ( n8298 , n8295 , n8297 );
buf ( n8299 , n8298 );
buf ( n8300 , n8299 );
nand ( n8301 , n8291 , n8300 );
buf ( n8302 , n8301 );
buf ( n8303 , n8302 );
xor ( n8304 , n8286 , n8303 );
xor ( n8305 , n6704 , n6714 );
and ( n8306 , n8305 , n6729 );
and ( n8307 , n6704 , n6714 );
or ( n8308 , n8306 , n8307 );
buf ( n8309 , n8308 );
buf ( n8310 , n8309 );
xor ( n8311 , n8304 , n8310 );
buf ( n8312 , n8311 );
buf ( n8313 , n8312 );
xor ( n8314 , n8250 , n8313 );
xor ( n8315 , n6732 , n6737 );
and ( n8316 , n8315 , n6744 );
and ( n8317 , n6732 , n6737 );
or ( n8318 , n8316 , n8317 );
buf ( n8319 , n8318 );
buf ( n8320 , n8319 );
xor ( n8321 , n8314 , n8320 );
buf ( n8322 , n8321 );
buf ( n8323 , n8322 );
xor ( n8324 , n8241 , n8323 );
buf ( n8325 , n8324 );
buf ( n8326 , n8325 );
xor ( n8327 , n8116 , n8326 );
buf ( n8328 , n8327 );
buf ( n8329 , n8328 );
xor ( n8330 , n8094 , n8329 );
buf ( n8331 , n8330 );
buf ( n8332 , n8331 );
xor ( n8333 , n6660 , n6666 );
and ( n8334 , n8333 , n6868 );
and ( n8335 , n6660 , n6666 );
or ( n8336 , n8334 , n8335 );
buf ( n8337 , n8336 );
buf ( n8338 , n8337 );
and ( n8339 , n8332 , n8338 );
buf ( n8340 , n8339 );
not ( n8341 , n8340 );
buf ( n8342 , n8331 );
not ( n8343 , n8342 );
buf ( n8344 , n8343 );
buf ( n8345 , n8344 );
buf ( n8346 , n8337 );
not ( n8347 , n8346 );
buf ( n8348 , n8347 );
buf ( n8349 , n8348 );
nand ( n8350 , n8345 , n8349 );
buf ( n8351 , n8350 );
nand ( n8352 , n8341 , n8351 );
not ( n8353 , n8352 );
and ( n8354 , n7827 , n8353 );
not ( n8355 , n7827 );
and ( n8356 , n8355 , n8352 );
nor ( n8357 , n8354 , n8356 );
not ( n8358 , n8357 );
xor ( n8359 , n6922 , n6992 );
and ( n8360 , n8359 , n7031 );
and ( n8361 , n6922 , n6992 );
or ( n8362 , n8360 , n8361 );
xor ( n8363 , n7169 , n7281 );
and ( n8364 , n8363 , n7298 );
and ( n8365 , n7169 , n7281 );
or ( n8366 , n8364 , n8365 );
xor ( n8367 , n8362 , n8366 );
not ( n8368 , n1596 );
not ( n8369 , n556 );
not ( n8370 , n7223 );
or ( n8371 , n8369 , n8370 );
not ( n8372 , n556 );
nand ( n8373 , n8372 , n7222 );
nand ( n8374 , n8371 , n8373 );
not ( n8375 , n8374 );
or ( n8376 , n8368 , n8375 );
and ( n8377 , n7124 , n3112 );
and ( n8378 , n7125 , n3109 );
nor ( n8379 , n8377 , n8378 );
nand ( n8380 , n8376 , n8379 );
xor ( n8381 , n7171 , n7188 );
and ( n8382 , n8381 , n7194 );
and ( n8383 , n7171 , n7188 );
or ( n8384 , n8382 , n8383 );
xor ( n8385 , n8380 , n8384 );
not ( n8386 , n3118 );
not ( n8387 , n554 );
not ( n8388 , n5247 );
or ( n8389 , n8387 , n8388 );
nand ( n8390 , n7147 , n1681 );
nand ( n8391 , n8389 , n8390 );
not ( n8392 , n8391 );
or ( n8393 , n8386 , n8392 );
nand ( n8394 , n6920 , n6906 );
nand ( n8395 , n8393 , n8394 );
xor ( n8396 , n8385 , n8395 );
not ( n8397 , n3068 );
and ( n8398 , n2981 , n3073 );
not ( n8399 , n2981 );
and ( n8400 , n8399 , n550 );
or ( n8401 , n8398 , n8400 );
not ( n8402 , n8401 );
or ( n8403 , n8397 , n8402 );
nand ( n8404 , n7009 , n5268 );
nand ( n8405 , n8403 , n8404 );
nand ( n8406 , n7020 , n3064 );
not ( n8407 , n3167 );
and ( n8408 , n2265 , n552 );
nand ( n8409 , n8407 , n8408 );
not ( n8410 , n552 );
nand ( n8411 , n8410 , n2265 , n3167 );
nand ( n8412 , n8406 , n8409 , n8411 );
xor ( n8413 , n8405 , n8412 );
not ( n8414 , n559 );
not ( n8415 , n558 );
nand ( n8416 , n7239 , n7231 );
nor ( n8417 , n7095 , n8416 );
not ( n8418 , n8417 );
not ( n8419 , n3033 );
or ( n8420 , n8418 , n8419 );
not ( n8421 , n8416 );
and ( n8422 , n7249 , n8421 );
nor ( n8423 , n577 , n561 );
not ( n8424 , n8423 );
or ( n8425 , n578 , n562 );
nand ( n8426 , n8424 , n8425 , n7116 );
or ( n8427 , n8423 , n7257 );
nand ( n8428 , n8426 , n8427 , n7232 );
nor ( n8429 , n8422 , n8428 );
nand ( n8430 , n8420 , n8429 );
nor ( n8431 , n560 , n576 );
not ( n8432 , n8431 );
nand ( n8433 , n560 , n576 );
nand ( n8434 , n8432 , n8433 );
and ( n8435 , n8430 , n8434 );
not ( n8436 , n8430 );
not ( n8437 , n8434 );
and ( n8438 , n8436 , n8437 );
nor ( n8439 , n8435 , n8438 );
not ( n8440 , n8439 );
not ( n8441 , n8440 );
not ( n8442 , n8441 );
or ( n8443 , n8415 , n8442 );
nand ( n8444 , n8440 , n1736 );
nand ( n8445 , n8443 , n8444 );
not ( n8446 , n8445 );
or ( n8447 , n8414 , n8446 );
nand ( n8448 , n7278 , n1739 );
nand ( n8449 , n8447 , n8448 );
xor ( n8450 , n8413 , n8449 );
xor ( n8451 , n8396 , n8450 );
xor ( n8452 , n7002 , n7011 );
and ( n8453 , n8452 , n7030 );
and ( n8454 , n7002 , n7011 );
or ( n8455 , n8453 , n8454 );
not ( n8456 , n6945 );
not ( n8457 , n546 );
not ( n8458 , n3049 );
or ( n8459 , n8457 , n8458 );
nand ( n8460 , n5261 , n6949 );
nand ( n8461 , n8459 , n8460 );
not ( n8462 , n8461 );
or ( n8463 , n8456 , n8462 );
xor ( n8464 , n546 , n547 );
not ( n8465 , n8464 );
nor ( n8466 , n8465 , n6945 );
nand ( n8467 , n7176 , n8466 );
nand ( n8468 , n8463 , n8467 );
or ( n8469 , n545 , n546 );
nand ( n8470 , n8469 , n1664 );
nand ( n8471 , n545 , n546 );
and ( n8472 , n8470 , n8471 , n544 );
not ( n8473 , n7170 );
not ( n8474 , n544 );
not ( n8475 , n1677 );
or ( n8476 , n8474 , n8475 );
not ( n8477 , n544 );
nand ( n8478 , n1680 , n8477 );
nand ( n8479 , n8476 , n8478 );
not ( n8480 , n8479 );
or ( n8481 , n8473 , n8480 );
not ( n8482 , n544 );
not ( n8483 , n1687 );
or ( n8484 , n8482 , n8483 );
nand ( n8485 , n1798 , n8477 );
nand ( n8486 , n8484 , n8485 );
xnor ( n8487 , n544 , n545 );
nor ( n8488 , n7170 , n8487 );
nand ( n8489 , n8486 , n8488 );
nand ( n8490 , n8481 , n8489 );
xor ( n8491 , n8472 , n8490 );
xor ( n8492 , n8468 , n8491 );
not ( n8493 , n6923 );
not ( n8494 , n548 );
not ( n8495 , n5304 );
or ( n8496 , n8494 , n8495 );
nand ( n8497 , n1772 , n5279 );
nand ( n8498 , n8496 , n8497 );
not ( n8499 , n8498 );
or ( n8500 , n8493 , n8499 );
nand ( n8501 , n6998 , n6939 );
nand ( n8502 , n8500 , n8501 );
xor ( n8503 , n8492 , n8502 );
xor ( n8504 , n8455 , n8503 );
xor ( n8505 , n7195 , n7205 );
and ( n8506 , n8505 , n7280 );
and ( n8507 , n7195 , n7205 );
or ( n8508 , n8506 , n8507 );
xor ( n8509 , n8504 , n8508 );
xor ( n8510 , n8451 , n8509 );
xor ( n8511 , n8367 , n8510 );
not ( n8512 , n8511 );
xor ( n8513 , n7032 , n7164 );
and ( n8514 , n8513 , n7299 );
and ( n8515 , n7032 , n7164 );
or ( n8516 , n8514 , n8515 );
not ( n8517 , n8516 );
nand ( n8518 , n8512 , n8517 );
buf ( n8519 , n8518 );
buf ( n8520 , n8511 );
nand ( n8521 , n8520 , n8516 );
nand ( n8522 , n8519 , n8521 );
not ( n8523 , n8522 );
or ( n8524 , n7362 , n7326 );
nand ( n8525 , n8524 , n7324 );
not ( n8526 , n8525 );
or ( n8527 , n8523 , n8526 );
or ( n8528 , n8522 , n8525 );
nand ( n8529 , n8527 , n8528 );
nor ( n8530 , n8358 , n8529 );
not ( n8531 , n8530 );
nand ( n8532 , n8358 , n8529 );
nand ( n8533 , n8531 , n8532 );
and ( n8534 , n7451 , n7369 );
nor ( n8535 , n8534 , n7372 );
nand ( n8536 , n7461 , n7369 , n7464 );
not ( n8537 , n7441 );
nor ( n8538 , n8537 , n7383 );
nand ( n8539 , n8538 , n7369 , n7464 );
nand ( n8540 , n8535 , n8536 , n8539 );
xor ( n8541 , n8533 , n8540 );
not ( n8542 , n8541 );
not ( n8543 , n8542 );
not ( n8544 , n8543 );
or ( n8545 , n7810 , n8544 );
nand ( n8546 , n8542 , n576 );
nand ( n8547 , n8545 , n8546 );
not ( n8548 , n8547 );
and ( n8549 , n7806 , n8548 );
not ( n8550 , n7806 );
and ( n8551 , n8550 , n8547 );
nor ( n8552 , n8549 , n8551 );
buf ( n8553 , n8552 );
not ( n8554 , n8553 );
and ( n8555 , n604 , n8554 );
not ( n8556 , n604 );
not ( n8557 , n8554 );
and ( n8558 , n8556 , n8557 );
or ( n8559 , n8555 , n8558 );
buf ( n8560 , n8559 );
not ( n8561 , n8560 );
or ( n8562 , n7792 , n8561 );
and ( n8563 , n604 , n7562 );
not ( n8564 , n604 );
and ( n8565 , n8564 , n7559 );
or ( n8566 , n8563 , n8565 );
buf ( n8567 , n8566 );
buf ( n8568 , n604 );
buf ( n8569 , n605 );
and ( n8570 , n8568 , n8569 );
buf ( n8571 , n7788 );
buf ( n8572 , n604 );
buf ( n8573 , n605 );
nor ( n8574 , n8572 , n8573 );
buf ( n8575 , n8574 );
buf ( n8576 , n8575 );
nor ( n8577 , n8570 , n8571 , n8576 );
buf ( n8578 , n8577 );
buf ( n8579 , n8578 );
buf ( n8580 , n8579 );
buf ( n8581 , n8580 );
buf ( n8582 , n8581 );
nand ( n8583 , n8567 , n8582 );
buf ( n8584 , n8583 );
buf ( n8585 , n8584 );
nand ( n8586 , n8562 , n8585 );
buf ( n8587 , n8586 );
buf ( n8588 , n8587 );
buf ( n8589 , n5550 );
not ( n8590 , n8589 );
buf ( n8591 , n598 );
not ( n8592 , n8591 );
buf ( n8593 , n5464 );
not ( n8594 , n8593 );
buf ( n8595 , n8594 );
buf ( n8596 , n8595 );
not ( n8597 , n8596 );
or ( n8598 , n8592 , n8597 );
buf ( n8599 , n5458 );
not ( n8600 , n8599 );
buf ( n8601 , n818 );
nand ( n8602 , n8600 , n8601 );
buf ( n8603 , n8602 );
buf ( n8604 , n8603 );
nand ( n8605 , n8598 , n8604 );
buf ( n8606 , n8605 );
buf ( n8607 , n8606 );
not ( n8608 , n8607 );
or ( n8609 , n8590 , n8608 );
buf ( n8610 , n598 );
not ( n8611 , n8610 );
buf ( n8612 , n2364 );
not ( n8613 , n8612 );
or ( n8614 , n8611 , n8613 );
buf ( n8615 , n2361 );
buf ( n8616 , n818 );
nand ( n8617 , n8615 , n8616 );
buf ( n8618 , n8617 );
buf ( n8619 , n8618 );
nand ( n8620 , n8614 , n8619 );
buf ( n8621 , n8620 );
buf ( n8622 , n8621 );
buf ( n8623 , n5631 );
nand ( n8624 , n8622 , n8623 );
buf ( n8625 , n8624 );
buf ( n8626 , n8625 );
nand ( n8627 , n8609 , n8626 );
buf ( n8628 , n8627 );
buf ( n8629 , n8628 );
xor ( n8630 , n2754 , n2758 );
xor ( n8631 , n8630 , n2897 );
buf ( n8632 , n8631 );
buf ( n8633 , n8632 );
xor ( n8634 , n8629 , n8633 );
buf ( n8635 , n2915 );
not ( n8636 , n8635 );
buf ( n8637 , n600 );
not ( n8638 , n8637 );
not ( n8639 , n5576 );
buf ( n8640 , n8639 );
not ( n8641 , n8640 );
or ( n8642 , n8638 , n8641 );
buf ( n8643 , n5576 );
buf ( n8644 , n5383 );
nand ( n8645 , n8643 , n8644 );
buf ( n8646 , n8645 );
buf ( n8647 , n8646 );
nand ( n8648 , n8642 , n8647 );
buf ( n8649 , n8648 );
buf ( n8650 , n8649 );
not ( n8651 , n8650 );
or ( n8652 , n8636 , n8651 );
buf ( n8653 , n600 );
not ( n8654 , n8653 );
buf ( n8655 , n5601 );
not ( n8656 , n8655 );
or ( n8657 , n8654 , n8656 );
buf ( n8658 , n7757 );
buf ( n8659 , n5382 );
nand ( n8660 , n8658 , n8659 );
buf ( n8661 , n8660 );
buf ( n8662 , n8661 );
nand ( n8663 , n8657 , n8662 );
buf ( n8664 , n8663 );
buf ( n8665 , n8664 );
buf ( n8666 , n5430 );
nand ( n8667 , n8665 , n8666 );
buf ( n8668 , n8667 );
buf ( n8669 , n8668 );
nand ( n8670 , n8652 , n8669 );
buf ( n8671 , n8670 );
buf ( n8672 , n8671 );
and ( n8673 , n8634 , n8672 );
and ( n8674 , n8629 , n8633 );
or ( n8675 , n8673 , n8674 );
buf ( n8676 , n8675 );
buf ( n8677 , n8676 );
buf ( n8678 , n5655 );
not ( n8679 , n8678 );
buf ( n8680 , n602 );
not ( n8681 , n8680 );
buf ( n8682 , n7648 );
not ( n8683 , n8682 );
buf ( n8684 , n8683 );
buf ( n8685 , n8684 );
not ( n8686 , n8685 );
or ( n8687 , n8681 , n8686 );
buf ( n8688 , n7648 );
buf ( n8689 , n2912 );
nand ( n8690 , n8688 , n8689 );
buf ( n8691 , n8690 );
buf ( n8692 , n8691 );
nand ( n8693 , n8687 , n8692 );
buf ( n8694 , n8693 );
buf ( n8695 , n8694 );
not ( n8696 , n8695 );
or ( n8697 , n8679 , n8696 );
buf ( n8698 , n602 );
not ( n8699 , n8698 );
buf ( n8700 , n5376 );
not ( n8701 , n8700 );
or ( n8702 , n8699 , n8701 );
buf ( n8703 , n5379 );
buf ( n8704 , n2912 );
nand ( n8705 , n8703 , n8704 );
buf ( n8706 , n8705 );
buf ( n8707 , n8706 );
nand ( n8708 , n8702 , n8707 );
buf ( n8709 , n8708 );
buf ( n8710 , n8709 );
buf ( n8711 , n7619 );
nand ( n8712 , n8710 , n8711 );
buf ( n8713 , n8712 );
buf ( n8714 , n8713 );
nand ( n8715 , n8697 , n8714 );
buf ( n8716 , n8715 );
buf ( n8717 , n8716 );
xor ( n8718 , n8677 , n8717 );
buf ( n8719 , n5550 );
not ( n8720 , n8719 );
buf ( n8721 , n5614 );
not ( n8722 , n8721 );
or ( n8723 , n8720 , n8722 );
buf ( n8724 , n8606 );
buf ( n8725 , n5631 );
nand ( n8726 , n8724 , n8725 );
buf ( n8727 , n8726 );
buf ( n8728 , n8727 );
nand ( n8729 , n8723 , n8728 );
buf ( n8730 , n8729 );
buf ( n8731 , n8730 );
buf ( n8732 , n2915 );
not ( n8733 , n8732 );
buf ( n8734 , n5418 );
not ( n8735 , n8734 );
or ( n8736 , n8733 , n8735 );
buf ( n8737 , n8649 );
buf ( n8738 , n5430 );
nand ( n8739 , n8737 , n8738 );
buf ( n8740 , n8739 );
buf ( n8741 , n8740 );
nand ( n8742 , n8736 , n8741 );
buf ( n8743 , n8742 );
buf ( n8744 , n8743 );
xor ( n8745 , n8731 , n8744 );
xor ( n8746 , n2411 , n2721 );
xor ( n8747 , n8746 , n2902 );
buf ( n8748 , n8747 );
buf ( n8749 , n8748 );
xor ( n8750 , n8745 , n8749 );
buf ( n8751 , n8750 );
buf ( n8752 , n8751 );
and ( n8753 , n8718 , n8752 );
and ( n8754 , n8677 , n8717 );
or ( n8755 , n8753 , n8754 );
buf ( n8756 , n8755 );
buf ( n8757 , n8756 );
xor ( n8758 , n8588 , n8757 );
xor ( n8759 , n8731 , n8744 );
and ( n8760 , n8759 , n8749 );
and ( n8761 , n8731 , n8744 );
or ( n8762 , n8760 , n8761 );
buf ( n8763 , n8762 );
buf ( n8764 , n8763 );
xor ( n8765 , n2907 , n5437 );
xor ( n8766 , n8765 , n5641 );
buf ( n8767 , n8766 );
buf ( n8768 , n8767 );
xor ( n8769 , n8764 , n8768 );
buf ( n8770 , n5655 );
not ( n8771 , n8770 );
buf ( n8772 , n7606 );
not ( n8773 , n8772 );
or ( n8774 , n8771 , n8773 );
buf ( n8775 , n8694 );
buf ( n8776 , n7619 );
nand ( n8777 , n8775 , n8776 );
buf ( n8778 , n8777 );
buf ( n8779 , n8778 );
nand ( n8780 , n8774 , n8779 );
buf ( n8781 , n8780 );
buf ( n8782 , n8781 );
xor ( n8783 , n8769 , n8782 );
buf ( n8784 , n8783 );
buf ( n8785 , n8784 );
and ( n8786 , n8758 , n8785 );
and ( n8787 , n8588 , n8757 );
or ( n8788 , n8786 , n8787 );
buf ( n8789 , n8788 );
buf ( n8790 , n8789 );
xor ( n8791 , n7787 , n8790 );
xor ( n8792 , n8764 , n8768 );
and ( n8793 , n8792 , n8782 );
and ( n8794 , n8764 , n8768 );
or ( n8795 , n8793 , n8794 );
buf ( n8796 , n8795 );
buf ( n8797 , n8796 );
buf ( n8798 , n7790 );
not ( n8799 , n8798 );
xor ( n8800 , n7999 , n8041 );
and ( n8801 , n8800 , n8063 );
and ( n8802 , n7999 , n8041 );
or ( n8803 , n8801 , n8802 );
buf ( n8804 , n8803 );
buf ( n8805 , n8804 );
buf ( n8806 , n8032 );
not ( n8807 , n8806 );
buf ( n8808 , n8014 );
nor ( n8809 , n8807 , n8808 );
buf ( n8810 , n8809 );
buf ( n8811 , n7967 );
not ( n8812 , n8811 );
buf ( n8813 , n7932 );
not ( n8814 , n8813 );
or ( n8815 , n8812 , n8814 );
buf ( n8816 , n7932 );
buf ( n8817 , n7967 );
or ( n8818 , n8816 , n8817 );
buf ( n8819 , n7948 );
nand ( n8820 , n8818 , n8819 );
buf ( n8821 , n8820 );
buf ( n8822 , n8821 );
nand ( n8823 , n8815 , n8822 );
buf ( n8824 , n8823 );
xor ( n8825 , n8810 , n8824 );
not ( n8826 , n7886 );
buf ( n8827 , n6504 );
not ( n8828 , n8827 );
buf ( n8829 , n4836 );
not ( n8830 , n8829 );
or ( n8831 , n8828 , n8830 );
buf ( n8832 , n7904 );
nand ( n8833 , n8831 , n8832 );
buf ( n8834 , n8833 );
not ( n8835 , n8834 );
or ( n8836 , n8826 , n8835 );
buf ( n8837 , n7886 );
buf ( n8838 , n8834 );
nor ( n8839 , n8837 , n8838 );
buf ( n8840 , n8839 );
or ( n8841 , n8840 , n7864 );
nand ( n8842 , n8836 , n8841 );
xor ( n8843 , n8825 , n8842 );
buf ( n8844 , n8843 );
xor ( n8845 , n8805 , n8844 );
not ( n8846 , n7915 );
not ( n8847 , n7841 );
or ( n8848 , n8846 , n8847 );
not ( n8849 , n7844 );
not ( n8850 , n7914 );
or ( n8851 , n8849 , n8850 );
nand ( n8852 , n8851 , n7970 );
nand ( n8853 , n8848 , n8852 );
buf ( n8854 , n8853 );
xor ( n8855 , n8845 , n8854 );
buf ( n8856 , n8855 );
xor ( n8857 , n7978 , n8066 );
and ( n8858 , n8857 , n8084 );
and ( n8859 , n7978 , n8066 );
or ( n8860 , n8858 , n8859 );
buf ( n8861 , n8860 );
xor ( n8862 , n8856 , n8861 );
buf ( n8863 , n574 );
buf ( n8864 , n575 );
and ( n8865 , n8863 , n8864 );
buf ( n8866 , n4953 );
buf ( n8867 , n8025 );
and ( n8868 , n8866 , n8867 );
nor ( n8869 , n8865 , n8868 );
buf ( n8870 , n8869 );
buf ( n8871 , n8870 );
not ( n8872 , n8871 );
buf ( n8873 , n8872 );
buf ( n8874 , n559 );
buf ( n8875 , n560 );
nand ( n8876 , n8874 , n8875 );
buf ( n8877 , n8876 );
and ( n8878 , n8873 , n8877 );
not ( n8879 , n8873 );
buf ( n8880 , n8877 );
not ( n8881 , n8880 );
buf ( n8882 , n8881 );
and ( n8883 , n8879 , n8882 );
or ( n8884 , n8878 , n8883 );
buf ( n8885 , n7926 );
not ( n8886 , n8885 );
buf ( n8887 , n1243 );
not ( n8888 , n8887 );
or ( n8889 , n8886 , n8888 );
buf ( n8890 , n888 );
buf ( n8891 , n545 );
buf ( n8892 , n572 );
xor ( n8893 , n8891 , n8892 );
buf ( n8894 , n8893 );
buf ( n8895 , n8894 );
nand ( n8896 , n8890 , n8895 );
buf ( n8897 , n8896 );
buf ( n8898 , n8897 );
nand ( n8899 , n8889 , n8898 );
buf ( n8900 , n8899 );
and ( n8901 , n8884 , n8900 );
not ( n8902 , n8884 );
not ( n8903 , n8900 );
and ( n8904 , n8902 , n8903 );
nor ( n8905 , n8901 , n8904 );
not ( n8906 , n8905 );
not ( n8907 , n8906 );
not ( n8908 , n7992 );
not ( n8909 , n6479 );
or ( n8910 , n8908 , n8909 );
buf ( n8911 , n5801 );
buf ( n8912 , n555 );
buf ( n8913 , n562 );
xor ( n8914 , n8912 , n8913 );
buf ( n8915 , n8914 );
buf ( n8916 , n8915 );
nand ( n8917 , n8911 , n8916 );
buf ( n8918 , n8917 );
nand ( n8919 , n8910 , n8918 );
buf ( n8920 , n7880 );
not ( n8921 , n8920 );
buf ( n8922 , n7872 );
not ( n8923 , n8922 );
or ( n8924 , n8921 , n8923 );
buf ( n8925 , n1979 );
buf ( n8926 , n547 );
buf ( n8927 , n570 );
xor ( n8928 , n8926 , n8927 );
buf ( n8929 , n8928 );
buf ( n8930 , n8929 );
nand ( n8931 , n8925 , n8930 );
buf ( n8932 , n8931 );
buf ( n8933 , n8932 );
nand ( n8934 , n8924 , n8933 );
buf ( n8935 , n8934 );
xor ( n8936 , n8919 , n8935 );
buf ( n8937 , n7901 );
not ( n8938 , n8937 );
buf ( n8939 , n5678 );
not ( n8940 , n8939 );
or ( n8941 , n8938 , n8940 );
buf ( n8942 , n4840 );
buf ( n8943 , n553 );
buf ( n8944 , n564 );
xor ( n8945 , n8943 , n8944 );
buf ( n8946 , n8945 );
buf ( n8947 , n8946 );
nand ( n8948 , n8942 , n8947 );
buf ( n8949 , n8948 );
buf ( n8950 , n8949 );
nand ( n8951 , n8941 , n8950 );
buf ( n8952 , n8951 );
xnor ( n8953 , n8936 , n8952 );
buf ( n8954 , n8953 );
not ( n8955 , n8954 );
buf ( n8956 , n8955 );
not ( n8957 , n8956 );
or ( n8958 , n8907 , n8957 );
buf ( n8959 , n8953 );
buf ( n8960 , n8905 );
nand ( n8961 , n8959 , n8960 );
buf ( n8962 , n8961 );
nand ( n8963 , n8958 , n8962 );
buf ( n8964 , n8963 );
not ( n8965 , n6595 );
and ( n8966 , n557 , n560 );
not ( n8967 , n557 );
and ( n8968 , n8967 , n7962 );
nor ( n8969 , n8966 , n8968 );
not ( n8970 , n8969 );
or ( n8971 , n8965 , n8970 );
nand ( n8972 , n7955 , n7964 );
nand ( n8973 , n8971 , n8972 );
buf ( n8974 , n8973 );
not ( n8975 , n7942 );
not ( n8976 , n4958 );
or ( n8977 , n8975 , n8976 );
and ( n8978 , n549 , n568 );
not ( n8979 , n549 );
and ( n8980 , n8979 , n3015 );
nor ( n8981 , n8978 , n8980 );
nand ( n8982 , n3436 , n8981 );
nand ( n8983 , n8977 , n8982 );
buf ( n8984 , n8983 );
xor ( n8985 , n8974 , n8984 );
buf ( n8986 , n7855 );
not ( n8987 , n8986 );
buf ( n8988 , n4380 );
not ( n8989 , n8988 );
or ( n8990 , n8987 , n8989 );
buf ( n8991 , n3743 );
buf ( n8992 , n551 );
buf ( n8993 , n566 );
xor ( n8994 , n8992 , n8993 );
buf ( n8995 , n8994 );
buf ( n8996 , n8995 );
nand ( n8997 , n8991 , n8996 );
buf ( n8998 , n8997 );
buf ( n8999 , n8998 );
nand ( n9000 , n8990 , n8999 );
buf ( n9001 , n9000 );
buf ( n9002 , n9001 );
xor ( n9003 , n8985 , n9002 );
buf ( n9004 , n9003 );
buf ( n9005 , n9004 );
xor ( n9006 , n8964 , n9005 );
buf ( n9007 , n9006 );
xor ( n9008 , n8862 , n9007 );
not ( n9009 , n9008 );
not ( n9010 , n9009 );
xor ( n9011 , n8109 , n8115 );
and ( n9012 , n9011 , n8326 );
and ( n9013 , n8109 , n8115 );
or ( n9014 , n9012 , n9013 );
buf ( n9015 , n9014 );
not ( n9016 , n9015 );
or ( n9017 , n9010 , n9016 );
not ( n9018 , n9015 );
nand ( n9019 , n9018 , n9008 );
nand ( n9020 , n9017 , n9019 );
xor ( n9021 , n8228 , n8240 );
and ( n9022 , n9021 , n8323 );
and ( n9023 , n8228 , n8240 );
or ( n9024 , n9022 , n9023 );
buf ( n9025 , n9024 );
buf ( n9026 , n7971 );
not ( n9027 , n9026 );
buf ( n9028 , n9027 );
buf ( n9029 , n9028 );
not ( n9030 , n9029 );
buf ( n9031 , n8086 );
not ( n9032 , n9031 );
or ( n9033 , n9030 , n9032 );
buf ( n9034 , n8086 );
buf ( n9035 , n9028 );
or ( n9036 , n9034 , n9035 );
buf ( n9037 , n7835 );
nand ( n9038 , n9036 , n9037 );
buf ( n9039 , n9038 );
buf ( n9040 , n9039 );
nand ( n9041 , n9033 , n9040 );
buf ( n9042 , n9041 );
xor ( n9043 , n9025 , n9042 );
buf ( n9044 , n8296 );
not ( n9045 , n9044 );
buf ( n9046 , n6349 );
buf ( n9047 , n6344 );
nor ( n9048 , n9046 , n9047 );
buf ( n9049 , n9048 );
buf ( n9050 , n9049 );
not ( n9051 , n9050 );
or ( n9052 , n9045 , n9051 );
buf ( n9053 , n5997 );
xor ( n9054 , n578 , n555 );
buf ( n9055 , n9054 );
nand ( n9056 , n9053 , n9055 );
buf ( n9057 , n9056 );
buf ( n9058 , n9057 );
nand ( n9059 , n9052 , n9058 );
buf ( n9060 , n9059 );
not ( n9061 , n8134 );
not ( n9062 , n1177 );
or ( n9063 , n9061 , n9062 );
buf ( n9064 , n1036 );
buf ( n9065 , n547 );
buf ( n9066 , n586 );
xor ( n9067 , n9065 , n9066 );
buf ( n9068 , n9067 );
buf ( n9069 , n9068 );
nand ( n9070 , n9064 , n9069 );
buf ( n9071 , n9070 );
nand ( n9072 , n9063 , n9071 );
xor ( n9073 , n9060 , n9072 );
not ( n9074 , n8121 );
not ( n9075 , n5060 );
or ( n9076 , n9074 , n9075 );
buf ( n9077 , n4544 );
xor ( n9078 , n580 , n553 );
buf ( n9079 , n9078 );
nand ( n9080 , n9077 , n9079 );
buf ( n9081 , n9080 );
nand ( n9082 , n9076 , n9081 );
xor ( n9083 , n9073 , n9082 );
buf ( n9084 , n8275 );
not ( n9085 , n9084 );
buf ( n9086 , n984 );
not ( n9087 , n9086 );
or ( n9088 , n9085 , n9087 );
buf ( n9089 , n590 );
buf ( n9090 , n591 );
nand ( n9091 , n9089 , n9090 );
buf ( n9092 , n9091 );
buf ( n9093 , n9092 );
nand ( n9094 , n9088 , n9093 );
buf ( n9095 , n9094 );
buf ( n9096 , n559 );
buf ( n9097 , n576 );
nand ( n9098 , n9096 , n9097 );
buf ( n9099 , n9098 );
xor ( n9100 , n9095 , n9099 );
buf ( n9101 , n8181 );
not ( n9102 , n9101 );
buf ( n9103 , n3639 );
not ( n9104 , n9103 );
or ( n9105 , n9102 , n9104 );
buf ( n9106 , n545 );
buf ( n9107 , n588 );
xor ( n9108 , n9106 , n9107 );
buf ( n9109 , n9108 );
buf ( n9110 , n9109 );
buf ( n9111 , n1071 );
nand ( n9112 , n9110 , n9111 );
buf ( n9113 , n9112 );
buf ( n9114 , n9113 );
nand ( n9115 , n9105 , n9114 );
buf ( n9116 , n9115 );
xor ( n9117 , n9100 , n9116 );
not ( n9118 , n9117 );
xor ( n9119 , n9083 , n9118 );
buf ( n9120 , n8203 );
not ( n9121 , n9120 );
buf ( n9122 , n8196 );
not ( n9123 , n9122 );
or ( n9124 , n9121 , n9123 );
buf ( n9125 , n6699 );
buf ( n9126 , n557 );
buf ( n9127 , n576 );
xor ( n9128 , n9126 , n9127 );
buf ( n9129 , n9128 );
buf ( n9130 , n9129 );
nand ( n9131 , n9125 , n9130 );
buf ( n9132 , n9131 );
buf ( n9133 , n9132 );
nand ( n9134 , n9124 , n9133 );
buf ( n9135 , n9134 );
buf ( n9136 , n9135 );
buf ( n9137 , n8149 );
not ( n9138 , n9137 );
buf ( n9139 , n4506 );
not ( n9140 , n9139 );
or ( n9141 , n9138 , n9140 );
buf ( n9142 , n3883 );
buf ( n9143 , n551 );
buf ( n9144 , n582 );
xor ( n9145 , n9143 , n9144 );
buf ( n9146 , n9145 );
buf ( n9147 , n9146 );
nand ( n9148 , n9142 , n9147 );
buf ( n9149 , n9148 );
buf ( n9150 , n9149 );
nand ( n9151 , n9141 , n9150 );
buf ( n9152 , n9151 );
buf ( n9153 , n9152 );
xor ( n9154 , n9136 , n9153 );
buf ( n9155 , n8216 );
not ( n9156 , n9155 );
buf ( n9157 , n3664 );
not ( n9158 , n9157 );
or ( n9159 , n9156 , n9158 );
buf ( n9160 , n4232 );
buf ( n9161 , n549 );
buf ( n9162 , n584 );
xor ( n9163 , n9161 , n9162 );
buf ( n9164 , n9163 );
buf ( n9165 , n9164 );
nand ( n9166 , n9160 , n9165 );
buf ( n9167 , n9166 );
buf ( n9168 , n9167 );
nand ( n9169 , n9159 , n9168 );
buf ( n9170 , n9169 );
buf ( n9171 , n9170 );
xnor ( n9172 , n9154 , n9171 );
buf ( n9173 , n9172 );
buf ( n9174 , n9173 );
not ( n9175 , n9174 );
buf ( n9176 , n9175 );
xor ( n9177 , n9119 , n9176 );
buf ( n9178 , n9177 );
xor ( n9179 , n8250 , n8313 );
and ( n9180 , n9179 , n8320 );
and ( n9181 , n8250 , n8313 );
or ( n9182 , n9180 , n9181 );
buf ( n9183 , n9182 );
buf ( n9184 , n9183 );
xor ( n9185 , n9178 , n9184 );
xor ( n9186 , n8286 , n8303 );
and ( n9187 , n9186 , n8310 );
and ( n9188 , n8286 , n8303 );
or ( n9189 , n9187 , n9188 );
buf ( n9190 , n9189 );
buf ( n9191 , n9190 );
buf ( n9192 , n8166 );
not ( n9193 , n9192 );
buf ( n9194 , n8221 );
not ( n9195 , n9194 );
or ( n9196 , n9193 , n9195 );
buf ( n9197 , n8156 );
nand ( n9198 , n9196 , n9197 );
buf ( n9199 , n9198 );
buf ( n9200 , n9199 );
buf ( n9201 , n8221 );
not ( n9202 , n9201 );
buf ( n9203 , n8165 );
nand ( n9204 , n9202 , n9203 );
buf ( n9205 , n9204 );
buf ( n9206 , n9205 );
nand ( n9207 , n9200 , n9206 );
buf ( n9208 , n9207 );
buf ( n9209 , n9208 );
xor ( n9210 , n9191 , n9209 );
and ( n9211 , n8266 , n8283 );
buf ( n9212 , n9211 );
buf ( n9213 , n9212 );
xor ( n9214 , n8125 , n8138 );
and ( n9215 , n9214 , n8155 );
and ( n9216 , n8125 , n8138 );
or ( n9217 , n9215 , n9216 );
buf ( n9218 , n9217 );
xor ( n9219 , n9213 , n9218 );
not ( n9220 , n8183 );
not ( n9221 , n8207 );
or ( n9222 , n9220 , n9221 );
or ( n9223 , n8183 , n8207 );
nand ( n9224 , n9223 , n8220 );
nand ( n9225 , n9222 , n9224 );
buf ( n9226 , n9225 );
xor ( n9227 , n9219 , n9226 );
buf ( n9228 , n9227 );
buf ( n9229 , n9228 );
xor ( n9230 , n9210 , n9229 );
buf ( n9231 , n9230 );
buf ( n9232 , n9231 );
xor ( n9233 , n9185 , n9232 );
buf ( n9234 , n9233 );
xor ( n9235 , n9043 , n9234 );
and ( n9236 , n9020 , n9235 );
not ( n9237 , n9020 );
not ( n9238 , n9235 );
and ( n9239 , n9237 , n9238 );
nor ( n9240 , n9236 , n9239 );
xor ( n9241 , n8088 , n8093 );
and ( n9242 , n9241 , n8329 );
and ( n9243 , n8088 , n8093 );
or ( n9244 , n9242 , n9243 );
buf ( n9245 , n9244 );
nor ( n9246 , n9240 , n9245 );
not ( n9247 , n9246 );
nand ( n9248 , n9245 , n9240 );
and ( n9249 , n9247 , n9248 );
not ( n9250 , n9249 );
not ( n9251 , n9250 );
buf ( n9252 , n6437 );
not ( n9253 , n9252 );
buf ( n9254 , n8331 );
buf ( n9255 , n8337 );
nor ( n9256 , n9254 , n9255 );
buf ( n9257 , n9256 );
buf ( n9258 , n9257 );
buf ( n9259 , n6879 );
nor ( n9260 , n9258 , n9259 );
buf ( n9261 , n9260 );
buf ( n9262 , n9261 );
not ( n9263 , n9262 );
or ( n9264 , n9253 , n9263 );
buf ( n9265 , n8351 );
buf ( n9266 , n6887 );
not ( n9267 , n9266 );
buf ( n9268 , n9267 );
buf ( n9269 , n9268 );
and ( n9270 , n9265 , n9269 );
buf ( n9271 , n8340 );
nor ( n9272 , n9270 , n9271 );
buf ( n9273 , n9272 );
buf ( n9274 , n9273 );
nand ( n9275 , n9264 , n9274 );
buf ( n9276 , n9275 );
buf ( n9277 , n9276 );
not ( n9278 , n9277 );
buf ( n9279 , n9278 );
buf ( n9280 , n9279 );
buf ( n9281 , n9257 );
buf ( n9282 , n6879 );
nor ( n9283 , n9281 , n9282 );
buf ( n9284 , n9283 );
nand ( n9285 , n6469 , n9284 , n6449 );
buf ( n9286 , n9285 );
buf ( n9287 , n6441 );
buf ( n9288 , n9284 );
buf ( n9289 , n6449 );
buf ( n9290 , n6454 );
nand ( n9291 , n9287 , n9288 , n9289 , n9290 );
buf ( n9292 , n9291 );
buf ( n9293 , n9292 );
and ( n9294 , n9280 , n9286 , n9293 );
buf ( n9295 , n9294 );
buf ( n9296 , n9295 );
buf ( n9297 , n9296 );
buf ( n9298 , n9297 );
buf ( n9299 , n9298 );
not ( n9300 , n9299 );
buf ( n9301 , n9300 );
not ( n9302 , n9301 );
or ( n9303 , n9251 , n9302 );
nand ( n9304 , n9249 , n9298 );
nand ( n9305 , n9303 , n9304 );
xor ( n9306 , n8405 , n8412 );
and ( n9307 , n9306 , n8449 );
and ( n9308 , n8405 , n8412 );
or ( n9309 , n9307 , n9308 );
and ( n9310 , n8472 , n8490 );
not ( n9311 , n3068 );
not ( n9312 , n3073 );
not ( n9313 , n3036 );
or ( n9314 , n9312 , n9313 );
nand ( n9315 , n3037 , n550 );
nand ( n9316 , n9314 , n9315 );
not ( n9317 , n9316 );
or ( n9318 , n9311 , n9317 );
not ( n9319 , n2981 );
not ( n9320 , n3073 );
or ( n9321 , n9319 , n9320 );
or ( n9322 , n3073 , n2981 );
nand ( n9323 , n9321 , n9322 );
nand ( n9324 , n9323 , n5268 );
nand ( n9325 , n9318 , n9324 );
xor ( n9326 , n9310 , n9325 );
buf ( n9327 , n3212 );
not ( n9328 , n9327 );
not ( n9329 , n548 );
not ( n9330 , n2252 );
or ( n9331 , n9329 , n9330 );
nand ( n9332 , n2251 , n5279 );
nand ( n9333 , n9331 , n9332 );
not ( n9334 , n9333 );
or ( n9335 , n9328 , n9334 );
nand ( n9336 , n8498 , n6939 );
nand ( n9337 , n9335 , n9336 );
xor ( n9338 , n9326 , n9337 );
xor ( n9339 , n9309 , n9338 );
xor ( n9340 , n8380 , n8384 );
and ( n9341 , n9340 , n8395 );
and ( n9342 , n8380 , n8384 );
or ( n9343 , n9341 , n9342 );
xor ( n9344 , n9339 , n9343 );
not ( n9345 , n3064 );
not ( n9346 , n552 );
not ( n9347 , n5201 );
or ( n9348 , n9346 , n9347 );
not ( n9349 , n552 );
nand ( n9350 , n9349 , n3167 );
nand ( n9351 , n9348 , n9350 );
not ( n9352 , n9351 );
or ( n9353 , n9345 , n9352 );
xor ( n9354 , n3264 , n552 );
nand ( n9355 , n9354 , n5299 );
nand ( n9356 , n9353 , n9355 );
not ( n9357 , n1739 );
not ( n9358 , n8445 );
or ( n9359 , n9357 , n9358 );
not ( n9360 , n1736 );
nor ( n9361 , n8431 , n7265 );
nand ( n9362 , n7253 , n9361 );
nor ( n9363 , n9362 , n7095 );
not ( n9364 , n9363 );
not ( n9365 , n3034 );
or ( n9366 , n9364 , n9365 );
and ( n9367 , n7253 , n9361 );
and ( n9368 , n7112 , n9367 );
not ( n9369 , n9361 );
not ( n9370 , n7258 );
or ( n9371 , n9369 , n9370 );
or ( n9372 , n8431 , n7232 );
nand ( n9373 , n9372 , n8433 );
not ( n9374 , n9373 );
nand ( n9375 , n9371 , n9374 );
nor ( n9376 , n9368 , n9375 );
nand ( n9377 , n9366 , n9376 );
not ( n9378 , n9377 );
not ( n9379 , n9378 );
not ( n9380 , n9379 );
or ( n9381 , n9360 , n9380 );
not ( n9382 , n9379 );
nand ( n9383 , n9382 , n558 );
nand ( n9384 , n9381 , n9383 );
nand ( n9385 , n559 , n9384 );
nand ( n9386 , n9359 , n9385 );
xor ( n9387 , n9356 , n9386 );
not ( n9388 , n8374 );
or ( n9389 , n9388 , n1658 );
and ( n9390 , n7276 , n1625 );
not ( n9391 , n7276 );
and ( n9392 , n9391 , n556 );
or ( n9393 , n9390 , n9392 );
not ( n9394 , n9393 );
or ( n9395 , n9394 , n1595 );
nand ( n9396 , n9389 , n9395 );
xor ( n9397 , n9387 , n9396 );
not ( n9398 , n6906 );
not ( n9399 , n8391 );
or ( n9400 , n9398 , n9399 );
not ( n9401 , n554 );
not ( n9402 , n7125 );
or ( n9403 , n9401 , n9402 );
nand ( n9404 , n7124 , n1681 );
nand ( n9405 , n9403 , n9404 );
nand ( n9406 , n9405 , n3118 );
nand ( n9407 , n9400 , n9406 );
nor ( n9408 , n1687 , n8477 );
buf ( n9409 , n7170 );
not ( n9410 , n9409 );
and ( n9411 , n1652 , n544 );
not ( n9412 , n1652 );
and ( n9413 , n9412 , n8477 );
or ( n9414 , n9411 , n9413 );
not ( n9415 , n9414 );
or ( n9416 , n9410 , n9415 );
nor ( n9417 , n8487 , n7170 );
nand ( n9418 , n8479 , n9417 );
nand ( n9419 , n9416 , n9418 );
xor ( n9420 , n9408 , n9419 );
not ( n9421 , n6945 );
and ( n9422 , n2220 , n546 );
not ( n9423 , n2220 );
and ( n9424 , n9423 , n6949 );
or ( n9425 , n9422 , n9424 );
not ( n9426 , n9425 );
or ( n9427 , n9421 , n9426 );
nand ( n9428 , n8461 , n8466 );
nand ( n9429 , n9427 , n9428 );
xor ( n9430 , n9420 , n9429 );
xor ( n9431 , n9407 , n9430 );
xor ( n9432 , n8468 , n8491 );
and ( n9433 , n9432 , n8502 );
and ( n9434 , n8468 , n8491 );
or ( n9435 , n9433 , n9434 );
xor ( n9436 , n9431 , n9435 );
xor ( n9437 , n9397 , n9436 );
xor ( n9438 , n8455 , n8503 );
and ( n9439 , n9438 , n8508 );
and ( n9440 , n8455 , n8503 );
or ( n9441 , n9439 , n9440 );
xor ( n9442 , n9437 , n9441 );
xor ( n9443 , n9344 , n9442 );
xor ( n9444 , n8396 , n8450 );
and ( n9445 , n9444 , n8509 );
and ( n9446 , n8396 , n8450 );
or ( n9447 , n9445 , n9446 );
xor ( n9448 , n9443 , n9447 );
xor ( n9449 , n8362 , n8366 );
and ( n9450 , n9449 , n8510 );
and ( n9451 , n8362 , n8366 );
or ( n9452 , n9450 , n9451 );
or ( n9453 , n9448 , n9452 );
nand ( n9454 , n9448 , n9452 );
nand ( n9455 , n9453 , n9454 );
not ( n9456 , n9455 );
not ( n9457 , n7300 );
not ( n9458 , n7323 );
and ( n9459 , n9457 , n9458 );
nor ( n9460 , n7352 , n7356 );
nor ( n9461 , n9459 , n9460 );
nand ( n9462 , n8518 , n7360 , n9461 );
or ( n9463 , n8520 , n8516 );
and ( n9464 , n7300 , n7323 );
nand ( n9465 , n9463 , n9464 );
nand ( n9466 , n9462 , n8521 , n9465 );
buf ( n9467 , n9466 );
not ( n9468 , n9467 );
not ( n9469 , n9468 );
or ( n9470 , n9456 , n9469 );
or ( n9471 , n9455 , n9468 );
nand ( n9472 , n9470 , n9471 );
nand ( n9473 , n9305 , n9472 );
buf ( n9474 , n9473 );
not ( n9475 , n9305 );
not ( n9476 , n9472 );
nand ( n9477 , n9475 , n9476 );
buf ( n9478 , n9477 );
nand ( n9479 , n9474 , n9478 );
not ( n9480 , n9479 );
not ( n9481 , n6903 );
not ( n9482 , n7367 );
and ( n9483 , n9481 , n9482 );
not ( n9484 , n8357 );
and ( n9485 , n8529 , n9484 );
nor ( n9486 , n9483 , n9485 );
nand ( n9487 , n9486 , n7440 , n7493 );
nand ( n9488 , n9486 , n7451 );
and ( n9489 , n8532 , n7372 );
nor ( n9490 , n9489 , n8530 );
nand ( n9491 , n9487 , n9488 , n9490 );
buf ( n9492 , n9491 );
not ( n9493 , n9492 );
or ( n9494 , n9480 , n9493 );
or ( n9495 , n9479 , n9492 );
nand ( n9496 , n9494 , n9495 );
buf ( n9497 , n9496 );
not ( n9498 , n9497 );
not ( n9499 , n9498 );
nand ( n9500 , n8541 , n7809 );
nand ( n9501 , n9500 , n7520 );
not ( n9502 , n9501 );
buf ( n9503 , n7795 );
buf ( n9504 , n7514 );
nand ( n9505 , n9502 , n9503 , n9504 );
not ( n9506 , n7554 );
not ( n9507 , n7795 );
not ( n9508 , n8541 );
nor ( n9509 , n9508 , n576 );
nor ( n9510 , n9507 , n9509 );
and ( n9511 , n9506 , n9510 );
nor ( n9512 , n8542 , n576 );
or ( n9513 , n9512 , n7800 );
nand ( n9514 , n9513 , n8546 );
nor ( n9515 , n9511 , n9514 );
nand ( n9516 , n9505 , n9515 );
buf ( n9517 , n9516 );
not ( n9518 , n9517 );
or ( n9519 , n9499 , n9518 );
not ( n9520 , n9516 );
not ( n9521 , n9520 );
or ( n9522 , n9521 , n9498 );
nand ( n9523 , n9519 , n9522 );
not ( n9524 , n9523 );
and ( n9525 , n604 , n9524 );
not ( n9526 , n604 );
buf ( n9527 , n9523 );
and ( n9528 , n9526 , n9527 );
or ( n9529 , n9525 , n9528 );
buf ( n9530 , n9529 );
not ( n9531 , n9530 );
or ( n9532 , n8799 , n9531 );
buf ( n9533 , n8559 );
buf ( n9534 , n8581 );
nand ( n9535 , n9533 , n9534 );
buf ( n9536 , n9535 );
buf ( n9537 , n9536 );
nand ( n9538 , n9532 , n9537 );
buf ( n9539 , n9538 );
buf ( n9540 , n9539 );
xor ( n9541 , n8797 , n9540 );
buf ( n9542 , n607 );
not ( n9543 , n9542 );
buf ( n9544 , n606 );
not ( n9545 , n9544 );
not ( n9546 , n9520 );
not ( n9547 , n9478 );
buf ( n9548 , n9491 );
not ( n9549 , n9548 );
or ( n9550 , n9547 , n9549 );
nand ( n9551 , n9550 , n9474 );
not ( n9552 , n9453 );
not ( n9553 , n9467 );
or ( n9554 , n9552 , n9553 );
nand ( n9555 , n9554 , n9454 );
xor ( n9556 , n9344 , n9442 );
and ( n9557 , n9556 , n9447 );
and ( n9558 , n9344 , n9442 );
or ( n9559 , n9557 , n9558 );
xor ( n9560 , n9356 , n9386 );
and ( n9561 , n9560 , n9396 );
and ( n9562 , n9356 , n9386 );
or ( n9563 , n9561 , n9562 );
not ( n9564 , n6939 );
not ( n9565 , n9333 );
or ( n9566 , n9564 , n9565 );
not ( n9567 , n548 );
not ( n9568 , n5186 );
or ( n9569 , n9567 , n9568 );
nand ( n9570 , n2981 , n5279 );
nand ( n9571 , n9569 , n9570 );
nand ( n9572 , n9571 , n3212 );
nand ( n9573 , n9566 , n9572 );
not ( n9574 , n9425 );
and ( n9575 , n7178 , n8464 );
not ( n9576 , n9575 );
or ( n9577 , n9574 , n9576 );
not ( n9578 , n5304 );
not ( n9579 , n6949 );
and ( n9580 , n9578 , n9579 );
and ( n9581 , n5304 , n6949 );
nor ( n9582 , n9580 , n9581 );
nand ( n9583 , n9582 , n6945 );
nand ( n9584 , n9577 , n9583 );
xor ( n9585 , n9573 , n9584 );
xnor ( n9586 , n5250 , n552 );
not ( n9587 , n5299 );
or ( n9588 , n9586 , n9587 );
nand ( n9589 , n9354 , n3064 );
nand ( n9590 , n9588 , n9589 );
xor ( n9591 , n9585 , n9590 );
xor ( n9592 , n9563 , n9591 );
nand ( n9593 , n8440 , n1625 , n7069 );
nand ( n9594 , n1659 , n9393 );
nand ( n9595 , n8441 , n7069 , n556 );
nand ( n9596 , n9593 , n9594 , n9595 );
not ( n9597 , n9316 );
not ( n9598 , n5268 );
or ( n9599 , n9597 , n9598 );
and ( n9600 , n3167 , n550 );
not ( n9601 , n3167 );
and ( n9602 , n9601 , n3073 );
nor ( n9603 , n9600 , n9602 );
not ( n9604 , n9603 );
not ( n9605 , n3068 );
or ( n9606 , n9604 , n9605 );
nand ( n9607 , n9599 , n9606 );
xor ( n9608 , n9596 , n9607 );
xor ( n9609 , n9408 , n9419 );
and ( n9610 , n9609 , n9429 );
and ( n9611 , n9408 , n9419 );
or ( n9612 , n9610 , n9611 );
xor ( n9613 , n9608 , n9612 );
xor ( n9614 , n9592 , n9613 );
not ( n9615 , n2276 );
not ( n9616 , n9405 );
or ( n9617 , n9615 , n9616 );
not ( n9618 , n3118 );
not ( n9619 , n9618 );
not ( n9620 , n554 );
not ( n9621 , n7223 );
or ( n9622 , n9620 , n9621 );
nand ( n9623 , n7222 , n1681 );
nand ( n9624 , n9622 , n9623 );
nand ( n9625 , n9619 , n9624 );
nand ( n9626 , n9617 , n9625 );
not ( n9627 , n9409 );
not ( n9628 , n544 );
not ( n9629 , n1621 );
or ( n9630 , n9628 , n9629 );
nand ( n9631 , n5261 , n8477 );
nand ( n9632 , n9630 , n9631 );
not ( n9633 , n9632 );
or ( n9634 , n9627 , n9633 );
nand ( n9635 , n9417 , n9414 );
nand ( n9636 , n9634 , n9635 );
not ( n9637 , n544 );
nor ( n9638 , n9637 , n1677 );
xor ( n9639 , n9636 , n9638 );
not ( n9640 , n1739 );
not ( n9641 , n9384 );
or ( n9642 , n9640 , n9641 );
nand ( n9643 , n9642 , n1774 );
xor ( n9644 , n9639 , n9643 );
xor ( n9645 , n9626 , n9644 );
xor ( n9646 , n9310 , n9325 );
and ( n9647 , n9646 , n9337 );
and ( n9648 , n9310 , n9325 );
or ( n9649 , n9647 , n9648 );
xor ( n9650 , n9645 , n9649 );
xor ( n9651 , n9407 , n9430 );
and ( n9652 , n9651 , n9435 );
and ( n9653 , n9407 , n9430 );
or ( n9654 , n9652 , n9653 );
xor ( n9655 , n9650 , n9654 );
xor ( n9656 , n9309 , n9338 );
and ( n9657 , n9656 , n9343 );
and ( n9658 , n9309 , n9338 );
or ( n9659 , n9657 , n9658 );
xor ( n9660 , n9655 , n9659 );
xor ( n9661 , n9614 , n9660 );
xor ( n9662 , n9397 , n9436 );
and ( n9663 , n9662 , n9441 );
and ( n9664 , n9397 , n9436 );
or ( n9665 , n9663 , n9664 );
xor ( n9666 , n9661 , n9665 );
nor ( n9667 , n9559 , n9666 );
not ( n9668 , n9667 );
not ( n9669 , n9666 );
not ( n9670 , n9559 );
nor ( n9671 , n9669 , n9670 );
not ( n9672 , n9671 );
and ( n9673 , n9668 , n9672 );
and ( n9674 , n9555 , n9673 );
not ( n9675 , n9555 );
not ( n9676 , n9673 );
and ( n9677 , n9675 , n9676 );
nor ( n9678 , n9674 , n9677 );
not ( n9679 , n9678 );
not ( n9680 , n9247 );
nand ( n9681 , n9279 , n9285 , n9292 );
not ( n9682 , n9681 );
or ( n9683 , n9680 , n9682 );
nand ( n9684 , n9683 , n9248 );
xor ( n9685 , n8805 , n8844 );
and ( n9686 , n9685 , n8854 );
and ( n9687 , n8805 , n8844 );
or ( n9688 , n9686 , n9687 );
buf ( n9689 , n9688 );
buf ( n9690 , n574 );
buf ( n9691 , n558 );
buf ( n9692 , n560 );
nand ( n9693 , n9691 , n9692 );
buf ( n9694 , n9693 );
buf ( n9695 , n9694 );
xor ( n9696 , n9690 , n9695 );
not ( n9697 , n6595 );
buf ( n9698 , n556 );
buf ( n9699 , n560 );
xor ( n9700 , n9698 , n9699 );
buf ( n9701 , n9700 );
not ( n9702 , n9701 );
or ( n9703 , n9697 , n9702 );
nand ( n9704 , n7964 , n8969 );
nand ( n9705 , n9703 , n9704 );
buf ( n9706 , n9705 );
xnor ( n9707 , n9696 , n9706 );
buf ( n9708 , n9707 );
buf ( n9709 , n9708 );
not ( n9710 , n9709 );
buf ( n9711 , n9710 );
buf ( n9712 , n9711 );
not ( n9713 , n9712 );
buf ( n9714 , n8894 );
not ( n9715 , n9714 );
buf ( n9716 , n1243 );
not ( n9717 , n9716 );
or ( n9718 , n9715 , n9717 );
buf ( n9719 , n888 );
buf ( n9720 , n544 );
buf ( n9721 , n572 );
xor ( n9722 , n9720 , n9721 );
buf ( n9723 , n9722 );
buf ( n9724 , n9723 );
nand ( n9725 , n9719 , n9724 );
buf ( n9726 , n9725 );
buf ( n9727 , n9726 );
nand ( n9728 , n9718 , n9727 );
buf ( n9729 , n9728 );
buf ( n9730 , n8929 );
not ( n9731 , n9730 );
buf ( n9732 , n1973 );
not ( n9733 , n9732 );
or ( n9734 , n9731 , n9733 );
buf ( n9735 , n1979 );
buf ( n9736 , n546 );
buf ( n9737 , n570 );
xor ( n9738 , n9736 , n9737 );
buf ( n9739 , n9738 );
buf ( n9740 , n9739 );
nand ( n9741 , n9735 , n9740 );
buf ( n9742 , n9741 );
buf ( n9743 , n9742 );
nand ( n9744 , n9734 , n9743 );
buf ( n9745 , n9744 );
xor ( n9746 , n9729 , n9745 );
buf ( n9747 , n8995 );
not ( n9748 , n9747 );
buf ( n9749 , n4380 );
not ( n9750 , n9749 );
or ( n9751 , n9748 , n9750 );
buf ( n9752 , n3743 );
xor ( n9753 , n566 , n550 );
buf ( n9754 , n9753 );
nand ( n9755 , n9752 , n9754 );
buf ( n9756 , n9755 );
buf ( n9757 , n9756 );
nand ( n9758 , n9751 , n9757 );
buf ( n9759 , n9758 );
not ( n9760 , n9759 );
and ( n9761 , n9746 , n9760 );
not ( n9762 , n9746 );
and ( n9763 , n9762 , n9759 );
nor ( n9764 , n9761 , n9763 );
buf ( n9765 , n9764 );
not ( n9766 , n9765 );
or ( n9767 , n9713 , n9766 );
not ( n9768 , n9764 );
nand ( n9769 , n9768 , n9708 );
buf ( n9770 , n9769 );
nand ( n9771 , n9767 , n9770 );
buf ( n9772 , n9771 );
buf ( n9773 , n9772 );
xor ( n9774 , n8810 , n8824 );
and ( n9775 , n9774 , n8842 );
and ( n9776 , n8810 , n8824 );
or ( n9777 , n9775 , n9776 );
buf ( n9778 , n9777 );
not ( n9779 , n9778 );
buf ( n9780 , n9779 );
buf ( n9781 , n9780 );
and ( n9782 , n9773 , n9781 );
not ( n9783 , n9773 );
buf ( n9784 , n9777 );
and ( n9785 , n9783 , n9784 );
nor ( n9786 , n9782 , n9785 );
buf ( n9787 , n9786 );
and ( n9788 , n9689 , n9787 );
not ( n9789 , n9689 );
buf ( n9790 , n9787 );
not ( n9791 , n9790 );
buf ( n9792 , n9791 );
and ( n9793 , n9789 , n9792 );
or ( n9794 , n9788 , n9793 );
buf ( n9795 , n8915 );
not ( n9796 , n9795 );
nor ( n9797 , n5813 , n5818 );
buf ( n9798 , n9797 );
buf ( n9799 , n9798 );
not ( n9800 , n9799 );
or ( n9801 , n9796 , n9800 );
buf ( n9802 , n5801 );
buf ( n9803 , n554 );
buf ( n9804 , n562 );
xor ( n9805 , n9803 , n9804 );
buf ( n9806 , n9805 );
buf ( n9807 , n9806 );
nand ( n9808 , n9802 , n9807 );
buf ( n9809 , n9808 );
buf ( n9810 , n9809 );
nand ( n9811 , n9801 , n9810 );
buf ( n9812 , n9811 );
buf ( n9813 , n8946 );
not ( n9814 , n9813 );
buf ( n9815 , n4836 );
not ( n9816 , n9815 );
or ( n9817 , n9814 , n9816 );
buf ( n9818 , n4840 );
buf ( n9819 , n552 );
buf ( n9820 , n564 );
xor ( n9821 , n9819 , n9820 );
buf ( n9822 , n9821 );
buf ( n9823 , n9822 );
nand ( n9824 , n9818 , n9823 );
buf ( n9825 , n9824 );
buf ( n9826 , n9825 );
nand ( n9827 , n9817 , n9826 );
buf ( n9828 , n9827 );
xor ( n9829 , n9812 , n9828 );
buf ( n9830 , n8981 );
not ( n9831 , n9830 );
buf ( n9832 , n3429 );
not ( n9833 , n9832 );
or ( n9834 , n9831 , n9833 );
buf ( n9835 , n3439 );
buf ( n9836 , n548 );
buf ( n9837 , n568 );
xor ( n9838 , n9836 , n9837 );
buf ( n9839 , n9838 );
buf ( n9840 , n9839 );
nand ( n9841 , n9835 , n9840 );
buf ( n9842 , n9841 );
buf ( n9843 , n9842 );
nand ( n9844 , n9834 , n9843 );
buf ( n9845 , n9844 );
xor ( n9846 , n9829 , n9845 );
buf ( n9847 , n8900 );
not ( n9848 , n9847 );
buf ( n9849 , n8870 );
buf ( n9850 , n8877 );
nand ( n9851 , n9849 , n9850 );
buf ( n9852 , n9851 );
buf ( n9853 , n9852 );
not ( n9854 , n9853 );
or ( n9855 , n9848 , n9854 );
buf ( n9856 , n8873 );
buf ( n9857 , n8882 );
nand ( n9858 , n9856 , n9857 );
buf ( n9859 , n9858 );
buf ( n9860 , n9859 );
nand ( n9861 , n9855 , n9860 );
buf ( n9862 , n9861 );
buf ( n9863 , n9862 );
or ( n9864 , n8919 , n8952 );
nand ( n9865 , n9864 , n8935 );
buf ( n9866 , n9865 );
nand ( n9867 , n8952 , n8919 );
buf ( n9868 , n9867 );
nand ( n9869 , n9866 , n9868 );
buf ( n9870 , n9869 );
buf ( n9871 , n9870 );
xor ( n9872 , n9863 , n9871 );
xor ( n9873 , n8974 , n8984 );
and ( n9874 , n9873 , n9002 );
and ( n9875 , n8974 , n8984 );
or ( n9876 , n9874 , n9875 );
buf ( n9877 , n9876 );
buf ( n9878 , n9877 );
xor ( n9879 , n9872 , n9878 );
buf ( n9880 , n9879 );
xor ( n9881 , n9846 , n9880 );
not ( n9882 , n8956 );
not ( n9883 , n8905 );
or ( n9884 , n9882 , n9883 );
not ( n9885 , n8906 );
not ( n9886 , n8953 );
or ( n9887 , n9885 , n9886 );
nand ( n9888 , n9887 , n9004 );
nand ( n9889 , n9884 , n9888 );
xnor ( n9890 , n9881 , n9889 );
buf ( n9891 , n9890 );
buf ( n9892 , n9891 );
buf ( n9893 , n9892 );
xor ( n9894 , n9794 , n9893 );
buf ( n9895 , n9894 );
buf ( n9896 , n9025 );
not ( n9897 , n9896 );
buf ( n9898 , n9042 );
not ( n9899 , n9898 );
or ( n9900 , n9897 , n9899 );
buf ( n9901 , n9042 );
buf ( n9902 , n9025 );
or ( n9903 , n9901 , n9902 );
buf ( n9904 , n9234 );
nand ( n9905 , n9903 , n9904 );
buf ( n9906 , n9905 );
buf ( n9907 , n9906 );
nand ( n9908 , n9900 , n9907 );
buf ( n9909 , n9908 );
buf ( n9910 , n9909 );
xor ( n9911 , n9895 , n9910 );
buf ( n9912 , n9007 );
not ( n9913 , n9912 );
buf ( n9914 , n8861 );
not ( n9915 , n9914 );
or ( n9916 , n9913 , n9915 );
buf ( n9917 , n8861 );
buf ( n9918 , n9007 );
or ( n9919 , n9917 , n9918 );
buf ( n9920 , n8856 );
nand ( n9921 , n9919 , n9920 );
buf ( n9922 , n9921 );
buf ( n9923 , n9922 );
nand ( n9924 , n9916 , n9923 );
buf ( n9925 , n9924 );
buf ( n9926 , n9925 );
xor ( n9927 , n9178 , n9184 );
and ( n9928 , n9927 , n9232 );
and ( n9929 , n9178 , n9184 );
or ( n9930 , n9928 , n9929 );
buf ( n9931 , n9930 );
buf ( n9932 , n9931 );
xor ( n9933 , n9926 , n9932 );
buf ( n9934 , n558 );
buf ( n9935 , n576 );
and ( n9936 , n9934 , n9935 );
buf ( n9937 , n9936 );
buf ( n9938 , n9937 );
buf ( n9939 , n1203 );
xor ( n9940 , n9938 , n9939 );
buf ( n9941 , n9129 );
not ( n9942 , n9941 );
buf ( n9943 , n8193 );
buf ( n9944 , n6699 );
nor ( n9945 , n9943 , n9944 );
buf ( n9946 , n9945 );
buf ( n9947 , n9946 );
not ( n9948 , n9947 );
or ( n9949 , n9942 , n9948 );
buf ( n9950 , n6699 );
buf ( n9951 , n9950 );
buf ( n9952 , n9951 );
buf ( n9953 , n9952 );
xor ( n9954 , n576 , n556 );
buf ( n9955 , n9954 );
nand ( n9956 , n9953 , n9955 );
buf ( n9957 , n9956 );
buf ( n9958 , n9957 );
nand ( n9959 , n9949 , n9958 );
buf ( n9960 , n9959 );
buf ( n9961 , n9960 );
xor ( n9962 , n9940 , n9961 );
buf ( n9963 , n9962 );
buf ( n9964 , n9963 );
buf ( n9965 , n9146 );
not ( n9966 , n9965 );
buf ( n9967 , n4205 );
not ( n9968 , n9967 );
or ( n9969 , n9966 , n9968 );
buf ( n9970 , n4211 );
xor ( n9971 , n582 , n550 );
buf ( n9972 , n9971 );
nand ( n9973 , n9970 , n9972 );
buf ( n9974 , n9973 );
buf ( n9975 , n9974 );
nand ( n9976 , n9969 , n9975 );
buf ( n9977 , n9976 );
buf ( n9978 , n9977 );
not ( n9979 , n9978 );
buf ( n9980 , n9979 );
buf ( n9981 , n9068 );
not ( n9982 , n9981 );
buf ( n9983 , n1177 );
not ( n9984 , n9983 );
or ( n9985 , n9982 , n9984 );
buf ( n9986 , n1036 );
buf ( n9987 , n546 );
buf ( n9988 , n586 );
xor ( n9989 , n9987 , n9988 );
buf ( n9990 , n9989 );
buf ( n9991 , n9990 );
nand ( n9992 , n9986 , n9991 );
buf ( n9993 , n9992 );
buf ( n9994 , n9993 );
nand ( n9995 , n9985 , n9994 );
buf ( n9996 , n9995 );
not ( n9997 , n9996 );
not ( n9998 , n9109 );
not ( n9999 , n1060 );
or ( n10000 , n9998 , n9999 );
buf ( n10001 , n544 );
buf ( n10002 , n588 );
xor ( n10003 , n10001 , n10002 );
buf ( n10004 , n10003 );
buf ( n10005 , n10004 );
buf ( n10006 , n1074 );
nand ( n10007 , n10005 , n10006 );
buf ( n10008 , n10007 );
nand ( n10009 , n10000 , n10008 );
not ( n10010 , n10009 );
not ( n10011 , n10010 );
or ( n10012 , n9997 , n10011 );
or ( n10013 , n10010 , n9996 );
nand ( n10014 , n10012 , n10013 );
xnor ( n10015 , n9980 , n10014 );
buf ( n10016 , n10015 );
xor ( n10017 , n9964 , n10016 );
xor ( n10018 , n9213 , n9218 );
and ( n10019 , n10018 , n9226 );
and ( n10020 , n9213 , n9218 );
or ( n10021 , n10019 , n10020 );
buf ( n10022 , n10021 );
buf ( n10023 , n10022 );
xor ( n10024 , n10017 , n10023 );
buf ( n10025 , n10024 );
buf ( n10026 , n10025 );
xor ( n10027 , n9191 , n9209 );
and ( n10028 , n10027 , n9229 );
and ( n10029 , n9191 , n9209 );
or ( n10030 , n10028 , n10029 );
buf ( n10031 , n10030 );
buf ( n10032 , n10031 );
xor ( n10033 , n10026 , n10032 );
buf ( n10034 , n9054 );
not ( n10035 , n10034 );
buf ( n10036 , n6350 );
not ( n10037 , n10036 );
or ( n10038 , n10035 , n10037 );
buf ( n10039 , n8294 );
xor ( n10040 , n578 , n554 );
buf ( n10041 , n10040 );
nand ( n10042 , n10039 , n10041 );
buf ( n10043 , n10042 );
buf ( n10044 , n10043 );
nand ( n10045 , n10038 , n10044 );
buf ( n10046 , n10045 );
buf ( n10047 , n10046 );
buf ( n10048 , n9078 );
not ( n10049 , n10048 );
buf ( n10050 , n5060 );
not ( n10051 , n10050 );
or ( n10052 , n10049 , n10051 );
buf ( n10053 , n5065 );
xor ( n10054 , n580 , n552 );
buf ( n10055 , n10054 );
nand ( n10056 , n10053 , n10055 );
buf ( n10057 , n10056 );
buf ( n10058 , n10057 );
nand ( n10059 , n10052 , n10058 );
buf ( n10060 , n10059 );
buf ( n10061 , n10060 );
xor ( n10062 , n10047 , n10061 );
buf ( n10063 , n9164 );
not ( n10064 , n10063 );
buf ( n10065 , n3664 );
not ( n10066 , n10065 );
or ( n10067 , n10064 , n10066 );
buf ( n10068 , n2123 );
xor ( n10069 , n584 , n548 );
buf ( n10070 , n10069 );
nand ( n10071 , n10068 , n10070 );
buf ( n10072 , n10071 );
buf ( n10073 , n10072 );
nand ( n10074 , n10067 , n10073 );
buf ( n10075 , n10074 );
buf ( n10076 , n10075 );
not ( n10077 , n10076 );
buf ( n10078 , n10077 );
buf ( n10079 , n10078 );
xor ( n10080 , n10062 , n10079 );
buf ( n10081 , n10080 );
buf ( n10082 , n10081 );
buf ( n10083 , n9117 );
not ( n10084 , n10083 );
buf ( n10085 , n9176 );
nand ( n10086 , n10084 , n10085 );
buf ( n10087 , n10086 );
buf ( n10088 , n10087 );
not ( n10089 , n9117 );
not ( n10090 , n9173 );
or ( n10091 , n10089 , n10090 );
nand ( n10092 , n10091 , n9083 );
buf ( n10093 , n10092 );
nand ( n10094 , n10088 , n10093 );
buf ( n10095 , n10094 );
buf ( n10096 , n10095 );
xor ( n10097 , n10082 , n10096 );
buf ( n10098 , n9116 );
not ( n10099 , n10098 );
buf ( n10100 , n9095 );
not ( n10101 , n10100 );
buf ( n10102 , n9099 );
nand ( n10103 , n10101 , n10102 );
buf ( n10104 , n10103 );
buf ( n10105 , n10104 );
not ( n10106 , n10105 );
or ( n10107 , n10099 , n10106 );
buf ( n10108 , n9099 );
not ( n10109 , n10108 );
buf ( n10110 , n9095 );
nand ( n10111 , n10109 , n10110 );
buf ( n10112 , n10111 );
buf ( n10113 , n10112 );
nand ( n10114 , n10107 , n10113 );
buf ( n10115 , n10114 );
buf ( n10116 , n10115 );
buf ( n10117 , n9060 );
buf ( n10118 , n9082 );
or ( n10119 , n10117 , n10118 );
buf ( n10120 , n9072 );
nand ( n10121 , n10119 , n10120 );
buf ( n10122 , n10121 );
buf ( n10123 , n10122 );
buf ( n10124 , n9060 );
buf ( n10125 , n9082 );
nand ( n10126 , n10124 , n10125 );
buf ( n10127 , n10126 );
buf ( n10128 , n10127 );
nand ( n10129 , n10123 , n10128 );
buf ( n10130 , n10129 );
buf ( n10131 , n10130 );
xor ( n10132 , n10116 , n10131 );
not ( n10133 , n9152 );
not ( n10134 , n9135 );
or ( n10135 , n10133 , n10134 );
buf ( n10136 , n9152 );
buf ( n10137 , n9135 );
nor ( n10138 , n10136 , n10137 );
buf ( n10139 , n10138 );
buf ( n10140 , n9170 );
not ( n10141 , n10140 );
buf ( n10142 , n10141 );
or ( n10143 , n10139 , n10142 );
nand ( n10144 , n10135 , n10143 );
buf ( n10145 , n10144 );
xor ( n10146 , n10132 , n10145 );
buf ( n10147 , n10146 );
buf ( n10148 , n10147 );
xor ( n10149 , n10097 , n10148 );
buf ( n10150 , n10149 );
buf ( n10151 , n10150 );
xor ( n10152 , n10033 , n10151 );
buf ( n10153 , n10152 );
buf ( n10154 , n10153 );
xor ( n10155 , n9933 , n10154 );
buf ( n10156 , n10155 );
buf ( n10157 , n10156 );
xor ( n10158 , n9911 , n10157 );
buf ( n10159 , n10158 );
not ( n10160 , n9235 );
not ( n10161 , n9015 );
nand ( n10162 , n10161 , n9009 );
not ( n10163 , n10162 );
or ( n10164 , n10160 , n10163 );
nand ( n10165 , n9008 , n9015 );
nand ( n10166 , n10164 , n10165 );
nor ( n10167 , n10159 , n10166 );
not ( n10168 , n10167 );
buf ( n10169 , n10159 );
buf ( n10170 , n10166 );
nand ( n10171 , n10169 , n10170 );
buf ( n10172 , n10171 );
nand ( n10173 , n10168 , n10172 );
xor ( n10174 , n9684 , n10173 );
not ( n10175 , n10174 );
nand ( n10176 , n9679 , n10175 );
nand ( n10177 , n9678 , n10174 );
and ( n10178 , n10176 , n10177 );
and ( n10179 , n9551 , n10178 );
not ( n10180 , n9551 );
not ( n10181 , n10178 );
and ( n10182 , n10180 , n10181 );
nor ( n10183 , n10179 , n10182 );
buf ( n10184 , n10183 );
nand ( n10185 , n10184 , n9497 );
not ( n10186 , n10185 );
nand ( n10187 , n9546 , n10186 );
nor ( n10188 , n9448 , n9452 );
nor ( n10189 , n9667 , n10188 );
not ( n10190 , n10189 );
not ( n10191 , n9466 );
or ( n10192 , n10190 , n10191 );
not ( n10193 , n9666 );
not ( n10194 , n9559 );
and ( n10195 , n10193 , n10194 );
nand ( n10196 , n9448 , n9452 );
nor ( n10197 , n10195 , n10196 );
nor ( n10198 , n10197 , n9671 );
nand ( n10199 , n10192 , n10198 );
not ( n10200 , n10199 );
xor ( n10201 , n9573 , n9584 );
and ( n10202 , n10201 , n9590 );
and ( n10203 , n9573 , n9584 );
or ( n10204 , n10202 , n10203 );
xor ( n10205 , n9596 , n9607 );
and ( n10206 , n10205 , n9612 );
and ( n10207 , n9596 , n9607 );
or ( n10208 , n10206 , n10207 );
xor ( n10209 , n10204 , n10208 );
not ( n10210 , n3109 );
not ( n10211 , n8439 );
not ( n10212 , n10211 );
not ( n10213 , n10212 );
or ( n10214 , n10210 , n10213 );
not ( n10215 , n556 );
not ( n10216 , n9378 );
or ( n10217 , n10215 , n10216 );
nand ( n10218 , n1625 , n9377 );
nand ( n10219 , n10217 , n10218 );
and ( n10220 , n10219 , n1594 );
and ( n10221 , n8440 , n3112 );
nor ( n10222 , n10220 , n10221 );
nand ( n10223 , n10214 , n10222 );
not ( n10224 , n5268 );
not ( n10225 , n9603 );
or ( n10226 , n10224 , n10225 );
and ( n10227 , n3264 , n550 );
not ( n10228 , n3264 );
and ( n10229 , n10228 , n3073 );
nor ( n10230 , n10227 , n10229 );
nand ( n10231 , n10230 , n3068 );
nand ( n10232 , n10226 , n10231 );
xor ( n10233 , n10223 , n10232 );
not ( n10234 , n2276 );
not ( n10235 , n9624 );
or ( n10236 , n10234 , n10235 );
xor ( n10237 , n554 , n7269 );
nand ( n10238 , n3118 , n10237 );
nand ( n10239 , n10236 , n10238 );
xor ( n10240 , n10233 , n10239 );
xor ( n10241 , n10209 , n10240 );
xor ( n10242 , n9650 , n9654 );
and ( n10243 , n10242 , n9659 );
and ( n10244 , n9650 , n9654 );
or ( n10245 , n10243 , n10244 );
xor ( n10246 , n10241 , n10245 );
xor ( n10247 , n9626 , n9644 );
and ( n10248 , n10247 , n9649 );
and ( n10249 , n9626 , n9644 );
or ( n10250 , n10248 , n10249 );
xor ( n10251 , n9636 , n9638 );
and ( n10252 , n10251 , n9643 );
and ( n10253 , n9636 , n9638 );
or ( n10254 , n10252 , n10253 );
not ( n10255 , n1740 );
nand ( n10256 , n10255 , n1774 );
not ( n10257 , n10256 );
not ( n10258 , n1652 );
nand ( n10259 , n10258 , n544 );
not ( n10260 , n10259 );
or ( n10261 , n10257 , n10260 );
or ( n10262 , n10259 , n10256 );
nand ( n10263 , n10261 , n10262 );
not ( n10264 , n9409 );
not ( n10265 , n2220 );
xor ( n10266 , n544 , n10265 );
not ( n10267 , n10266 );
or ( n10268 , n10264 , n10267 );
nand ( n10269 , n9632 , n9417 );
nand ( n10270 , n10268 , n10269 );
xor ( n10271 , n10263 , n10270 );
xor ( n10272 , n10254 , n10271 );
not ( n10273 , n6939 );
not ( n10274 , n9571 );
or ( n10275 , n10273 , n10274 );
not ( n10276 , n548 );
not ( n10277 , n3037 );
or ( n10278 , n10276 , n10277 );
nand ( n10279 , n3036 , n5279 );
nand ( n10280 , n10278 , n10279 );
nand ( n10281 , n10280 , n3212 );
nand ( n10282 , n10275 , n10281 );
not ( n10283 , n546 );
not ( n10284 , n3195 );
or ( n10285 , n10283 , n10284 );
nand ( n10286 , n2251 , n6949 );
nand ( n10287 , n10285 , n10286 );
not ( n10288 , n10287 );
not ( n10289 , n6945 );
or ( n10290 , n10288 , n10289 );
nand ( n10291 , n9582 , n9575 );
nand ( n10292 , n10290 , n10291 );
xor ( n10293 , n10282 , n10292 );
and ( n10294 , n552 , n7125 );
not ( n10295 , n552 );
and ( n10296 , n10295 , n7124 );
or ( n10297 , n10294 , n10296 );
not ( n10298 , n10297 );
not ( n10299 , n2265 );
or ( n10300 , n10298 , n10299 );
not ( n10301 , n9586 );
nand ( n10302 , n10301 , n3064 );
nand ( n10303 , n10300 , n10302 );
xor ( n10304 , n10293 , n10303 );
xor ( n10305 , n10272 , n10304 );
xor ( n10306 , n10250 , n10305 );
xor ( n10307 , n9563 , n9591 );
and ( n10308 , n10307 , n9613 );
and ( n10309 , n9563 , n9591 );
or ( n10310 , n10308 , n10309 );
xor ( n10311 , n10306 , n10310 );
xor ( n10312 , n10246 , n10311 );
xor ( n10313 , n9614 , n9660 );
and ( n10314 , n10313 , n9665 );
and ( n10315 , n9614 , n9660 );
or ( n10316 , n10314 , n10315 );
nor ( n10317 , n10312 , n10316 );
not ( n10318 , n10317 );
nand ( n10319 , n10312 , n10316 );
buf ( n10320 , n10319 );
nand ( n10321 , n10318 , n10320 );
and ( n10322 , n10200 , n10321 );
not ( n10323 , n10200 );
not ( n10324 , n10321 );
and ( n10325 , n10323 , n10324 );
nor ( n10326 , n10322 , n10325 );
not ( n10327 , n10326 );
nor ( n10328 , n10167 , n9246 );
not ( n10329 , n10328 );
not ( n10330 , n9681 );
or ( n10331 , n10329 , n10330 );
or ( n10332 , n9248 , n10167 );
nand ( n10333 , n10332 , n10172 );
buf ( n10334 , n10333 );
not ( n10335 , n10334 );
buf ( n10336 , n10335 );
nand ( n10337 , n10331 , n10336 );
buf ( n10338 , n557 );
buf ( n10339 , n560 );
and ( n10340 , n10338 , n10339 );
buf ( n10341 , n10340 );
buf ( n10342 , n10341 );
buf ( n10343 , n9753 );
not ( n10344 , n10343 );
buf ( n10345 , n4044 );
not ( n10346 , n10345 );
or ( n10347 , n10344 , n10346 );
buf ( n10348 , n3743 );
xor ( n10349 , n566 , n549 );
buf ( n10350 , n10349 );
nand ( n10351 , n10348 , n10350 );
buf ( n10352 , n10351 );
buf ( n10353 , n10352 );
nand ( n10354 , n10347 , n10353 );
buf ( n10355 , n10354 );
buf ( n10356 , n10355 );
xor ( n10357 , n10342 , n10356 );
buf ( n10358 , n9739 );
not ( n10359 , n10358 );
buf ( n10360 , n850 );
not ( n10361 , n10360 );
or ( n10362 , n10359 , n10361 );
buf ( n10363 , n856 );
buf ( n10364 , n545 );
buf ( n10365 , n570 );
xor ( n10366 , n10364 , n10365 );
buf ( n10367 , n10366 );
buf ( n10368 , n10367 );
nand ( n10369 , n10363 , n10368 );
buf ( n10370 , n10369 );
buf ( n10371 , n10370 );
nand ( n10372 , n10362 , n10371 );
buf ( n10373 , n10372 );
buf ( n10374 , n10373 );
xor ( n10375 , n10357 , n10374 );
buf ( n10376 , n10375 );
buf ( n10377 , n10376 );
buf ( n10378 , n9701 );
not ( n10379 , n10378 );
buf ( n10380 , n7964 );
buf ( n10381 , n10380 );
not ( n10382 , n10381 );
or ( n10383 , n10379 , n10382 );
buf ( n10384 , n6595 );
buf ( n10385 , n555 );
buf ( n10386 , n560 );
xor ( n10387 , n10385 , n10386 );
buf ( n10388 , n10387 );
buf ( n10389 , n10388 );
nand ( n10390 , n10384 , n10389 );
buf ( n10391 , n10390 );
buf ( n10392 , n10391 );
nand ( n10393 , n10383 , n10392 );
buf ( n10394 , n10393 );
buf ( n10395 , n10394 );
buf ( n10396 , n9845 );
xor ( n10397 , n10395 , n10396 );
buf ( n10398 , n9723 );
not ( n10399 , n10398 );
buf ( n10400 , n884 );
not ( n10401 , n10400 );
or ( n10402 , n10399 , n10401 );
buf ( n10403 , n572 );
buf ( n10404 , n888 );
nand ( n10405 , n10403 , n10404 );
buf ( n10406 , n10405 );
buf ( n10407 , n10406 );
nand ( n10408 , n10402 , n10407 );
buf ( n10409 , n10408 );
buf ( n10410 , n10409 );
not ( n10411 , n10410 );
buf ( n10412 , n10411 );
buf ( n10413 , n10412 );
xor ( n10414 , n10397 , n10413 );
buf ( n10415 , n10414 );
buf ( n10416 , n10415 );
xor ( n10417 , n10377 , n10416 );
xor ( n10418 , n9863 , n9871 );
and ( n10419 , n10418 , n9878 );
and ( n10420 , n9863 , n9871 );
or ( n10421 , n10419 , n10420 );
buf ( n10422 , n10421 );
buf ( n10423 , n10422 );
xor ( n10424 , n10417 , n10423 );
buf ( n10425 , n10424 );
buf ( n10426 , n10425 );
buf ( n10427 , n9846 );
not ( n10428 , n10427 );
buf ( n10429 , n9880 );
not ( n10430 , n10429 );
buf ( n10431 , n10430 );
buf ( n10432 , n10431 );
not ( n10433 , n10432 );
or ( n10434 , n10428 , n10433 );
buf ( n10435 , n9889 );
nand ( n10436 , n10434 , n10435 );
buf ( n10437 , n10436 );
buf ( n10438 , n10437 );
buf ( n10439 , n9846 );
not ( n10440 , n10439 );
buf ( n10441 , n9880 );
nand ( n10442 , n10440 , n10441 );
buf ( n10443 , n10442 );
buf ( n10444 , n10443 );
nand ( n10445 , n10438 , n10444 );
buf ( n10446 , n10445 );
buf ( n10447 , n10446 );
xor ( n10448 , n10426 , n10447 );
buf ( n10449 , n9828 );
buf ( n10450 , n9812 );
nor ( n10451 , n10449 , n10450 );
buf ( n10452 , n10451 );
buf ( n10453 , n10452 );
buf ( n10454 , n9845 );
or ( n10455 , n10453 , n10454 );
buf ( n10456 , n9828 );
buf ( n10457 , n9812 );
nand ( n10458 , n10456 , n10457 );
buf ( n10459 , n10458 );
buf ( n10460 , n10459 );
nand ( n10461 , n10455 , n10460 );
buf ( n10462 , n10461 );
buf ( n10463 , n10462 );
buf ( n10464 , n9694 );
buf ( n10465 , n574 );
nand ( n10466 , n10464 , n10465 );
buf ( n10467 , n10466 );
not ( n10468 , n10467 );
not ( n10469 , n9705 );
or ( n10470 , n10468 , n10469 );
or ( n10471 , n9694 , n574 );
nand ( n10472 , n10470 , n10471 );
buf ( n10473 , n10472 );
buf ( n10474 , n9745 );
not ( n10475 , n10474 );
buf ( n10476 , n9729 );
not ( n10477 , n10476 );
or ( n10478 , n10475 , n10477 );
or ( n10479 , n9745 , n9729 );
nand ( n10480 , n10479 , n9759 );
buf ( n10481 , n10480 );
nand ( n10482 , n10478 , n10481 );
buf ( n10483 , n10482 );
buf ( n10484 , n10483 );
xor ( n10485 , n10473 , n10484 );
buf ( n10486 , n9822 );
not ( n10487 , n10486 );
buf ( n10488 , n5678 );
not ( n10489 , n10488 );
or ( n10490 , n10487 , n10489 );
xor ( n10491 , n551 , n564 );
nand ( n10492 , n4840 , n10491 );
buf ( n10493 , n10492 );
nand ( n10494 , n10490 , n10493 );
buf ( n10495 , n10494 );
buf ( n10496 , n10495 );
buf ( n10497 , n9806 );
not ( n10498 , n10497 );
buf ( n10499 , n9797 );
not ( n10500 , n10499 );
or ( n10501 , n10498 , n10500 );
buf ( n10502 , n5801 );
buf ( n10503 , n553 );
buf ( n10504 , n562 );
xor ( n10505 , n10503 , n10504 );
buf ( n10506 , n10505 );
buf ( n10507 , n10506 );
nand ( n10508 , n10502 , n10507 );
buf ( n10509 , n10508 );
buf ( n10510 , n10509 );
nand ( n10511 , n10501 , n10510 );
buf ( n10512 , n10511 );
buf ( n10513 , n10512 );
xor ( n10514 , n10496 , n10513 );
buf ( n10515 , n9839 );
not ( n10516 , n10515 );
buf ( n10517 , n3429 );
not ( n10518 , n10517 );
or ( n10519 , n10516 , n10518 );
buf ( n10520 , n3772 );
buf ( n10521 , n547 );
buf ( n10522 , n568 );
xor ( n10523 , n10521 , n10522 );
buf ( n10524 , n10523 );
buf ( n10525 , n10524 );
nand ( n10526 , n10520 , n10525 );
buf ( n10527 , n10526 );
buf ( n10528 , n10527 );
nand ( n10529 , n10519 , n10528 );
buf ( n10530 , n10529 );
buf ( n10531 , n10530 );
xor ( n10532 , n10514 , n10531 );
buf ( n10533 , n10532 );
buf ( n10534 , n10533 );
xor ( n10535 , n10485 , n10534 );
buf ( n10536 , n10535 );
buf ( n10537 , n10536 );
xor ( n10538 , n10463 , n10537 );
or ( n10539 , n9777 , n9711 );
nand ( n10540 , n10539 , n9768 );
buf ( n10541 , n10540 );
buf ( n10542 , n9777 );
buf ( n10543 , n9711 );
nand ( n10544 , n10542 , n10543 );
buf ( n10545 , n10544 );
buf ( n10546 , n10545 );
nand ( n10547 , n10541 , n10546 );
buf ( n10548 , n10547 );
buf ( n10549 , n10548 );
xor ( n10550 , n10538 , n10549 );
buf ( n10551 , n10550 );
buf ( n10552 , n10551 );
xor ( n10553 , n10448 , n10552 );
buf ( n10554 , n10553 );
buf ( n10555 , n10554 );
xor ( n10556 , n9926 , n9932 );
and ( n10557 , n10556 , n10154 );
and ( n10558 , n9926 , n9932 );
or ( n10559 , n10557 , n10558 );
buf ( n10560 , n10559 );
buf ( n10561 , n10560 );
xor ( n10562 , n10555 , n10561 );
not ( n10563 , n9890 );
buf ( n10564 , n9689 );
not ( n10565 , n10564 );
buf ( n10566 , n10565 );
nand ( n10567 , n10566 , n9787 );
not ( n10568 , n10567 );
or ( n10569 , n10563 , n10568 );
nand ( n10570 , n9792 , n9689 );
nand ( n10571 , n10569 , n10570 );
buf ( n10572 , n10571 );
xor ( n10573 , n10026 , n10032 );
and ( n10574 , n10573 , n10151 );
and ( n10575 , n10026 , n10032 );
or ( n10576 , n10574 , n10575 );
buf ( n10577 , n10576 );
buf ( n10578 , n10577 );
xor ( n10579 , n10572 , n10578 );
buf ( n10580 , n9990 );
not ( n10581 , n10580 );
buf ( n10582 , n1177 );
not ( n10583 , n10582 );
or ( n10584 , n10581 , n10583 );
buf ( n10585 , n1036 );
buf ( n10586 , n545 );
buf ( n10587 , n586 );
xor ( n10588 , n10586 , n10587 );
buf ( n10589 , n10588 );
buf ( n10590 , n10589 );
nand ( n10591 , n10585 , n10590 );
buf ( n10592 , n10591 );
buf ( n10593 , n10592 );
nand ( n10594 , n10584 , n10593 );
buf ( n10595 , n10594 );
buf ( n10596 , n10595 );
buf ( n10597 , n557 );
buf ( n10598 , n576 );
nand ( n10599 , n10597 , n10598 );
buf ( n10600 , n10599 );
buf ( n10601 , n10600 );
not ( n10602 , n10601 );
buf ( n10603 , n10602 );
buf ( n10604 , n10603 );
and ( n10605 , n10596 , n10604 );
not ( n10606 , n10596 );
buf ( n10607 , n10600 );
and ( n10608 , n10606 , n10607 );
nor ( n10609 , n10605 , n10608 );
buf ( n10610 , n10609 );
buf ( n10611 , n9971 );
not ( n10612 , n10611 );
buf ( n10613 , n4205 );
not ( n10614 , n10613 );
or ( n10615 , n10612 , n10614 );
buf ( n10616 , n3883 );
xor ( n10617 , n582 , n549 );
buf ( n10618 , n10617 );
nand ( n10619 , n10616 , n10618 );
buf ( n10620 , n10619 );
buf ( n10621 , n10620 );
nand ( n10622 , n10615 , n10621 );
buf ( n10623 , n10622 );
xor ( n10624 , n10610 , n10623 );
buf ( n10625 , n10624 );
buf ( n10626 , n9954 );
not ( n10627 , n10626 );
buf ( n10628 , n9946 );
not ( n10629 , n10628 );
or ( n10630 , n10627 , n10629 );
buf ( n10631 , n9952 );
buf ( n10632 , n555 );
buf ( n10633 , n576 );
xor ( n10634 , n10632 , n10633 );
buf ( n10635 , n10634 );
buf ( n10636 , n10635 );
nand ( n10637 , n10631 , n10636 );
buf ( n10638 , n10637 );
buf ( n10639 , n10638 );
nand ( n10640 , n10630 , n10639 );
buf ( n10641 , n10640 );
buf ( n10642 , n10641 );
buf ( n10643 , n10004 );
not ( n10644 , n10643 );
buf ( n10645 , n1060 );
not ( n10646 , n10645 );
or ( n10647 , n10644 , n10646 );
buf ( n10648 , n588 );
buf ( n10649 , n1074 );
nand ( n10650 , n10648 , n10649 );
buf ( n10651 , n10650 );
buf ( n10652 , n10651 );
nand ( n10653 , n10647 , n10652 );
buf ( n10654 , n10653 );
buf ( n10655 , n10654 );
not ( n10656 , n10655 );
buf ( n10657 , n10656 );
buf ( n10658 , n10657 );
xor ( n10659 , n10642 , n10658 );
buf ( n10660 , n10075 );
xor ( n10661 , n10659 , n10660 );
buf ( n10662 , n10661 );
buf ( n10663 , n10662 );
xor ( n10664 , n10625 , n10663 );
xor ( n10665 , n10116 , n10131 );
and ( n10666 , n10665 , n10145 );
and ( n10667 , n10116 , n10131 );
or ( n10668 , n10666 , n10667 );
buf ( n10669 , n10668 );
buf ( n10670 , n10669 );
xor ( n10671 , n10664 , n10670 );
buf ( n10672 , n10671 );
buf ( n10673 , n10672 );
xor ( n10674 , n10082 , n10096 );
and ( n10675 , n10674 , n10148 );
and ( n10676 , n10082 , n10096 );
or ( n10677 , n10675 , n10676 );
buf ( n10678 , n10677 );
buf ( n10679 , n10678 );
xor ( n10680 , n10673 , n10679 );
xor ( n10681 , n10047 , n10061 );
and ( n10682 , n10681 , n10079 );
and ( n10683 , n10047 , n10061 );
or ( n10684 , n10682 , n10683 );
buf ( n10685 , n10684 );
buf ( n10686 , n10685 );
xor ( n10687 , n9938 , n9939 );
and ( n10688 , n10687 , n9961 );
and ( n10689 , n9938 , n9939 );
or ( n10690 , n10688 , n10689 );
buf ( n10691 , n10690 );
buf ( n10692 , n10691 );
buf ( n10693 , n9977 );
not ( n10694 , n10693 );
buf ( n10695 , n10009 );
not ( n10696 , n10695 );
or ( n10697 , n10694 , n10696 );
buf ( n10698 , n9980 );
not ( n10699 , n10698 );
buf ( n10700 , n10010 );
not ( n10701 , n10700 );
or ( n10702 , n10699 , n10701 );
buf ( n10703 , n9996 );
nand ( n10704 , n10702 , n10703 );
buf ( n10705 , n10704 );
buf ( n10706 , n10705 );
nand ( n10707 , n10697 , n10706 );
buf ( n10708 , n10707 );
buf ( n10709 , n10708 );
xor ( n10710 , n10692 , n10709 );
buf ( n10711 , n551 );
buf ( n10712 , n580 );
xor ( n10713 , n10711 , n10712 );
buf ( n10714 , n10713 );
not ( n10715 , n10714 );
not ( n10716 , n4544 );
or ( n10717 , n10715 , n10716 );
nand ( n10718 , n5058 , n4541 , n10054 );
nand ( n10719 , n10717 , n10718 );
buf ( n10720 , n10719 );
buf ( n10721 , n10040 );
not ( n10722 , n10721 );
buf ( n10723 , n6350 );
not ( n10724 , n10723 );
or ( n10725 , n10722 , n10724 );
buf ( n10726 , n5997 );
buf ( n10727 , n553 );
buf ( n10728 , n578 );
xor ( n10729 , n10727 , n10728 );
buf ( n10730 , n10729 );
buf ( n10731 , n10730 );
nand ( n10732 , n10726 , n10731 );
buf ( n10733 , n10732 );
buf ( n10734 , n10733 );
nand ( n10735 , n10725 , n10734 );
buf ( n10736 , n10735 );
buf ( n10737 , n10736 );
xor ( n10738 , n10720 , n10737 );
buf ( n10739 , n10069 );
not ( n10740 , n10739 );
buf ( n10741 , n3664 );
not ( n10742 , n10741 );
or ( n10743 , n10740 , n10742 );
buf ( n10744 , n2135 );
xor ( n10745 , n584 , n547 );
buf ( n10746 , n10745 );
nand ( n10747 , n10744 , n10746 );
buf ( n10748 , n10747 );
buf ( n10749 , n10748 );
nand ( n10750 , n10743 , n10749 );
buf ( n10751 , n10750 );
buf ( n10752 , n10751 );
xor ( n10753 , n10738 , n10752 );
buf ( n10754 , n10753 );
buf ( n10755 , n10754 );
xor ( n10756 , n10710 , n10755 );
buf ( n10757 , n10756 );
buf ( n10758 , n10757 );
xor ( n10759 , n10686 , n10758 );
xor ( n10760 , n9964 , n10016 );
and ( n10761 , n10760 , n10023 );
and ( n10762 , n9964 , n10016 );
or ( n10763 , n10761 , n10762 );
buf ( n10764 , n10763 );
buf ( n10765 , n10764 );
xor ( n10766 , n10759 , n10765 );
buf ( n10767 , n10766 );
buf ( n10768 , n10767 );
xor ( n10769 , n10680 , n10768 );
buf ( n10770 , n10769 );
buf ( n10771 , n10770 );
xor ( n10772 , n10579 , n10771 );
buf ( n10773 , n10772 );
buf ( n10774 , n10773 );
xor ( n10775 , n10562 , n10774 );
buf ( n10776 , n10775 );
xor ( n10777 , n9895 , n9910 );
and ( n10778 , n10777 , n10157 );
and ( n10779 , n9895 , n9910 );
or ( n10780 , n10778 , n10779 );
buf ( n10781 , n10780 );
or ( n10782 , n10776 , n10781 );
buf ( n10783 , n10776 );
buf ( n10784 , n10781 );
nand ( n10785 , n10783 , n10784 );
buf ( n10786 , n10785 );
nand ( n10787 , n10782 , n10786 );
and ( n10788 , n10337 , n10787 );
not ( n10789 , n10337 );
not ( n10790 , n10787 );
and ( n10791 , n10789 , n10790 );
nor ( n10792 , n10788 , n10791 );
not ( n10793 , n10792 );
nand ( n10794 , n10327 , n10793 );
not ( n10795 , n10794 );
not ( n10796 , n10326 );
nor ( n10797 , n10796 , n10793 );
or ( n10798 , n10795 , n10797 );
not ( n10799 , n10798 );
not ( n10800 , n9678 );
not ( n10801 , n10174 );
or ( n10802 , n10800 , n10801 );
nand ( n10803 , n10802 , n9477 );
not ( n10804 , n10803 );
nand ( n10805 , n10804 , n9548 );
not ( n10806 , n9473 );
not ( n10807 , n10806 );
not ( n10808 , n10177 );
or ( n10809 , n10807 , n10808 );
nand ( n10810 , n10809 , n10176 );
buf ( n10811 , n10810 );
not ( n10812 , n10811 );
nand ( n10813 , n10805 , n10812 );
not ( n10814 , n10813 );
or ( n10815 , n10799 , n10814 );
nor ( n10816 , n10798 , n10811 );
nand ( n10817 , n10805 , n10816 );
nand ( n10818 , n10815 , n10817 );
buf ( n10819 , n10818 );
buf ( n10820 , n10819 );
buf ( n10821 , n10820 );
buf ( n10822 , n10821 );
buf ( n10823 , n10822 );
not ( n10824 , n10823 );
and ( n10825 , n10187 , n10824 );
not ( n10826 , n10187 );
and ( n10827 , n10826 , n10823 );
nor ( n10828 , n10825 , n10827 );
buf ( n10829 , n10828 );
buf ( n10830 , n10829 );
not ( n10831 , n10830 );
buf ( n10832 , n10831 );
not ( n10833 , n10832 );
or ( n10834 , n9545 , n10833 );
buf ( n10835 , n10829 );
not ( n10836 , n606 );
buf ( n10837 , n10836 );
nand ( n10838 , n10835 , n10837 );
buf ( n10839 , n10838 );
buf ( n10840 , n10839 );
nand ( n10841 , n10834 , n10840 );
buf ( n10842 , n10841 );
buf ( n10843 , n10842 );
not ( n10844 , n10843 );
or ( n10845 , n9543 , n10844 );
buf ( n10846 , n606 );
not ( n10847 , n10846 );
not ( n10848 , n9505 );
not ( n10849 , n9515 );
or ( n10850 , n10848 , n10849 );
nand ( n10851 , n10850 , n9497 );
buf ( n10852 , n10184 );
buf ( n10853 , n10852 );
buf ( n10854 , n10853 );
or ( n10855 , n10851 , n10854 );
nand ( n10856 , n10854 , n10851 );
nand ( n10857 , n10855 , n10856 );
buf ( n10858 , n10857 );
buf ( n10859 , n10858 );
not ( n10860 , n10859 );
buf ( n10861 , n10860 );
buf ( n10862 , n10861 );
not ( n10863 , n10862 );
or ( n10864 , n10847 , n10863 );
buf ( n10865 , n10858 );
buf ( n10866 , n10836 );
nand ( n10867 , n10865 , n10866 );
buf ( n10868 , n10867 );
buf ( n10869 , n10868 );
nand ( n10870 , n10864 , n10869 );
buf ( n10871 , n10870 );
buf ( n10872 , n10871 );
buf ( n10873 , n10836 );
buf ( n10874 , n607 );
nor ( n10875 , n10873 , n10874 );
buf ( n10876 , n10875 );
buf ( n10877 , n10876 );
buf ( n10878 , n10877 );
buf ( n10879 , n10878 );
buf ( n10880 , n10879 );
buf ( n10881 , n10880 );
buf ( n10882 , n10881 );
buf ( n10883 , n10882 );
nand ( n10884 , n10872 , n10883 );
buf ( n10885 , n10884 );
buf ( n10886 , n10885 );
nand ( n10887 , n10845 , n10886 );
buf ( n10888 , n10887 );
buf ( n10889 , n10888 );
xor ( n10890 , n9541 , n10889 );
buf ( n10891 , n10890 );
buf ( n10892 , n10891 );
xor ( n10893 , n8791 , n10892 );
buf ( n10894 , n10893 );
buf ( n10895 , n10894 );
not ( n10896 , n10895 );
buf ( n10897 , n607 );
not ( n10898 , n10897 );
buf ( n10899 , n10871 );
not ( n10900 , n10899 );
or ( n10901 , n10898 , n10900 );
not ( n10902 , n9527 );
and ( n10903 , n10902 , n10836 );
not ( n10904 , n10902 );
and ( n10905 , n10904 , n606 );
nor ( n10906 , n10903 , n10905 );
buf ( n10907 , n10906 );
buf ( n10908 , n10882 );
nand ( n10909 , n10907 , n10908 );
buf ( n10910 , n10909 );
buf ( n10911 , n10910 );
nand ( n10912 , n10901 , n10911 );
buf ( n10913 , n10912 );
buf ( n10914 , n10913 );
buf ( n10915 , n5549 );
not ( n10916 , n10915 );
buf ( n10917 , n8621 );
not ( n10918 , n10917 );
or ( n10919 , n10916 , n10918 );
buf ( n10920 , n5631 );
buf ( n10921 , n598 );
not ( n10922 , n10921 );
buf ( n10923 , n5487 );
not ( n10924 , n10923 );
or ( n10925 , n10922 , n10924 );
buf ( n10926 , n2390 );
buf ( n10927 , n818 );
nand ( n10928 , n10926 , n10927 );
buf ( n10929 , n10928 );
buf ( n10930 , n10929 );
nand ( n10931 , n10925 , n10930 );
buf ( n10932 , n10931 );
buf ( n10933 , n10932 );
nand ( n10934 , n10920 , n10933 );
buf ( n10935 , n10934 );
buf ( n10936 , n10935 );
nand ( n10937 , n10919 , n10936 );
buf ( n10938 , n10937 );
buf ( n10939 , n10938 );
xor ( n10940 , n2763 , n2788 );
xor ( n10941 , n10940 , n2892 );
buf ( n10942 , n10941 );
buf ( n10943 , n10942 );
xor ( n10944 , n10939 , n10943 );
buf ( n10945 , n2914 );
buf ( n10946 , n10945 );
not ( n10947 , n10946 );
buf ( n10948 , n8664 );
not ( n10949 , n10948 );
or ( n10950 , n10947 , n10949 );
and ( n10951 , n5458 , n600 );
not ( n10952 , n5458 );
and ( n10953 , n10952 , n5382 );
or ( n10954 , n10951 , n10953 );
buf ( n10955 , n10954 );
buf ( n10956 , n5430 );
nand ( n10957 , n10955 , n10956 );
buf ( n10958 , n10957 );
buf ( n10959 , n10958 );
nand ( n10960 , n10950 , n10959 );
buf ( n10961 , n10960 );
buf ( n10962 , n10961 );
and ( n10963 , n10944 , n10962 );
and ( n10964 , n10939 , n10943 );
or ( n10965 , n10963 , n10964 );
buf ( n10966 , n10965 );
buf ( n10967 , n10966 );
not ( n10968 , n5655 );
not ( n10969 , n8709 );
or ( n10970 , n10968 , n10969 );
buf ( n10971 , n602 );
not ( n10972 , n10971 );
buf ( n10973 , n5407 );
not ( n10974 , n10973 );
or ( n10975 , n10972 , n10974 );
buf ( n10976 , n5411 );
buf ( n10977 , n2912 );
nand ( n10978 , n10976 , n10977 );
buf ( n10979 , n10978 );
buf ( n10980 , n10979 );
nand ( n10981 , n10975 , n10980 );
buf ( n10982 , n10981 );
buf ( n10983 , n10982 );
buf ( n10984 , n7619 );
nand ( n10985 , n10983 , n10984 );
buf ( n10986 , n10985 );
nand ( n10987 , n10970 , n10986 );
buf ( n10988 , n10987 );
xor ( n10989 , n10967 , n10988 );
xor ( n10990 , n8629 , n8633 );
xor ( n10991 , n10990 , n8672 );
buf ( n10992 , n10991 );
buf ( n10993 , n10992 );
and ( n10994 , n10989 , n10993 );
and ( n10995 , n10967 , n10988 );
or ( n10996 , n10994 , n10995 );
buf ( n10997 , n10996 );
buf ( n10998 , n10997 );
buf ( n10999 , n7789 );
not ( n11000 , n10999 );
buf ( n11001 , n8566 );
not ( n11002 , n11001 );
or ( n11003 , n11000 , n11002 );
not ( n11004 , n7589 );
not ( n11005 , n7586 );
or ( n11006 , n11004 , n11005 );
nand ( n11007 , n7585 , n7588 );
nand ( n11008 , n11006 , n11007 );
buf ( n11009 , n11008 );
not ( n11010 , n11009 );
buf ( n11011 , n11010 );
and ( n11012 , n604 , n11011 );
not ( n11013 , n604 );
and ( n11014 , n11013 , n11008 );
or ( n11015 , n11012 , n11014 );
buf ( n11016 , n11015 );
buf ( n11017 , n8581 );
nand ( n11018 , n11016 , n11017 );
buf ( n11019 , n11018 );
buf ( n11020 , n11019 );
nand ( n11021 , n11003 , n11020 );
buf ( n11022 , n11021 );
buf ( n11023 , n11022 );
xor ( n11024 , n10998 , n11023 );
xor ( n11025 , n8677 , n8717 );
xor ( n11026 , n11025 , n8752 );
buf ( n11027 , n11026 );
buf ( n11028 , n11027 );
and ( n11029 , n11024 , n11028 );
and ( n11030 , n10998 , n11023 );
or ( n11031 , n11029 , n11030 );
buf ( n11032 , n11031 );
buf ( n11033 , n11032 );
xor ( n11034 , n10914 , n11033 );
xor ( n11035 , n8588 , n8757 );
xor ( n11036 , n11035 , n8785 );
buf ( n11037 , n11036 );
buf ( n11038 , n11037 );
and ( n11039 , n11034 , n11038 );
and ( n11040 , n10914 , n11033 );
or ( n11041 , n11039 , n11040 );
buf ( n11042 , n11041 );
buf ( n11043 , n11042 );
not ( n11044 , n11043 );
buf ( n11045 , n11044 );
buf ( n11046 , n11045 );
nand ( n11047 , n10896 , n11046 );
buf ( n11048 , n11047 );
not ( n11049 , n11048 );
buf ( n11050 , n607 );
not ( n11051 , n11050 );
buf ( n11052 , n606 );
not ( n11053 , n11052 );
buf ( n11054 , n8554 );
not ( n11055 , n11054 );
or ( n11056 , n11053 , n11055 );
buf ( n11057 , n8557 );
buf ( n11058 , n10836 );
nand ( n11059 , n11057 , n11058 );
buf ( n11060 , n11059 );
buf ( n11061 , n11060 );
nand ( n11062 , n11056 , n11061 );
buf ( n11063 , n11062 );
buf ( n11064 , n11063 );
not ( n11065 , n11064 );
or ( n11066 , n11051 , n11065 );
buf ( n11067 , n606 );
not ( n11068 , n11067 );
buf ( n11069 , n7562 );
not ( n11070 , n11069 );
or ( n11071 , n11068 , n11070 );
buf ( n11072 , n7559 );
buf ( n11073 , n10836 );
nand ( n11074 , n11072 , n11073 );
buf ( n11075 , n11074 );
buf ( n11076 , n11075 );
nand ( n11077 , n11071 , n11076 );
buf ( n11078 , n11077 );
buf ( n11079 , n11078 );
buf ( n11080 , n10882 );
nand ( n11081 , n11079 , n11080 );
buf ( n11082 , n11081 );
buf ( n11083 , n11082 );
nand ( n11084 , n11066 , n11083 );
buf ( n11085 , n11084 );
buf ( n11086 , n11085 );
buf ( n11087 , n10945 );
not ( n11088 , n11087 );
buf ( n11089 , n10954 );
not ( n11090 , n11089 );
or ( n11091 , n11088 , n11090 );
buf ( n11092 , n600 );
not ( n11093 , n11092 );
buf ( n11094 , n2358 );
not ( n11095 , n11094 );
buf ( n11096 , n11095 );
buf ( n11097 , n11096 );
not ( n11098 , n11097 );
or ( n11099 , n11093 , n11098 );
buf ( n11100 , n11096 );
not ( n11101 , n11100 );
buf ( n11102 , n11101 );
buf ( n11103 , n11102 );
buf ( n11104 , n5382 );
nand ( n11105 , n11103 , n11104 );
buf ( n11106 , n11105 );
buf ( n11107 , n11106 );
nand ( n11108 , n11099 , n11107 );
buf ( n11109 , n11108 );
buf ( n11110 , n11109 );
buf ( n11111 , n5430 );
nand ( n11112 , n11110 , n11111 );
buf ( n11113 , n11112 );
buf ( n11114 , n11113 );
nand ( n11115 , n11091 , n11114 );
buf ( n11116 , n11115 );
buf ( n11117 , n11116 );
buf ( n11118 , n5549 );
not ( n11119 , n11118 );
buf ( n11120 , n10932 );
not ( n11121 , n11120 );
or ( n11122 , n11119 , n11121 );
buf ( n11123 , n598 );
not ( n11124 , n11123 );
buf ( n11125 , n2738 );
not ( n11126 , n11125 );
or ( n11127 , n11124 , n11126 );
buf ( n11128 , n7719 );
buf ( n11129 , n818 );
nand ( n11130 , n11128 , n11129 );
buf ( n11131 , n11130 );
buf ( n11132 , n11131 );
nand ( n11133 , n11127 , n11132 );
buf ( n11134 , n11133 );
buf ( n11135 , n11134 );
buf ( n11136 , n5631 );
nand ( n11137 , n11135 , n11136 );
buf ( n11138 , n11137 );
buf ( n11139 , n11138 );
nand ( n11140 , n11122 , n11139 );
buf ( n11141 , n11140 );
buf ( n11142 , n11141 );
xor ( n11143 , n2800 , n2825 );
xor ( n11144 , n11143 , n2887 );
buf ( n11145 , n11144 );
buf ( n11146 , n11145 );
xor ( n11147 , n11142 , n11146 );
xor ( n11148 , n2831 , n2869 );
xor ( n11149 , n11148 , n2883 );
buf ( n11150 , n11149 );
buf ( n11151 , n11150 );
buf ( n11152 , n5549 );
not ( n11153 , n11152 );
buf ( n11154 , n11134 );
not ( n11155 , n11154 );
or ( n11156 , n11153 , n11155 );
buf ( n11157 , n598 );
not ( n11158 , n11157 );
buf ( n11159 , n2576 );
not ( n11160 , n11159 );
or ( n11161 , n11158 , n11160 );
buf ( n11162 , n818 );
buf ( n11163 , n2570 );
nand ( n11164 , n11162 , n11163 );
buf ( n11165 , n11164 );
buf ( n11166 , n11165 );
nand ( n11167 , n11161 , n11166 );
buf ( n11168 , n11167 );
buf ( n11169 , n11168 );
buf ( n11170 , n5630 );
nand ( n11171 , n11169 , n11170 );
buf ( n11172 , n11171 );
buf ( n11173 , n11172 );
nand ( n11174 , n11156 , n11173 );
buf ( n11175 , n11174 );
buf ( n11176 , n11175 );
xor ( n11177 , n11151 , n11176 );
buf ( n11178 , n2865 );
not ( n11179 , n11178 );
buf ( n11180 , n2848 );
not ( n11181 , n11180 );
or ( n11182 , n11179 , n11181 );
buf ( n11183 , n2848 );
buf ( n11184 , n2865 );
or ( n11185 , n11183 , n11184 );
nand ( n11186 , n11182 , n11185 );
buf ( n11187 , n11186 );
buf ( n11188 , n11187 );
buf ( n11189 , n5549 );
not ( n11190 , n11189 );
buf ( n11191 , n11168 );
not ( n11192 , n11191 );
or ( n11193 , n11190 , n11192 );
buf ( n11194 , n598 );
not ( n11195 , n11194 );
buf ( n11196 , n2612 );
not ( n11197 , n11196 );
or ( n11198 , n11195 , n11197 );
buf ( n11199 , n2510 );
buf ( n11200 , n818 );
nand ( n11201 , n11199 , n11200 );
buf ( n11202 , n11201 );
buf ( n11203 , n11202 );
nand ( n11204 , n11198 , n11203 );
buf ( n11205 , n11204 );
buf ( n11206 , n11205 );
buf ( n11207 , n5630 );
nand ( n11208 , n11206 , n11207 );
buf ( n11209 , n11208 );
buf ( n11210 , n11209 );
nand ( n11211 , n11193 , n11210 );
buf ( n11212 , n11211 );
buf ( n11213 , n11212 );
xor ( n11214 , n11188 , n11213 );
buf ( n11215 , n2412 );
buf ( n11216 , n825 );
not ( n11217 , n11216 );
buf ( n11218 , n11217 );
buf ( n11219 , n11218 );
nor ( n11220 , n11215 , n11219 );
buf ( n11221 , n11220 );
buf ( n11222 , n11221 );
not ( n11223 , n5549 );
not ( n11224 , n598 );
not ( n11225 , n2431 );
or ( n11226 , n11224 , n11225 );
buf ( n11227 , n2425 );
buf ( n11228 , n818 );
nand ( n11229 , n11227 , n11228 );
buf ( n11230 , n11229 );
nand ( n11231 , n11226 , n11230 );
not ( n11232 , n11231 );
or ( n11233 , n11223 , n11232 );
buf ( n11234 , n5630 );
buf ( n11235 , n598 );
nand ( n11236 , n11234 , n11235 );
buf ( n11237 , n11236 );
buf ( n11238 , n11237 );
not ( n11239 , n11238 );
buf ( n11240 , n2466 );
not ( n11241 , n11240 );
and ( n11242 , n11239 , n11241 );
buf ( n11243 , n2466 );
buf ( n11244 , n5630 );
buf ( n11245 , n598 );
not ( n11246 , n11245 );
and ( n11247 , n11244 , n11246 );
buf ( n11248 , n11247 );
buf ( n11249 , n11248 );
and ( n11250 , n11243 , n11249 );
nor ( n11251 , n11242 , n11250 );
buf ( n11252 , n11251 );
nand ( n11253 , n11233 , n11252 );
buf ( n11254 , n11253 );
buf ( n11255 , n599 );
buf ( n11256 , n600 );
or ( n11257 , n11255 , n11256 );
buf ( n11258 , n2466 );
nand ( n11259 , n11257 , n11258 );
buf ( n11260 , n11259 );
buf ( n11261 , n11260 );
buf ( n11262 , n599 );
buf ( n11263 , n600 );
and ( n11264 , n11262 , n11263 );
buf ( n11265 , n818 );
nor ( n11266 , n11264 , n11265 );
buf ( n11267 , n11266 );
buf ( n11268 , n11267 );
nand ( n11269 , n11261 , n11268 );
buf ( n11270 , n11269 );
buf ( n11271 , n11270 );
not ( n11272 , n11271 );
and ( n11273 , n11254 , n11272 );
buf ( n11274 , n11273 );
buf ( n11275 , n11274 );
xor ( n11276 , n11222 , n11275 );
buf ( n11277 , n5549 );
not ( n11278 , n11277 );
buf ( n11279 , n11205 );
not ( n11280 , n11279 );
or ( n11281 , n11278 , n11280 );
nand ( n11282 , n11231 , n5630 );
buf ( n11283 , n11282 );
nand ( n11284 , n11281 , n11283 );
buf ( n11285 , n11284 );
buf ( n11286 , n11285 );
and ( n11287 , n11276 , n11286 );
or ( n11288 , n11287 , C0 );
buf ( n11289 , n11288 );
buf ( n11290 , n11289 );
and ( n11291 , n11214 , n11290 );
and ( n11292 , n11188 , n11213 );
or ( n11293 , n11291 , n11292 );
buf ( n11294 , n11293 );
buf ( n11295 , n11294 );
and ( n11296 , n11177 , n11295 );
and ( n11297 , n11151 , n11176 );
or ( n11298 , n11296 , n11297 );
buf ( n11299 , n11298 );
buf ( n11300 , n11299 );
xor ( n11301 , n11147 , n11300 );
buf ( n11302 , n11301 );
buf ( n11303 , n11302 );
xor ( n11304 , n11117 , n11303 );
buf ( n11305 , n5655 );
not ( n11306 , n11305 );
buf ( n11307 , n602 );
not ( n11308 , n11307 );
buf ( n11309 , n5572 );
not ( n11310 , n11309 );
or ( n11311 , n11308 , n11310 );
buf ( n11312 , n5576 );
buf ( n11313 , n2912 );
nand ( n11314 , n11312 , n11313 );
buf ( n11315 , n11314 );
buf ( n11316 , n11315 );
nand ( n11317 , n11311 , n11316 );
buf ( n11318 , n11317 );
buf ( n11319 , n11318 );
not ( n11320 , n11319 );
or ( n11321 , n11306 , n11320 );
buf ( n11322 , n602 );
not ( n11323 , n11322 );
buf ( n11324 , n5601 );
not ( n11325 , n11324 );
or ( n11326 , n11323 , n11325 );
buf ( n11327 , n7757 );
buf ( n11328 , n2912 );
nand ( n11329 , n11327 , n11328 );
buf ( n11330 , n11329 );
buf ( n11331 , n11330 );
nand ( n11332 , n11326 , n11331 );
buf ( n11333 , n11332 );
buf ( n11334 , n11333 );
buf ( n11335 , n7619 );
nand ( n11336 , n11334 , n11335 );
buf ( n11337 , n11336 );
buf ( n11338 , n11337 );
nand ( n11339 , n11321 , n11338 );
buf ( n11340 , n11339 );
buf ( n11341 , n11340 );
and ( n11342 , n11304 , n11341 );
and ( n11343 , n11117 , n11303 );
or ( n11344 , n11342 , n11343 );
buf ( n11345 , n11344 );
buf ( n11346 , n11345 );
buf ( n11347 , n7790 );
not ( n11348 , n11347 );
buf ( n11349 , n604 );
buf ( n11350 , n7648 );
and ( n11351 , n11349 , n11350 );
not ( n11352 , n11349 );
buf ( n11353 , n8684 );
and ( n11354 , n11352 , n11353 );
nor ( n11355 , n11351 , n11354 );
buf ( n11356 , n11355 );
buf ( n11357 , n11356 );
not ( n11358 , n11357 );
or ( n11359 , n11348 , n11358 );
and ( n11360 , n604 , n5369 );
not ( n11361 , n604 );
buf ( n11362 , n5373 );
buf ( n11363 , n11362 );
buf ( n11364 , n11363 );
and ( n11365 , n11361 , n11364 );
or ( n11366 , n11360 , n11365 );
buf ( n11367 , n11366 );
buf ( n11368 , n8581 );
nand ( n11369 , n11367 , n11368 );
buf ( n11370 , n11369 );
buf ( n11371 , n11370 );
nand ( n11372 , n11359 , n11371 );
buf ( n11373 , n11372 );
buf ( n11374 , n11373 );
xor ( n11375 , n11346 , n11374 );
xor ( n11376 , n11142 , n11146 );
and ( n11377 , n11376 , n11300 );
and ( n11378 , n11142 , n11146 );
or ( n11379 , n11377 , n11378 );
buf ( n11380 , n11379 );
buf ( n11381 , n11380 );
buf ( n11382 , n5655 );
not ( n11383 , n11382 );
buf ( n11384 , n10982 );
not ( n11385 , n11384 );
or ( n11386 , n11383 , n11385 );
buf ( n11387 , n11318 );
buf ( n11388 , n7619 );
nand ( n11389 , n11387 , n11388 );
buf ( n11390 , n11389 );
buf ( n11391 , n11390 );
nand ( n11392 , n11386 , n11391 );
buf ( n11393 , n11392 );
buf ( n11394 , n11393 );
xor ( n11395 , n11381 , n11394 );
xor ( n11396 , n10939 , n10943 );
xor ( n11397 , n11396 , n10962 );
buf ( n11398 , n11397 );
buf ( n11399 , n11398 );
xor ( n11400 , n11395 , n11399 );
buf ( n11401 , n11400 );
buf ( n11402 , n11401 );
and ( n11403 , n11375 , n11402 );
and ( n11404 , n11346 , n11374 );
or ( n11405 , n11403 , n11404 );
buf ( n11406 , n11405 );
buf ( n11407 , n11406 );
xor ( n11408 , n11086 , n11407 );
xor ( n11409 , n11381 , n11394 );
and ( n11410 , n11409 , n11399 );
and ( n11411 , n11381 , n11394 );
or ( n11412 , n11410 , n11411 );
buf ( n11413 , n11412 );
buf ( n11414 , n11413 );
xor ( n11415 , n10967 , n10988 );
xor ( n11416 , n11415 , n10993 );
buf ( n11417 , n11416 );
buf ( n11418 , n11417 );
xor ( n11419 , n11414 , n11418 );
buf ( n11420 , n7789 );
not ( n11421 , n11420 );
buf ( n11422 , n11015 );
not ( n11423 , n11422 );
or ( n11424 , n11421 , n11423 );
buf ( n11425 , n11356 );
buf ( n11426 , n8581 );
nand ( n11427 , n11425 , n11426 );
buf ( n11428 , n11427 );
buf ( n11429 , n11428 );
nand ( n11430 , n11424 , n11429 );
buf ( n11431 , n11430 );
buf ( n11432 , n11431 );
xor ( n11433 , n11419 , n11432 );
buf ( n11434 , n11433 );
buf ( n11435 , n11434 );
xor ( n11436 , n11408 , n11435 );
buf ( n11437 , n11436 );
buf ( n11438 , n11437 );
buf ( n11439 , n2915 );
not ( n11440 , n11439 );
buf ( n11441 , n11109 );
not ( n11442 , n11441 );
or ( n11443 , n11440 , n11442 );
buf ( n11444 , n600 );
not ( n11445 , n11444 );
buf ( n11446 , n5487 );
not ( n11447 , n11446 );
or ( n11448 , n11445 , n11447 );
buf ( n11449 , n5382 );
buf ( n11450 , n2389 );
nand ( n11451 , n11449 , n11450 );
buf ( n11452 , n11451 );
buf ( n11453 , n11452 );
nand ( n11454 , n11448 , n11453 );
buf ( n11455 , n11454 );
buf ( n11456 , n11455 );
buf ( n11457 , n5430 );
nand ( n11458 , n11456 , n11457 );
buf ( n11459 , n11458 );
buf ( n11460 , n11459 );
nand ( n11461 , n11443 , n11460 );
buf ( n11462 , n11461 );
buf ( n11463 , n11462 );
xor ( n11464 , n11151 , n11176 );
xor ( n11465 , n11464 , n11295 );
buf ( n11466 , n11465 );
buf ( n11467 , n11466 );
xor ( n11468 , n11463 , n11467 );
buf ( n11469 , n2915 );
not ( n11470 , n11469 );
buf ( n11471 , n11455 );
not ( n11472 , n11471 );
or ( n11473 , n11470 , n11472 );
buf ( n11474 , n600 );
not ( n11475 , n11474 );
buf ( n11476 , n2555 );
not ( n11477 , n11476 );
or ( n11478 , n11475 , n11477 );
buf ( n11479 , n7719 );
buf ( n11480 , n5382 );
nand ( n11481 , n11479 , n11480 );
buf ( n11482 , n11481 );
buf ( n11483 , n11482 );
nand ( n11484 , n11478 , n11483 );
buf ( n11485 , n11484 );
buf ( n11486 , n11485 );
buf ( n11487 , n5430 );
nand ( n11488 , n11486 , n11487 );
buf ( n11489 , n11488 );
buf ( n11490 , n11489 );
nand ( n11491 , n11473 , n11490 );
buf ( n11492 , n11491 );
buf ( n11493 , n11492 );
xor ( n11494 , n11188 , n11213 );
xor ( n11495 , n11494 , n11290 );
buf ( n11496 , n11495 );
buf ( n11497 , n11496 );
xor ( n11498 , n11493 , n11497 );
xor ( n11499 , n11222 , n11275 );
xor ( n11500 , n11499 , n11286 );
buf ( n11501 , n11500 );
buf ( n11502 , n11501 );
buf ( n11503 , n2915 );
not ( n11504 , n11503 );
buf ( n11505 , n11485 );
not ( n11506 , n11505 );
or ( n11507 , n11504 , n11506 );
buf ( n11508 , n600 );
not ( n11509 , n11508 );
buf ( n11510 , n2576 );
not ( n11511 , n11510 );
or ( n11512 , n11509 , n11511 );
buf ( n11513 , n2570 );
buf ( n11514 , n5382 );
nand ( n11515 , n11513 , n11514 );
buf ( n11516 , n11515 );
buf ( n11517 , n11516 );
nand ( n11518 , n11512 , n11517 );
buf ( n11519 , n11518 );
buf ( n11520 , n11519 );
buf ( n11521 , n5430 );
nand ( n11522 , n11520 , n11521 );
buf ( n11523 , n11522 );
buf ( n11524 , n11523 );
nand ( n11525 , n11507 , n11524 );
buf ( n11526 , n11525 );
buf ( n11527 , n11526 );
xor ( n11528 , n11502 , n11527 );
buf ( n11529 , n11270 );
not ( n11530 , n11529 );
buf ( n11531 , n11253 );
not ( n11532 , n11531 );
or ( n11533 , n11530 , n11532 );
buf ( n11534 , n11253 );
buf ( n11535 , n11270 );
or ( n11536 , n11534 , n11535 );
nand ( n11537 , n11533 , n11536 );
buf ( n11538 , n11537 );
buf ( n11539 , n11538 );
buf ( n11540 , n2412 );
buf ( n11541 , n5618 );
nor ( n11542 , n11540 , n11541 );
buf ( n11543 , n11542 );
buf ( n11544 , n11543 );
buf ( n11545 , n2915 );
not ( n11546 , n11545 );
buf ( n11547 , n11546 );
not ( n11548 , n600 );
nor ( n11549 , n11547 , n11548 );
not ( n11550 , n11549 );
not ( n11551 , n2431 );
or ( n11552 , n11550 , n11551 );
buf ( n11553 , n2428 );
nor ( n11554 , n11547 , n600 );
and ( n11555 , n11553 , n11554 );
buf ( n11556 , n2466 );
buf ( n11557 , n5430 );
buf ( n11558 , n600 );
not ( n11559 , n11558 );
and ( n11560 , n11557 , n11559 );
buf ( n11561 , n11560 );
buf ( n11562 , n11561 );
and ( n11563 , n11556 , n11562 );
buf ( n11564 , n2412 );
buf ( n11565 , n5430 );
buf ( n11566 , n600 );
nand ( n11567 , n11565 , n11566 );
buf ( n11568 , n11567 );
buf ( n11569 , n11568 );
not ( n11570 , n11569 );
buf ( n11571 , n11570 );
buf ( n11572 , n11571 );
and ( n11573 , n11564 , n11572 );
nor ( n11574 , n11563 , n11573 );
buf ( n11575 , n11574 );
not ( n11576 , n11575 );
nor ( n11577 , n11555 , n11576 );
nand ( n11578 , n11552 , n11577 );
buf ( n11579 , n11578 );
not ( n11580 , n11579 );
buf ( n11581 , n601 );
buf ( n11582 , n602 );
or ( n11583 , n11581 , n11582 );
buf ( n11584 , n2466 );
nand ( n11585 , n11583 , n11584 );
buf ( n11586 , n11585 );
buf ( n11587 , n11586 );
buf ( n11588 , n601 );
buf ( n11589 , n602 );
nand ( n11590 , n11588 , n11589 );
buf ( n11591 , n11590 );
buf ( n11592 , n11591 );
buf ( n11593 , n600 );
nand ( n11594 , n11587 , n11592 , n11593 );
buf ( n11595 , n11594 );
buf ( n11596 , n11595 );
nor ( n11597 , n11580 , n11596 );
buf ( n11598 , n11597 );
buf ( n11599 , n11598 );
xor ( n11600 , n11544 , n11599 );
not ( n11601 , n2915 );
not ( n11602 , n2504 );
not ( n11603 , n600 );
and ( n11604 , C1 , n11603 );
or ( n11605 , C0 , n11604 );
and ( n11606 , n11602 , n11605 );
not ( n11607 , n11602 );
not ( n11608 , n5382 );
and ( n11609 , C1 , n11608 );
or ( n11610 , n11609 , C0 );
and ( n11611 , n11607 , n11610 );
or ( n11612 , n11606 , n11611 );
not ( n11613 , n11612 );
or ( n11614 , n11601 , n11613 );
or ( n11615 , n600 , n11553 );
or ( n11616 , n2431 , n11548 );
nand ( n11617 , n11615 , n11616 , n5430 );
nand ( n11618 , n11614 , n11617 );
buf ( n11619 , n11618 );
and ( n11620 , n11600 , n11619 );
or ( n11621 , n11620 , C0 );
buf ( n11622 , n11621 );
buf ( n11623 , n11622 );
xor ( n11624 , n11539 , n11623 );
buf ( n11625 , n2915 );
not ( n11626 , n11625 );
buf ( n11627 , n11519 );
not ( n11628 , n11627 );
or ( n11629 , n11626 , n11628 );
nand ( n11630 , n11612 , n5430 );
buf ( n11631 , n11630 );
nand ( n11632 , n11629 , n11631 );
buf ( n11633 , n11632 );
buf ( n11634 , n11633 );
and ( n11635 , n11624 , n11634 );
and ( n11636 , n11539 , n11623 );
or ( n11637 , n11635 , n11636 );
buf ( n11638 , n11637 );
buf ( n11639 , n11638 );
and ( n11640 , n11528 , n11639 );
and ( n11641 , n11502 , n11527 );
or ( n11642 , n11640 , n11641 );
buf ( n11643 , n11642 );
buf ( n11644 , n11643 );
and ( n11645 , n11498 , n11644 );
and ( n11646 , n11493 , n11497 );
or ( n11647 , n11645 , n11646 );
buf ( n11648 , n11647 );
buf ( n11649 , n11648 );
and ( n11650 , n11468 , n11649 );
and ( n11651 , n11463 , n11467 );
or ( n11652 , n11650 , n11651 );
buf ( n11653 , n11652 );
buf ( n11654 , n11653 );
buf ( n11655 , n7790 );
not ( n11656 , n11655 );
buf ( n11657 , n11366 );
not ( n11658 , n11657 );
or ( n11659 , n11656 , n11658 );
buf ( n11660 , n8581 );
and ( n11661 , n604 , n5411 );
not ( n11662 , n604 );
and ( n11663 , n11662 , n5407 );
nor ( n11664 , n11661 , n11663 );
buf ( n11665 , n11664 );
nand ( n11666 , n11660 , n11665 );
buf ( n11667 , n11666 );
buf ( n11668 , n11667 );
nand ( n11669 , n11659 , n11668 );
buf ( n11670 , n11669 );
buf ( n11671 , n11670 );
xor ( n11672 , n11654 , n11671 );
xor ( n11673 , n11117 , n11303 );
xor ( n11674 , n11673 , n11341 );
buf ( n11675 , n11674 );
buf ( n11676 , n11675 );
and ( n11677 , n11672 , n11676 );
and ( n11678 , n11654 , n11671 );
or ( n11679 , n11677 , n11678 );
buf ( n11680 , n11679 );
buf ( n11681 , n11680 );
buf ( n11682 , n607 );
not ( n11683 , n11682 );
buf ( n11684 , n11078 );
not ( n11685 , n11684 );
or ( n11686 , n11683 , n11685 );
buf ( n11687 , n606 );
not ( n11688 , n11687 );
buf ( n11689 , n7593 );
not ( n11690 , n11689 );
or ( n11691 , n11688 , n11690 );
buf ( n11692 , n7599 );
buf ( n11693 , n10836 );
nand ( n11694 , n11692 , n11693 );
buf ( n11695 , n11694 );
buf ( n11696 , n11695 );
nand ( n11697 , n11691 , n11696 );
buf ( n11698 , n11697 );
buf ( n11699 , n11698 );
buf ( n11700 , n10879 );
nand ( n11701 , n11699 , n11700 );
buf ( n11702 , n11701 );
buf ( n11703 , n11702 );
nand ( n11704 , n11686 , n11703 );
buf ( n11705 , n11704 );
buf ( n11706 , n11705 );
xor ( n11707 , n11681 , n11706 );
xor ( n11708 , n11346 , n11374 );
xor ( n11709 , n11708 , n11402 );
buf ( n11710 , n11709 );
buf ( n11711 , n11710 );
and ( n11712 , n11707 , n11711 );
and ( n11713 , n11681 , n11706 );
or ( n11714 , n11712 , n11713 );
buf ( n11715 , n11714 );
buf ( n11716 , n11715 );
nor ( n11717 , n11438 , n11716 );
buf ( n11718 , n11717 );
buf ( n11719 , n11718 );
not ( n11720 , n11719 );
buf ( n11721 , n11720 );
not ( n11722 , n11721 );
xor ( n11723 , n11681 , n11706 );
xor ( n11724 , n11723 , n11711 );
buf ( n11725 , n11724 );
buf ( n11726 , n11725 );
buf ( n11727 , n5655 );
not ( n11728 , n11727 );
buf ( n11729 , n11333 );
not ( n11730 , n11729 );
or ( n11731 , n11728 , n11730 );
buf ( n11732 , n602 );
not ( n11733 , n11732 );
buf ( n11734 , n5458 );
not ( n11735 , n11734 );
or ( n11736 , n11733 , n11735 );
buf ( n11737 , n2912 );
buf ( n11738 , n5464 );
nand ( n11739 , n11737 , n11738 );
buf ( n11740 , n11739 );
buf ( n11741 , n11740 );
nand ( n11742 , n11736 , n11741 );
buf ( n11743 , n11742 );
buf ( n11744 , n11743 );
buf ( n11745 , n7619 );
nand ( n11746 , n11744 , n11745 );
buf ( n11747 , n11746 );
buf ( n11748 , n11747 );
nand ( n11749 , n11731 , n11748 );
buf ( n11750 , n11749 );
buf ( n11751 , n11750 );
buf ( n11752 , n7790 );
not ( n11753 , n11752 );
buf ( n11754 , n11664 );
not ( n11755 , n11754 );
or ( n11756 , n11753 , n11755 );
buf ( n11757 , n604 );
not ( n11758 , n11757 );
not ( n11759 , n5571 );
buf ( n11760 , n11759 );
not ( n11761 , n11760 );
or ( n11762 , n11758 , n11761 );
buf ( n11763 , n604 );
not ( n11764 , n11763 );
buf ( n11765 , n5571 );
nand ( n11766 , n11764 , n11765 );
buf ( n11767 , n11766 );
buf ( n11768 , n11767 );
nand ( n11769 , n11762 , n11768 );
buf ( n11770 , n11769 );
buf ( n11771 , n11770 );
buf ( n11772 , n8578 );
nand ( n11773 , n11771 , n11772 );
buf ( n11774 , n11773 );
buf ( n11775 , n11774 );
nand ( n11776 , n11756 , n11775 );
buf ( n11777 , n11776 );
buf ( n11778 , n11777 );
xor ( n11779 , n11751 , n11778 );
xor ( n11780 , n11463 , n11467 );
xor ( n11781 , n11780 , n11649 );
buf ( n11782 , n11781 );
buf ( n11783 , n11782 );
and ( n11784 , n11779 , n11783 );
and ( n11785 , n11751 , n11778 );
or ( n11786 , n11784 , n11785 );
buf ( n11787 , n11786 );
buf ( n11788 , n11787 );
xor ( n11789 , n11654 , n11671 );
xor ( n11790 , n11789 , n11676 );
buf ( n11791 , n11790 );
buf ( n11792 , n11791 );
xor ( n11793 , n11788 , n11792 );
buf ( n11794 , n607 );
not ( n11795 , n11794 );
buf ( n11796 , n11698 );
not ( n11797 , n11796 );
or ( n11798 , n11795 , n11797 );
not ( n11799 , n7648 );
not ( n11800 , n10836 );
or ( n11801 , n11799 , n11800 );
not ( n11802 , n7648 );
nand ( n11803 , n11802 , n606 );
nand ( n11804 , n11801 , n11803 );
buf ( n11805 , n11804 );
buf ( n11806 , n10879 );
nand ( n11807 , n11805 , n11806 );
buf ( n11808 , n11807 );
buf ( n11809 , n11808 );
nand ( n11810 , n11798 , n11809 );
buf ( n11811 , n11810 );
buf ( n11812 , n11811 );
and ( n11813 , n11793 , n11812 );
and ( n11814 , n11788 , n11792 );
or ( n11815 , n11813 , n11814 );
buf ( n11816 , n11815 );
buf ( n11817 , n11816 );
nor ( n11818 , n11726 , n11817 );
buf ( n11819 , n11818 );
not ( n11820 , n11819 );
not ( n11821 , n11820 );
buf ( n11822 , n5655 );
not ( n11823 , n11822 );
buf ( n11824 , n602 );
not ( n11825 , n11824 );
buf ( n11826 , n5487 );
not ( n11827 , n11826 );
or ( n11828 , n11825 , n11827 );
buf ( n11829 , n2912 );
buf ( n11830 , n2389 );
nand ( n11831 , n11829 , n11830 );
buf ( n11832 , n11831 );
buf ( n11833 , n11832 );
nand ( n11834 , n11828 , n11833 );
buf ( n11835 , n11834 );
buf ( n11836 , n11835 );
not ( n11837 , n11836 );
or ( n11838 , n11823 , n11837 );
buf ( n11839 , n602 );
not ( n11840 , n11839 );
buf ( n11841 , n2738 );
not ( n11842 , n11841 );
or ( n11843 , n11840 , n11842 );
buf ( n11844 , n7719 );
buf ( n11845 , n2912 );
nand ( n11846 , n11844 , n11845 );
buf ( n11847 , n11846 );
buf ( n11848 , n11847 );
nand ( n11849 , n11843 , n11848 );
buf ( n11850 , n11849 );
buf ( n11851 , n11850 );
buf ( n11852 , n7619 );
nand ( n11853 , n11851 , n11852 );
buf ( n11854 , n11853 );
buf ( n11855 , n11854 );
nand ( n11856 , n11838 , n11855 );
buf ( n11857 , n11856 );
buf ( n11858 , n11857 );
xor ( n11859 , n11539 , n11623 );
xor ( n11860 , n11859 , n11634 );
buf ( n11861 , n11860 );
buf ( n11862 , n11861 );
xor ( n11863 , n11858 , n11862 );
xor ( n11864 , n11544 , n11599 );
xor ( n11865 , n11864 , n11619 );
buf ( n11866 , n11865 );
buf ( n11867 , n11866 );
buf ( n11868 , n5655 );
not ( n11869 , n11868 );
buf ( n11870 , n11850 );
not ( n11871 , n11870 );
or ( n11872 , n11869 , n11871 );
buf ( n11873 , n2912 );
not ( n11874 , n11873 );
buf ( n11875 , n2570 );
not ( n11876 , n11875 );
or ( n11877 , n11874 , n11876 );
not ( n11878 , n2570 );
nand ( n11879 , n11878 , n602 );
buf ( n11880 , n11879 );
nand ( n11881 , n11877 , n11880 );
buf ( n11882 , n11881 );
buf ( n11883 , n11882 );
buf ( n11884 , n7619 );
nand ( n11885 , n11883 , n11884 );
buf ( n11886 , n11885 );
buf ( n11887 , n11886 );
nand ( n11888 , n11872 , n11887 );
buf ( n11889 , n11888 );
buf ( n11890 , n11889 );
xor ( n11891 , n11867 , n11890 );
buf ( n11892 , n11595 );
not ( n11893 , n11892 );
buf ( n11894 , n11578 );
not ( n11895 , n11894 );
or ( n11896 , n11893 , n11895 );
buf ( n11897 , n11578 );
buf ( n11898 , n11595 );
or ( n11899 , n11897 , n11898 );
nand ( n11900 , n11896 , n11899 );
buf ( n11901 , n11900 );
buf ( n11902 , n11901 );
buf ( n11903 , n2412 );
buf ( n11904 , n11547 );
nor ( n11905 , n11903 , n11904 );
buf ( n11906 , n11905 );
buf ( n11907 , n11906 );
buf ( n11908 , n2912 );
buf ( n11909 , n2425 );
and ( n11910 , n11908 , n11909 );
not ( n11911 , n11908 );
buf ( n11912 , n2437 );
and ( n11913 , n11911 , n11912 );
nor ( n11914 , n11910 , n11913 );
buf ( n11915 , n11914 );
buf ( n11916 , n11915 );
buf ( n11917 , n5652 );
or ( n11918 , n11916 , n11917 );
buf ( n11919 , n2466 );
buf ( n11920 , n7619 );
buf ( n11921 , n2912 );
and ( n11922 , n11920 , n11921 );
buf ( n11923 , n11922 );
buf ( n11924 , n11923 );
and ( n11925 , n11919 , n11924 );
buf ( n11926 , n2412 );
buf ( n11927 , n7619 );
buf ( n11928 , n602 );
and ( n11929 , n11927 , n11928 );
buf ( n11930 , n11929 );
buf ( n11931 , n11930 );
and ( n11932 , n11926 , n11931 );
nor ( n11933 , n11925 , n11932 );
buf ( n11934 , n11933 );
buf ( n11935 , n11934 );
nand ( n11936 , n11918 , n11935 );
buf ( n11937 , n11936 );
buf ( n11938 , n11937 );
not ( n11939 , n11938 );
buf ( n11940 , n603 );
buf ( n11941 , n604 );
or ( n11942 , n11940 , n11941 );
buf ( n11943 , n2466 );
nand ( n11944 , n11942 , n11943 );
buf ( n11945 , n11944 );
buf ( n11946 , n11945 );
buf ( n11947 , n5651 );
buf ( n11948 , n602 );
nand ( n11949 , n11946 , n11947 , n11948 );
buf ( n11950 , n11949 );
buf ( n11951 , n11950 );
nor ( n11952 , n11939 , n11951 );
buf ( n11953 , n11952 );
buf ( n11954 , n11953 );
xor ( n11955 , n11907 , n11954 );
or ( n11956 , n5652 , n2912 );
nor ( n11957 , n11956 , n2510 );
not ( n11958 , n7619 );
nor ( n11959 , n11958 , n11915 );
nor ( n11960 , n11957 , n11959 );
not ( n11961 , n5652 );
nand ( n11962 , n11961 , n2510 , n2912 );
nand ( n11963 , n11960 , n11962 );
buf ( n11964 , n11963 );
and ( n11965 , n11955 , n11964 );
or ( n11966 , n11965 , C0 );
buf ( n11967 , n11966 );
buf ( n11968 , n11967 );
xor ( n11969 , n11902 , n11968 );
buf ( n11970 , n5655 );
not ( n11971 , n11970 );
buf ( n11972 , n11882 );
not ( n11973 , n11972 );
or ( n11974 , n11971 , n11973 );
xnor ( n11975 , n2912 , n2510 );
nand ( n11976 , n11975 , n7619 );
buf ( n11977 , n11976 );
nand ( n11978 , n11974 , n11977 );
buf ( n11979 , n11978 );
buf ( n11980 , n11979 );
and ( n11981 , n11969 , n11980 );
and ( n11982 , n11902 , n11968 );
or ( n11983 , n11981 , n11982 );
buf ( n11984 , n11983 );
buf ( n11985 , n11984 );
and ( n11986 , n11891 , n11985 );
and ( n11987 , n11867 , n11890 );
or ( n11988 , n11986 , n11987 );
buf ( n11989 , n11988 );
buf ( n11990 , n11989 );
and ( n11991 , n11863 , n11990 );
and ( n11992 , n11858 , n11862 );
or ( n11993 , n11991 , n11992 );
buf ( n11994 , n11993 );
buf ( n11995 , n11994 );
buf ( n11996 , n607 );
not ( n11997 , n11996 );
buf ( n11998 , n606 );
buf ( n11999 , n5411 );
and ( n12000 , n11998 , n11999 );
not ( n12001 , n11998 );
buf ( n12002 , n5407 );
and ( n12003 , n12001 , n12002 );
nor ( n12004 , n12000 , n12003 );
buf ( n12005 , n12004 );
buf ( n12006 , n12005 );
not ( n12007 , n12006 );
or ( n12008 , n11997 , n12007 );
buf ( n12009 , n606 );
not ( n12010 , n12009 );
buf ( n12011 , n11759 );
not ( n12012 , n12011 );
or ( n12013 , n12010 , n12012 );
buf ( n12014 , n10836 );
buf ( n12015 , n5571 );
nand ( n12016 , n12014 , n12015 );
buf ( n12017 , n12016 );
buf ( n12018 , n12017 );
nand ( n12019 , n12013 , n12018 );
buf ( n12020 , n12019 );
buf ( n12021 , n12020 );
buf ( n12022 , n10879 );
nand ( n12023 , n12021 , n12022 );
buf ( n12024 , n12023 );
buf ( n12025 , n12024 );
nand ( n12026 , n12008 , n12025 );
buf ( n12027 , n12026 );
buf ( n12028 , n12027 );
xor ( n12029 , n11995 , n12028 );
buf ( n12030 , n5655 );
not ( n12031 , n12030 );
buf ( n12032 , n602 );
not ( n12033 , n12032 );
buf ( n12034 , n11096 );
not ( n12035 , n12034 );
or ( n12036 , n12033 , n12035 );
buf ( n12037 , n11102 );
buf ( n12038 , n2912 );
nand ( n12039 , n12037 , n12038 );
buf ( n12040 , n12039 );
buf ( n12041 , n12040 );
nand ( n12042 , n12036 , n12041 );
buf ( n12043 , n12042 );
buf ( n12044 , n12043 );
not ( n12045 , n12044 );
or ( n12046 , n12031 , n12045 );
buf ( n12047 , n11835 );
buf ( n12048 , n7619 );
nand ( n12049 , n12047 , n12048 );
buf ( n12050 , n12049 );
buf ( n12051 , n12050 );
nand ( n12052 , n12046 , n12051 );
buf ( n12053 , n12052 );
buf ( n12054 , n12053 );
xor ( n12055 , n11502 , n11527 );
xor ( n12056 , n12055 , n11639 );
buf ( n12057 , n12056 );
buf ( n12058 , n12057 );
xor ( n12059 , n12054 , n12058 );
buf ( n12060 , n7789 );
not ( n12061 , n12060 );
buf ( n12062 , n604 );
not ( n12063 , n12062 );
buf ( n12064 , n5598 );
not ( n12065 , n12064 );
or ( n12066 , n12063 , n12065 );
buf ( n12067 , n604 );
not ( n12068 , n12067 );
buf ( n12069 , n7751 );
nand ( n12070 , n12068 , n12069 );
buf ( n12071 , n12070 );
buf ( n12072 , n12071 );
nand ( n12073 , n12066 , n12072 );
buf ( n12074 , n12073 );
buf ( n12075 , n12074 );
not ( n12076 , n12075 );
or ( n12077 , n12061 , n12076 );
not ( n12078 , n604 );
not ( n12079 , n5458 );
or ( n12080 , n12078 , n12079 );
buf ( n12081 , n604 );
not ( n12082 , n12081 );
buf ( n12083 , n5455 );
nand ( n12084 , n12082 , n12083 );
buf ( n12085 , n12084 );
nand ( n12086 , n12080 , n12085 );
buf ( n12087 , n12086 );
buf ( n12088 , n8578 );
nand ( n12089 , n12087 , n12088 );
buf ( n12090 , n12089 );
buf ( n12091 , n12090 );
nand ( n12092 , n12077 , n12091 );
buf ( n12093 , n12092 );
buf ( n12094 , n12093 );
xor ( n12095 , n12059 , n12094 );
buf ( n12096 , n12095 );
buf ( n12097 , n12096 );
xor ( n12098 , n12029 , n12097 );
buf ( n12099 , n12098 );
buf ( n12100 , n12099 );
not ( n12101 , n12100 );
not ( n12102 , n7789 );
not ( n12103 , n12086 );
or ( n12104 , n12102 , n12103 );
xor ( n12105 , n604 , n2361 );
nand ( n12106 , n12105 , n8578 );
nand ( n12107 , n12104 , n12106 );
buf ( n12108 , n12107 );
xor ( n12109 , n11858 , n11862 );
xor ( n12110 , n12109 , n11990 );
buf ( n12111 , n12110 );
buf ( n12112 , n12111 );
xor ( n12113 , n12108 , n12112 );
buf ( n12114 , n607 );
not ( n12115 , n12114 );
buf ( n12116 , n12020 );
not ( n12117 , n12116 );
or ( n12118 , n12115 , n12117 );
buf ( n12119 , n606 );
not ( n12120 , n12119 );
buf ( n12121 , n5598 );
not ( n12122 , n12121 );
or ( n12123 , n12120 , n12122 );
not ( n12124 , n5598 );
nand ( n12125 , n12124 , n10836 );
buf ( n12126 , n12125 );
nand ( n12127 , n12123 , n12126 );
buf ( n12128 , n12127 );
buf ( n12129 , n12128 );
buf ( n12130 , n10879 );
nand ( n12131 , n12129 , n12130 );
buf ( n12132 , n12131 );
buf ( n12133 , n12132 );
nand ( n12134 , n12118 , n12133 );
buf ( n12135 , n12134 );
buf ( n12136 , n12135 );
and ( n12137 , n12113 , n12136 );
and ( n12138 , n12108 , n12112 );
or ( n12139 , n12137 , n12138 );
buf ( n12140 , n12139 );
buf ( n12141 , n12140 );
not ( n12142 , n12141 );
buf ( n12143 , n12142 );
buf ( n12144 , n12143 );
nand ( n12145 , n12101 , n12144 );
buf ( n12146 , n12145 );
not ( n12147 , n12146 );
buf ( n12148 , n7789 );
not ( n12149 , n12148 );
buf ( n12150 , n12105 );
not ( n12151 , n12150 );
or ( n12152 , n12149 , n12151 );
not ( n12153 , n2389 );
and ( n12154 , n604 , n12153 );
not ( n12155 , n604 );
and ( n12156 , n12155 , n2389 );
or ( n12157 , n12154 , n12156 );
buf ( n12158 , n12157 );
buf ( n12159 , n8578 );
nand ( n12160 , n12158 , n12159 );
buf ( n12161 , n12160 );
buf ( n12162 , n12161 );
nand ( n12163 , n12152 , n12162 );
buf ( n12164 , n12163 );
buf ( n12165 , n12164 );
xor ( n12166 , n11867 , n11890 );
xor ( n12167 , n12166 , n11985 );
buf ( n12168 , n12167 );
buf ( n12169 , n12168 );
xor ( n12170 , n12165 , n12169 );
buf ( n12171 , n607 );
not ( n12172 , n12171 );
buf ( n12173 , n12128 );
not ( n12174 , n12173 );
or ( n12175 , n12172 , n12174 );
buf ( n12176 , n606 );
buf ( n12177 , n5455 );
xor ( n12178 , n12176 , n12177 );
buf ( n12179 , n12178 );
buf ( n12180 , n12179 );
buf ( n12181 , n10879 );
nand ( n12182 , n12180 , n12181 );
buf ( n12183 , n12182 );
buf ( n12184 , n12183 );
nand ( n12185 , n12175 , n12184 );
buf ( n12186 , n12185 );
buf ( n12187 , n12186 );
and ( n12188 , n12170 , n12187 );
and ( n12189 , n12165 , n12169 );
or ( n12190 , n12188 , n12189 );
buf ( n12191 , n12190 );
xor ( n12192 , n12108 , n12112 );
xor ( n12193 , n12192 , n12136 );
buf ( n12194 , n12193 );
xor ( n12195 , n12191 , n12194 );
buf ( n12196 , n7789 );
not ( n12197 , n12196 );
buf ( n12198 , n12157 );
not ( n12199 , n12198 );
or ( n12200 , n12197 , n12199 );
buf ( n12201 , n604 );
not ( n12202 , n12201 );
buf ( n12203 , n2555 );
not ( n12204 , n12203 );
or ( n12205 , n12202 , n12204 );
buf ( n12206 , n604 );
not ( n12207 , n12206 );
buf ( n12208 , n2552 );
nand ( n12209 , n12207 , n12208 );
buf ( n12210 , n12209 );
buf ( n12211 , n12210 );
nand ( n12212 , n12205 , n12211 );
buf ( n12213 , n12212 );
buf ( n12214 , n12213 );
buf ( n12215 , n8578 );
nand ( n12216 , n12214 , n12215 );
buf ( n12217 , n12216 );
buf ( n12218 , n12217 );
nand ( n12219 , n12200 , n12218 );
buf ( n12220 , n12219 );
buf ( n12221 , n12220 );
xor ( n12222 , n11902 , n11968 );
xor ( n12223 , n12222 , n11980 );
buf ( n12224 , n12223 );
buf ( n12225 , n12224 );
xor ( n12226 , n12221 , n12225 );
xor ( n12227 , n11907 , n11954 );
xor ( n12228 , n12227 , n11964 );
buf ( n12229 , n12228 );
buf ( n12230 , n12229 );
buf ( n12231 , n7789 );
not ( n12232 , n12231 );
buf ( n12233 , n12213 );
not ( n12234 , n12233 );
or ( n12235 , n12232 , n12234 );
not ( n12236 , n604 );
not ( n12237 , n11878 );
or ( n12238 , n12236 , n12237 );
or ( n12239 , n11878 , n604 );
nand ( n12240 , n12238 , n12239 );
buf ( n12241 , n12240 );
buf ( n12242 , n8578 );
nand ( n12243 , n12241 , n12242 );
buf ( n12244 , n12243 );
buf ( n12245 , n12244 );
nand ( n12246 , n12235 , n12245 );
buf ( n12247 , n12246 );
buf ( n12248 , n12247 );
xor ( n12249 , n12230 , n12248 );
buf ( n12250 , n11950 );
not ( n12251 , n12250 );
buf ( n12252 , n11937 );
not ( n12253 , n12252 );
or ( n12254 , n12251 , n12253 );
buf ( n12255 , n11937 );
buf ( n12256 , n11950 );
or ( n12257 , n12255 , n12256 );
nand ( n12258 , n12254 , n12257 );
buf ( n12259 , n12258 );
buf ( n12260 , n12259 );
buf ( n12261 , n7789 );
not ( n12262 , n12261 );
buf ( n12263 , n12240 );
not ( n12264 , n12263 );
or ( n12265 , n12262 , n12264 );
and ( n12266 , n604 , n2612 );
not ( n12267 , n604 );
and ( n12268 , n12267 , n2510 );
or ( n12269 , n12266 , n12268 );
buf ( n12270 , n12269 );
buf ( n12271 , n8578 );
nand ( n12272 , n12270 , n12271 );
buf ( n12273 , n12272 );
buf ( n12274 , n12273 );
nand ( n12275 , n12265 , n12274 );
buf ( n12276 , n12275 );
buf ( n12277 , n12276 );
xor ( n12278 , n12260 , n12277 );
buf ( n12279 , n2412 );
buf ( n12280 , n5652 );
nor ( n12281 , n12279 , n12280 );
buf ( n12282 , n12281 );
buf ( n12283 , n12282 );
buf ( n12284 , n7789 );
not ( n12285 , n12284 );
buf ( n12286 , n604 );
not ( n12287 , n12286 );
buf ( n12288 , n2424 );
not ( n12289 , n12288 );
or ( n12290 , n12287 , n12289 );
buf ( n12291 , n604 );
not ( n12292 , n12291 );
buf ( n12293 , n2425 );
nand ( n12294 , n12292 , n12293 );
buf ( n12295 , n12294 );
buf ( n12296 , n12295 );
nand ( n12297 , n12290 , n12296 );
buf ( n12298 , n12297 );
buf ( n12299 , n12298 );
not ( n12300 , n12299 );
or ( n12301 , n12285 , n12300 );
buf ( n12302 , n604 );
buf ( n12303 , n2466 );
and ( n12304 , n12302 , n12303 );
not ( n12305 , n12302 );
buf ( n12306 , n2412 );
and ( n12307 , n12305 , n12306 );
nor ( n12308 , n12304 , n12307 );
buf ( n12309 , n12308 );
buf ( n12310 , n12309 );
buf ( n12311 , n8578 );
nand ( n12312 , n12310 , n12311 );
buf ( n12313 , n12312 );
buf ( n12314 , n12313 );
nand ( n12315 , n12301 , n12314 );
buf ( n12316 , n12315 );
buf ( n12317 , n12316 );
not ( n12318 , n12317 );
buf ( n12319 , n605 );
buf ( n12320 , n606 );
or ( n12321 , n12319 , n12320 );
buf ( n12322 , n2466 );
nand ( n12323 , n12321 , n12322 );
buf ( n12324 , n12323 );
buf ( n12325 , n12324 );
buf ( n12326 , n605 );
buf ( n12327 , n606 );
and ( n12328 , n12326 , n12327 );
not ( n12329 , n604 );
buf ( n12330 , n12329 );
nor ( n12331 , n12328 , n12330 );
buf ( n12332 , n12331 );
buf ( n12333 , n12332 );
nand ( n12334 , n12325 , n12333 );
buf ( n12335 , n12334 );
buf ( n12336 , n12335 );
nor ( n12337 , n12318 , n12336 );
buf ( n12338 , n12337 );
buf ( n12339 , n12338 );
xor ( n12340 , n12283 , n12339 );
buf ( n12341 , n7789 );
not ( n12342 , n12341 );
buf ( n12343 , n12269 );
not ( n12344 , n12343 );
or ( n12345 , n12342 , n12344 );
buf ( n12346 , n12298 );
buf ( n12347 , n8578 );
nand ( n12348 , n12346 , n12347 );
buf ( n12349 , n12348 );
buf ( n12350 , n12349 );
nand ( n12351 , n12345 , n12350 );
buf ( n12352 , n12351 );
buf ( n12353 , n12352 );
and ( n12354 , n12340 , n12353 );
or ( n12355 , n12354 , C0 );
buf ( n12356 , n12355 );
buf ( n12357 , n12356 );
and ( n12358 , n12278 , n12357 );
and ( n12359 , n12260 , n12277 );
or ( n12360 , n12358 , n12359 );
buf ( n12361 , n12360 );
buf ( n12362 , n12361 );
and ( n12363 , n12249 , n12362 );
and ( n12364 , n12230 , n12248 );
or ( n12365 , n12363 , n12364 );
buf ( n12366 , n12365 );
buf ( n12367 , n12366 );
and ( n12368 , n12226 , n12367 );
and ( n12369 , n12221 , n12225 );
or ( n12370 , n12368 , n12369 );
buf ( n12371 , n12370 );
xor ( n12372 , n12165 , n12169 );
xor ( n12373 , n12372 , n12187 );
buf ( n12374 , n12373 );
xor ( n12375 , n12371 , n12374 );
xor ( n12376 , n12230 , n12248 );
xor ( n12377 , n12376 , n12362 );
buf ( n12378 , n12377 );
not ( n12379 , n12378 );
buf ( n12380 , n607 );
not ( n12381 , n12380 );
buf ( n12382 , n606 );
buf ( n12383 , n2361 );
and ( n12384 , n12382 , n12383 );
not ( n12385 , n12382 );
buf ( n12386 , n11096 );
and ( n12387 , n12385 , n12386 );
nor ( n12388 , n12384 , n12387 );
buf ( n12389 , n12388 );
buf ( n12390 , n12389 );
not ( n12391 , n12390 );
or ( n12392 , n12381 , n12391 );
not ( n12393 , n606 );
not ( n12394 , n5487 );
or ( n12395 , n12393 , n12394 );
buf ( n12396 , n2389 );
buf ( n12397 , n10836 );
nand ( n12398 , n12396 , n12397 );
buf ( n12399 , n12398 );
nand ( n12400 , n12395 , n12399 );
buf ( n12401 , n12400 );
buf ( n12402 , n10879 );
nand ( n12403 , n12401 , n12402 );
buf ( n12404 , n12403 );
buf ( n12405 , n12404 );
nand ( n12406 , n12392 , n12405 );
buf ( n12407 , n12406 );
not ( n12408 , n12407 );
nand ( n12409 , n12379 , n12408 );
not ( n12410 , n607 );
not ( n12411 , n12399 );
not ( n12412 , n12411 );
or ( n12413 , n12410 , n12412 );
and ( n12414 , n607 , n606 );
and ( n12415 , n12153 , n12414 );
and ( n12416 , n2549 , n10836 );
not ( n12417 , n2549 );
and ( n12418 , n12417 , n606 );
or ( n12419 , n12416 , n12418 );
and ( n12420 , n12419 , n10879 );
nor ( n12421 , n12415 , n12420 );
nand ( n12422 , n12413 , n12421 );
buf ( n12423 , n12422 );
xor ( n12424 , n12260 , n12277 );
xor ( n12425 , n12424 , n12357 );
buf ( n12426 , n12425 );
buf ( n12427 , n12426 );
xor ( n12428 , n12423 , n12427 );
buf ( n12429 , n12335 );
not ( n12430 , n12429 );
buf ( n12431 , n12316 );
not ( n12432 , n12431 );
or ( n12433 , n12430 , n12432 );
buf ( n12434 , n12316 );
buf ( n12435 , n12335 );
or ( n12436 , n12434 , n12435 );
nand ( n12437 , n12433 , n12436 );
buf ( n12438 , n12437 );
buf ( n12439 , n12438 );
buf ( n12440 , n2412 );
buf ( n12441 , n7789 );
not ( n12442 , n12441 );
buf ( n12443 , n12442 );
buf ( n12444 , n12443 );
nor ( n12445 , n12440 , n12444 );
buf ( n12446 , n12445 );
buf ( n12447 , n12446 );
buf ( n12448 , n606 );
not ( n12449 , n12448 );
buf ( n12450 , n2424 );
not ( n12451 , n12450 );
or ( n12452 , n12449 , n12451 );
buf ( n12453 , n2425 );
buf ( n12454 , n10836 );
nand ( n12455 , n12453 , n12454 );
buf ( n12456 , n12455 );
buf ( n12457 , n12456 );
nand ( n12458 , n12452 , n12457 );
buf ( n12459 , n12458 );
buf ( n12460 , n12459 );
buf ( n12461 , n607 );
and ( n12462 , n12460 , n12461 );
buf ( n12463 , n10876 );
not ( n12464 , n12463 );
buf ( n12465 , n2466 );
nor ( n12466 , n12464 , n12465 );
buf ( n12467 , n12466 );
buf ( n12468 , n12467 );
nor ( n12469 , n12462 , n12468 );
buf ( n12470 , n12469 );
buf ( n12471 , n12470 );
buf ( n12472 , n2412 );
buf ( n12473 , n607 );
not ( n12474 , n12473 );
buf ( n12475 , n12474 );
buf ( n12476 , n12475 );
nor ( n12477 , n12472 , n12476 );
buf ( n12478 , n12477 );
buf ( n12479 , n12478 );
buf ( n12480 , n12479 );
buf ( n12481 , n12480 );
buf ( n12482 , n12481 );
buf ( n12483 , n10836 );
or ( n12484 , n12482 , n12483 );
buf ( n12485 , n12484 );
buf ( n12486 , n12485 );
nor ( n12487 , n12471 , n12486 );
buf ( n12488 , n12487 );
buf ( n12489 , n12488 );
xor ( n12490 , n12447 , n12489 );
xor ( n12491 , n2506 , n10836 );
buf ( n12492 , n12491 );
buf ( n12493 , n12475 );
or ( n12494 , n12492 , n12493 );
buf ( n12495 , n10876 );
buf ( n12496 , n12459 );
nand ( n12497 , n12495 , n12496 );
buf ( n12498 , n12497 );
buf ( n12499 , n12498 );
nand ( n12500 , n12494 , n12499 );
buf ( n12501 , n12500 );
buf ( n12502 , n12501 );
and ( n12503 , n12490 , n12502 );
or ( n12504 , n12503 , C0 );
buf ( n12505 , n12504 );
buf ( n12506 , n12505 );
xor ( n12507 , n12439 , n12506 );
not ( n12508 , n10836 );
not ( n12509 , n11878 );
or ( n12510 , n12508 , n12509 );
nand ( n12511 , n2570 , n606 );
nand ( n12512 , n12510 , n12511 );
buf ( n12513 , n12512 );
buf ( n12514 , n12475 );
or ( n12515 , n12513 , n12514 );
buf ( n12516 , n12491 );
not ( n12517 , n12516 );
buf ( n12518 , n10879 );
nand ( n12519 , n12517 , n12518 );
buf ( n12520 , n12519 );
buf ( n12521 , n12520 );
nand ( n12522 , n12515 , n12521 );
buf ( n12523 , n12522 );
buf ( n12524 , n12523 );
and ( n12525 , n12507 , n12524 );
and ( n12526 , n12439 , n12506 );
or ( n12527 , n12525 , n12526 );
buf ( n12528 , n12527 );
not ( n12529 , n12528 );
buf ( n12530 , n607 );
not ( n12531 , n12530 );
buf ( n12532 , n12419 );
not ( n12533 , n12532 );
or ( n12534 , n12531 , n12533 );
buf ( n12535 , n12512 );
not ( n12536 , n12535 );
buf ( n12537 , n10879 );
nand ( n12538 , n12536 , n12537 );
buf ( n12539 , n12538 );
buf ( n12540 , n12539 );
nand ( n12541 , n12534 , n12540 );
buf ( n12542 , n12541 );
xor ( n12543 , n12283 , n12339 );
xor ( n12544 , n12543 , n12353 );
buf ( n12545 , n12544 );
nor ( n12546 , n12542 , n12545 );
or ( n12547 , n12529 , n12546 );
nand ( n12548 , n12545 , n12542 );
nand ( n12549 , n12547 , n12548 );
buf ( n12550 , n12549 );
and ( n12551 , n12428 , n12550 );
and ( n12552 , n12423 , n12427 );
or ( n12553 , n12551 , n12552 );
buf ( n12554 , n12553 );
and ( n12555 , n12409 , n12554 );
and ( n12556 , n12378 , n12407 );
nor ( n12557 , n12555 , n12556 );
buf ( n12558 , n12557 );
xor ( n12559 , n12221 , n12225 );
xor ( n12560 , n12559 , n12367 );
buf ( n12561 , n12560 );
buf ( n12562 , n12561 );
not ( n12563 , n12389 );
not ( n12564 , n10879 );
or ( n12565 , n12563 , n12564 );
buf ( n12566 , n12179 );
not ( n12567 , n12566 );
buf ( n12568 , n12567 );
or ( n12569 , n12568 , n12475 );
nand ( n12570 , n12565 , n12569 );
buf ( n12571 , n12570 );
nor ( n12572 , n12562 , n12571 );
buf ( n12573 , n12572 );
buf ( n12574 , n12573 );
or ( n12575 , n12558 , n12574 );
buf ( n12576 , n12561 );
buf ( n12577 , n12570 );
nand ( n12578 , n12576 , n12577 );
buf ( n12579 , n12578 );
buf ( n12580 , n12579 );
nand ( n12581 , n12575 , n12580 );
buf ( n12582 , n12581 );
and ( n12583 , n12375 , n12582 );
and ( n12584 , n12371 , n12374 );
or ( n12585 , n12583 , n12584 );
and ( n12586 , n12195 , n12585 );
and ( n12587 , n12191 , n12194 );
or ( n12588 , n12586 , n12587 );
not ( n12589 , n12588 );
or ( n12590 , n12147 , n12589 );
buf ( n12591 , n12099 );
buf ( n12592 , n12140 );
nand ( n12593 , n12591 , n12592 );
buf ( n12594 , n12593 );
nand ( n12595 , n12590 , n12594 );
buf ( n12596 , n12595 );
not ( n12597 , n12596 );
xor ( n12598 , n11995 , n12028 );
and ( n12599 , n12598 , n12097 );
and ( n12600 , n11995 , n12028 );
or ( n12601 , n12599 , n12600 );
buf ( n12602 , n12601 );
not ( n12603 , n12602 );
buf ( n12604 , n607 );
not ( n12605 , n12604 );
and ( n12606 , n606 , n5369 );
not ( n12607 , n606 );
and ( n12608 , n12607 , n5373 );
or ( n12609 , n12606 , n12608 );
buf ( n12610 , n12609 );
not ( n12611 , n12610 );
or ( n12612 , n12605 , n12611 );
buf ( n12613 , n12005 );
buf ( n12614 , n10879 );
nand ( n12615 , n12613 , n12614 );
buf ( n12616 , n12615 );
buf ( n12617 , n12616 );
nand ( n12618 , n12612 , n12617 );
buf ( n12619 , n12618 );
buf ( n12620 , n12619 );
xor ( n12621 , n12054 , n12058 );
and ( n12622 , n12621 , n12094 );
and ( n12623 , n12054 , n12058 );
or ( n12624 , n12622 , n12623 );
buf ( n12625 , n12624 );
buf ( n12626 , n12625 );
xor ( n12627 , n12620 , n12626 );
buf ( n12628 , n5655 );
not ( n12629 , n12628 );
buf ( n12630 , n11743 );
not ( n12631 , n12630 );
or ( n12632 , n12629 , n12631 );
buf ( n12633 , n12043 );
buf ( n12634 , n7619 );
nand ( n12635 , n12633 , n12634 );
buf ( n12636 , n12635 );
buf ( n12637 , n12636 );
nand ( n12638 , n12632 , n12637 );
buf ( n12639 , n12638 );
buf ( n12640 , n12639 );
xor ( n12641 , n11493 , n11497 );
xor ( n12642 , n12641 , n11644 );
buf ( n12643 , n12642 );
buf ( n12644 , n12643 );
xor ( n12645 , n12640 , n12644 );
buf ( n12646 , n7789 );
not ( n12647 , n12646 );
buf ( n12648 , n11770 );
not ( n12649 , n12648 );
or ( n12650 , n12647 , n12649 );
buf ( n12651 , n12074 );
buf ( n12652 , n12651 );
buf ( n12653 , n12652 );
buf ( n12654 , n12653 );
buf ( n12655 , n8578 );
nand ( n12656 , n12654 , n12655 );
buf ( n12657 , n12656 );
buf ( n12658 , n12657 );
nand ( n12659 , n12650 , n12658 );
buf ( n12660 , n12659 );
buf ( n12661 , n12660 );
xor ( n12662 , n12645 , n12661 );
buf ( n12663 , n12662 );
buf ( n12664 , n12663 );
xor ( n12665 , n12627 , n12664 );
buf ( n12666 , n12665 );
buf ( n12667 , n12666 );
not ( n12668 , n12667 );
buf ( n12669 , n12668 );
nand ( n12670 , n12603 , n12669 );
buf ( n12671 , n12670 );
not ( n12672 , n12671 );
or ( n12673 , n12597 , n12672 );
buf ( n12674 , n12669 );
not ( n12675 , n12674 );
buf ( n12676 , n12602 );
nand ( n12677 , n12675 , n12676 );
buf ( n12678 , n12677 );
buf ( n12679 , n12678 );
nand ( n12680 , n12673 , n12679 );
buf ( n12681 , n12680 );
buf ( n12682 , n12681 );
not ( n12683 , n12682 );
xor ( n12684 , n12640 , n12644 );
and ( n12685 , n12684 , n12661 );
and ( n12686 , n12640 , n12644 );
or ( n12687 , n12685 , n12686 );
buf ( n12688 , n12687 );
buf ( n12689 , n12688 );
xor ( n12690 , n11751 , n11778 );
xor ( n12691 , n12690 , n11783 );
buf ( n12692 , n12691 );
buf ( n12693 , n12692 );
xor ( n12694 , n12689 , n12693 );
buf ( n12695 , n607 );
not ( n12696 , n12695 );
buf ( n12697 , n11804 );
not ( n12698 , n12697 );
or ( n12699 , n12696 , n12698 );
buf ( n12700 , n12609 );
buf ( n12701 , n10879 );
nand ( n12702 , n12700 , n12701 );
buf ( n12703 , n12702 );
buf ( n12704 , n12703 );
nand ( n12705 , n12699 , n12704 );
buf ( n12706 , n12705 );
buf ( n12707 , n12706 );
xor ( n12708 , n12694 , n12707 );
buf ( n12709 , n12708 );
buf ( n12710 , n12709 );
xor ( n12711 , n12620 , n12626 );
and ( n12712 , n12711 , n12664 );
and ( n12713 , n12620 , n12626 );
or ( n12714 , n12712 , n12713 );
buf ( n12715 , n12714 );
buf ( n12716 , n12715 );
nor ( n12717 , n12710 , n12716 );
buf ( n12718 , n12717 );
buf ( n12719 , n12718 );
not ( n12720 , n12719 );
buf ( n12721 , n12720 );
buf ( n12722 , n12721 );
not ( n12723 , n12722 );
or ( n12724 , n12683 , n12723 );
buf ( n12725 , n12709 );
buf ( n12726 , n12715 );
nand ( n12727 , n12725 , n12726 );
buf ( n12728 , n12727 );
buf ( n12729 , n12728 );
nand ( n12730 , n12724 , n12729 );
buf ( n12731 , n12730 );
not ( n12732 , n12731 );
xor ( n12733 , n11788 , n11792 );
xor ( n12734 , n12733 , n11812 );
buf ( n12735 , n12734 );
buf ( n12736 , n12735 );
not ( n12737 , n12736 );
xor ( n12738 , n12689 , n12693 );
and ( n12739 , n12738 , n12707 );
and ( n12740 , n12689 , n12693 );
or ( n12741 , n12739 , n12740 );
buf ( n12742 , n12741 );
buf ( n12743 , n12742 );
not ( n12744 , n12743 );
buf ( n12745 , n12744 );
buf ( n12746 , n12745 );
nand ( n12747 , n12737 , n12746 );
buf ( n12748 , n12747 );
not ( n12749 , n12748 );
or ( n12750 , n12732 , n12749 );
buf ( n12751 , n12735 );
buf ( n12752 , n12742 );
nand ( n12753 , n12751 , n12752 );
buf ( n12754 , n12753 );
nand ( n12755 , n12750 , n12754 );
not ( n12756 , n12755 );
or ( n12757 , n11821 , n12756 );
nand ( n12758 , n11725 , n11816 );
nand ( n12759 , n12757 , n12758 );
not ( n12760 , n12759 );
or ( n12761 , n11722 , n12760 );
buf ( n12762 , n11437 );
buf ( n12763 , n11715 );
nand ( n12764 , n12762 , n12763 );
buf ( n12765 , n12764 );
nand ( n12766 , n12761 , n12765 );
buf ( n12767 , n12766 );
not ( n12768 , n12767 );
buf ( n12769 , n12768 );
xor ( n12770 , n11414 , n11418 );
and ( n12771 , n12770 , n11432 );
and ( n12772 , n11414 , n11418 );
or ( n12773 , n12771 , n12772 );
buf ( n12774 , n12773 );
buf ( n12775 , n12774 );
not ( n12776 , n607 );
not ( n12777 , n10906 );
or ( n12778 , n12776 , n12777 );
nand ( n12779 , n11063 , n10882 );
nand ( n12780 , n12778 , n12779 );
buf ( n12781 , n12780 );
xor ( n12782 , n12775 , n12781 );
xor ( n12783 , n10998 , n11023 );
xor ( n12784 , n12783 , n11028 );
buf ( n12785 , n12784 );
buf ( n12786 , n12785 );
xor ( n12787 , n12782 , n12786 );
buf ( n12788 , n12787 );
buf ( n12789 , n12788 );
xor ( n12790 , n11086 , n11407 );
and ( n12791 , n12790 , n11435 );
and ( n12792 , n11086 , n11407 );
or ( n12793 , n12791 , n12792 );
buf ( n12794 , n12793 );
buf ( n12795 , n12794 );
nor ( n12796 , n12789 , n12795 );
buf ( n12797 , n12796 );
or ( n12798 , n12769 , n12797 );
buf ( n12799 , n12788 );
buf ( n12800 , n12794 );
nand ( n12801 , n12799 , n12800 );
buf ( n12802 , n12801 );
nand ( n12803 , n12798 , n12802 );
not ( n12804 , n12803 );
xor ( n12805 , n10914 , n11033 );
xor ( n12806 , n12805 , n11038 );
buf ( n12807 , n12806 );
buf ( n12808 , n12807 );
not ( n12809 , n12808 );
xor ( n12810 , n12775 , n12781 );
and ( n12811 , n12810 , n12786 );
and ( n12812 , n12775 , n12781 );
or ( n12813 , n12811 , n12812 );
buf ( n12814 , n12813 );
buf ( n12815 , n12814 );
not ( n12816 , n12815 );
buf ( n12817 , n12816 );
buf ( n12818 , n12817 );
nand ( n12819 , n12809 , n12818 );
buf ( n12820 , n12819 );
not ( n12821 , n12820 );
or ( n12822 , n12804 , n12821 );
buf ( n12823 , n12807 );
buf ( n12824 , n12814 );
nand ( n12825 , n12823 , n12824 );
buf ( n12826 , n12825 );
nand ( n12827 , n12822 , n12826 );
not ( n12828 , n12827 );
or ( n12829 , n11049 , n12828 );
nand ( n12830 , n10894 , n11042 );
buf ( n12831 , n12830 );
nand ( n12832 , n12829 , n12831 );
xor ( n12833 , n7633 , n7655 );
and ( n12834 , n12833 , n7781 );
and ( n12835 , n7633 , n7655 );
or ( n12836 , n12834 , n12835 );
buf ( n12837 , n12836 );
buf ( n12838 , n12837 );
buf ( n12839 , n5655 );
not ( n12840 , n12839 );
buf ( n12841 , n602 );
not ( n12842 , n12841 );
buf ( n12843 , n8554 );
not ( n12844 , n12843 );
or ( n12845 , n12842 , n12844 );
buf ( n12846 , n8557 );
buf ( n12847 , n2912 );
nand ( n12848 , n12846 , n12847 );
buf ( n12849 , n12848 );
buf ( n12850 , n12849 );
nand ( n12851 , n12845 , n12850 );
buf ( n12852 , n12851 );
buf ( n12853 , n12852 );
not ( n12854 , n12853 );
or ( n12855 , n12840 , n12854 );
buf ( n12856 , n7572 );
buf ( n12857 , n7619 );
nand ( n12858 , n12856 , n12857 );
buf ( n12859 , n12858 );
buf ( n12860 , n12859 );
nand ( n12861 , n12855 , n12860 );
buf ( n12862 , n12861 );
buf ( n12863 , n12862 );
xor ( n12864 , n12838 , n12863 );
xor ( n12865 , n7662 , n7687 );
and ( n12866 , n12865 , n7778 );
and ( n12867 , n7662 , n7687 );
or ( n12868 , n12866 , n12867 );
buf ( n12869 , n12868 );
buf ( n12870 , n12869 );
buf ( n12871 , n2915 );
not ( n12872 , n12871 );
buf ( n12873 , n600 );
not ( n12874 , n12873 );
buf ( n12875 , n7593 );
not ( n12876 , n12875 );
or ( n12877 , n12874 , n12876 );
buf ( n12878 , n7650 );
buf ( n12879 , n11008 );
nand ( n12880 , n12878 , n12879 );
buf ( n12881 , n12880 );
buf ( n12882 , n12881 );
nand ( n12883 , n12877 , n12882 );
buf ( n12884 , n12883 );
buf ( n12885 , n12884 );
not ( n12886 , n12885 );
or ( n12887 , n12872 , n12886 );
nand ( n12888 , n7652 , n5430 );
buf ( n12889 , n12888 );
nand ( n12890 , n12887 , n12889 );
buf ( n12891 , n12890 );
buf ( n12892 , n12891 );
xor ( n12893 , n12870 , n12892 );
xor ( n12894 , n7705 , n7742 );
and ( n12895 , n12894 , n7775 );
and ( n12896 , n7705 , n7742 );
or ( n12897 , n12895 , n12896 );
buf ( n12898 , n12897 );
buf ( n12899 , n12898 );
not ( n12900 , n5549 );
not ( n12901 , n598 );
not ( n12902 , n5376 );
or ( n12903 , n12901 , n12902 );
buf ( n12904 , n11364 );
buf ( n12905 , n818 );
nand ( n12906 , n12904 , n12905 );
buf ( n12907 , n12906 );
nand ( n12908 , n12903 , n12907 );
not ( n12909 , n12908 );
or ( n12910 , n12900 , n12909 );
nand ( n12911 , n7676 , n5631 );
nand ( n12912 , n12910 , n12911 );
buf ( n12913 , n12912 );
xor ( n12914 , n12899 , n12913 );
not ( n12915 , n2541 );
not ( n12916 , n5464 );
not ( n12917 , n2481 );
or ( n12918 , n12916 , n12917 );
nand ( n12919 , n594 , n5458 );
nand ( n12920 , n12918 , n12919 );
not ( n12921 , n12920 );
or ( n12922 , n12915 , n12921 );
buf ( n12923 , n7694 );
buf ( n12924 , n2592 );
nand ( n12925 , n12923 , n12924 );
buf ( n12926 , n12925 );
nand ( n12927 , n12922 , n12926 );
buf ( n12928 , n12927 );
buf ( n12929 , n2573 );
buf ( n12930 , n592 );
and ( n12931 , n12929 , n12930 );
buf ( n12932 , n12931 );
buf ( n12933 , n12932 );
buf ( n12934 , n2452 );
not ( n12935 , n12934 );
buf ( n12936 , n592 );
not ( n12937 , n5487 );
buf ( n12938 , n12937 );
xor ( n12939 , n12936 , n12938 );
buf ( n12940 , n12939 );
buf ( n12941 , n12940 );
not ( n12942 , n12941 );
or ( n12943 , n12935 , n12942 );
buf ( n12944 , n7726 );
buf ( n12945 , n2460 );
nand ( n12946 , n12944 , n12945 );
buf ( n12947 , n12946 );
buf ( n12948 , n12947 );
nand ( n12949 , n12943 , n12948 );
buf ( n12950 , n12949 );
buf ( n12951 , n12950 );
xor ( n12952 , n12933 , n12951 );
xor ( n12953 , n7710 , n7732 );
and ( n12954 , n12953 , n7739 );
and ( n12955 , n7710 , n7732 );
or ( n12956 , n12954 , n12955 );
buf ( n12957 , n12956 );
buf ( n12958 , n12957 );
xor ( n12959 , n12952 , n12958 );
buf ( n12960 , n12959 );
buf ( n12961 , n12960 );
xor ( n12962 , n12928 , n12961 );
buf ( n12963 , n825 );
not ( n12964 , n12963 );
buf ( n12965 , n596 );
not ( n12966 , n12965 );
buf ( n12967 , n8639 );
not ( n12968 , n12967 );
or ( n12969 , n12966 , n12968 );
buf ( n12970 , n5576 );
buf ( n12971 , n2371 );
nand ( n12972 , n12970 , n12971 );
buf ( n12973 , n12972 );
buf ( n12974 , n12973 );
nand ( n12975 , n12969 , n12974 );
buf ( n12976 , n12975 );
buf ( n12977 , n12976 );
not ( n12978 , n12977 );
or ( n12979 , n12964 , n12978 );
buf ( n12980 , n7764 );
buf ( n12981 , n2404 );
nand ( n12982 , n12980 , n12981 );
buf ( n12983 , n12982 );
buf ( n12984 , n12983 );
nand ( n12985 , n12979 , n12984 );
buf ( n12986 , n12985 );
buf ( n12987 , n12986 );
xor ( n12988 , n12962 , n12987 );
buf ( n12989 , n12988 );
buf ( n12990 , n12989 );
xor ( n12991 , n12914 , n12990 );
buf ( n12992 , n12991 );
buf ( n12993 , n12992 );
xor ( n12994 , n12893 , n12993 );
buf ( n12995 , n12994 );
buf ( n12996 , n12995 );
xor ( n12997 , n12864 , n12996 );
buf ( n12998 , n12997 );
buf ( n12999 , n12998 );
xor ( n13000 , n8797 , n9540 );
and ( n13001 , n13000 , n10889 );
and ( n13002 , n8797 , n9540 );
or ( n13003 , n13001 , n13002 );
buf ( n13004 , n13003 );
buf ( n13005 , n13004 );
xor ( n13006 , n12999 , n13005 );
xor ( n13007 , n5646 , n7626 );
and ( n13008 , n13007 , n7784 );
and ( n13009 , n5646 , n7626 );
or ( n13010 , n13008 , n13009 );
buf ( n13011 , n13010 );
buf ( n13012 , n13011 );
buf ( n13013 , n7790 );
not ( n13014 , n13013 );
and ( n13015 , n604 , n10861 );
not ( n13016 , n604 );
and ( n13017 , n13016 , n10858 );
or ( n13018 , n13015 , n13017 );
buf ( n13019 , n13018 );
not ( n13020 , n13019 );
or ( n13021 , n13014 , n13020 );
buf ( n13022 , n9529 );
buf ( n13023 , n8581 );
nand ( n13024 , n13022 , n13023 );
buf ( n13025 , n13024 );
buf ( n13026 , n13025 );
nand ( n13027 , n13021 , n13026 );
buf ( n13028 , n13027 );
buf ( n13029 , n13028 );
xor ( n13030 , n13012 , n13029 );
buf ( n13031 , n607 );
not ( n13032 , n13031 );
buf ( n13033 , n606 );
not ( n13034 , n13033 );
nor ( n13035 , n10803 , n10797 );
not ( n13036 , n13035 );
not ( n13037 , n9491 );
or ( n13038 , n13036 , n13037 );
not ( n13039 , n9679 );
not ( n13040 , n10175 );
and ( n13041 , n13039 , n13040 );
nor ( n13042 , n13041 , n10797 );
nand ( n13043 , n10176 , n9473 );
and ( n13044 , n13042 , n13043 );
nor ( n13045 , n13044 , n10795 );
nand ( n13046 , n13038 , n13045 );
xor ( n13047 , n10395 , n10396 );
and ( n13048 , n13047 , n10413 );
and ( n13049 , n10395 , n10396 );
or ( n13050 , n13048 , n13049 );
buf ( n13051 , n13050 );
buf ( n13052 , n13051 );
buf ( n13053 , n556 );
buf ( n13054 , n560 );
and ( n13055 , n13053 , n13054 );
buf ( n13056 , n13055 );
buf ( n13057 , n13056 );
buf ( n13058 , n10491 );
not ( n13059 , n13058 );
buf ( n13060 , n4836 );
not ( n13061 , n13060 );
or ( n13062 , n13059 , n13061 );
buf ( n13063 , n4840 );
buf ( n13064 , n550 );
buf ( n13065 , n564 );
xor ( n13066 , n13064 , n13065 );
buf ( n13067 , n13066 );
buf ( n13068 , n13067 );
nand ( n13069 , n13063 , n13068 );
buf ( n13070 , n13069 );
buf ( n13071 , n13070 );
nand ( n13072 , n13062 , n13071 );
buf ( n13073 , n13072 );
buf ( n13074 , n13073 );
xor ( n13075 , n13057 , n13074 );
buf ( n13076 , n10524 );
not ( n13077 , n13076 );
buf ( n13078 , n3429 );
not ( n13079 , n13078 );
or ( n13080 , n13077 , n13079 );
buf ( n13081 , n3439 );
xor ( n13082 , n568 , n546 );
buf ( n13083 , n13082 );
nand ( n13084 , n13081 , n13083 );
buf ( n13085 , n13084 );
buf ( n13086 , n13085 );
nand ( n13087 , n13080 , n13086 );
buf ( n13088 , n13087 );
buf ( n13089 , n13088 );
xor ( n13090 , n13075 , n13089 );
buf ( n13091 , n13090 );
buf ( n13092 , n13091 );
xor ( n13093 , n13052 , n13092 );
not ( n13094 , n10506 );
not ( n13095 , n9798 );
or ( n13096 , n13094 , n13095 );
buf ( n13097 , n5801 );
buf ( n13098 , n552 );
buf ( n13099 , n562 );
xor ( n13100 , n13098 , n13099 );
buf ( n13101 , n13100 );
buf ( n13102 , n13101 );
nand ( n13103 , n13097 , n13102 );
buf ( n13104 , n13103 );
nand ( n13105 , n13096 , n13104 );
not ( n13106 , n13105 );
buf ( n13107 , n10388 );
not ( n13108 , n13107 );
buf ( n13109 , n10380 );
not ( n13110 , n13109 );
or ( n13111 , n13108 , n13110 );
buf ( n13112 , n6595 );
buf ( n13113 , n554 );
buf ( n13114 , n560 );
xor ( n13115 , n13113 , n13114 );
buf ( n13116 , n13115 );
buf ( n13117 , n13116 );
nand ( n13118 , n13112 , n13117 );
buf ( n13119 , n13118 );
buf ( n13120 , n13119 );
nand ( n13121 , n13111 , n13120 );
buf ( n13122 , n13121 );
and ( n13123 , n13106 , n13122 );
not ( n13124 , n13106 );
not ( n13125 , n13122 );
and ( n13126 , n13124 , n13125 );
nor ( n13127 , n13123 , n13126 );
and ( n13128 , n13127 , n10412 );
not ( n13129 , n13127 );
and ( n13130 , n13129 , n10409 );
nor ( n13131 , n13128 , n13130 );
buf ( n13132 , n13131 );
xor ( n13133 , n13093 , n13132 );
buf ( n13134 , n13133 );
buf ( n13135 , n13134 );
xor ( n13136 , n10463 , n10537 );
and ( n13137 , n13136 , n10549 );
and ( n13138 , n10463 , n10537 );
or ( n13139 , n13137 , n13138 );
buf ( n13140 , n13139 );
buf ( n13141 , n13140 );
xor ( n13142 , n13135 , n13141 );
xor ( n13143 , n10473 , n10484 );
and ( n13144 , n13143 , n10534 );
and ( n13145 , n10473 , n10484 );
or ( n13146 , n13144 , n13145 );
buf ( n13147 , n13146 );
buf ( n13148 , n13147 );
xor ( n13149 , n10342 , n10356 );
and ( n13150 , n13149 , n10374 );
and ( n13151 , n10342 , n10356 );
or ( n13152 , n13150 , n13151 );
buf ( n13153 , n13152 );
buf ( n13154 , n13153 );
xor ( n13155 , n10496 , n10513 );
and ( n13156 , n13155 , n10531 );
and ( n13157 , n10496 , n10513 );
or ( n13158 , n13156 , n13157 );
buf ( n13159 , n13158 );
buf ( n13160 , n13159 );
xor ( n13161 , n13154 , n13160 );
buf ( n13162 , n10367 );
not ( n13163 , n13162 );
buf ( n13164 , n7872 );
not ( n13165 , n13164 );
or ( n13166 , n13163 , n13165 );
buf ( n13167 , n1979 );
buf ( n13168 , n544 );
buf ( n13169 , n570 );
xor ( n13170 , n13168 , n13169 );
buf ( n13171 , n13170 );
buf ( n13172 , n13171 );
nand ( n13173 , n13167 , n13172 );
buf ( n13174 , n13173 );
buf ( n13175 , n13174 );
nand ( n13176 , n13166 , n13175 );
buf ( n13177 , n13176 );
buf ( n13178 , n13177 );
or ( n13179 , n888 , n4434 );
nand ( n13180 , n13179 , n572 );
buf ( n13181 , n13180 );
xor ( n13182 , n13178 , n13181 );
buf ( n13183 , n10349 );
not ( n13184 , n13183 );
buf ( n13185 , n4380 );
not ( n13186 , n13185 );
or ( n13187 , n13184 , n13186 );
buf ( n13188 , n3743 );
buf ( n13189 , n548 );
buf ( n13190 , n566 );
xor ( n13191 , n13189 , n13190 );
buf ( n13192 , n13191 );
buf ( n13193 , n13192 );
nand ( n13194 , n13188 , n13193 );
buf ( n13195 , n13194 );
buf ( n13196 , n13195 );
nand ( n13197 , n13187 , n13196 );
buf ( n13198 , n13197 );
buf ( n13199 , n13198 );
xor ( n13200 , n13182 , n13199 );
buf ( n13201 , n13200 );
buf ( n13202 , n13201 );
xor ( n13203 , n13161 , n13202 );
buf ( n13204 , n13203 );
buf ( n13205 , n13204 );
xor ( n13206 , n13148 , n13205 );
xor ( n13207 , n10377 , n10416 );
and ( n13208 , n13207 , n10423 );
and ( n13209 , n10377 , n10416 );
or ( n13210 , n13208 , n13209 );
buf ( n13211 , n13210 );
buf ( n13212 , n13211 );
xor ( n13213 , n13206 , n13212 );
buf ( n13214 , n13213 );
buf ( n13215 , n13214 );
xor ( n13216 , n13142 , n13215 );
buf ( n13217 , n13216 );
buf ( n13218 , n13217 );
xor ( n13219 , n10572 , n10578 );
and ( n13220 , n13219 , n10771 );
and ( n13221 , n10572 , n10578 );
or ( n13222 , n13220 , n13221 );
buf ( n13223 , n13222 );
buf ( n13224 , n13223 );
xor ( n13225 , n13218 , n13224 );
xor ( n13226 , n10426 , n10447 );
and ( n13227 , n13226 , n10552 );
and ( n13228 , n10426 , n10447 );
or ( n13229 , n13227 , n13228 );
buf ( n13230 , n13229 );
buf ( n13231 , n13230 );
xor ( n13232 , n10673 , n10679 );
and ( n13233 , n13232 , n10768 );
and ( n13234 , n10673 , n10679 );
or ( n13235 , n13233 , n13234 );
buf ( n13236 , n13235 );
buf ( n13237 , n13236 );
xor ( n13238 , n13231 , n13237 );
xor ( n13239 , n10642 , n10658 );
and ( n13240 , n13239 , n10660 );
and ( n13241 , n10642 , n10658 );
or ( n13242 , n13240 , n13241 );
buf ( n13243 , n13242 );
buf ( n13244 , n13243 );
buf ( n13245 , n556 );
buf ( n13246 , n576 );
and ( n13247 , n13245 , n13246 );
buf ( n13248 , n13247 );
buf ( n13249 , n13248 );
not ( n13250 , n10714 );
not ( n13251 , n5059 );
not ( n13252 , n13251 );
or ( n13253 , n13250 , n13252 );
not ( n13254 , n550 );
not ( n13255 , n7240 );
or ( n13256 , n13254 , n13255 );
nand ( n13257 , n6311 , n580 );
nand ( n13258 , n13256 , n13257 );
nand ( n13259 , n4538 , n13258 );
nand ( n13260 , n13253 , n13259 );
buf ( n13261 , n13260 );
xor ( n13262 , n13249 , n13261 );
buf ( n13263 , n10745 );
not ( n13264 , n13263 );
buf ( n13265 , n3664 );
not ( n13266 , n13265 );
or ( n13267 , n13264 , n13266 );
buf ( n13268 , n2123 );
xor ( n13269 , n584 , n546 );
buf ( n13270 , n13269 );
nand ( n13271 , n13268 , n13270 );
buf ( n13272 , n13271 );
buf ( n13273 , n13272 );
nand ( n13274 , n13267 , n13273 );
buf ( n13275 , n13274 );
buf ( n13276 , n13275 );
xor ( n13277 , n13262 , n13276 );
buf ( n13278 , n13277 );
buf ( n13279 , n13278 );
xor ( n13280 , n13244 , n13279 );
buf ( n13281 , n10635 );
not ( n13282 , n13281 );
buf ( n13283 , n9946 );
not ( n13284 , n13283 );
or ( n13285 , n13282 , n13284 );
buf ( n13286 , n9952 );
buf ( n13287 , n554 );
buf ( n13288 , n576 );
xor ( n13289 , n13287 , n13288 );
buf ( n13290 , n13289 );
buf ( n13291 , n13290 );
nand ( n13292 , n13286 , n13291 );
buf ( n13293 , n13292 );
buf ( n13294 , n13293 );
nand ( n13295 , n13285 , n13294 );
buf ( n13296 , n13295 );
buf ( n13297 , n13296 );
buf ( n13298 , n10730 );
not ( n13299 , n13298 );
buf ( n13300 , n9049 );
not ( n13301 , n13300 );
or ( n13302 , n13299 , n13301 );
buf ( n13303 , n5997 );
xor ( n13304 , n578 , n552 );
buf ( n13305 , n13304 );
nand ( n13306 , n13303 , n13305 );
buf ( n13307 , n13306 );
buf ( n13308 , n13307 );
nand ( n13309 , n13302 , n13308 );
buf ( n13310 , n13309 );
buf ( n13311 , n13310 );
xor ( n13312 , n13297 , n13311 );
buf ( n13313 , n13312 );
buf ( n13314 , n13313 );
buf ( n13315 , n10654 );
xor ( n13316 , n13314 , n13315 );
buf ( n13317 , n13316 );
buf ( n13318 , n13317 );
xor ( n13319 , n13280 , n13318 );
buf ( n13320 , n13319 );
buf ( n13321 , n13320 );
xor ( n13322 , n10686 , n10758 );
and ( n13323 , n13322 , n10765 );
and ( n13324 , n10686 , n10758 );
or ( n13325 , n13323 , n13324 );
buf ( n13326 , n13325 );
buf ( n13327 , n13326 );
xor ( n13328 , n13321 , n13327 );
xor ( n13329 , n10692 , n10709 );
and ( n13330 , n13329 , n10755 );
and ( n13331 , n10692 , n10709 );
or ( n13332 , n13330 , n13331 );
buf ( n13333 , n13332 );
buf ( n13334 , n13333 );
buf ( n13335 , n10623 );
buf ( n13336 , n10603 );
or ( n13337 , n13335 , n13336 );
buf ( n13338 , n10595 );
nand ( n13339 , n13337 , n13338 );
buf ( n13340 , n13339 );
buf ( n13341 , n13340 );
buf ( n13342 , n10623 );
buf ( n13343 , n10603 );
nand ( n13344 , n13342 , n13343 );
buf ( n13345 , n13344 );
buf ( n13346 , n13345 );
nand ( n13347 , n13341 , n13346 );
buf ( n13348 , n13347 );
buf ( n13349 , n13348 );
xor ( n13350 , n10720 , n10737 );
and ( n13351 , n13350 , n10752 );
and ( n13352 , n10720 , n10737 );
or ( n13353 , n13351 , n13352 );
buf ( n13354 , n13353 );
buf ( n13355 , n13354 );
xor ( n13356 , n13349 , n13355 );
buf ( n13357 , n10617 );
not ( n13358 , n13357 );
buf ( n13359 , n4205 );
not ( n13360 , n13359 );
or ( n13361 , n13358 , n13360 );
buf ( n13362 , n4211 );
buf ( n13363 , n548 );
buf ( n13364 , n582 );
xor ( n13365 , n13363 , n13364 );
buf ( n13366 , n13365 );
buf ( n13367 , n13366 );
nand ( n13368 , n13362 , n13367 );
buf ( n13369 , n13368 );
buf ( n13370 , n13369 );
nand ( n13371 , n13361 , n13370 );
buf ( n13372 , n13371 );
buf ( n13373 , n10589 );
not ( n13374 , n13373 );
buf ( n13375 , n3616 );
not ( n13376 , n13375 );
or ( n13377 , n13374 , n13376 );
buf ( n13378 , n1036 );
buf ( n13379 , n544 );
buf ( n13380 , n586 );
xor ( n13381 , n13379 , n13380 );
buf ( n13382 , n13381 );
buf ( n13383 , n13382 );
nand ( n13384 , n13378 , n13383 );
buf ( n13385 , n13384 );
buf ( n13386 , n13385 );
nand ( n13387 , n13377 , n13386 );
buf ( n13388 , n13387 );
xor ( n13389 , n13372 , n13388 );
not ( n13390 , n1071 );
buf ( n13391 , n13390 );
not ( n13392 , n13391 );
buf ( n13393 , n3636 );
not ( n13394 , n13393 );
or ( n13395 , n13392 , n13394 );
buf ( n13396 , n588 );
nand ( n13397 , n13395 , n13396 );
buf ( n13398 , n13397 );
xor ( n13399 , n13389 , n13398 );
buf ( n13400 , n13399 );
xor ( n13401 , n13356 , n13400 );
buf ( n13402 , n13401 );
buf ( n13403 , n13402 );
xor ( n13404 , n13334 , n13403 );
xor ( n13405 , n10625 , n10663 );
and ( n13406 , n13405 , n10670 );
and ( n13407 , n10625 , n10663 );
or ( n13408 , n13406 , n13407 );
buf ( n13409 , n13408 );
buf ( n13410 , n13409 );
xor ( n13411 , n13404 , n13410 );
buf ( n13412 , n13411 );
buf ( n13413 , n13412 );
xor ( n13414 , n13328 , n13413 );
buf ( n13415 , n13414 );
buf ( n13416 , n13415 );
xor ( n13417 , n13238 , n13416 );
buf ( n13418 , n13417 );
buf ( n13419 , n13418 );
xor ( n13420 , n13225 , n13419 );
buf ( n13421 , n13420 );
xor ( n13422 , n10555 , n10561 );
and ( n13423 , n13422 , n10774 );
and ( n13424 , n10555 , n10561 );
or ( n13425 , n13423 , n13424 );
buf ( n13426 , n13425 );
nor ( n13427 , n13421 , n13426 );
buf ( n13428 , n13427 );
buf ( n13429 , n13421 );
buf ( n13430 , n13426 );
and ( n13431 , n13429 , n13430 );
buf ( n13432 , n13431 );
nor ( n13433 , n13428 , n13432 );
not ( n13434 , n13433 );
not ( n13435 , n13434 );
buf ( n13436 , n10333 );
not ( n13437 , n13436 );
buf ( n13438 , n10782 );
not ( n13439 , n13438 );
or ( n13440 , n13437 , n13439 );
buf ( n13441 , n10786 );
nand ( n13442 , n13440 , n13441 );
buf ( n13443 , n13442 );
buf ( n13444 , n13443 );
not ( n13445 , n13444 );
buf ( n13446 , n13445 );
and ( n13447 , n10782 , n10328 );
nand ( n13448 , n13447 , n9681 );
nand ( n13449 , n13446 , n13448 );
not ( n13450 , n13449 );
or ( n13451 , n13435 , n13450 );
nand ( n13452 , n13446 , n13448 , n13433 );
nand ( n13453 , n13451 , n13452 );
not ( n13454 , n13453 );
not ( n13455 , n10318 );
not ( n13456 , n10199 );
or ( n13457 , n13455 , n13456 );
nand ( n13458 , n13457 , n10320 );
xor ( n13459 , n10241 , n10245 );
and ( n13460 , n13459 , n10311 );
and ( n13461 , n10241 , n10245 );
or ( n13462 , n13460 , n13461 );
not ( n13463 , n13462 );
not ( n13464 , n8466 );
not ( n13465 , n10287 );
or ( n13466 , n13464 , n13465 );
not ( n13467 , n7178 );
and ( n13468 , n2981 , n6949 );
not ( n13469 , n2981 );
and ( n13470 , n13469 , n546 );
or ( n13471 , n13468 , n13470 );
nand ( n13472 , n13467 , n13471 );
nand ( n13473 , n13466 , n13472 );
not ( n13474 , n9409 );
not ( n13475 , n2944 );
nand ( n13476 , n13475 , n8477 );
nand ( n13477 , n5304 , n544 );
nand ( n13478 , n13476 , n13477 );
not ( n13479 , n13478 );
or ( n13480 , n13474 , n13479 );
nand ( n13481 , n10266 , n9417 );
nand ( n13482 , n13480 , n13481 );
xor ( n13483 , n13473 , n13482 );
not ( n13484 , n3068 );
not ( n13485 , n3073 );
not ( n13486 , n7147 );
or ( n13487 , n13485 , n13486 );
nand ( n13488 , n550 , n5247 );
nand ( n13489 , n13487 , n13488 );
not ( n13490 , n13489 );
or ( n13491 , n13484 , n13490 );
nand ( n13492 , n10230 , n5268 );
nand ( n13493 , n13491 , n13492 );
xor ( n13494 , n13483 , n13493 );
xor ( n13495 , n10282 , n10292 );
and ( n13496 , n13495 , n10303 );
and ( n13497 , n10282 , n10292 );
or ( n13498 , n13496 , n13497 );
xor ( n13499 , n13494 , n13498 );
not ( n13500 , n3118 );
not ( n13501 , n554 );
not ( n13502 , n8439 );
or ( n13503 , n13501 , n13502 );
not ( n13504 , n8439 );
nand ( n13505 , n13504 , n1681 );
nand ( n13506 , n13503 , n13505 );
not ( n13507 , n13506 );
or ( n13508 , n13500 , n13507 );
nand ( n13509 , n10237 , n2276 );
nand ( n13510 , n13508 , n13509 );
not ( n13511 , n6923 );
not ( n13512 , n548 );
not ( n13513 , n3168 );
or ( n13514 , n13512 , n13513 );
nand ( n13515 , n3167 , n5279 );
nand ( n13516 , n13514 , n13515 );
not ( n13517 , n13516 );
or ( n13518 , n13511 , n13517 );
nand ( n13519 , n10280 , n6939 );
nand ( n13520 , n13518 , n13519 );
xor ( n13521 , n13510 , n13520 );
not ( n13522 , n3064 );
not ( n13523 , n10297 );
or ( n13524 , n13522 , n13523 );
and ( n13525 , n552 , n7223 );
not ( n13526 , n552 );
and ( n13527 , n13526 , n7222 );
or ( n13528 , n13525 , n13527 );
nand ( n13529 , n13528 , n2265 );
nand ( n13530 , n13524 , n13529 );
xor ( n13531 , n13521 , n13530 );
xor ( n13532 , n13499 , n13531 );
and ( n13533 , n10270 , n10263 );
not ( n13534 , n1659 );
not ( n13535 , n10219 );
or ( n13536 , n13534 , n13535 );
nand ( n13537 , n13536 , n7199 );
not ( n13538 , n544 );
not ( n13539 , n10258 );
or ( n13540 , n13538 , n13539 );
nand ( n13541 , n13540 , n10256 );
xor ( n13542 , n13537 , n13541 );
not ( n13543 , n3049 );
nand ( n13544 , n13543 , n544 );
xor ( n13545 , n13542 , n13544 );
xor ( n13546 , n13533 , n13545 );
xor ( n13547 , n10223 , n10232 );
and ( n13548 , n13547 , n10239 );
and ( n13549 , n10223 , n10232 );
or ( n13550 , n13548 , n13549 );
xor ( n13551 , n13546 , n13550 );
xor ( n13552 , n10254 , n10271 );
and ( n13553 , n13552 , n10304 );
and ( n13554 , n10254 , n10271 );
or ( n13555 , n13553 , n13554 );
xor ( n13556 , n13551 , n13555 );
xor ( n13557 , n10204 , n10208 );
and ( n13558 , n13557 , n10240 );
and ( n13559 , n10204 , n10208 );
or ( n13560 , n13558 , n13559 );
xor ( n13561 , n13556 , n13560 );
xor ( n13562 , n13532 , n13561 );
xor ( n13563 , n10250 , n10305 );
and ( n13564 , n13563 , n10310 );
and ( n13565 , n10250 , n10305 );
or ( n13566 , n13564 , n13565 );
xor ( n13567 , n13562 , n13566 );
buf ( n13568 , n13567 );
not ( n13569 , n13568 );
or ( n13570 , n13463 , n13569 );
nor ( n13571 , n13567 , n13462 );
not ( n13572 , n13571 );
nand ( n13573 , n13570 , n13572 );
not ( n13574 , n13573 );
and ( n13575 , n13458 , n13574 );
not ( n13576 , n13458 );
and ( n13577 , n13576 , n13573 );
nor ( n13578 , n13575 , n13577 );
nor ( n13579 , n13454 , n13578 );
not ( n13580 , n13579 );
nand ( n13581 , n13578 , n13454 );
buf ( n13582 , n13581 );
nand ( n13583 , n13580 , n13582 );
and ( n13584 , n13046 , n13583 );
not ( n13585 , n13046 );
not ( n13586 , n13583 );
and ( n13587 , n13585 , n13586 );
nor ( n13588 , n13584 , n13587 );
not ( n13589 , n13588 );
buf ( n13590 , n13589 );
buf ( n13591 , n13590 );
buf ( n13592 , n13591 );
not ( n13593 , n13592 );
not ( n13594 , n10822 );
nor ( n13595 , n13594 , n10185 );
nand ( n13596 , n9517 , n13595 );
not ( n13597 , n13596 );
or ( n13598 , n13593 , n13597 );
not ( n13599 , n13596 );
not ( n13600 , n13592 );
nand ( n13601 , n13599 , n13600 );
nand ( n13602 , n13598 , n13601 );
buf ( n13603 , n13602 );
not ( n13604 , n13603 );
buf ( n13605 , n13604 );
buf ( n13606 , n13605 );
not ( n13607 , n13606 );
or ( n13608 , n13034 , n13607 );
buf ( n13609 , n13602 );
buf ( n13610 , n13609 );
buf ( n13611 , n13610 );
buf ( n13612 , n13611 );
buf ( n13613 , n10836 );
nand ( n13614 , n13612 , n13613 );
buf ( n13615 , n13614 );
buf ( n13616 , n13615 );
nand ( n13617 , n13608 , n13616 );
buf ( n13618 , n13617 );
buf ( n13619 , n13618 );
not ( n13620 , n13619 );
or ( n13621 , n13032 , n13620 );
buf ( n13622 , n10842 );
buf ( n13623 , n10882 );
nand ( n13624 , n13622 , n13623 );
buf ( n13625 , n13624 );
buf ( n13626 , n13625 );
nand ( n13627 , n13621 , n13626 );
buf ( n13628 , n13627 );
buf ( n13629 , n13628 );
xor ( n13630 , n13030 , n13629 );
buf ( n13631 , n13630 );
buf ( n13632 , n13631 );
xor ( n13633 , n13006 , n13632 );
buf ( n13634 , n13633 );
xor ( n13635 , n7787 , n8790 );
and ( n13636 , n13635 , n10892 );
and ( n13637 , n7787 , n8790 );
or ( n13638 , n13636 , n13637 );
buf ( n13639 , n13638 );
or ( n13640 , n13634 , n13639 );
buf ( n13641 , n13640 );
buf ( n13642 , n13634 );
buf ( n13643 , n13639 );
nand ( n13644 , n13642 , n13643 );
buf ( n13645 , n13644 );
buf ( n13646 , n13645 );
buf ( n13647 , n13646 );
buf ( n13648 , n13647 );
buf ( n13649 , n13648 );
nand ( n13650 , n13641 , n13649 );
buf ( n13651 , n13650 );
xnor ( n13652 , n12832 , n13651 );
buf ( n13653 , n13652 );
not ( n13654 , n12807 );
not ( n13655 , n12814 );
or ( n13656 , n13654 , n13655 );
nand ( n13657 , n13656 , n12820 );
buf ( n13658 , n12803 );
buf ( n13659 , n13658 );
buf ( n13660 , n13659 );
xnor ( n13661 , n13657 , n13660 );
buf ( n13662 , n13661 );
not ( n13663 , n5558 );
buf ( n13664 , n2314 );
buf ( n13665 , n4793 );
buf ( n13666 , n2343 );
buf ( n13667 , n2174 );
buf ( n13668 , n6394 );
buf ( n13669 , n6146 );
buf ( n13670 , n5146 );
buf ( n13671 , n4595 );
buf ( n13672 , n4001 );
buf ( n13673 , n8087 );
buf ( n13674 , n5939 );
buf ( n13675 , n1086 );
buf ( n13676 , n3516 );
buf ( n13677 , n2038 );
buf ( n13678 , n934 );
buf ( n13679 , n8114 );
buf ( n13680 , n1224 );
buf ( n13681 , n3684 );
buf ( n13682 , n6180 );
buf ( n13683 , n5945 );
buf ( n13684 , n4477 );
buf ( n13685 , n4314 );
buf ( n13686 , n10770 );
not ( n13687 , n10810 );
nand ( n13688 , n10792 , n10326 );
and ( n13689 , n13581 , n13688 );
not ( n13690 , n13689 );
or ( n13691 , n13687 , n13690 );
not ( n13692 , n13453 );
nand ( n13693 , n13692 , n13578 );
and ( n13694 , n13693 , n10795 );
nor ( n13695 , n13694 , n13579 );
nand ( n13696 , n13691 , n13695 );
not ( n13697 , n13696 );
nand ( n13698 , n10804 , n13689 );
not ( n13699 , n13698 );
nand ( n13700 , n13699 , n9548 );
nand ( n13701 , n13697 , n13700 );
nor ( n13702 , n13571 , n10317 );
not ( n13703 , n13702 );
not ( n13704 , n10199 );
or ( n13705 , n13703 , n13704 );
not ( n13706 , n13462 );
not ( n13707 , n13567 );
or ( n13708 , n13706 , n13707 );
nand ( n13709 , n13708 , n10319 );
nand ( n13710 , n13709 , n13572 );
nand ( n13711 , n13705 , n13710 );
buf ( n13712 , n13711 );
xor ( n13713 , n13510 , n13520 );
and ( n13714 , n13713 , n13530 );
and ( n13715 , n13510 , n13520 );
or ( n13716 , n13714 , n13715 );
xor ( n13717 , n13473 , n13482 );
and ( n13718 , n13717 , n13493 );
and ( n13719 , n13473 , n13482 );
or ( n13720 , n13718 , n13719 );
xor ( n13721 , n13716 , n13720 );
not ( n13722 , n2276 );
not ( n13723 , n13506 );
or ( n13724 , n13722 , n13723 );
buf ( n13725 , n9379 );
and ( n13726 , n554 , n13725 );
not ( n13727 , n554 );
not ( n13728 , n9379 );
and ( n13729 , n13727 , n13728 );
nor ( n13730 , n13726 , n13729 );
nand ( n13731 , n13730 , n3118 );
nand ( n13732 , n13724 , n13731 );
not ( n13733 , n6939 );
not ( n13734 , n13516 );
or ( n13735 , n13733 , n13734 );
and ( n13736 , n3264 , n548 );
not ( n13737 , n3264 );
and ( n13738 , n13737 , n5279 );
nor ( n13739 , n13736 , n13738 );
buf ( n13740 , n13739 );
nand ( n13741 , n13740 , n9327 );
nand ( n13742 , n13735 , n13741 );
xor ( n13743 , n13732 , n13742 );
not ( n13744 , n3064 );
not ( n13745 , n13528 );
or ( n13746 , n13744 , n13745 );
and ( n13747 , n552 , n7270 );
not ( n13748 , n552 );
and ( n13749 , n13748 , n7269 );
or ( n13750 , n13747 , n13749 );
nand ( n13751 , n13750 , n5299 );
nand ( n13752 , n13746 , n13751 );
xor ( n13753 , n13743 , n13752 );
xor ( n13754 , n13721 , n13753 );
xor ( n13755 , n13533 , n13545 );
and ( n13756 , n13755 , n13550 );
and ( n13757 , n13533 , n13545 );
or ( n13758 , n13756 , n13757 );
xor ( n13759 , n13537 , n13541 );
and ( n13760 , n13759 , n13544 );
and ( n13761 , n13537 , n13541 );
or ( n13762 , n13760 , n13761 );
not ( n13763 , n1595 );
not ( n13764 , n1658 );
or ( n13765 , n13763 , n13764 );
nand ( n13766 , n13765 , n556 );
and ( n13767 , n544 , n10265 );
xor ( n13768 , n13766 , n13767 );
not ( n13769 , n13544 );
xor ( n13770 , n13768 , n13769 );
xor ( n13771 , n13762 , n13770 );
not ( n13772 , n6945 );
not ( n13773 , n546 );
not ( n13774 , n7015 );
or ( n13775 , n13773 , n13774 );
nand ( n13776 , n6949 , n3036 );
nand ( n13777 , n13775 , n13776 );
not ( n13778 , n13777 );
or ( n13779 , n13772 , n13778 );
nand ( n13780 , n13471 , n9575 );
nand ( n13781 , n13779 , n13780 );
not ( n13782 , n9409 );
xor ( n13783 , n544 , n2251 );
not ( n13784 , n13783 );
or ( n13785 , n13782 , n13784 );
not ( n13786 , n13476 );
not ( n13787 , n13477 );
or ( n13788 , n13786 , n13787 );
nand ( n13789 , n13788 , n9417 );
nand ( n13790 , n13785 , n13789 );
xor ( n13791 , n13781 , n13790 );
not ( n13792 , n3068 );
not ( n13793 , n550 );
not ( n13794 , n7125 );
or ( n13795 , n13793 , n13794 );
nand ( n13796 , n7124 , n3073 );
nand ( n13797 , n13795 , n13796 );
not ( n13798 , n13797 );
or ( n13799 , n13792 , n13798 );
nand ( n13800 , n13489 , n5268 );
nand ( n13801 , n13799 , n13800 );
xor ( n13802 , n13791 , n13801 );
xor ( n13803 , n13771 , n13802 );
xor ( n13804 , n13758 , n13803 );
xor ( n13805 , n13494 , n13498 );
and ( n13806 , n13805 , n13531 );
and ( n13807 , n13494 , n13498 );
or ( n13808 , n13806 , n13807 );
xor ( n13809 , n13804 , n13808 );
xor ( n13810 , n13754 , n13809 );
xor ( n13811 , n13551 , n13555 );
and ( n13812 , n13811 , n13560 );
and ( n13813 , n13551 , n13555 );
or ( n13814 , n13812 , n13813 );
xor ( n13815 , n13810 , n13814 );
xor ( n13816 , n13532 , n13561 );
and ( n13817 , n13816 , n13566 );
and ( n13818 , n13532 , n13561 );
or ( n13819 , n13817 , n13818 );
nor ( n13820 , n13815 , n13819 );
buf ( n13821 , n13820 );
not ( n13822 , n13821 );
nand ( n13823 , n13815 , n13819 );
nand ( n13824 , n13822 , n13823 );
not ( n13825 , n13824 );
and ( n13826 , n13712 , n13825 );
not ( n13827 , n13712 );
and ( n13828 , n13827 , n13824 );
nor ( n13829 , n13826 , n13828 );
xor ( n13830 , n13052 , n13092 );
and ( n13831 , n13830 , n13132 );
and ( n13832 , n13052 , n13092 );
or ( n13833 , n13831 , n13832 );
buf ( n13834 , n13833 );
buf ( n13835 , n13834 );
xor ( n13836 , n13148 , n13205 );
and ( n13837 , n13836 , n13212 );
and ( n13838 , n13148 , n13205 );
or ( n13839 , n13837 , n13838 );
buf ( n13840 , n13839 );
buf ( n13841 , n13840 );
xor ( n13842 , n13835 , n13841 );
xor ( n13843 , n13154 , n13160 );
and ( n13844 , n13843 , n13202 );
and ( n13845 , n13154 , n13160 );
or ( n13846 , n13844 , n13845 );
buf ( n13847 , n13846 );
buf ( n13848 , n13847 );
buf ( n13849 , n13171 );
not ( n13850 , n13849 );
buf ( n13851 , n850 );
not ( n13852 , n13851 );
or ( n13853 , n13850 , n13852 );
buf ( n13854 , n570 );
buf ( n13855 , n856 );
nand ( n13856 , n13854 , n13855 );
buf ( n13857 , n13856 );
buf ( n13858 , n13857 );
nand ( n13859 , n13853 , n13858 );
buf ( n13860 , n13859 );
buf ( n13861 , n13860 );
not ( n13862 , n13861 );
buf ( n13863 , n13862 );
buf ( n13864 , n13863 );
xor ( n13865 , n13057 , n13074 );
and ( n13866 , n13865 , n13089 );
and ( n13867 , n13057 , n13074 );
or ( n13868 , n13866 , n13867 );
buf ( n13869 , n13868 );
buf ( n13870 , n13869 );
xor ( n13871 , n13864 , n13870 );
xor ( n13872 , n13178 , n13181 );
and ( n13873 , n13872 , n13199 );
and ( n13874 , n13178 , n13181 );
or ( n13875 , n13873 , n13874 );
buf ( n13876 , n13875 );
buf ( n13877 , n13876 );
xor ( n13878 , n13871 , n13877 );
buf ( n13879 , n13878 );
buf ( n13880 , n13879 );
xor ( n13881 , n13848 , n13880 );
buf ( n13882 , n13125 );
not ( n13883 , n13882 );
buf ( n13884 , n13106 );
not ( n13885 , n13884 );
or ( n13886 , n13883 , n13885 );
buf ( n13887 , n10409 );
nand ( n13888 , n13886 , n13887 );
buf ( n13889 , n13888 );
buf ( n13890 , n13889 );
buf ( n13891 , n13105 );
buf ( n13892 , n13122 );
nand ( n13893 , n13891 , n13892 );
buf ( n13894 , n13893 );
buf ( n13895 , n13894 );
nand ( n13896 , n13890 , n13895 );
buf ( n13897 , n13896 );
buf ( n13898 , n13897 );
buf ( n13899 , n555 );
buf ( n13900 , n560 );
and ( n13901 , n13899 , n13900 );
buf ( n13902 , n13901 );
buf ( n13903 , n13902 );
buf ( n13904 , n13116 );
not ( n13905 , n13904 );
buf ( n13906 , n10380 );
not ( n13907 , n13906 );
or ( n13908 , n13905 , n13907 );
buf ( n13909 , n6595 );
buf ( n13910 , n553 );
buf ( n13911 , n560 );
xor ( n13912 , n13910 , n13911 );
buf ( n13913 , n13912 );
buf ( n13914 , n13913 );
nand ( n13915 , n13909 , n13914 );
buf ( n13916 , n13915 );
buf ( n13917 , n13916 );
nand ( n13918 , n13908 , n13917 );
buf ( n13919 , n13918 );
buf ( n13920 , n13919 );
xor ( n13921 , n13903 , n13920 );
buf ( n13922 , n13192 );
not ( n13923 , n13922 );
buf ( n13924 , n4380 );
buf ( n13925 , n13924 );
buf ( n13926 , n13925 );
buf ( n13927 , n13926 );
not ( n13928 , n13927 );
or ( n13929 , n13923 , n13928 );
buf ( n13930 , n3743 );
buf ( n13931 , n547 );
buf ( n13932 , n566 );
xor ( n13933 , n13931 , n13932 );
buf ( n13934 , n13933 );
buf ( n13935 , n13934 );
nand ( n13936 , n13930 , n13935 );
buf ( n13937 , n13936 );
buf ( n13938 , n13937 );
nand ( n13939 , n13929 , n13938 );
buf ( n13940 , n13939 );
buf ( n13941 , n13940 );
xor ( n13942 , n13921 , n13941 );
buf ( n13943 , n13942 );
buf ( n13944 , n13943 );
xor ( n13945 , n13898 , n13944 );
buf ( n13946 , n13067 );
not ( n13947 , n13946 );
buf ( n13948 , n4836 );
not ( n13949 , n13948 );
or ( n13950 , n13947 , n13949 );
buf ( n13951 , n4840 );
buf ( n13952 , n549 );
buf ( n13953 , n564 );
xor ( n13954 , n13952 , n13953 );
buf ( n13955 , n13954 );
buf ( n13956 , n13955 );
nand ( n13957 , n13951 , n13956 );
buf ( n13958 , n13957 );
buf ( n13959 , n13958 );
nand ( n13960 , n13950 , n13959 );
buf ( n13961 , n13960 );
buf ( n13962 , n13961 );
buf ( n13963 , n13101 );
not ( n13964 , n13963 );
buf ( n13965 , n9798 );
not ( n13966 , n13965 );
or ( n13967 , n13964 , n13966 );
buf ( n13968 , n5801 );
buf ( n13969 , n551 );
buf ( n13970 , n562 );
xor ( n13971 , n13969 , n13970 );
buf ( n13972 , n13971 );
buf ( n13973 , n13972 );
nand ( n13974 , n13968 , n13973 );
buf ( n13975 , n13974 );
buf ( n13976 , n13975 );
nand ( n13977 , n13967 , n13976 );
buf ( n13978 , n13977 );
buf ( n13979 , n13978 );
xor ( n13980 , n13962 , n13979 );
buf ( n13981 , n13082 );
not ( n13982 , n13981 );
buf ( n13983 , n3429 );
not ( n13984 , n13983 );
or ( n13985 , n13982 , n13984 );
buf ( n13986 , n3439 );
buf ( n13987 , n545 );
buf ( n13988 , n568 );
xor ( n13989 , n13987 , n13988 );
buf ( n13990 , n13989 );
buf ( n13991 , n13990 );
nand ( n13992 , n13986 , n13991 );
buf ( n13993 , n13992 );
buf ( n13994 , n13993 );
nand ( n13995 , n13985 , n13994 );
buf ( n13996 , n13995 );
buf ( n13997 , n13996 );
xor ( n13998 , n13980 , n13997 );
buf ( n13999 , n13998 );
buf ( n14000 , n13999 );
xor ( n14001 , n13945 , n14000 );
buf ( n14002 , n14001 );
buf ( n14003 , n14002 );
xor ( n14004 , n13881 , n14003 );
buf ( n14005 , n14004 );
buf ( n14006 , n14005 );
xor ( n14007 , n13842 , n14006 );
buf ( n14008 , n14007 );
buf ( n14009 , n14008 );
xor ( n14010 , n13231 , n13237 );
and ( n14011 , n14010 , n13416 );
and ( n14012 , n13231 , n13237 );
or ( n14013 , n14011 , n14012 );
buf ( n14014 , n14013 );
buf ( n14015 , n14014 );
xor ( n14016 , n14009 , n14015 );
xor ( n14017 , n13135 , n13141 );
and ( n14018 , n14017 , n13215 );
and ( n14019 , n13135 , n13141 );
or ( n14020 , n14018 , n14019 );
buf ( n14021 , n14020 );
buf ( n14022 , n14021 );
xor ( n14023 , n13321 , n13327 );
and ( n14024 , n14023 , n13413 );
and ( n14025 , n13321 , n13327 );
or ( n14026 , n14024 , n14025 );
buf ( n14027 , n14026 );
buf ( n14028 , n14027 );
xor ( n14029 , n14022 , n14028 );
xor ( n14030 , n13244 , n13279 );
and ( n14031 , n14030 , n13318 );
and ( n14032 , n13244 , n13279 );
or ( n14033 , n14031 , n14032 );
buf ( n14034 , n14033 );
buf ( n14035 , n14034 );
buf ( n14036 , n13382 );
not ( n14037 , n14036 );
buf ( n14038 , n1177 );
not ( n14039 , n14038 );
or ( n14040 , n14037 , n14039 );
buf ( n14041 , n1036 );
buf ( n14042 , n586 );
nand ( n14043 , n14041 , n14042 );
buf ( n14044 , n14043 );
buf ( n14045 , n14044 );
nand ( n14046 , n14040 , n14045 );
buf ( n14047 , n14046 );
buf ( n14048 , n14047 );
not ( n14049 , n14048 );
buf ( n14050 , n14049 );
buf ( n14051 , n14050 );
xor ( n14052 , n13249 , n13261 );
and ( n14053 , n14052 , n13276 );
and ( n14054 , n13249 , n13261 );
or ( n14055 , n14053 , n14054 );
buf ( n14056 , n14055 );
buf ( n14057 , n14056 );
xor ( n14058 , n14051 , n14057 );
buf ( n14059 , n13398 );
buf ( n14060 , n13388 );
or ( n14061 , n14059 , n14060 );
buf ( n14062 , n13372 );
nand ( n14063 , n14061 , n14062 );
buf ( n14064 , n14063 );
buf ( n14065 , n14064 );
buf ( n14066 , n13398 );
buf ( n14067 , n13388 );
nand ( n14068 , n14066 , n14067 );
buf ( n14069 , n14068 );
buf ( n14070 , n14069 );
nand ( n14071 , n14065 , n14070 );
buf ( n14072 , n14071 );
buf ( n14073 , n14072 );
xor ( n14074 , n14058 , n14073 );
buf ( n14075 , n14074 );
buf ( n14076 , n14075 );
xor ( n14077 , n13349 , n13355 );
and ( n14078 , n14077 , n13400 );
and ( n14079 , n13349 , n13355 );
or ( n14080 , n14078 , n14079 );
buf ( n14081 , n14080 );
buf ( n14082 , n14081 );
xor ( n14083 , n14076 , n14082 );
buf ( n14084 , n13310 );
not ( n14085 , n14084 );
buf ( n14086 , n10654 );
not ( n14087 , n14086 );
or ( n14088 , n14085 , n14087 );
buf ( n14089 , n10654 );
buf ( n14090 , n13310 );
or ( n14091 , n14089 , n14090 );
buf ( n14092 , n13296 );
nand ( n14093 , n14091 , n14092 );
buf ( n14094 , n14093 );
buf ( n14095 , n14094 );
nand ( n14096 , n14088 , n14095 );
buf ( n14097 , n14096 );
buf ( n14098 , n14097 );
nand ( n14099 , n555 , n576 );
not ( n14100 , n9946 );
not ( n14101 , n13290 );
or ( n14102 , n14100 , n14101 );
buf ( n14103 , n6699 );
buf ( n14104 , n553 );
buf ( n14105 , n576 );
xor ( n14106 , n14104 , n14105 );
buf ( n14107 , n14106 );
buf ( n14108 , n14107 );
nand ( n14109 , n14103 , n14108 );
buf ( n14110 , n14109 );
nand ( n14111 , n14102 , n14110 );
xor ( n14112 , n14099 , n14111 );
not ( n14113 , n13366 );
not ( n14114 , n4205 );
or ( n14115 , n14113 , n14114 );
buf ( n14116 , n4211 );
buf ( n14117 , n547 );
buf ( n14118 , n582 );
xor ( n14119 , n14117 , n14118 );
buf ( n14120 , n14119 );
buf ( n14121 , n14120 );
nand ( n14122 , n14116 , n14121 );
buf ( n14123 , n14122 );
nand ( n14124 , n14115 , n14123 );
xnor ( n14125 , n14112 , n14124 );
buf ( n14126 , n14125 );
xor ( n14127 , n14098 , n14126 );
not ( n14128 , n13304 );
not ( n14129 , n9049 );
or ( n14130 , n14128 , n14129 );
buf ( n14131 , n5997 );
buf ( n14132 , n551 );
buf ( n14133 , n578 );
xor ( n14134 , n14132 , n14133 );
buf ( n14135 , n14134 );
buf ( n14136 , n14135 );
nand ( n14137 , n14131 , n14136 );
buf ( n14138 , n14137 );
nand ( n14139 , n14130 , n14138 );
buf ( n14140 , n13269 );
not ( n14141 , n14140 );
buf ( n14142 , n6758 );
not ( n14143 , n14142 );
or ( n14144 , n14141 , n14143 );
buf ( n14145 , n2123 );
xor ( n14146 , n584 , n545 );
buf ( n14147 , n14146 );
nand ( n14148 , n14145 , n14147 );
buf ( n14149 , n14148 );
buf ( n14150 , n14149 );
nand ( n14151 , n14144 , n14150 );
buf ( n14152 , n14151 );
xor ( n14153 , n14139 , n14152 );
buf ( n14154 , n549 );
buf ( n14155 , n580 );
xor ( n14156 , n14154 , n14155 );
buf ( n14157 , n14156 );
not ( n14158 , n14157 );
not ( n14159 , n5065 );
or ( n14160 , n14158 , n14159 );
nand ( n14161 , n13258 , n5060 );
nand ( n14162 , n14160 , n14161 );
xor ( n14163 , n14153 , n14162 );
buf ( n14164 , n14163 );
xor ( n14165 , n14127 , n14164 );
buf ( n14166 , n14165 );
buf ( n14167 , n14166 );
xor ( n14168 , n14083 , n14167 );
buf ( n14169 , n14168 );
buf ( n14170 , n14169 );
xor ( n14171 , n14035 , n14170 );
xor ( n14172 , n13334 , n13403 );
and ( n14173 , n14172 , n13410 );
and ( n14174 , n13334 , n13403 );
or ( n14175 , n14173 , n14174 );
buf ( n14176 , n14175 );
buf ( n14177 , n14176 );
xor ( n14178 , n14171 , n14177 );
buf ( n14179 , n14178 );
buf ( n14180 , n14179 );
xor ( n14181 , n14029 , n14180 );
buf ( n14182 , n14181 );
buf ( n14183 , n14182 );
xor ( n14184 , n14016 , n14183 );
buf ( n14185 , n14184 );
buf ( n14186 , n14185 );
not ( n14187 , n14186 );
buf ( n14188 , n14187 );
buf ( n14189 , n14188 );
xor ( n14190 , n13218 , n13224 );
and ( n14191 , n14190 , n13419 );
and ( n14192 , n13218 , n13224 );
or ( n14193 , n14191 , n14192 );
buf ( n14194 , n14193 );
buf ( n14195 , n14194 );
not ( n14196 , n14195 );
buf ( n14197 , n14196 );
buf ( n14198 , n14197 );
nand ( n14199 , n14189 , n14198 );
buf ( n14200 , n14199 );
buf ( n14201 , n14200 );
buf ( n14202 , n14201 );
buf ( n14203 , n14202 );
not ( n14204 , n14197 );
nand ( n14205 , n14204 , n14185 );
and ( n14206 , n14203 , n14205 );
not ( n14207 , n13427 );
not ( n14208 , n10167 );
nand ( n14209 , n14207 , n14208 , n10782 , n9247 );
buf ( n14210 , n14209 );
not ( n14211 , n14210 );
buf ( n14212 , n14211 );
not ( n14213 , n14212 );
not ( n14214 , n9301 );
or ( n14215 , n14213 , n14214 );
not ( n14216 , n10776 );
not ( n14217 , n10781 );
and ( n14218 , n14216 , n14217 );
nor ( n14219 , n14218 , n13427 );
not ( n14220 , n14219 );
not ( n14221 , n10333 );
or ( n14222 , n14220 , n14221 );
buf ( n14223 , n13427 );
not ( n14224 , n14223 );
buf ( n14225 , n10786 );
not ( n14226 , n14225 );
and ( n14227 , n14224 , n14226 );
buf ( n14228 , n13432 );
nor ( n14229 , n14227 , n14228 );
buf ( n14230 , n14229 );
nand ( n14231 , n14222 , n14230 );
buf ( n14232 , n14231 );
not ( n14233 , n14232 );
buf ( n14234 , n14233 );
nand ( n14235 , n14215 , n14234 );
and ( n14236 , n14206 , n14235 );
not ( n14237 , n14206 );
not ( n14238 , n14234 );
nor ( n14239 , n9298 , n14209 );
nor ( n14240 , n14238 , n14239 );
and ( n14241 , n14237 , n14240 );
nor ( n14242 , n14236 , n14241 );
not ( n14243 , n14242 );
nor ( n14244 , n13829 , n14243 );
not ( n14245 , n14244 );
not ( n14246 , n14242 );
nand ( n14247 , n14246 , n13829 );
buf ( n14248 , n14247 );
and ( n14249 , n14245 , n14248 );
and ( n14250 , n13701 , n14249 );
not ( n14251 , n13701 );
not ( n14252 , n14249 );
and ( n14253 , n14251 , n14252 );
nor ( n14254 , n14250 , n14253 );
nand ( n14255 , n14254 , n10819 , n13589 );
nand ( n14256 , n10184 , n9497 );
nor ( n14257 , n14255 , n14256 );
not ( n14258 , n13822 );
not ( n14259 , n13711 );
or ( n14260 , n14258 , n14259 );
buf ( n14261 , n13823 );
nand ( n14262 , n14260 , n14261 );
not ( n14263 , n9409 );
not ( n14264 , n544 );
not ( n14265 , n5186 );
or ( n14266 , n14264 , n14265 );
nand ( n14267 , n2981 , n8477 );
nand ( n14268 , n14266 , n14267 );
not ( n14269 , n14268 );
or ( n14270 , n14263 , n14269 );
nand ( n14271 , n13783 , n9417 );
nand ( n14272 , n14270 , n14271 );
buf ( n14273 , n1772 );
and ( n14274 , n14273 , n544 );
xor ( n14275 , n14272 , n14274 );
not ( n14276 , n5299 );
and ( n14277 , n552 , n8441 );
not ( n14278 , n552 );
and ( n14279 , n14278 , n10211 );
or ( n14280 , n14277 , n14279 );
not ( n14281 , n14280 );
or ( n14282 , n14276 , n14281 );
nand ( n14283 , n13750 , n3064 );
nand ( n14284 , n14282 , n14283 );
xor ( n14285 , n14275 , n14284 );
xor ( n14286 , n13732 , n13742 );
and ( n14287 , n14286 , n13752 );
and ( n14288 , n13732 , n13742 );
or ( n14289 , n14287 , n14288 );
xor ( n14290 , n14285 , n14289 );
not ( n14291 , n3212 );
not ( n14292 , n548 );
not ( n14293 , n5247 );
or ( n14294 , n14292 , n14293 );
nand ( n14295 , n5240 , n5221 );
not ( n14296 , n14295 );
not ( n14297 , n5245 );
or ( n14298 , n14296 , n14297 );
nand ( n14299 , n14298 , n5279 );
nand ( n14300 , n14294 , n14299 );
not ( n14301 , n14300 );
or ( n14302 , n14291 , n14301 );
nand ( n14303 , n13739 , n6939 );
nand ( n14304 , n14302 , n14303 );
not ( n14305 , n6945 );
not ( n14306 , n546 );
not ( n14307 , n5201 );
or ( n14308 , n14306 , n14307 );
nand ( n14309 , n3167 , n6949 );
nand ( n14310 , n14308 , n14309 );
not ( n14311 , n14310 );
or ( n14312 , n14305 , n14311 );
nand ( n14313 , n13777 , n9575 );
nand ( n14314 , n14312 , n14313 );
xor ( n14315 , n14304 , n14314 );
not ( n14316 , n3068 );
not ( n14317 , n550 );
not ( n14318 , n7223 );
or ( n14319 , n14317 , n14318 );
nand ( n14320 , n7222 , n3073 );
nand ( n14321 , n14319 , n14320 );
not ( n14322 , n14321 );
or ( n14323 , n14316 , n14322 );
nand ( n14324 , n13797 , n5268 );
nand ( n14325 , n14323 , n14324 );
xor ( n14326 , n14315 , n14325 );
xor ( n14327 , n14290 , n14326 );
xor ( n14328 , n13762 , n13770 );
and ( n14329 , n14328 , n13802 );
and ( n14330 , n13762 , n13770 );
or ( n14331 , n14329 , n14330 );
buf ( n14332 , n13730 );
and ( n14333 , n14332 , n6906 );
nor ( n14334 , n9618 , n1681 );
nor ( n14335 , n14333 , n14334 );
xor ( n14336 , n13766 , n13767 );
and ( n14337 , n14336 , n13769 );
and ( n14338 , n13766 , n13767 );
or ( n14339 , n14337 , n14338 );
xor ( n14340 , n14335 , n14339 );
xor ( n14341 , n13781 , n13790 );
and ( n14342 , n14341 , n13801 );
and ( n14343 , n13781 , n13790 );
or ( n14344 , n14342 , n14343 );
xor ( n14345 , n14340 , n14344 );
xor ( n14346 , n14331 , n14345 );
xor ( n14347 , n13716 , n13720 );
and ( n14348 , n14347 , n13753 );
and ( n14349 , n13716 , n13720 );
or ( n14350 , n14348 , n14349 );
xor ( n14351 , n14346 , n14350 );
xor ( n14352 , n14327 , n14351 );
xor ( n14353 , n13758 , n13803 );
and ( n14354 , n14353 , n13808 );
and ( n14355 , n13758 , n13803 );
or ( n14356 , n14354 , n14355 );
xor ( n14357 , n14352 , n14356 );
xor ( n14358 , n13754 , n13809 );
and ( n14359 , n14358 , n13814 );
and ( n14360 , n13754 , n13809 );
or ( n14361 , n14359 , n14360 );
nand ( n14362 , n14357 , n14361 );
not ( n14363 , n14357 );
not ( n14364 , n14361 );
nand ( n14365 , n14363 , n14364 );
nand ( n14366 , n14362 , n14365 );
not ( n14367 , n14366 );
and ( n14368 , n14262 , n14367 );
not ( n14369 , n14262 );
and ( n14370 , n14369 , n14366 );
nor ( n14371 , n14368 , n14370 );
buf ( n14372 , n9301 );
not ( n14373 , n14372 );
buf ( n14374 , n14203 );
not ( n14375 , n14374 );
buf ( n14376 , n14209 );
nor ( n14377 , n14375 , n14376 );
buf ( n14378 , n14377 );
buf ( n14379 , n14378 );
not ( n14380 , n14379 );
or ( n14381 , n14373 , n14380 );
not ( n14382 , n14203 );
not ( n14383 , n14231 );
or ( n14384 , n14382 , n14383 );
nand ( n14385 , n14384 , n14205 );
buf ( n14386 , n14385 );
not ( n14387 , n14386 );
buf ( n14388 , n14387 );
buf ( n14389 , n14388 );
nand ( n14390 , n14381 , n14389 );
buf ( n14391 , n14390 );
xor ( n14392 , n13903 , n13920 );
and ( n14393 , n14392 , n13941 );
and ( n14394 , n13903 , n13920 );
or ( n14395 , n14393 , n14394 );
buf ( n14396 , n14395 );
buf ( n14397 , n14396 );
buf ( n14398 , n13990 );
not ( n14399 , n14398 );
buf ( n14400 , n3429 );
not ( n14401 , n14400 );
or ( n14402 , n14399 , n14401 );
buf ( n14403 , n3439 );
buf ( n14404 , n544 );
buf ( n14405 , n568 );
xor ( n14406 , n14404 , n14405 );
buf ( n14407 , n14406 );
buf ( n14408 , n14407 );
nand ( n14409 , n14403 , n14408 );
buf ( n14410 , n14409 );
buf ( n14411 , n14410 );
nand ( n14412 , n14402 , n14411 );
buf ( n14413 , n14412 );
buf ( n14414 , n14413 );
buf ( n14415 , n13955 );
not ( n14416 , n14415 );
buf ( n14417 , n4836 );
buf ( n14418 , n14417 );
buf ( n14419 , n14418 );
buf ( n14420 , n14419 );
not ( n14421 , n14420 );
or ( n14422 , n14416 , n14421 );
buf ( n14423 , n4840 );
buf ( n14424 , n548 );
buf ( n14425 , n564 );
xor ( n14426 , n14424 , n14425 );
buf ( n14427 , n14426 );
buf ( n14428 , n14427 );
nand ( n14429 , n14423 , n14428 );
buf ( n14430 , n14429 );
buf ( n14431 , n14430 );
nand ( n14432 , n14422 , n14431 );
buf ( n14433 , n14432 );
buf ( n14434 , n14433 );
xor ( n14435 , n14414 , n14434 );
buf ( n14436 , n856 );
buf ( n14437 , n850 );
or ( n14438 , n14436 , n14437 );
buf ( n14439 , n570 );
nand ( n14440 , n14438 , n14439 );
buf ( n14441 , n14440 );
buf ( n14442 , n14441 );
xor ( n14443 , n14435 , n14442 );
buf ( n14444 , n14443 );
buf ( n14445 , n14444 );
xor ( n14446 , n14397 , n14445 );
buf ( n14447 , n13913 );
not ( n14448 , n14447 );
buf ( n14449 , n10380 );
not ( n14450 , n14449 );
or ( n14451 , n14448 , n14450 );
buf ( n14452 , n6595 );
buf ( n14453 , n552 );
buf ( n14454 , n560 );
xor ( n14455 , n14453 , n14454 );
buf ( n14456 , n14455 );
buf ( n14457 , n14456 );
nand ( n14458 , n14452 , n14457 );
buf ( n14459 , n14458 );
buf ( n14460 , n14459 );
nand ( n14461 , n14451 , n14460 );
buf ( n14462 , n14461 );
buf ( n14463 , n14462 );
buf ( n14464 , n13972 );
not ( n14465 , n14464 );
buf ( n14466 , n9798 );
not ( n14467 , n14466 );
or ( n14468 , n14465 , n14467 );
buf ( n14469 , n5801 );
buf ( n14470 , n550 );
buf ( n14471 , n562 );
xor ( n14472 , n14470 , n14471 );
buf ( n14473 , n14472 );
buf ( n14474 , n14473 );
nand ( n14475 , n14469 , n14474 );
buf ( n14476 , n14475 );
buf ( n14477 , n14476 );
nand ( n14478 , n14468 , n14477 );
buf ( n14479 , n14478 );
buf ( n14480 , n14479 );
xor ( n14481 , n14463 , n14480 );
buf ( n14482 , n13934 );
not ( n14483 , n14482 );
buf ( n14484 , n13926 );
not ( n14485 , n14484 );
or ( n14486 , n14483 , n14485 );
buf ( n14487 , n3743 );
buf ( n14488 , n546 );
buf ( n14489 , n566 );
xor ( n14490 , n14488 , n14489 );
buf ( n14491 , n14490 );
buf ( n14492 , n14491 );
nand ( n14493 , n14487 , n14492 );
buf ( n14494 , n14493 );
buf ( n14495 , n14494 );
nand ( n14496 , n14486 , n14495 );
buf ( n14497 , n14496 );
buf ( n14498 , n14497 );
xor ( n14499 , n14481 , n14498 );
buf ( n14500 , n14499 );
buf ( n14501 , n14500 );
xor ( n14502 , n14446 , n14501 );
buf ( n14503 , n14502 );
buf ( n14504 , n14503 );
xor ( n14505 , n13848 , n13880 );
and ( n14506 , n14505 , n14003 );
and ( n14507 , n13848 , n13880 );
or ( n14508 , n14506 , n14507 );
buf ( n14509 , n14508 );
buf ( n14510 , n14509 );
xor ( n14511 , n14504 , n14510 );
buf ( n14512 , n554 );
buf ( n14513 , n560 );
and ( n14514 , n14512 , n14513 );
buf ( n14515 , n14514 );
buf ( n14516 , n14515 );
buf ( n14517 , n13860 );
xor ( n14518 , n14516 , n14517 );
xor ( n14519 , n13962 , n13979 );
and ( n14520 , n14519 , n13997 );
and ( n14521 , n13962 , n13979 );
or ( n14522 , n14520 , n14521 );
buf ( n14523 , n14522 );
buf ( n14524 , n14523 );
xor ( n14525 , n14518 , n14524 );
buf ( n14526 , n14525 );
buf ( n14527 , n14526 );
xor ( n14528 , n13864 , n13870 );
and ( n14529 , n14528 , n13877 );
and ( n14530 , n13864 , n13870 );
or ( n14531 , n14529 , n14530 );
buf ( n14532 , n14531 );
buf ( n14533 , n14532 );
xor ( n14534 , n14527 , n14533 );
xor ( n14535 , n13898 , n13944 );
and ( n14536 , n14535 , n14000 );
and ( n14537 , n13898 , n13944 );
or ( n14538 , n14536 , n14537 );
buf ( n14539 , n14538 );
buf ( n14540 , n14539 );
xor ( n14541 , n14534 , n14540 );
buf ( n14542 , n14541 );
buf ( n14543 , n14542 );
xor ( n14544 , n14511 , n14543 );
buf ( n14545 , n14544 );
not ( n14546 , n14099 );
not ( n14547 , n14111 );
not ( n14548 , n14547 );
or ( n14549 , n14546 , n14548 );
nand ( n14550 , n14549 , n14124 );
not ( n14551 , n14099 );
nand ( n14552 , n14551 , n14111 );
nand ( n14553 , n14550 , n14552 );
buf ( n14554 , n14553 );
buf ( n14555 , n1036 );
buf ( n14556 , n3616 );
or ( n14557 , n14555 , n14556 );
buf ( n14558 , n586 );
nand ( n14559 , n14557 , n14558 );
buf ( n14560 , n14559 );
buf ( n14561 , n14560 );
buf ( n14562 , n14146 );
not ( n14563 , n14562 );
buf ( n14564 , n6758 );
not ( n14565 , n14564 );
or ( n14566 , n14563 , n14565 );
xor ( n14567 , n584 , n544 );
nand ( n14568 , n2123 , n14567 );
buf ( n14569 , n14568 );
nand ( n14570 , n14566 , n14569 );
buf ( n14571 , n14570 );
buf ( n14572 , n14571 );
xor ( n14573 , n14561 , n14572 );
buf ( n14574 , n14157 );
not ( n14575 , n14574 );
buf ( n14576 , n5060 );
not ( n14577 , n14576 );
or ( n14578 , n14575 , n14577 );
buf ( n14579 , n5065 );
buf ( n14580 , n548 );
buf ( n14581 , n580 );
xor ( n14582 , n14580 , n14581 );
buf ( n14583 , n14582 );
buf ( n14584 , n14583 );
nand ( n14585 , n14579 , n14584 );
buf ( n14586 , n14585 );
buf ( n14587 , n14586 );
nand ( n14588 , n14578 , n14587 );
buf ( n14589 , n14588 );
buf ( n14590 , n14589 );
xor ( n14591 , n14573 , n14590 );
buf ( n14592 , n14591 );
buf ( n14593 , n14592 );
xor ( n14594 , n14554 , n14593 );
buf ( n14595 , n14120 );
not ( n14596 , n14595 );
buf ( n14597 , n4205 );
not ( n14598 , n14597 );
or ( n14599 , n14596 , n14598 );
buf ( n14600 , n4211 );
buf ( n14601 , n546 );
buf ( n14602 , n582 );
xor ( n14603 , n14601 , n14602 );
buf ( n14604 , n14603 );
buf ( n14605 , n14604 );
nand ( n14606 , n14600 , n14605 );
buf ( n14607 , n14606 );
buf ( n14608 , n14607 );
nand ( n14609 , n14599 , n14608 );
buf ( n14610 , n14609 );
buf ( n14611 , n14610 );
buf ( n14612 , n14107 );
not ( n14613 , n14612 );
buf ( n14614 , n9946 );
buf ( n14615 , n14614 );
buf ( n14616 , n14615 );
buf ( n14617 , n14616 );
not ( n14618 , n14617 );
or ( n14619 , n14613 , n14618 );
buf ( n14620 , n9952 );
buf ( n14621 , n552 );
buf ( n14622 , n576 );
xor ( n14623 , n14621 , n14622 );
buf ( n14624 , n14623 );
buf ( n14625 , n14624 );
nand ( n14626 , n14620 , n14625 );
buf ( n14627 , n14626 );
buf ( n14628 , n14627 );
nand ( n14629 , n14619 , n14628 );
buf ( n14630 , n14629 );
buf ( n14631 , n14630 );
xor ( n14632 , n14611 , n14631 );
buf ( n14633 , n14135 );
not ( n14634 , n14633 );
buf ( n14635 , n6350 );
buf ( n14636 , n14635 );
buf ( n14637 , n14636 );
buf ( n14638 , n14637 );
not ( n14639 , n14638 );
or ( n14640 , n14634 , n14639 );
buf ( n14641 , n8294 );
buf ( n14642 , n550 );
buf ( n14643 , n578 );
xor ( n14644 , n14642 , n14643 );
buf ( n14645 , n14644 );
buf ( n14646 , n14645 );
nand ( n14647 , n14641 , n14646 );
buf ( n14648 , n14647 );
buf ( n14649 , n14648 );
nand ( n14650 , n14640 , n14649 );
buf ( n14651 , n14650 );
buf ( n14652 , n14651 );
xor ( n14653 , n14632 , n14652 );
buf ( n14654 , n14653 );
buf ( n14655 , n14654 );
xor ( n14656 , n14594 , n14655 );
buf ( n14657 , n14656 );
buf ( n14658 , n14657 );
buf ( n14659 , n554 );
buf ( n14660 , n576 );
nand ( n14661 , n14659 , n14660 );
buf ( n14662 , n14661 );
xor ( n14663 , n14047 , n14662 );
not ( n14664 , n14139 );
not ( n14665 , n14152 );
or ( n14666 , n14664 , n14665 );
or ( n14667 , n14139 , n14152 );
nand ( n14668 , n14667 , n14162 );
nand ( n14669 , n14666 , n14668 );
xnor ( n14670 , n14663 , n14669 );
buf ( n14671 , n14670 );
xor ( n14672 , n14051 , n14057 );
and ( n14673 , n14672 , n14073 );
and ( n14674 , n14051 , n14057 );
or ( n14675 , n14673 , n14674 );
buf ( n14676 , n14675 );
buf ( n14677 , n14676 );
xor ( n14678 , n14671 , n14677 );
xor ( n14679 , n14098 , n14126 );
and ( n14680 , n14679 , n14164 );
and ( n14681 , n14098 , n14126 );
or ( n14682 , n14680 , n14681 );
buf ( n14683 , n14682 );
buf ( n14684 , n14683 );
xor ( n14685 , n14678 , n14684 );
buf ( n14686 , n14685 );
buf ( n14687 , n14686 );
xor ( n14688 , n14658 , n14687 );
xor ( n14689 , n14076 , n14082 );
and ( n14690 , n14689 , n14167 );
and ( n14691 , n14076 , n14082 );
or ( n14692 , n14690 , n14691 );
buf ( n14693 , n14692 );
buf ( n14694 , n14693 );
xor ( n14695 , n14688 , n14694 );
buf ( n14696 , n14695 );
xor ( n14697 , n13835 , n13841 );
and ( n14698 , n14697 , n14006 );
and ( n14699 , n13835 , n13841 );
or ( n14700 , n14698 , n14699 );
buf ( n14701 , n14700 );
xor ( n14702 , n14696 , n14701 );
xor ( n14703 , n14035 , n14170 );
and ( n14704 , n14703 , n14177 );
and ( n14705 , n14035 , n14170 );
or ( n14706 , n14704 , n14705 );
buf ( n14707 , n14706 );
xor ( n14708 , n14702 , n14707 );
xor ( n14709 , n14545 , n14708 );
xor ( n14710 , n14022 , n14028 );
and ( n14711 , n14710 , n14180 );
and ( n14712 , n14022 , n14028 );
or ( n14713 , n14711 , n14712 );
buf ( n14714 , n14713 );
xor ( n14715 , n14709 , n14714 );
buf ( n14716 , n14715 );
not ( n14717 , n14716 );
buf ( n14718 , n14717 );
buf ( n14719 , n14718 );
xor ( n14720 , n14009 , n14015 );
and ( n14721 , n14720 , n14183 );
and ( n14722 , n14009 , n14015 );
or ( n14723 , n14721 , n14722 );
buf ( n14724 , n14723 );
buf ( n14725 , n14724 );
not ( n14726 , n14725 );
buf ( n14727 , n14726 );
buf ( n14728 , n14727 );
nand ( n14729 , n14719 , n14728 );
buf ( n14730 , n14729 );
buf ( n14731 , n14730 );
buf ( n14732 , n14731 );
buf ( n14733 , n14732 );
not ( n14734 , n14718 );
nand ( n14735 , n14734 , n14724 );
buf ( n14736 , n14735 );
buf ( n14737 , n14736 );
buf ( n14738 , n14737 );
nand ( n14739 , n14733 , n14738 );
and ( n14740 , n14391 , n14739 );
not ( n14741 , n14391 );
and ( n14742 , n14733 , n14738 );
and ( n14743 , n14741 , n14742 );
nor ( n14744 , n14740 , n14743 );
nand ( n14745 , n14371 , n14744 );
nand ( n14746 , n14745 , n14247 );
not ( n14747 , n14746 );
not ( n14748 , n14747 );
not ( n14749 , n14748 );
buf ( n14750 , n9295 );
not ( n14751 , n14750 );
buf ( n14752 , n14751 );
nand ( n14753 , n14752 , n14212 );
buf ( n14754 , n14730 );
buf ( n14755 , n14200 );
and ( n14756 , n14754 , n14755 );
buf ( n14757 , n14756 );
buf ( n14758 , n14757 );
buf ( n14759 , n14758 );
buf ( n14760 , n14759 );
not ( n14761 , n14760 );
or ( n14762 , n14753 , n14761 );
buf ( n14763 , n14757 );
not ( n14764 , n14763 );
buf ( n14765 , n14231 );
not ( n14766 , n14765 );
or ( n14767 , n14764 , n14766 );
nand ( n14768 , n14735 , n14205 );
buf ( n14769 , n14768 );
buf ( n14770 , n14733 );
nand ( n14771 , n14769 , n14770 );
buf ( n14772 , n14771 );
buf ( n14773 , n14772 );
nand ( n14774 , n14767 , n14773 );
buf ( n14775 , n14774 );
not ( n14776 , n14775 );
nand ( n14777 , n14762 , n14776 );
not ( n14778 , n14777 );
xor ( n14779 , n14545 , n14708 );
and ( n14780 , n14779 , n14714 );
and ( n14781 , n14545 , n14708 );
or ( n14782 , n14780 , n14781 );
buf ( n14783 , n553 );
buf ( n14784 , n560 );
and ( n14785 , n14783 , n14784 );
buf ( n14786 , n14785 );
buf ( n14787 , n14786 );
buf ( n14788 , n14427 );
not ( n14789 , n14788 );
buf ( n14790 , n14419 );
not ( n14791 , n14790 );
or ( n14792 , n14789 , n14791 );
buf ( n14793 , n4840 );
buf ( n14794 , n547 );
buf ( n14795 , n564 );
xor ( n14796 , n14794 , n14795 );
buf ( n14797 , n14796 );
buf ( n14798 , n14797 );
nand ( n14799 , n14793 , n14798 );
buf ( n14800 , n14799 );
buf ( n14801 , n14800 );
nand ( n14802 , n14792 , n14801 );
buf ( n14803 , n14802 );
buf ( n14804 , n14803 );
xor ( n14805 , n14787 , n14804 );
buf ( n14806 , n13926 );
buf ( n14807 , n14491 );
and ( n14808 , n14806 , n14807 );
buf ( n14809 , n3743 );
buf ( n14810 , n545 );
buf ( n14811 , n566 );
xor ( n14812 , n14810 , n14811 );
buf ( n14813 , n14812 );
buf ( n14814 , n14813 );
and ( n14815 , n14809 , n14814 );
nor ( n14816 , n14808 , n14815 );
buf ( n14817 , n14816 );
buf ( n14818 , n14817 );
xor ( n14819 , n14805 , n14818 );
buf ( n14820 , n14819 );
buf ( n14821 , n14820 );
xor ( n14822 , n14516 , n14517 );
and ( n14823 , n14822 , n14524 );
and ( n14824 , n14516 , n14517 );
or ( n14825 , n14823 , n14824 );
buf ( n14826 , n14825 );
buf ( n14827 , n14826 );
xor ( n14828 , n14821 , n14827 );
xor ( n14829 , n14397 , n14445 );
and ( n14830 , n14829 , n14501 );
and ( n14831 , n14397 , n14445 );
or ( n14832 , n14830 , n14831 );
buf ( n14833 , n14832 );
buf ( n14834 , n14833 );
xor ( n14835 , n14828 , n14834 );
buf ( n14836 , n14835 );
xor ( n14837 , n14463 , n14480 );
and ( n14838 , n14837 , n14498 );
and ( n14839 , n14463 , n14480 );
or ( n14840 , n14838 , n14839 );
buf ( n14841 , n14840 );
buf ( n14842 , n14841 );
buf ( n14843 , n14407 );
not ( n14844 , n14843 );
buf ( n14845 , n3429 );
not ( n14846 , n14845 );
or ( n14847 , n14844 , n14846 );
buf ( n14848 , n3439 );
buf ( n14849 , n568 );
nand ( n14850 , n14848 , n14849 );
buf ( n14851 , n14850 );
buf ( n14852 , n14851 );
nand ( n14853 , n14847 , n14852 );
buf ( n14854 , n14853 );
buf ( n14855 , n14473 );
not ( n14856 , n14855 );
buf ( n14857 , n9798 );
not ( n14858 , n14857 );
or ( n14859 , n14856 , n14858 );
buf ( n14860 , n5801 );
xor ( n14861 , n549 , n562 );
buf ( n14862 , n14861 );
nand ( n14863 , n14860 , n14862 );
buf ( n14864 , n14863 );
buf ( n14865 , n14864 );
nand ( n14866 , n14859 , n14865 );
buf ( n14867 , n14866 );
xor ( n14868 , n14854 , n14867 );
buf ( n14869 , n14456 );
not ( n14870 , n14869 );
buf ( n14871 , n10380 );
not ( n14872 , n14871 );
or ( n14873 , n14870 , n14872 );
buf ( n14874 , n6595 );
buf ( n14875 , n551 );
buf ( n14876 , n560 );
xor ( n14877 , n14875 , n14876 );
buf ( n14878 , n14877 );
buf ( n14879 , n14878 );
nand ( n14880 , n14874 , n14879 );
buf ( n14881 , n14880 );
buf ( n14882 , n14881 );
nand ( n14883 , n14873 , n14882 );
buf ( n14884 , n14883 );
xor ( n14885 , n14868 , n14884 );
buf ( n14886 , n14885 );
xor ( n14887 , n14842 , n14886 );
xor ( n14888 , n14414 , n14434 );
and ( n14889 , n14888 , n14442 );
and ( n14890 , n14414 , n14434 );
or ( n14891 , n14889 , n14890 );
buf ( n14892 , n14891 );
buf ( n14893 , n14892 );
xor ( n14894 , n14887 , n14893 );
buf ( n14895 , n14894 );
buf ( n14896 , n14895 );
xor ( n14897 , n14527 , n14533 );
and ( n14898 , n14897 , n14540 );
and ( n14899 , n14527 , n14533 );
or ( n14900 , n14898 , n14899 );
buf ( n14901 , n14900 );
nand ( n14902 , n14836 , n14896 , n14901 );
not ( n14903 , n14836 );
not ( n14904 , n14896 );
nand ( n14905 , n14903 , n14901 , n14904 );
not ( n14906 , n14901 );
nand ( n14907 , n14906 , n14836 , n14904 );
not ( n14908 , n14836 );
nand ( n14909 , n14908 , n14906 , n14896 );
nand ( n14910 , n14902 , n14905 , n14907 , n14909 );
xor ( n14911 , n14696 , n14701 );
and ( n14912 , n14911 , n14707 );
and ( n14913 , n14696 , n14701 );
or ( n14914 , n14912 , n14913 );
xor ( n14915 , n14910 , n14914 );
xor ( n14916 , n14658 , n14687 );
and ( n14917 , n14916 , n14694 );
and ( n14918 , n14658 , n14687 );
or ( n14919 , n14917 , n14918 );
buf ( n14920 , n14919 );
xor ( n14921 , n14611 , n14631 );
and ( n14922 , n14921 , n14652 );
and ( n14923 , n14611 , n14631 );
or ( n14924 , n14922 , n14923 );
buf ( n14925 , n14924 );
buf ( n14926 , n14925 );
xor ( n14927 , n14561 , n14572 );
and ( n14928 , n14927 , n14590 );
and ( n14929 , n14561 , n14572 );
or ( n14930 , n14928 , n14929 );
buf ( n14931 , n14930 );
buf ( n14932 , n14931 );
xor ( n14933 , n14926 , n14932 );
not ( n14934 , n14567 );
not ( n14935 , n3664 );
or ( n14936 , n14934 , n14935 );
nand ( n14937 , n4232 , n584 );
nand ( n14938 , n14936 , n14937 );
not ( n14939 , n14938 );
buf ( n14940 , n14624 );
not ( n14941 , n14940 );
buf ( n14942 , n14616 );
not ( n14943 , n14942 );
or ( n14944 , n14941 , n14943 );
buf ( n14945 , n9952 );
buf ( n14946 , n551 );
buf ( n14947 , n576 );
xor ( n14948 , n14946 , n14947 );
buf ( n14949 , n14948 );
buf ( n14950 , n14949 );
nand ( n14951 , n14945 , n14950 );
buf ( n14952 , n14951 );
buf ( n14953 , n14952 );
nand ( n14954 , n14944 , n14953 );
buf ( n14955 , n14954 );
not ( n14956 , n14955 );
not ( n14957 , n14956 );
or ( n14958 , n14939 , n14957 );
not ( n14959 , n14938 );
nand ( n14960 , n14959 , n14955 );
nand ( n14961 , n14958 , n14960 );
buf ( n14962 , n14645 );
not ( n14963 , n14962 );
buf ( n14964 , n14637 );
not ( n14965 , n14964 );
or ( n14966 , n14963 , n14965 );
buf ( n14967 , n8294 );
buf ( n14968 , n549 );
buf ( n14969 , n578 );
xor ( n14970 , n14968 , n14969 );
buf ( n14971 , n14970 );
buf ( n14972 , n14971 );
nand ( n14973 , n14967 , n14972 );
buf ( n14974 , n14973 );
buf ( n14975 , n14974 );
nand ( n14976 , n14966 , n14975 );
buf ( n14977 , n14976 );
and ( n14978 , n14961 , n14977 );
not ( n14979 , n14961 );
not ( n14980 , n14977 );
and ( n14981 , n14979 , n14980 );
nor ( n14982 , n14978 , n14981 );
buf ( n14983 , n14982 );
xor ( n14984 , n14933 , n14983 );
buf ( n14985 , n14984 );
buf ( n14986 , n14985 );
buf ( n14987 , n553 );
buf ( n14988 , n576 );
and ( n14989 , n14987 , n14988 );
buf ( n14990 , n14989 );
buf ( n14991 , n14990 );
buf ( n14992 , n14583 );
not ( n14993 , n14992 );
buf ( n14994 , n5060 );
not ( n14995 , n14994 );
or ( n14996 , n14993 , n14995 );
buf ( n14997 , n5065 );
buf ( n14998 , n547 );
buf ( n14999 , n580 );
xor ( n15000 , n14998 , n14999 );
buf ( n15001 , n15000 );
buf ( n15002 , n15001 );
nand ( n15003 , n14997 , n15002 );
buf ( n15004 , n15003 );
buf ( n15005 , n15004 );
nand ( n15006 , n14996 , n15005 );
buf ( n15007 , n15006 );
buf ( n15008 , n15007 );
xor ( n15009 , n14991 , n15008 );
not ( n15010 , n14604 );
not ( n15011 , n4205 );
or ( n15012 , n15010 , n15011 );
buf ( n15013 , n4211 );
buf ( n15014 , n545 );
buf ( n15015 , n582 );
xor ( n15016 , n15014 , n15015 );
buf ( n15017 , n15016 );
buf ( n15018 , n15017 );
nand ( n15019 , n15013 , n15018 );
buf ( n15020 , n15019 );
nand ( n15021 , n15012 , n15020 );
buf ( n15022 , n15021 );
not ( n15023 , n15022 );
buf ( n15024 , n15023 );
buf ( n15025 , n15024 );
xor ( n15026 , n15009 , n15025 );
buf ( n15027 , n15026 );
buf ( n15028 , n15027 );
buf ( n15029 , n14050 );
buf ( n15030 , n14662 );
nand ( n15031 , n15029 , n15030 );
buf ( n15032 , n15031 );
buf ( n15033 , n15032 );
not ( n15034 , n15033 );
buf ( n15035 , n14669 );
not ( n15036 , n15035 );
or ( n15037 , n15034 , n15036 );
buf ( n15038 , n14662 );
not ( n15039 , n15038 );
buf ( n15040 , n14047 );
nand ( n15041 , n15039 , n15040 );
buf ( n15042 , n15041 );
buf ( n15043 , n15042 );
nand ( n15044 , n15037 , n15043 );
buf ( n15045 , n15044 );
buf ( n15046 , n15045 );
xor ( n15047 , n15028 , n15046 );
xor ( n15048 , n14554 , n14593 );
and ( n15049 , n15048 , n14655 );
and ( n15050 , n14554 , n14593 );
or ( n15051 , n15049 , n15050 );
buf ( n15052 , n15051 );
buf ( n15053 , n15052 );
xor ( n15054 , n15047 , n15053 );
buf ( n15055 , n15054 );
buf ( n15056 , n15055 );
xor ( n15057 , n14986 , n15056 );
xor ( n15058 , n14671 , n14677 );
and ( n15059 , n15058 , n14684 );
and ( n15060 , n14671 , n14677 );
or ( n15061 , n15059 , n15060 );
buf ( n15062 , n15061 );
buf ( n15063 , n15062 );
xor ( n15064 , n15057 , n15063 );
buf ( n15065 , n15064 );
xor ( n15066 , n14920 , n15065 );
xor ( n15067 , n14504 , n14510 );
and ( n15068 , n15067 , n14543 );
and ( n15069 , n14504 , n14510 );
or ( n15070 , n15068 , n15069 );
buf ( n15071 , n15070 );
xor ( n15072 , n15066 , n15071 );
xor ( n15073 , n14915 , n15072 );
nor ( n15074 , n14782 , n15073 );
buf ( n15075 , n15074 );
not ( n15076 , n15075 );
buf ( n15077 , n15076 );
nand ( n15078 , n15073 , n14782 );
nand ( n15079 , n15077 , n15078 );
buf ( n15080 , n15079 );
not ( n15081 , n15080 );
and ( n15082 , n14778 , n15081 );
and ( n15083 , n14777 , n15080 );
nor ( n15084 , n15082 , n15083 );
nor ( n15085 , n14357 , n14361 );
nor ( n15086 , n13819 , n13815 );
nor ( n15087 , n15085 , n15086 );
nand ( n15088 , n15087 , n13702 );
not ( n15089 , n15088 );
not ( n15090 , n15089 );
not ( n15091 , n10199 );
or ( n15092 , n15090 , n15091 );
not ( n15093 , n13709 );
nor ( n15094 , n13567 , n13462 );
nor ( n15095 , n13820 , n15094 );
not ( n15096 , n15095 );
or ( n15097 , n15093 , n15096 );
nand ( n15098 , n13815 , n13819 );
and ( n15099 , n14362 , n15098 );
nand ( n15100 , n15097 , n15099 );
buf ( n15101 , n14365 );
nand ( n15102 , n15100 , n15101 );
nand ( n15103 , n15092 , n15102 );
buf ( n15104 , n15103 );
xor ( n15105 , n14304 , n14314 );
and ( n15106 , n15105 , n14325 );
and ( n15107 , n14304 , n14314 );
or ( n15108 , n15106 , n15107 );
not ( n15109 , n9618 );
not ( n15110 , n6905 );
or ( n15111 , n15109 , n15110 );
nand ( n15112 , n15111 , n554 );
not ( n15113 , n9417 );
not ( n15114 , n14268 );
or ( n15115 , n15113 , n15114 );
not ( n15116 , n544 );
not ( n15117 , n3036 );
not ( n15118 , n15117 );
or ( n15119 , n15116 , n15118 );
nand ( n15120 , n3036 , n8477 );
nand ( n15121 , n15119 , n15120 );
nand ( n15122 , n15121 , n9409 );
nand ( n15123 , n15115 , n15122 );
xor ( n15124 , n15112 , n15123 );
and ( n15125 , n544 , n2251 );
xor ( n15126 , n15124 , n15125 );
xor ( n15127 , n15108 , n15126 );
not ( n15128 , n3064 );
not ( n15129 , n14280 );
or ( n15130 , n15128 , n15129 );
and ( n15131 , n552 , n13728 );
not ( n15132 , n552 );
and ( n15133 , n15132 , n13725 );
or ( n15134 , n15131 , n15133 );
nand ( n15135 , n15134 , n5299 );
nand ( n15136 , n15130 , n15135 );
not ( n15137 , n9327 );
not ( n15138 , n548 );
not ( n15139 , n7125 );
or ( n15140 , n15138 , n15139 );
nand ( n15141 , n7124 , n5279 );
nand ( n15142 , n15140 , n15141 );
not ( n15143 , n15142 );
or ( n15144 , n15137 , n15143 );
nand ( n15145 , n14300 , n6939 );
nand ( n15146 , n15144 , n15145 );
xor ( n15147 , n15136 , n15146 );
not ( n15148 , n14335 );
xor ( n15149 , n15147 , n15148 );
xor ( n15150 , n15127 , n15149 );
xor ( n15151 , n14335 , n14339 );
and ( n15152 , n15151 , n14344 );
and ( n15153 , n14335 , n14339 );
or ( n15154 , n15152 , n15153 );
not ( n15155 , n9575 );
not ( n15156 , n14310 );
or ( n15157 , n15155 , n15156 );
and ( n15158 , n6918 , n6949 );
not ( n15159 , n6918 );
and ( n15160 , n15159 , n546 );
or ( n15161 , n15158 , n15160 );
nand ( n15162 , n15161 , n6945 );
nand ( n15163 , n15157 , n15162 );
not ( n15164 , n5268 );
not ( n15165 , n14321 );
or ( n15166 , n15164 , n15165 );
not ( n15167 , n550 );
not ( n15168 , n7270 );
or ( n15169 , n15167 , n15168 );
nand ( n15170 , n7269 , n3073 );
nand ( n15171 , n15169 , n15170 );
nand ( n15172 , n15171 , n3068 );
nand ( n15173 , n15166 , n15172 );
xor ( n15174 , n15163 , n15173 );
xor ( n15175 , n14272 , n14274 );
and ( n15176 , n15175 , n14284 );
and ( n15177 , n14272 , n14274 );
or ( n15178 , n15176 , n15177 );
xor ( n15179 , n15174 , n15178 );
xor ( n15180 , n15154 , n15179 );
xor ( n15181 , n14285 , n14289 );
and ( n15182 , n15181 , n14326 );
and ( n15183 , n14285 , n14289 );
or ( n15184 , n15182 , n15183 );
xor ( n15185 , n15180 , n15184 );
xor ( n15186 , n15150 , n15185 );
xor ( n15187 , n14331 , n14345 );
and ( n15188 , n15187 , n14350 );
and ( n15189 , n14331 , n14345 );
or ( n15190 , n15188 , n15189 );
xor ( n15191 , n15186 , n15190 );
buf ( n15192 , n15191 );
not ( n15193 , n15192 );
xor ( n15194 , n14327 , n14351 );
and ( n15195 , n15194 , n14356 );
and ( n15196 , n14327 , n14351 );
or ( n15197 , n15195 , n15196 );
not ( n15198 , n15197 );
nand ( n15199 , n15193 , n15198 );
nand ( n15200 , n15191 , n15197 );
nand ( n15201 , n15199 , n15200 );
not ( n15202 , n15201 );
and ( n15203 , n15104 , n15202 );
not ( n15204 , n15104 );
and ( n15205 , n15204 , n15201 );
nor ( n15206 , n15203 , n15205 );
nand ( n15207 , n15084 , n15206 );
and ( n15208 , n13699 , n15207 );
nand ( n15209 , n14749 , n15208 , n9492 );
and ( n15210 , n14747 , n15207 );
not ( n15211 , n13696 );
not ( n15212 , n15211 );
and ( n15213 , n15210 , n15212 );
not ( n15214 , n15207 );
not ( n15215 , n14745 );
not ( n15216 , n14244 );
or ( n15217 , n15215 , n15216 );
not ( n15218 , n14371 );
not ( n15219 , n14744 );
nand ( n15220 , n15218 , n15219 );
nand ( n15221 , n15217 , n15220 );
not ( n15222 , n15221 );
or ( n15223 , n15214 , n15222 );
nor ( n15224 , n15084 , n15206 );
not ( n15225 , n15224 );
nand ( n15226 , n15223 , n15225 );
nor ( n15227 , n15213 , n15226 );
nand ( n15228 , n15209 , n15227 );
not ( n15229 , n15199 );
not ( n15230 , n15103 );
or ( n15231 , n15229 , n15230 );
buf ( n15232 , n15200 );
nand ( n15233 , n15231 , n15232 );
xor ( n15234 , n15112 , n15123 );
and ( n15235 , n15234 , n15125 );
and ( n15236 , n15112 , n15123 );
or ( n15237 , n15235 , n15236 );
xor ( n15238 , n15136 , n15146 );
and ( n15239 , n15238 , n15148 );
and ( n15240 , n15136 , n15146 );
or ( n15241 , n15239 , n15240 );
xor ( n15242 , n15237 , n15241 );
not ( n15243 , n9409 );
xor ( n15244 , n544 , n6908 );
not ( n15245 , n15244 );
or ( n15246 , n15243 , n15245 );
nand ( n15247 , n15121 , n9417 );
nand ( n15248 , n15246 , n15247 );
not ( n15249 , n6939 );
not ( n15250 , n15142 );
or ( n15251 , n15249 , n15250 );
not ( n15252 , n548 );
not ( n15253 , n7223 );
or ( n15254 , n15252 , n15253 );
nand ( n15255 , n7222 , n5279 );
nand ( n15256 , n15254 , n15255 );
nand ( n15257 , n15256 , n9327 );
nand ( n15258 , n15251 , n15257 );
xor ( n15259 , n15248 , n15258 );
and ( n15260 , n15134 , n3064 );
nor ( n15261 , n15260 , n8408 );
xor ( n15262 , n15259 , n15261 );
xor ( n15263 , n15242 , n15262 );
not ( n15264 , n544 );
buf ( n15265 , n2982 );
nor ( n15266 , n15264 , n15265 );
not ( n15267 , n3068 );
not ( n15268 , n550 );
buf ( n15269 , n8440 );
not ( n15270 , n15269 );
not ( n15271 , n15270 );
or ( n15272 , n15268 , n15271 );
nand ( n15273 , n15269 , n3073 );
nand ( n15274 , n15272 , n15273 );
not ( n15275 , n15274 );
or ( n15276 , n15267 , n15275 );
nand ( n15277 , n15171 , n5268 );
nand ( n15278 , n15276 , n15277 );
xor ( n15279 , n15266 , n15278 );
not ( n15280 , n9575 );
not ( n15281 , n15161 );
or ( n15282 , n15280 , n15281 );
not ( n15283 , n546 );
not ( n15284 , n7150 );
or ( n15285 , n15283 , n15284 );
nand ( n15286 , n7147 , n6949 );
nand ( n15287 , n15285 , n15286 );
nand ( n15288 , n15287 , n7179 );
nand ( n15289 , n15282 , n15288 );
xor ( n15290 , n15279 , n15289 );
xor ( n15291 , n15163 , n15173 );
and ( n15292 , n15291 , n15178 );
and ( n15293 , n15163 , n15173 );
or ( n15294 , n15292 , n15293 );
xor ( n15295 , n15290 , n15294 );
xor ( n15296 , n15108 , n15126 );
and ( n15297 , n15296 , n15149 );
and ( n15298 , n15108 , n15126 );
or ( n15299 , n15297 , n15298 );
xor ( n15300 , n15295 , n15299 );
xor ( n15301 , n15263 , n15300 );
xor ( n15302 , n15154 , n15179 );
and ( n15303 , n15302 , n15184 );
and ( n15304 , n15154 , n15179 );
or ( n15305 , n15303 , n15304 );
xor ( n15306 , n15301 , n15305 );
xor ( n15307 , n15150 , n15185 );
and ( n15308 , n15307 , n15190 );
and ( n15309 , n15150 , n15185 );
or ( n15310 , n15308 , n15309 );
nor ( n15311 , n15306 , n15310 );
not ( n15312 , n15311 );
buf ( n15313 , n15306 );
nand ( n15314 , n15313 , n15310 );
nand ( n15315 , n15312 , n15314 );
not ( n15316 , n15315 );
and ( n15317 , n15233 , n15316 );
not ( n15318 , n15233 );
and ( n15319 , n15318 , n15315 );
nor ( n15320 , n15317 , n15319 );
buf ( n15321 , n14757 );
buf ( n15322 , n15077 );
and ( n15323 , n15321 , n15322 );
buf ( n15324 , n15323 );
not ( n15325 , n15324 );
not ( n15326 , n14212 );
not ( n15327 , n14752 );
or ( n15328 , n15326 , n15327 );
nand ( n15329 , n15328 , n14234 );
not ( n15330 , n15329 );
or ( n15331 , n15325 , n15330 );
nand ( n15332 , n14768 , n15077 , n14733 );
nand ( n15333 , n15332 , n15078 );
xor ( n15334 , n14910 , n14914 );
and ( n15335 , n15334 , n15072 );
and ( n15336 , n14910 , n14914 );
or ( n15337 , n15335 , n15336 );
buf ( n15338 , n15337 );
xor ( n15339 , n14842 , n14886 );
and ( n15340 , n15339 , n14893 );
and ( n15341 , n14842 , n14886 );
or ( n15342 , n15340 , n15341 );
buf ( n15343 , n15342 );
buf ( n15344 , n15343 );
buf ( n15345 , n14817 );
not ( n15346 , n15345 );
buf ( n15347 , n15346 );
buf ( n15348 , n15347 );
buf ( n15349 , n14884 );
not ( n15350 , n15349 );
buf ( n15351 , n14854 );
not ( n15352 , n15351 );
or ( n15353 , n15350 , n15352 );
buf ( n15354 , n14854 );
buf ( n15355 , n14884 );
or ( n15356 , n15354 , n15355 );
buf ( n15357 , n14867 );
nand ( n15358 , n15356 , n15357 );
buf ( n15359 , n15358 );
buf ( n15360 , n15359 );
nand ( n15361 , n15353 , n15360 );
buf ( n15362 , n15361 );
buf ( n15363 , n15362 );
xor ( n15364 , n15348 , n15363 );
buf ( n15365 , n552 );
buf ( n15366 , n560 );
and ( n15367 , n15365 , n15366 );
buf ( n15368 , n15367 );
buf ( n15369 , n15368 );
buf ( n15370 , n14878 );
not ( n15371 , n15370 );
buf ( n15372 , n10380 );
not ( n15373 , n15372 );
or ( n15374 , n15371 , n15373 );
buf ( n15375 , n6595 );
buf ( n15376 , n550 );
buf ( n15377 , n560 );
xor ( n15378 , n15376 , n15377 );
buf ( n15379 , n15378 );
buf ( n15380 , n15379 );
nand ( n15381 , n15375 , n15380 );
buf ( n15382 , n15381 );
buf ( n15383 , n15382 );
nand ( n15384 , n15374 , n15383 );
buf ( n15385 , n15384 );
buf ( n15386 , n15385 );
xor ( n15387 , n15369 , n15386 );
buf ( n15388 , n14797 );
not ( n15389 , n15388 );
buf ( n15390 , n14419 );
not ( n15391 , n15390 );
or ( n15392 , n15389 , n15391 );
buf ( n15393 , n4840 );
buf ( n15394 , n546 );
buf ( n15395 , n564 );
xor ( n15396 , n15394 , n15395 );
buf ( n15397 , n15396 );
buf ( n15398 , n15397 );
nand ( n15399 , n15393 , n15398 );
buf ( n15400 , n15399 );
buf ( n15401 , n15400 );
nand ( n15402 , n15392 , n15401 );
buf ( n15403 , n15402 );
buf ( n15404 , n15403 );
xor ( n15405 , n15387 , n15404 );
buf ( n15406 , n15405 );
buf ( n15407 , n15406 );
xor ( n15408 , n15364 , n15407 );
buf ( n15409 , n15408 );
buf ( n15410 , n14813 );
not ( n15411 , n15410 );
buf ( n15412 , n13926 );
not ( n15413 , n15412 );
or ( n15414 , n15411 , n15413 );
buf ( n15415 , n3743 );
buf ( n15416 , n544 );
buf ( n15417 , n566 );
xor ( n15418 , n15416 , n15417 );
buf ( n15419 , n15418 );
buf ( n15420 , n15419 );
nand ( n15421 , n15415 , n15420 );
buf ( n15422 , n15421 );
buf ( n15423 , n15422 );
nand ( n15424 , n15414 , n15423 );
buf ( n15425 , n15424 );
buf ( n15426 , n15425 );
not ( n15427 , n15426 );
buf ( n15428 , n3429 );
buf ( n15429 , n3439 );
or ( n15430 , n15428 , n15429 );
buf ( n15431 , n568 );
nand ( n15432 , n15430 , n15431 );
buf ( n15433 , n15432 );
buf ( n15434 , n15433 );
not ( n15435 , n15434 );
buf ( n15436 , n15435 );
buf ( n15437 , n15436 );
not ( n15438 , n15437 );
or ( n15439 , n15427 , n15438 );
buf ( n15440 , n15425 );
buf ( n15441 , n15436 );
or ( n15442 , n15440 , n15441 );
nand ( n15443 , n15439 , n15442 );
buf ( n15444 , n15443 );
buf ( n15445 , n15444 );
buf ( n15446 , n548 );
buf ( n15447 , n562 );
xor ( n15448 , n15446 , n15447 );
buf ( n15449 , n15448 );
and ( n15450 , n5801 , n15449 );
nand ( n15451 , n14861 , n9797 );
not ( n15452 , n15451 );
nor ( n15453 , n15450 , n15452 );
buf ( n15454 , n15453 );
and ( n15455 , n15445 , n15454 );
not ( n15456 , n15445 );
not ( n15457 , n15449 );
not ( n15458 , n5801 );
or ( n15459 , n15457 , n15458 );
nand ( n15460 , n15459 , n15451 );
buf ( n15461 , n15460 );
and ( n15462 , n15456 , n15461 );
nor ( n15463 , n15455 , n15462 );
buf ( n15464 , n15463 );
buf ( n15465 , n15464 );
not ( n15466 , n15465 );
buf ( n15467 , n15466 );
xor ( n15468 , n14787 , n14804 );
and ( n15469 , n15468 , n14818 );
and ( n15470 , n14787 , n14804 );
or ( n15471 , n15469 , n15470 );
buf ( n15472 , n15471 );
buf ( n15473 , n15472 );
not ( n15474 , n15473 );
buf ( n15475 , n15474 );
xor ( n15476 , n15467 , n15475 );
xnor ( n15477 , n15409 , n15476 );
buf ( n15478 , n15477 );
xor ( n15479 , n15344 , n15478 );
xor ( n15480 , n14821 , n14827 );
and ( n15481 , n15480 , n14834 );
and ( n15482 , n14821 , n14827 );
or ( n15483 , n15481 , n15482 );
buf ( n15484 , n15483 );
buf ( n15485 , n15484 );
xor ( n15486 , n15479 , n15485 );
buf ( n15487 , n15486 );
buf ( n15488 , n15487 );
xor ( n15489 , n14920 , n15065 );
and ( n15490 , n15489 , n15071 );
and ( n15491 , n14920 , n15065 );
or ( n15492 , n15490 , n15491 );
buf ( n15493 , n15492 );
xor ( n15494 , n15488 , n15493 );
xor ( n15495 , n14986 , n15056 );
and ( n15496 , n15495 , n15063 );
and ( n15497 , n14986 , n15056 );
or ( n15498 , n15496 , n15497 );
buf ( n15499 , n15498 );
buf ( n15500 , n15499 );
xor ( n15501 , n14926 , n14932 );
and ( n15502 , n15501 , n14983 );
and ( n15503 , n14926 , n14932 );
or ( n15504 , n15502 , n15503 );
buf ( n15505 , n15504 );
buf ( n15506 , n15505 );
xor ( n15507 , n15028 , n15046 );
and ( n15508 , n15507 , n15053 );
and ( n15509 , n15028 , n15046 );
or ( n15510 , n15508 , n15509 );
buf ( n15511 , n15510 );
buf ( n15512 , n15511 );
xor ( n15513 , n15506 , n15512 );
xor ( n15514 , n14991 , n15008 );
and ( n15515 , n15514 , n15025 );
and ( n15516 , n14991 , n15008 );
or ( n15517 , n15515 , n15516 );
buf ( n15518 , n15517 );
buf ( n15519 , n15518 );
buf ( n15520 , n15017 );
not ( n15521 , n15520 );
buf ( n15522 , n4205 );
not ( n15523 , n15522 );
or ( n15524 , n15521 , n15523 );
buf ( n15525 , n4211 );
buf ( n15526 , n544 );
buf ( n15527 , n582 );
xor ( n15528 , n15526 , n15527 );
buf ( n15529 , n15528 );
buf ( n15530 , n15529 );
nand ( n15531 , n15525 , n15530 );
buf ( n15532 , n15531 );
buf ( n15533 , n15532 );
nand ( n15534 , n15524 , n15533 );
buf ( n15535 , n15534 );
buf ( n15536 , n15535 );
not ( n15537 , n2132 );
not ( n15538 , n3663 );
or ( n15539 , n15537 , n15538 );
nand ( n15540 , n15539 , n584 );
buf ( n15541 , n15540 );
xor ( n15542 , n15536 , n15541 );
buf ( n15543 , n14971 );
not ( n15544 , n15543 );
buf ( n15545 , n14637 );
not ( n15546 , n15545 );
or ( n15547 , n15544 , n15546 );
buf ( n15548 , n8294 );
buf ( n15549 , n548 );
buf ( n15550 , n578 );
xor ( n15551 , n15549 , n15550 );
buf ( n15552 , n15551 );
buf ( n15553 , n15552 );
nand ( n15554 , n15548 , n15553 );
buf ( n15555 , n15554 );
buf ( n15556 , n15555 );
nand ( n15557 , n15547 , n15556 );
buf ( n15558 , n15557 );
buf ( n15559 , n15558 );
xor ( n15560 , n15542 , n15559 );
buf ( n15561 , n15560 );
buf ( n15562 , n15561 );
xor ( n15563 , n15519 , n15562 );
not ( n15564 , n14955 );
not ( n15565 , n14977 );
or ( n15566 , n15564 , n15565 );
or ( n15567 , n14977 , n14955 );
nand ( n15568 , n15567 , n14938 );
nand ( n15569 , n15566 , n15568 );
xor ( n15570 , n15021 , n15569 );
buf ( n15571 , n552 );
buf ( n15572 , n576 );
and ( n15573 , n15571 , n15572 );
buf ( n15574 , n15573 );
buf ( n15575 , n15001 );
not ( n15576 , n15575 );
buf ( n15577 , n5060 );
not ( n15578 , n15577 );
or ( n15579 , n15576 , n15578 );
buf ( n15580 , n5065 );
buf ( n15581 , n546 );
buf ( n15582 , n580 );
xor ( n15583 , n15581 , n15582 );
buf ( n15584 , n15583 );
buf ( n15585 , n15584 );
nand ( n15586 , n15580 , n15585 );
buf ( n15587 , n15586 );
buf ( n15588 , n15587 );
nand ( n15589 , n15579 , n15588 );
buf ( n15590 , n15589 );
xor ( n15591 , n15574 , n15590 );
buf ( n15592 , n14949 );
not ( n15593 , n15592 );
buf ( n15594 , n14616 );
not ( n15595 , n15594 );
or ( n15596 , n15593 , n15595 );
buf ( n15597 , n9952 );
buf ( n15598 , n550 );
buf ( n15599 , n576 );
xor ( n15600 , n15598 , n15599 );
buf ( n15601 , n15600 );
buf ( n15602 , n15601 );
nand ( n15603 , n15597 , n15602 );
buf ( n15604 , n15603 );
buf ( n15605 , n15604 );
nand ( n15606 , n15596 , n15605 );
buf ( n15607 , n15606 );
xor ( n15608 , n15591 , n15607 );
xor ( n15609 , n15570 , n15608 );
buf ( n15610 , n15609 );
xor ( n15611 , n15563 , n15610 );
buf ( n15612 , n15611 );
buf ( n15613 , n15612 );
xor ( n15614 , n15513 , n15613 );
buf ( n15615 , n15614 );
buf ( n15616 , n15615 );
xor ( n15617 , n15500 , n15616 );
not ( n15618 , n14836 );
not ( n15619 , n14896 );
or ( n15620 , n15618 , n15619 );
or ( n15621 , n14836 , n14896 );
nand ( n15622 , n15621 , n14901 );
nand ( n15623 , n15620 , n15622 );
buf ( n15624 , n15623 );
xor ( n15625 , n15617 , n15624 );
buf ( n15626 , n15625 );
buf ( n15627 , n15626 );
xor ( n15628 , n15494 , n15627 );
buf ( n15629 , n15628 );
buf ( n15630 , n15629 );
nor ( n15631 , n15338 , n15630 );
buf ( n15632 , n15631 );
buf ( n15633 , n15632 );
buf ( n15634 , n15633 );
buf ( n15635 , n15634 );
not ( n15636 , n15635 );
buf ( n15637 , n15337 );
buf ( n15638 , n15629 );
nand ( n15639 , n15637 , n15638 );
buf ( n15640 , n15639 );
nand ( n15641 , n15636 , n15640 );
nor ( n15642 , n15333 , n15641 );
nand ( n15643 , n15331 , n15642 );
nand ( n15644 , n15333 , n15641 );
nand ( n15645 , n15329 , n15641 , n15324 );
nand ( n15646 , n15643 , n15644 , n15645 );
not ( n15647 , n15646 );
nand ( n15648 , n15320 , n15647 );
buf ( n15649 , n15648 );
not ( n15650 , n15320 );
buf ( n15651 , n15646 );
nand ( n15652 , n15650 , n15651 );
buf ( n15653 , n15652 );
nand ( n15654 , n15649 , n15653 );
xnor ( n15655 , n15228 , n15654 );
nand ( n15656 , n15225 , n15207 );
not ( n15657 , n15656 );
not ( n15658 , n15657 );
nand ( n15659 , n13696 , n14747 );
not ( n15660 , n15221 );
nand ( n15661 , n14747 , n13699 , n9492 );
nand ( n15662 , n15659 , n15660 , n15661 );
not ( n15663 , n15662 );
not ( n15664 , n15663 );
or ( n15665 , n15658 , n15664 );
nand ( n15666 , n15662 , n15656 );
nand ( n15667 , n15665 , n15666 );
and ( n15668 , n15220 , n14745 );
not ( n15669 , n13045 );
and ( n15670 , n14247 , n13582 );
and ( n15671 , n15669 , n15670 );
not ( n15672 , n13579 );
not ( n15673 , n14247 );
or ( n15674 , n15672 , n15673 );
nand ( n15675 , n15674 , n14245 );
nor ( n15676 , n15671 , n15675 );
nand ( n15677 , n14248 , n9492 , n13699 );
nand ( n15678 , n15676 , n15677 );
xor ( n15679 , n15668 , n15678 );
buf ( n15680 , n15679 );
nand ( n15681 , n14257 , n15655 , n15667 , n15680 );
not ( n15682 , n15681 );
not ( n15683 , n15682 );
not ( n15684 , n15683 );
not ( n15685 , n15084 );
not ( n15686 , n15206 );
or ( n15687 , n15685 , n15686 );
nand ( n15688 , n15687 , n15648 );
not ( n15689 , n15688 );
and ( n15690 , n14745 , n14247 );
nand ( n15691 , n15689 , n15690 );
not ( n15692 , n15691 );
buf ( n15693 , n15692 );
not ( n15694 , n15211 );
and ( n15695 , n15693 , n15694 );
not ( n15696 , n15689 );
not ( n15697 , n15221 );
or ( n15698 , n15696 , n15697 );
not ( n15699 , n15224 );
not ( n15700 , n15648 );
or ( n15701 , n15699 , n15700 );
nand ( n15702 , n15701 , n15652 );
not ( n15703 , n15702 );
nand ( n15704 , n15698 , n15703 );
nor ( n15705 , n15695 , n15704 );
nand ( n15706 , n15692 , n13699 );
not ( n15707 , n15706 );
nand ( n15708 , n9492 , n15707 );
nand ( n15709 , n15705 , n15708 );
not ( n15710 , n15709 );
xor ( n15711 , n15263 , n15300 );
and ( n15712 , n15711 , n15305 );
and ( n15713 , n15263 , n15300 );
or ( n15714 , n15712 , n15713 );
not ( n15715 , n15714 );
xor ( n15716 , n15237 , n15241 );
and ( n15717 , n15716 , n15262 );
and ( n15718 , n15237 , n15241 );
or ( n15719 , n15717 , n15718 );
not ( n15720 , n9587 );
not ( n15721 , n7028 );
or ( n15722 , n15720 , n15721 );
nand ( n15723 , n15722 , n552 );
not ( n15724 , n544 );
nor ( n15725 , n15724 , n15117 );
xor ( n15726 , n15723 , n15725 );
not ( n15727 , n5268 );
not ( n15728 , n15274 );
or ( n15729 , n15727 , n15728 );
not ( n15730 , n3073 );
buf ( n15731 , n13725 );
not ( n15732 , n15731 );
or ( n15733 , n15730 , n15732 );
not ( n15734 , n15731 );
nand ( n15735 , n15734 , n550 );
nand ( n15736 , n15733 , n15735 );
nand ( n15737 , n15736 , n3068 );
nand ( n15738 , n15729 , n15737 );
xor ( n15739 , n15726 , n15738 );
not ( n15740 , n9575 );
not ( n15741 , n15287 );
or ( n15742 , n15740 , n15741 );
not ( n15743 , n546 );
not ( n15744 , n7125 );
or ( n15745 , n15743 , n15744 );
nand ( n15746 , n7124 , n6949 );
nand ( n15747 , n15745 , n15746 );
nand ( n15748 , n15747 , n7179 );
nand ( n15749 , n15742 , n15748 );
not ( n15750 , n9417 );
not ( n15751 , n15244 );
or ( n15752 , n15750 , n15751 );
xor ( n15753 , n544 , n6918 );
nand ( n15754 , n15753 , n9409 );
nand ( n15755 , n15752 , n15754 );
xor ( n15756 , n15749 , n15755 );
not ( n15757 , n6939 );
not ( n15758 , n15256 );
or ( n15759 , n15757 , n15758 );
not ( n15760 , n548 );
not ( n15761 , n7270 );
or ( n15762 , n15760 , n15761 );
not ( n15763 , n7270 );
nand ( n15764 , n15763 , n5279 );
nand ( n15765 , n15762 , n15764 );
nand ( n15766 , n15765 , n9327 );
nand ( n15767 , n15759 , n15766 );
xor ( n15768 , n15756 , n15767 );
xor ( n15769 , n15739 , n15768 );
not ( n15770 , n15261 );
xor ( n15771 , n15266 , n15278 );
and ( n15772 , n15771 , n15289 );
and ( n15773 , n15266 , n15278 );
or ( n15774 , n15772 , n15773 );
xor ( n15775 , n15770 , n15774 );
xor ( n15776 , n15248 , n15258 );
and ( n15777 , n15776 , n15261 );
and ( n15778 , n15248 , n15258 );
or ( n15779 , n15777 , n15778 );
xor ( n15780 , n15775 , n15779 );
xor ( n15781 , n15769 , n15780 );
xor ( n15782 , n15719 , n15781 );
xor ( n15783 , n15290 , n15294 );
and ( n15784 , n15783 , n15299 );
and ( n15785 , n15290 , n15294 );
or ( n15786 , n15784 , n15785 );
xor ( n15787 , n15782 , n15786 );
not ( n15788 , n15787 );
nand ( n15789 , n15715 , n15788 );
nand ( n15790 , n15714 , n15787 );
nand ( n15791 , n15789 , n15790 );
not ( n15792 , n15791 );
not ( n15793 , n15792 );
nor ( n15794 , n15192 , n15197 );
nor ( n15795 , n15311 , n15794 );
not ( n15796 , n15795 );
not ( n15797 , n15104 );
or ( n15798 , n15796 , n15797 );
nor ( n15799 , n15310 , n15306 );
or ( n15800 , n15799 , n15200 );
nand ( n15801 , n15306 , n15310 );
nand ( n15802 , n15800 , n15801 );
buf ( n15803 , n15802 );
not ( n15804 , n15803 );
nand ( n15805 , n15798 , n15804 );
not ( n15806 , n15805 );
not ( n15807 , n15806 );
or ( n15808 , n15793 , n15807 );
nand ( n15809 , n15805 , n15791 );
nand ( n15810 , n15808 , n15809 );
xor ( n15811 , n15344 , n15478 );
and ( n15812 , n15811 , n15485 );
and ( n15813 , n15344 , n15478 );
or ( n15814 , n15812 , n15813 );
buf ( n15815 , n15814 );
buf ( n15816 , n15815 );
xor ( n15817 , n15021 , n15569 );
and ( n15818 , n15817 , n15608 );
and ( n15819 , n15021 , n15569 );
or ( n15820 , n15818 , n15819 );
buf ( n15821 , n15820 );
buf ( n15822 , n551 );
buf ( n15823 , n576 );
and ( n15824 , n15822 , n15823 );
buf ( n15825 , n15824 );
not ( n15826 , n15529 );
not ( n15827 , n4205 );
or ( n15828 , n15826 , n15827 );
buf ( n15829 , n4211 );
buf ( n15830 , n582 );
nand ( n15831 , n15829 , n15830 );
buf ( n15832 , n15831 );
nand ( n15833 , n15828 , n15832 );
xor ( n15834 , n15825 , n15833 );
buf ( n15835 , n15601 );
not ( n15836 , n15835 );
buf ( n15837 , n14616 );
not ( n15838 , n15837 );
or ( n15839 , n15836 , n15838 );
buf ( n15840 , n9952 );
buf ( n15841 , n549 );
buf ( n15842 , n576 );
xor ( n15843 , n15841 , n15842 );
buf ( n15844 , n15843 );
buf ( n15845 , n15844 );
nand ( n15846 , n15840 , n15845 );
buf ( n15847 , n15846 );
buf ( n15848 , n15847 );
nand ( n15849 , n15839 , n15848 );
buf ( n15850 , n15849 );
xor ( n15851 , n15834 , n15850 );
buf ( n15852 , n15851 );
xor ( n15853 , n15536 , n15541 );
and ( n15854 , n15853 , n15559 );
and ( n15855 , n15536 , n15541 );
or ( n15856 , n15854 , n15855 );
buf ( n15857 , n15856 );
buf ( n15858 , n15857 );
xor ( n15859 , n15852 , n15858 );
buf ( n15860 , n15552 );
not ( n15861 , n15860 );
buf ( n15862 , n14637 );
not ( n15863 , n15862 );
or ( n15864 , n15861 , n15863 );
buf ( n15865 , n8294 );
buf ( n15866 , n547 );
buf ( n15867 , n578 );
xor ( n15868 , n15866 , n15867 );
buf ( n15869 , n15868 );
buf ( n15870 , n15869 );
nand ( n15871 , n15865 , n15870 );
buf ( n15872 , n15871 );
buf ( n15873 , n15872 );
nand ( n15874 , n15864 , n15873 );
buf ( n15875 , n15874 );
buf ( n15876 , n15875 );
buf ( n15877 , n15584 );
not ( n15878 , n15877 );
buf ( n15879 , n5060 );
buf ( n15880 , n15879 );
buf ( n15881 , n15880 );
buf ( n15882 , n15881 );
not ( n15883 , n15882 );
or ( n15884 , n15878 , n15883 );
buf ( n15885 , n5065 );
buf ( n15886 , n545 );
buf ( n15887 , n580 );
xor ( n15888 , n15886 , n15887 );
buf ( n15889 , n15888 );
buf ( n15890 , n15889 );
nand ( n15891 , n15885 , n15890 );
buf ( n15892 , n15891 );
buf ( n15893 , n15892 );
nand ( n15894 , n15884 , n15893 );
buf ( n15895 , n15894 );
buf ( n15896 , n15895 );
not ( n15897 , n15896 );
buf ( n15898 , n15897 );
buf ( n15899 , n15898 );
xor ( n15900 , n15876 , n15899 );
not ( n15901 , n15607 );
or ( n15902 , n15590 , n15574 );
not ( n15903 , n15902 );
or ( n15904 , n15901 , n15903 );
nand ( n15905 , n15590 , n15574 );
nand ( n15906 , n15904 , n15905 );
buf ( n15907 , n15906 );
xor ( n15908 , n15900 , n15907 );
buf ( n15909 , n15908 );
buf ( n15910 , n15909 );
xor ( n15911 , n15859 , n15910 );
buf ( n15912 , n15911 );
buf ( n15913 , n15912 );
xor ( n15914 , n15821 , n15913 );
xor ( n15915 , n15519 , n15562 );
and ( n15916 , n15915 , n15610 );
and ( n15917 , n15519 , n15562 );
or ( n15918 , n15916 , n15917 );
buf ( n15919 , n15918 );
buf ( n15920 , n15919 );
xor ( n15921 , n15914 , n15920 );
buf ( n15922 , n15921 );
buf ( n15923 , n15922 );
not ( n15924 , n15923 );
buf ( n15925 , n15924 );
buf ( n15926 , n15925 );
and ( n15927 , n15816 , n15926 );
not ( n15928 , n15816 );
buf ( n15929 , n15922 );
and ( n15930 , n15928 , n15929 );
nor ( n15931 , n15927 , n15930 );
buf ( n15932 , n15931 );
xor ( n15933 , n15506 , n15512 );
and ( n15934 , n15933 , n15613 );
and ( n15935 , n15506 , n15512 );
or ( n15936 , n15934 , n15935 );
buf ( n15937 , n15936 );
not ( n15938 , n15937 );
and ( n15939 , n15932 , n15938 );
not ( n15940 , n15932 );
and ( n15941 , n15940 , n15937 );
nor ( n15942 , n15939 , n15941 );
not ( n15943 , n15942 );
not ( n15944 , n15943 );
xor ( n15945 , n15500 , n15616 );
and ( n15946 , n15945 , n15624 );
and ( n15947 , n15500 , n15616 );
or ( n15948 , n15946 , n15947 );
buf ( n15949 , n15948 );
xor ( n15950 , n15348 , n15363 );
and ( n15951 , n15950 , n15407 );
and ( n15952 , n15348 , n15363 );
or ( n15953 , n15951 , n15952 );
buf ( n15954 , n15953 );
buf ( n15955 , n15954 );
buf ( n15956 , n551 );
buf ( n15957 , n560 );
and ( n15958 , n15956 , n15957 );
buf ( n15959 , n15958 );
buf ( n15960 , n15959 );
buf ( n15961 , n15379 );
not ( n15962 , n15961 );
buf ( n15963 , n10380 );
not ( n15964 , n15963 );
or ( n15965 , n15962 , n15964 );
buf ( n15966 , n6595 );
buf ( n15967 , n549 );
buf ( n15968 , n560 );
xor ( n15969 , n15967 , n15968 );
buf ( n15970 , n15969 );
buf ( n15971 , n15970 );
nand ( n15972 , n15966 , n15971 );
buf ( n15973 , n15972 );
buf ( n15974 , n15973 );
nand ( n15975 , n15965 , n15974 );
buf ( n15976 , n15975 );
buf ( n15977 , n15976 );
xor ( n15978 , n15960 , n15977 );
buf ( n15979 , n15419 );
not ( n15980 , n15979 );
buf ( n15981 , n13926 );
not ( n15982 , n15981 );
or ( n15983 , n15980 , n15982 );
buf ( n15984 , n3743 );
buf ( n15985 , n566 );
nand ( n15986 , n15984 , n15985 );
buf ( n15987 , n15986 );
buf ( n15988 , n15987 );
nand ( n15989 , n15983 , n15988 );
buf ( n15990 , n15989 );
buf ( n15991 , n15990 );
xor ( n15992 , n15978 , n15991 );
buf ( n15993 , n15992 );
buf ( n15994 , n15993 );
buf ( n15995 , n15453 );
not ( n15996 , n15995 );
buf ( n15997 , n15436 );
not ( n15998 , n15997 );
or ( n15999 , n15996 , n15998 );
buf ( n16000 , n15425 );
nand ( n16001 , n15999 , n16000 );
buf ( n16002 , n16001 );
buf ( n16003 , n16002 );
buf ( n16004 , n15433 );
buf ( n16005 , n15460 );
nand ( n16006 , n16004 , n16005 );
buf ( n16007 , n16006 );
buf ( n16008 , n16007 );
nand ( n16009 , n16003 , n16008 );
buf ( n16010 , n16009 );
buf ( n16011 , n16010 );
xor ( n16012 , n15994 , n16011 );
buf ( n16013 , n15449 );
not ( n16014 , n16013 );
buf ( n16015 , n9798 );
not ( n16016 , n16015 );
or ( n16017 , n16014 , n16016 );
buf ( n16018 , n5801 );
buf ( n16019 , n547 );
buf ( n16020 , n562 );
xor ( n16021 , n16019 , n16020 );
buf ( n16022 , n16021 );
buf ( n16023 , n16022 );
nand ( n16024 , n16018 , n16023 );
buf ( n16025 , n16024 );
buf ( n16026 , n16025 );
nand ( n16027 , n16017 , n16026 );
buf ( n16028 , n16027 );
buf ( n16029 , n16028 );
buf ( n16030 , n15397 );
not ( n16031 , n16030 );
buf ( n16032 , n14419 );
not ( n16033 , n16032 );
or ( n16034 , n16031 , n16033 );
buf ( n16035 , n4840 );
buf ( n16036 , n545 );
buf ( n16037 , n564 );
xor ( n16038 , n16036 , n16037 );
buf ( n16039 , n16038 );
buf ( n16040 , n16039 );
nand ( n16041 , n16035 , n16040 );
buf ( n16042 , n16041 );
buf ( n16043 , n16042 );
nand ( n16044 , n16034 , n16043 );
buf ( n16045 , n16044 );
buf ( n16046 , n16045 );
not ( n16047 , n16046 );
buf ( n16048 , n16047 );
buf ( n16049 , n16048 );
xor ( n16050 , n16029 , n16049 );
xor ( n16051 , n15369 , n15386 );
and ( n16052 , n16051 , n15404 );
and ( n16053 , n15369 , n15386 );
or ( n16054 , n16052 , n16053 );
buf ( n16055 , n16054 );
buf ( n16056 , n16055 );
xor ( n16057 , n16050 , n16056 );
buf ( n16058 , n16057 );
buf ( n16059 , n16058 );
xor ( n16060 , n16012 , n16059 );
buf ( n16061 , n16060 );
buf ( n16062 , n16061 );
xor ( n16063 , n15955 , n16062 );
buf ( n16064 , n15464 );
buf ( n16065 , n15475 );
nand ( n16066 , n16064 , n16065 );
buf ( n16067 , n16066 );
buf ( n16068 , n16067 );
not ( n16069 , n16068 );
buf ( n16070 , n15409 );
not ( n16071 , n16070 );
or ( n16072 , n16069 , n16071 );
buf ( n16073 , n15467 );
buf ( n16074 , n15472 );
nand ( n16075 , n16073 , n16074 );
buf ( n16076 , n16075 );
buf ( n16077 , n16076 );
nand ( n16078 , n16072 , n16077 );
buf ( n16079 , n16078 );
buf ( n16080 , n16079 );
xor ( n16081 , n16063 , n16080 );
buf ( n16082 , n16081 );
buf ( n16083 , n16082 );
not ( n16084 , n16083 );
buf ( n16085 , n16084 );
and ( n16086 , n15949 , n16085 );
not ( n16087 , n15949 );
and ( n16088 , n16087 , n16082 );
nor ( n16089 , n16086 , n16088 );
not ( n16090 , n16089 );
not ( n16091 , n16090 );
or ( n16092 , n15944 , n16091 );
nand ( n16093 , n16089 , n15942 );
nand ( n16094 , n16092 , n16093 );
buf ( n16095 , n16094 );
xor ( n16096 , n15488 , n15493 );
and ( n16097 , n16096 , n15627 );
and ( n16098 , n15488 , n15493 );
or ( n16099 , n16097 , n16098 );
buf ( n16100 , n16099 );
buf ( n16101 , n16100 );
nor ( n16102 , n16095 , n16101 );
buf ( n16103 , n16102 );
buf ( n16104 , n16103 );
not ( n16105 , n16104 );
buf ( n16106 , n16105 );
buf ( n16107 , n16106 );
buf ( n16108 , n16094 );
buf ( n16109 , n16100 );
nand ( n16110 , n16108 , n16109 );
buf ( n16111 , n16110 );
buf ( n16112 , n16111 );
nand ( n16113 , n16107 , n16112 );
buf ( n16114 , n16113 );
not ( n16115 , n16114 );
buf ( n16116 , n9298 );
not ( n16117 , n16116 );
buf ( n16118 , n16117 );
not ( n16119 , n16118 );
buf ( n16120 , n14757 );
buf ( n16121 , n15074 );
buf ( n16122 , n15632 );
nor ( n16123 , n16121 , n16122 );
buf ( n16124 , n16123 );
buf ( n16125 , n16124 );
and ( n16126 , n16120 , n16125 );
buf ( n16127 , n16126 );
nand ( n16128 , n16127 , n14212 );
not ( n16129 , n16128 );
not ( n16130 , n16129 );
or ( n16131 , n16119 , n16130 );
not ( n16132 , n14231 );
not ( n16133 , n16127 );
or ( n16134 , n16132 , n16133 );
and ( n16135 , n15078 , n15640 );
not ( n16136 , n16135 );
not ( n16137 , n15332 );
or ( n16138 , n16136 , n16137 );
buf ( n16139 , n15635 );
not ( n16140 , n16139 );
buf ( n16141 , n16140 );
nand ( n16142 , n16138 , n16141 );
nand ( n16143 , n16134 , n16142 );
not ( n16144 , n16143 );
nand ( n16145 , n16131 , n16144 );
not ( n16146 , n16145 );
not ( n16147 , n16146 );
or ( n16148 , n16115 , n16147 );
buf ( n16149 , n16114 );
not ( n16150 , n16149 );
buf ( n16151 , n16150 );
not ( n16152 , n16151 );
or ( n16153 , n16152 , n16146 );
nand ( n16154 , n16148 , n16153 );
nand ( n16155 , n15810 , n16154 );
not ( n16156 , n14235 );
not ( n16157 , n14760 );
buf ( n16158 , n16124 );
buf ( n16159 , n16106 );
nand ( n16160 , n16158 , n16159 );
buf ( n16161 , n16160 );
nor ( n16162 , n16157 , n16161 );
not ( n16163 , n16162 );
or ( n16164 , n16156 , n16163 );
not ( n16165 , n16161 );
not ( n16166 , n14772 );
and ( n16167 , n16165 , n16166 );
not ( n16168 , n15640 );
nor ( n16169 , n15635 , n15078 );
nor ( n16170 , n16168 , n16169 );
buf ( n16171 , n16170 );
buf ( n16172 , n16103 );
or ( n16173 , n16171 , n16172 );
buf ( n16174 , n16111 );
nand ( n16175 , n16173 , n16174 );
buf ( n16176 , n16175 );
nor ( n16177 , n16167 , n16176 );
nand ( n16178 , n16164 , n16177 );
buf ( n16179 , n15943 );
buf ( n16180 , n16085 );
nand ( n16181 , n16179 , n16180 );
buf ( n16182 , n16181 );
buf ( n16183 , n16182 );
buf ( n16184 , n15949 );
buf ( n16185 , n16184 );
and ( n16186 , n16183 , n16185 );
buf ( n16187 , n15943 );
buf ( n16188 , n16085 );
nor ( n16189 , n16187 , n16188 );
buf ( n16190 , n16189 );
buf ( n16191 , n16190 );
nor ( n16192 , n16186 , n16191 );
buf ( n16193 , n16192 );
buf ( n16194 , n16193 );
not ( n16195 , n16194 );
buf ( n16196 , n16195 );
buf ( n16197 , n16196 );
xor ( n16198 , n15955 , n16062 );
and ( n16199 , n16198 , n16080 );
and ( n16200 , n15955 , n16062 );
or ( n16201 , n16199 , n16200 );
buf ( n16202 , n16201 );
buf ( n16203 , n16202 );
xor ( n16204 , n15876 , n15899 );
and ( n16205 , n16204 , n15907 );
and ( n16206 , n15876 , n15899 );
or ( n16207 , n16205 , n16206 );
buf ( n16208 , n16207 );
buf ( n16209 , n16208 );
xor ( n16210 , n15825 , n15833 );
and ( n16211 , n16210 , n15850 );
and ( n16212 , n15825 , n15833 );
or ( n16213 , n16211 , n16212 );
not ( n16214 , n16213 );
buf ( n16215 , n550 );
buf ( n16216 , n576 );
and ( n16217 , n16215 , n16216 );
buf ( n16218 , n16217 );
buf ( n16219 , n16218 );
buf ( n16220 , n15895 );
xor ( n16221 , n16219 , n16220 );
buf ( n16222 , n15869 );
not ( n16223 , n16222 );
buf ( n16224 , n14637 );
not ( n16225 , n16224 );
or ( n16226 , n16223 , n16225 );
buf ( n16227 , n8294 );
buf ( n16228 , n546 );
buf ( n16229 , n578 );
xor ( n16230 , n16228 , n16229 );
buf ( n16231 , n16230 );
buf ( n16232 , n16231 );
nand ( n16233 , n16227 , n16232 );
buf ( n16234 , n16233 );
buf ( n16235 , n16234 );
nand ( n16236 , n16226 , n16235 );
buf ( n16237 , n16236 );
buf ( n16238 , n16237 );
xor ( n16239 , n16221 , n16238 );
buf ( n16240 , n16239 );
not ( n16241 , n16240 );
and ( n16242 , n16214 , n16241 );
not ( n16243 , n16214 );
not ( n16244 , n16241 );
and ( n16245 , n16243 , n16244 );
nor ( n16246 , n16242 , n16245 );
buf ( n16247 , n4211 );
not ( n16248 , n16247 );
buf ( n16249 , n16248 );
buf ( n16250 , n16249 );
not ( n16251 , n16250 );
buf ( n16252 , n4202 );
not ( n16253 , n16252 );
or ( n16254 , n16251 , n16253 );
buf ( n16255 , n582 );
nand ( n16256 , n16254 , n16255 );
buf ( n16257 , n16256 );
buf ( n16258 , n15844 );
not ( n16259 , n16258 );
buf ( n16260 , n14616 );
not ( n16261 , n16260 );
or ( n16262 , n16259 , n16261 );
buf ( n16263 , n9952 );
buf ( n16264 , n548 );
buf ( n16265 , n576 );
xor ( n16266 , n16264 , n16265 );
buf ( n16267 , n16266 );
buf ( n16268 , n16267 );
nand ( n16269 , n16263 , n16268 );
buf ( n16270 , n16269 );
buf ( n16271 , n16270 );
nand ( n16272 , n16262 , n16271 );
buf ( n16273 , n16272 );
not ( n16274 , n16273 );
and ( n16275 , n16257 , n16274 );
not ( n16276 , n16257 );
not ( n16277 , n16274 );
and ( n16278 , n16276 , n16277 );
or ( n16279 , n16275 , n16278 );
buf ( n16280 , n15889 );
not ( n16281 , n16280 );
buf ( n16282 , n15881 );
not ( n16283 , n16282 );
or ( n16284 , n16281 , n16283 );
buf ( n16285 , n5065 );
buf ( n16286 , n544 );
buf ( n16287 , n580 );
xor ( n16288 , n16286 , n16287 );
buf ( n16289 , n16288 );
buf ( n16290 , n16289 );
nand ( n16291 , n16285 , n16290 );
buf ( n16292 , n16291 );
buf ( n16293 , n16292 );
nand ( n16294 , n16284 , n16293 );
buf ( n16295 , n16294 );
not ( n16296 , n16295 );
not ( n16297 , n16296 );
xor ( n16298 , n16279 , n16297 );
and ( n16299 , n16246 , n16298 );
not ( n16300 , n16246 );
not ( n16301 , n16298 );
and ( n16302 , n16300 , n16301 );
nor ( n16303 , n16299 , n16302 );
buf ( n16304 , n16303 );
xor ( n16305 , n16209 , n16304 );
xor ( n16306 , n15852 , n15858 );
and ( n16307 , n16306 , n15910 );
and ( n16308 , n15852 , n15858 );
or ( n16309 , n16307 , n16308 );
buf ( n16310 , n16309 );
buf ( n16311 , n16310 );
xor ( n16312 , n16305 , n16311 );
buf ( n16313 , n16312 );
buf ( n16314 , n16313 );
xor ( n16315 , n15821 , n15913 );
and ( n16316 , n16315 , n15920 );
and ( n16317 , n15821 , n15913 );
or ( n16318 , n16316 , n16317 );
buf ( n16319 , n16318 );
buf ( n16320 , n16319 );
xor ( n16321 , n16314 , n16320 );
xor ( n16322 , n16029 , n16049 );
and ( n16323 , n16322 , n16056 );
and ( n16324 , n16029 , n16049 );
or ( n16325 , n16323 , n16324 );
buf ( n16326 , n16325 );
buf ( n16327 , n16326 );
xor ( n16328 , n15960 , n15977 );
and ( n16329 , n16328 , n15991 );
and ( n16330 , n15960 , n15977 );
or ( n16331 , n16329 , n16330 );
buf ( n16332 , n16331 );
buf ( n16333 , n16332 );
buf ( n16334 , n550 );
buf ( n16335 , n560 );
and ( n16336 , n16334 , n16335 );
buf ( n16337 , n16336 );
buf ( n16338 , n16337 );
buf ( n16339 , n16045 );
xor ( n16340 , n16338 , n16339 );
buf ( n16341 , n16022 );
not ( n16342 , n16341 );
buf ( n16343 , n9798 );
not ( n16344 , n16343 );
or ( n16345 , n16342 , n16344 );
buf ( n16346 , n5801 );
buf ( n16347 , n546 );
buf ( n16348 , n562 );
xor ( n16349 , n16347 , n16348 );
buf ( n16350 , n16349 );
buf ( n16351 , n16350 );
nand ( n16352 , n16346 , n16351 );
buf ( n16353 , n16352 );
buf ( n16354 , n16353 );
nand ( n16355 , n16345 , n16354 );
buf ( n16356 , n16355 );
buf ( n16357 , n16356 );
xor ( n16358 , n16340 , n16357 );
buf ( n16359 , n16358 );
buf ( n16360 , n16359 );
xor ( n16361 , n16333 , n16360 );
buf ( n16362 , n15970 );
not ( n16363 , n16362 );
buf ( n16364 , n10380 );
not ( n16365 , n16364 );
or ( n16366 , n16363 , n16365 );
buf ( n16367 , n6595 );
buf ( n16368 , n548 );
buf ( n16369 , n560 );
xor ( n16370 , n16368 , n16369 );
buf ( n16371 , n16370 );
buf ( n16372 , n16371 );
nand ( n16373 , n16367 , n16372 );
buf ( n16374 , n16373 );
buf ( n16375 , n16374 );
nand ( n16376 , n16366 , n16375 );
buf ( n16377 , n16376 );
buf ( n16378 , n16377 );
buf ( n16379 , n16039 );
not ( n16380 , n16379 );
buf ( n16381 , n14419 );
not ( n16382 , n16381 );
or ( n16383 , n16380 , n16382 );
buf ( n16384 , n4840 );
xor ( n16385 , n564 , n544 );
buf ( n16386 , n16385 );
nand ( n16387 , n16384 , n16386 );
buf ( n16388 , n16387 );
buf ( n16389 , n16388 );
nand ( n16390 , n16383 , n16389 );
buf ( n16391 , n16390 );
buf ( n16392 , n16391 );
xor ( n16393 , n16378 , n16392 );
buf ( n16394 , n3743 );
buf ( n16395 , n13926 );
or ( n16396 , n16394 , n16395 );
buf ( n16397 , n566 );
nand ( n16398 , n16396 , n16397 );
buf ( n16399 , n16398 );
buf ( n16400 , n16399 );
xor ( n16401 , n16393 , n16400 );
buf ( n16402 , n16401 );
buf ( n16403 , n16402 );
xor ( n16404 , n16361 , n16403 );
buf ( n16405 , n16404 );
buf ( n16406 , n16405 );
xor ( n16407 , n16327 , n16406 );
xor ( n16408 , n15994 , n16011 );
and ( n16409 , n16408 , n16059 );
and ( n16410 , n15994 , n16011 );
or ( n16411 , n16409 , n16410 );
buf ( n16412 , n16411 );
buf ( n16413 , n16412 );
xor ( n16414 , n16407 , n16413 );
buf ( n16415 , n16414 );
buf ( n16416 , n16415 );
xor ( n16417 , n16321 , n16416 );
buf ( n16418 , n16417 );
buf ( n16419 , n16418 );
xor ( n16420 , n16203 , n16419 );
buf ( n16421 , n15937 );
not ( n16422 , n16421 );
buf ( n16423 , n15815 );
not ( n16424 , n16423 );
or ( n16425 , n16422 , n16424 );
buf ( n16426 , n15815 );
buf ( n16427 , n15937 );
or ( n16428 , n16426 , n16427 );
buf ( n16429 , n15922 );
nand ( n16430 , n16428 , n16429 );
buf ( n16431 , n16430 );
buf ( n16432 , n16431 );
nand ( n16433 , n16425 , n16432 );
buf ( n16434 , n16433 );
buf ( n16435 , n16434 );
xor ( n16436 , n16420 , n16435 );
buf ( n16437 , n16436 );
buf ( n16438 , n16437 );
nor ( n16439 , n16197 , n16438 );
buf ( n16440 , n16439 );
not ( n16441 , n16440 );
buf ( n16442 , n16437 );
buf ( n16443 , n16196 );
nand ( n16444 , n16442 , n16443 );
buf ( n16445 , n16444 );
nand ( n16446 , n16441 , n16445 );
and ( n16447 , n16178 , n16446 );
not ( n16448 , n16178 );
not ( n16449 , n16446 );
and ( n16450 , n16448 , n16449 );
nor ( n16451 , n16447 , n16450 );
nand ( n16452 , n15795 , n15789 );
not ( n16453 , n16452 );
nand ( n16454 , n15104 , n16453 );
not ( n16455 , n16454 );
not ( n16456 , n15714 );
nand ( n16457 , n16456 , n15788 );
not ( n16458 , n16457 );
not ( n16459 , n15802 );
or ( n16460 , n16458 , n16459 );
nand ( n16461 , n16460 , n15790 );
not ( n16462 , n16461 );
buf ( n16463 , n16462 );
not ( n16464 , n16463 );
or ( n16465 , n16455 , n16464 );
and ( n16466 , n544 , n6908 );
not ( n16467 , n6945 );
not ( n16468 , n546 );
buf ( n16469 , n7223 );
not ( n16470 , n16469 );
or ( n16471 , n16468 , n16470 );
not ( n16472 , n16469 );
nand ( n16473 , n16472 , n6949 );
nand ( n16474 , n16471 , n16473 );
not ( n16475 , n16474 );
or ( n16476 , n16467 , n16475 );
nand ( n16477 , n15747 , n9575 );
nand ( n16478 , n16476 , n16477 );
xor ( n16479 , n16466 , n16478 );
xor ( n16480 , n15749 , n15755 );
and ( n16481 , n16480 , n15767 );
and ( n16482 , n15749 , n15755 );
or ( n16483 , n16481 , n16482 );
xor ( n16484 , n16479 , n16483 );
xor ( n16485 , n15723 , n15725 );
and ( n16486 , n16485 , n15738 );
and ( n16487 , n15723 , n15725 );
or ( n16488 , n16486 , n16487 );
not ( n16489 , n9327 );
not ( n16490 , n548 );
not ( n16491 , n15270 );
or ( n16492 , n16490 , n16491 );
nand ( n16493 , n15269 , n5279 );
nand ( n16494 , n16492 , n16493 );
not ( n16495 , n16494 );
or ( n16496 , n16489 , n16495 );
nand ( n16497 , n15765 , n6939 );
nand ( n16498 , n16496 , n16497 );
not ( n16499 , n15736 );
not ( n16500 , n16499 );
not ( n16501 , n5268 );
not ( n16502 , n16501 );
and ( n16503 , n16500 , n16502 );
and ( n16504 , n3068 , n550 );
nor ( n16505 , n16503 , n16504 );
xor ( n16506 , n16498 , n16505 );
not ( n16507 , n9409 );
xor ( n16508 , n544 , n7147 );
not ( n16509 , n16508 );
or ( n16510 , n16507 , n16509 );
nand ( n16511 , n15753 , n9417 );
nand ( n16512 , n16510 , n16511 );
xor ( n16513 , n16506 , n16512 );
xor ( n16514 , n16488 , n16513 );
xor ( n16515 , n15770 , n15774 );
and ( n16516 , n16515 , n15779 );
and ( n16517 , n15770 , n15774 );
or ( n16518 , n16516 , n16517 );
xor ( n16519 , n16514 , n16518 );
xor ( n16520 , n16484 , n16519 );
xor ( n16521 , n15739 , n15768 );
and ( n16522 , n16521 , n15780 );
and ( n16523 , n15739 , n15768 );
or ( n16524 , n16522 , n16523 );
xor ( n16525 , n16520 , n16524 );
xor ( n16526 , n15719 , n15781 );
and ( n16527 , n16526 , n15786 );
and ( n16528 , n15719 , n15781 );
or ( n16529 , n16527 , n16528 );
xor ( n16530 , n16525 , n16529 );
nand ( n16531 , n16465 , n16530 );
nor ( n16532 , n16529 , n16525 );
not ( n16533 , n16532 );
nand ( n16534 , n16529 , n16525 );
nand ( n16535 , n16533 , n16534 );
nand ( n16536 , n16454 , n16463 , n16535 );
nand ( n16537 , n16451 , n16531 , n16536 );
and ( n16538 , n16155 , n16537 );
xor ( n16539 , n16327 , n16406 );
and ( n16540 , n16539 , n16413 );
and ( n16541 , n16327 , n16406 );
or ( n16542 , n16540 , n16541 );
buf ( n16543 , n16542 );
buf ( n16544 , n16543 );
xor ( n16545 , n16314 , n16320 );
and ( n16546 , n16545 , n16416 );
and ( n16547 , n16314 , n16320 );
or ( n16548 , n16546 , n16547 );
buf ( n16549 , n16548 );
buf ( n16550 , n16549 );
xor ( n16551 , n16544 , n16550 );
xor ( n16552 , n16338 , n16339 );
and ( n16553 , n16552 , n16357 );
and ( n16554 , n16338 , n16339 );
or ( n16555 , n16553 , n16554 );
buf ( n16556 , n16555 );
buf ( n16557 , n16556 );
buf ( n16558 , n16385 );
not ( n16559 , n16558 );
buf ( n16560 , n14419 );
not ( n16561 , n16560 );
or ( n16562 , n16559 , n16561 );
buf ( n16563 , n4840 );
buf ( n16564 , n564 );
nand ( n16565 , n16563 , n16564 );
buf ( n16566 , n16565 );
buf ( n16567 , n16566 );
nand ( n16568 , n16562 , n16567 );
buf ( n16569 , n16568 );
buf ( n16570 , n16569 );
not ( n16571 , n16570 );
buf ( n16572 , n16571 );
buf ( n16573 , n16572 );
xor ( n16574 , n16378 , n16392 );
and ( n16575 , n16574 , n16400 );
and ( n16576 , n16378 , n16392 );
or ( n16577 , n16575 , n16576 );
buf ( n16578 , n16577 );
buf ( n16579 , n16578 );
xor ( n16580 , n16573 , n16579 );
buf ( n16581 , n549 );
buf ( n16582 , n560 );
and ( n16583 , n16581 , n16582 );
buf ( n16584 , n16583 );
buf ( n16585 , n16584 );
buf ( n16586 , n16371 );
not ( n16587 , n16586 );
buf ( n16588 , n10380 );
not ( n16589 , n16588 );
or ( n16590 , n16587 , n16589 );
buf ( n16591 , n6595 );
xor ( n16592 , n560 , n547 );
buf ( n16593 , n16592 );
nand ( n16594 , n16591 , n16593 );
buf ( n16595 , n16594 );
buf ( n16596 , n16595 );
nand ( n16597 , n16590 , n16596 );
buf ( n16598 , n16597 );
buf ( n16599 , n16598 );
xor ( n16600 , n16585 , n16599 );
buf ( n16601 , n16350 );
not ( n16602 , n16601 );
buf ( n16603 , n9798 );
not ( n16604 , n16603 );
or ( n16605 , n16602 , n16604 );
buf ( n16606 , n5801 );
buf ( n16607 , n545 );
buf ( n16608 , n562 );
xor ( n16609 , n16607 , n16608 );
buf ( n16610 , n16609 );
buf ( n16611 , n16610 );
nand ( n16612 , n16606 , n16611 );
buf ( n16613 , n16612 );
buf ( n16614 , n16613 );
nand ( n16615 , n16605 , n16614 );
buf ( n16616 , n16615 );
buf ( n16617 , n16616 );
xor ( n16618 , n16600 , n16617 );
buf ( n16619 , n16618 );
buf ( n16620 , n16619 );
xor ( n16621 , n16580 , n16620 );
buf ( n16622 , n16621 );
buf ( n16623 , n16622 );
xor ( n16624 , n16557 , n16623 );
xor ( n16625 , n16333 , n16360 );
and ( n16626 , n16625 , n16403 );
and ( n16627 , n16333 , n16360 );
or ( n16628 , n16626 , n16627 );
buf ( n16629 , n16628 );
buf ( n16630 , n16629 );
xor ( n16631 , n16624 , n16630 );
buf ( n16632 , n16631 );
buf ( n16633 , n16632 );
xor ( n16634 , n16219 , n16220 );
and ( n16635 , n16634 , n16238 );
and ( n16636 , n16219 , n16220 );
or ( n16637 , n16635 , n16636 );
buf ( n16638 , n16637 );
not ( n16639 , n16214 );
not ( n16640 , n16241 );
or ( n16641 , n16639 , n16640 );
nand ( n16642 , n16641 , n16298 );
not ( n16643 , n16214 );
nand ( n16644 , n16643 , n16244 );
nand ( n16645 , n16642 , n16644 );
xor ( n16646 , n16638 , n16645 );
not ( n16647 , n16289 );
not ( n16648 , n15881 );
or ( n16649 , n16647 , n16648 );
buf ( n16650 , n5065 );
buf ( n16651 , n580 );
nand ( n16652 , n16650 , n16651 );
buf ( n16653 , n16652 );
nand ( n16654 , n16649 , n16653 );
not ( n16655 , n16654 );
not ( n16656 , n16296 );
nand ( n16657 , n16656 , n16277 );
not ( n16658 , n16274 );
not ( n16659 , n16296 );
or ( n16660 , n16658 , n16659 );
nand ( n16661 , n16660 , n16257 );
nand ( n16662 , n16657 , n16661 );
xor ( n16663 , n16655 , n16662 );
buf ( n16664 , n549 );
buf ( n16665 , n576 );
and ( n16666 , n16664 , n16665 );
buf ( n16667 , n16666 );
buf ( n16668 , n16231 );
not ( n16669 , n16668 );
buf ( n16670 , n14637 );
not ( n16671 , n16670 );
or ( n16672 , n16669 , n16671 );
buf ( n16673 , n8294 );
buf ( n16674 , n545 );
buf ( n16675 , n578 );
xor ( n16676 , n16674 , n16675 );
buf ( n16677 , n16676 );
buf ( n16678 , n16677 );
nand ( n16679 , n16673 , n16678 );
buf ( n16680 , n16679 );
buf ( n16681 , n16680 );
nand ( n16682 , n16672 , n16681 );
buf ( n16683 , n16682 );
xor ( n16684 , n16667 , n16683 );
buf ( n16685 , n16267 );
not ( n16686 , n16685 );
buf ( n16687 , n14616 );
not ( n16688 , n16687 );
or ( n16689 , n16686 , n16688 );
buf ( n16690 , n9952 );
buf ( n16691 , n576 );
buf ( n16692 , n547 );
xor ( n16693 , n16691 , n16692 );
buf ( n16694 , n16693 );
buf ( n16695 , n16694 );
nand ( n16696 , n16690 , n16695 );
buf ( n16697 , n16696 );
buf ( n16698 , n16697 );
nand ( n16699 , n16689 , n16698 );
buf ( n16700 , n16699 );
xor ( n16701 , n16684 , n16700 );
xor ( n16702 , n16663 , n16701 );
xor ( n16703 , n16646 , n16702 );
buf ( n16704 , n16703 );
xor ( n16705 , n16633 , n16704 );
xor ( n16706 , n16209 , n16304 );
and ( n16707 , n16706 , n16311 );
and ( n16708 , n16209 , n16304 );
or ( n16709 , n16707 , n16708 );
buf ( n16710 , n16709 );
buf ( n16711 , n16710 );
xor ( n16712 , n16705 , n16711 );
buf ( n16713 , n16712 );
buf ( n16714 , n16713 );
xor ( n16715 , n16551 , n16714 );
buf ( n16716 , n16715 );
buf ( n16717 , n16716 );
xor ( n16718 , n16203 , n16419 );
and ( n16719 , n16718 , n16435 );
and ( n16720 , n16203 , n16419 );
or ( n16721 , n16719 , n16720 );
buf ( n16722 , n16721 );
buf ( n16723 , n16722 );
and ( n16724 , n16717 , n16723 );
buf ( n16725 , n16724 );
buf ( n16726 , n16725 );
not ( n16727 , n16726 );
buf ( n16728 , n16727 );
buf ( n16729 , n16722 );
buf ( n16730 , n16716 );
nor ( n16731 , n16729 , n16730 );
buf ( n16732 , n16731 );
buf ( n16733 , n16732 );
not ( n16734 , n16733 );
buf ( n16735 , n16734 );
nand ( n16736 , n16728 , n16735 );
not ( n16737 , n16736 );
buf ( n16738 , n16127 );
buf ( n16739 , n16103 );
buf ( n16740 , n16440 );
nor ( n16741 , n16739 , n16740 );
buf ( n16742 , n16741 );
buf ( n16743 , n16742 );
buf ( n16744 , n16743 );
buf ( n16745 , n16744 );
nand ( n16746 , n16118 , n14212 , n16738 , n16745 );
nand ( n16747 , n16143 , n16745 );
buf ( n16748 , n16440 );
buf ( n16749 , n16111 );
or ( n16750 , n16748 , n16749 );
buf ( n16751 , n16445 );
nand ( n16752 , n16750 , n16751 );
buf ( n16753 , n16752 );
buf ( n16754 , n16753 );
not ( n16755 , n16754 );
nand ( n16756 , n16746 , n16747 , n16755 );
not ( n16757 , n16756 );
or ( n16758 , n16737 , n16757 );
nor ( n16759 , n16754 , n16736 );
nand ( n16760 , n16747 , n16759 , n16746 );
nand ( n16761 , n16758 , n16760 );
not ( n16762 , n16761 );
not ( n16763 , n16762 );
or ( n16764 , n16529 , n16525 );
not ( n16765 , n16764 );
not ( n16766 , n16461 );
or ( n16767 , n16765 , n16766 );
nand ( n16768 , n16767 , n16534 );
not ( n16769 , n16768 );
not ( n16770 , n15102 );
nand ( n16771 , n10199 , n15089 );
not ( n16772 , n16771 );
or ( n16773 , n16770 , n16772 );
nor ( n16774 , n16452 , n16532 );
nand ( n16775 , n16773 , n16774 );
nand ( n16776 , n16769 , n16775 );
buf ( n16777 , n16776 );
xor ( n16778 , n16484 , n16519 );
and ( n16779 , n16778 , n16524 );
and ( n16780 , n16484 , n16519 );
or ( n16781 , n16779 , n16780 );
xor ( n16782 , n16466 , n16478 );
and ( n16783 , n16782 , n16483 );
and ( n16784 , n16466 , n16478 );
or ( n16785 , n16783 , n16784 );
xor ( n16786 , n16498 , n16505 );
and ( n16787 , n16786 , n16512 );
and ( n16788 , n16498 , n16505 );
or ( n16789 , n16787 , n16788 );
not ( n16790 , n9605 );
not ( n16791 , n16501 );
or ( n16792 , n16790 , n16791 );
nand ( n16793 , n16792 , n550 );
not ( n16794 , n6939 );
not ( n16795 , n16494 );
or ( n16796 , n16794 , n16795 );
not ( n16797 , n548 );
not ( n16798 , n15734 );
or ( n16799 , n16797 , n16798 );
nand ( n16800 , n15731 , n5279 );
nand ( n16801 , n16799 , n16800 );
nand ( n16802 , n16801 , n9327 );
nand ( n16803 , n16796 , n16802 );
xor ( n16804 , n16793 , n16803 );
not ( n16805 , n9417 );
not ( n16806 , n16508 );
or ( n16807 , n16805 , n16806 );
buf ( n16808 , n7124 );
xor ( n16809 , n544 , n16808 );
nand ( n16810 , n16809 , n9409 );
nand ( n16811 , n16807 , n16810 );
xor ( n16812 , n16804 , n16811 );
xor ( n16813 , n16789 , n16812 );
and ( n16814 , n544 , n6918 );
not ( n16815 , n9575 );
not ( n16816 , n16474 );
or ( n16817 , n16815 , n16816 );
not ( n16818 , n546 );
not ( n16819 , n7270 );
or ( n16820 , n16818 , n16819 );
nand ( n16821 , n15763 , n6949 );
nand ( n16822 , n16820 , n16821 );
nand ( n16823 , n16822 , n7179 );
nand ( n16824 , n16817 , n16823 );
xor ( n16825 , n16814 , n16824 );
not ( n16826 , n16505 );
xor ( n16827 , n16825 , n16826 );
xor ( n16828 , n16813 , n16827 );
xor ( n16829 , n16785 , n16828 );
xor ( n16830 , n16488 , n16513 );
and ( n16831 , n16830 , n16518 );
and ( n16832 , n16488 , n16513 );
or ( n16833 , n16831 , n16832 );
xor ( n16834 , n16829 , n16833 );
not ( n16835 , n16834 );
not ( n16836 , n16835 );
and ( n16837 , n16781 , n16836 );
not ( n16838 , n16781 );
and ( n16839 , n16838 , n16835 );
nor ( n16840 , n16837 , n16839 );
and ( n16841 , n16777 , n16840 );
not ( n16842 , n16777 );
not ( n16843 , n16840 );
and ( n16844 , n16842 , n16843 );
nor ( n16845 , n16841 , n16844 );
not ( n16846 , n16845 );
or ( n16847 , n16763 , n16846 );
not ( n16848 , n16781 );
nand ( n16849 , n16848 , n16835 );
not ( n16850 , n16849 );
not ( n16851 , n16776 );
or ( n16852 , n16850 , n16851 );
nand ( n16853 , n16781 , n16836 );
nand ( n16854 , n16852 , n16853 );
not ( n16855 , n16854 );
xor ( n16856 , n16785 , n16828 );
and ( n16857 , n16856 , n16833 );
and ( n16858 , n16785 , n16828 );
or ( n16859 , n16857 , n16858 );
not ( n16860 , n16859 );
not ( n16861 , n16860 );
and ( n16862 , n544 , n7147 );
not ( n16863 , n6945 );
not ( n16864 , n546 );
not ( n16865 , n15270 );
or ( n16866 , n16864 , n16865 );
nand ( n16867 , n15269 , n6949 );
nand ( n16868 , n16866 , n16867 );
not ( n16869 , n16868 );
or ( n16870 , n16863 , n16869 );
nand ( n16871 , n16822 , n9575 );
nand ( n16872 , n16870 , n16871 );
xor ( n16873 , n16862 , n16872 );
and ( n16874 , n16801 , n6939 );
not ( n16875 , n9327 );
nor ( n16876 , n16875 , n5279 );
nor ( n16877 , n16874 , n16876 );
xor ( n16878 , n16873 , n16877 );
not ( n16879 , n9409 );
xor ( n16880 , n544 , n16472 );
not ( n16881 , n16880 );
or ( n16882 , n16879 , n16881 );
nand ( n16883 , n16809 , n9417 );
nand ( n16884 , n16882 , n16883 );
xor ( n16885 , n16814 , n16824 );
and ( n16886 , n16885 , n16826 );
and ( n16887 , n16814 , n16824 );
or ( n16888 , n16886 , n16887 );
xor ( n16889 , n16884 , n16888 );
xor ( n16890 , n16793 , n16803 );
and ( n16891 , n16890 , n16811 );
and ( n16892 , n16793 , n16803 );
or ( n16893 , n16891 , n16892 );
xor ( n16894 , n16889 , n16893 );
xor ( n16895 , n16878 , n16894 );
xor ( n16896 , n16789 , n16812 );
and ( n16897 , n16896 , n16827 );
and ( n16898 , n16789 , n16812 );
or ( n16899 , n16897 , n16898 );
xor ( n16900 , n16895 , n16899 );
not ( n16901 , n16900 );
not ( n16902 , n16901 );
or ( n16903 , n16861 , n16902 );
nand ( n16904 , n16859 , n16900 );
nand ( n16905 , n16903 , n16904 );
nand ( n16906 , n16855 , n16905 );
xor ( n16907 , n16544 , n16550 );
and ( n16908 , n16907 , n16714 );
and ( n16909 , n16544 , n16550 );
or ( n16910 , n16908 , n16909 );
buf ( n16911 , n16910 );
buf ( n16912 , n16911 );
xor ( n16913 , n16557 , n16623 );
and ( n16914 , n16913 , n16630 );
and ( n16915 , n16557 , n16623 );
or ( n16916 , n16914 , n16915 );
buf ( n16917 , n16916 );
buf ( n16918 , n16917 );
buf ( n16919 , n548 );
buf ( n16920 , n560 );
and ( n16921 , n16919 , n16920 );
buf ( n16922 , n16921 );
buf ( n16923 , n16922 );
buf ( n16924 , n16610 );
not ( n16925 , n16924 );
buf ( n16926 , n9798 );
not ( n16927 , n16926 );
or ( n16928 , n16925 , n16927 );
buf ( n16929 , n5801 );
and ( n16930 , n562 , n544 );
not ( n16931 , n562 );
and ( n16932 , n16931 , n8477 );
nor ( n16933 , n16930 , n16932 );
buf ( n16934 , n16933 );
nand ( n16935 , n16929 , n16934 );
buf ( n16936 , n16935 );
buf ( n16937 , n16936 );
nand ( n16938 , n16928 , n16937 );
buf ( n16939 , n16938 );
buf ( n16940 , n16939 );
xor ( n16941 , n16923 , n16940 );
buf ( n16942 , n4840 );
buf ( n16943 , n14419 );
or ( n16944 , n16942 , n16943 );
buf ( n16945 , n564 );
nand ( n16946 , n16944 , n16945 );
buf ( n16947 , n16946 );
buf ( n16948 , n16947 );
xor ( n16949 , n16941 , n16948 );
buf ( n16950 , n16949 );
buf ( n16951 , n16950 );
buf ( n16952 , n16569 );
buf ( n16953 , n16592 );
not ( n16954 , n16953 );
buf ( n16955 , n10380 );
not ( n16956 , n16955 );
or ( n16957 , n16954 , n16956 );
buf ( n16958 , n6595 );
buf ( n16959 , n560 );
buf ( n16960 , n546 );
xor ( n16961 , n16959 , n16960 );
buf ( n16962 , n16961 );
buf ( n16963 , n16962 );
nand ( n16964 , n16958 , n16963 );
buf ( n16965 , n16964 );
buf ( n16966 , n16965 );
nand ( n16967 , n16957 , n16966 );
buf ( n16968 , n16967 );
buf ( n16969 , n16968 );
xor ( n16970 , n16952 , n16969 );
xor ( n16971 , n16585 , n16599 );
and ( n16972 , n16971 , n16617 );
and ( n16973 , n16585 , n16599 );
or ( n16974 , n16972 , n16973 );
buf ( n16975 , n16974 );
buf ( n16976 , n16975 );
xor ( n16977 , n16970 , n16976 );
buf ( n16978 , n16977 );
buf ( n16979 , n16978 );
xor ( n16980 , n16951 , n16979 );
xor ( n16981 , n16573 , n16579 );
and ( n16982 , n16981 , n16620 );
and ( n16983 , n16573 , n16579 );
or ( n16984 , n16982 , n16983 );
buf ( n16985 , n16984 );
buf ( n16986 , n16985 );
xor ( n16987 , n16980 , n16986 );
buf ( n16988 , n16987 );
buf ( n16989 , n16988 );
or ( n16990 , n16667 , n16700 );
nand ( n16991 , n16990 , n16683 );
nand ( n16992 , n16700 , n16667 );
nand ( n16993 , n16991 , n16992 );
buf ( n16994 , n16694 );
not ( n16995 , n16994 );
buf ( n16996 , n14616 );
not ( n16997 , n16996 );
or ( n16998 , n16995 , n16997 );
buf ( n16999 , n9952 );
buf ( n17000 , n576 );
buf ( n17001 , n546 );
xor ( n17002 , n17000 , n17001 );
buf ( n17003 , n17002 );
buf ( n17004 , n17003 );
nand ( n17005 , n16999 , n17004 );
buf ( n17006 , n17005 );
buf ( n17007 , n17006 );
nand ( n17008 , n16998 , n17007 );
buf ( n17009 , n17008 );
and ( n17010 , n16654 , n17009 );
not ( n17011 , n16654 );
not ( n17012 , n17009 );
and ( n17013 , n17011 , n17012 );
nor ( n17014 , n17010 , n17013 );
xor ( n17015 , n16993 , n17014 );
xor ( n17016 , n16655 , n16662 );
and ( n17017 , n17016 , n16701 );
and ( n17018 , n16655 , n16662 );
or ( n17019 , n17017 , n17018 );
xor ( n17020 , n17015 , n17019 );
buf ( n17021 , n548 );
buf ( n17022 , n576 );
and ( n17023 , n17021 , n17022 );
buf ( n17024 , n17023 );
buf ( n17025 , n17024 );
buf ( n17026 , n16677 );
not ( n17027 , n17026 );
buf ( n17028 , n14637 );
not ( n17029 , n17028 );
or ( n17030 , n17027 , n17029 );
buf ( n17031 , n8294 );
buf ( n17032 , n544 );
buf ( n17033 , n578 );
xor ( n17034 , n17032 , n17033 );
buf ( n17035 , n17034 );
buf ( n17036 , n17035 );
nand ( n17037 , n17031 , n17036 );
buf ( n17038 , n17037 );
buf ( n17039 , n17038 );
nand ( n17040 , n17030 , n17039 );
buf ( n17041 , n17040 );
buf ( n17042 , n17041 );
xor ( n17043 , n17025 , n17042 );
buf ( n17044 , n5065 );
buf ( n17045 , n15881 );
or ( n17046 , n17044 , n17045 );
buf ( n17047 , n580 );
nand ( n17048 , n17046 , n17047 );
buf ( n17049 , n17048 );
buf ( n17050 , n17049 );
xor ( n17051 , n17043 , n17050 );
buf ( n17052 , n17051 );
xor ( n17053 , n17020 , n17052 );
buf ( n17054 , n17053 );
xor ( n17055 , n16989 , n17054 );
xor ( n17056 , n16638 , n16645 );
and ( n17057 , n17056 , n16702 );
and ( n17058 , n16638 , n16645 );
or ( n17059 , n17057 , n17058 );
buf ( n17060 , n17059 );
xor ( n17061 , n17055 , n17060 );
buf ( n17062 , n17061 );
buf ( n17063 , n17062 );
xor ( n17064 , n16918 , n17063 );
xor ( n17065 , n16633 , n16704 );
and ( n17066 , n17065 , n16711 );
and ( n17067 , n16633 , n16704 );
or ( n17068 , n17066 , n17067 );
buf ( n17069 , n17068 );
buf ( n17070 , n17069 );
xor ( n17071 , n17064 , n17070 );
buf ( n17072 , n17071 );
buf ( n17073 , n17072 );
and ( n17074 , n16912 , n17073 );
buf ( n17075 , n17074 );
buf ( n17076 , n16911 );
buf ( n17077 , n17072 );
nor ( n17078 , n17076 , n17077 );
buf ( n17079 , n17078 );
nor ( n17080 , n17075 , n17079 );
not ( n17081 , n17080 );
and ( n17082 , n16742 , n16735 );
nand ( n17083 , n16143 , n17082 );
nand ( n17084 , n16129 , n17082 , n16118 );
buf ( n17085 , n16735 );
not ( n17086 , n17085 );
buf ( n17087 , n16753 );
not ( n17088 , n17087 );
or ( n17089 , n17086 , n17088 );
buf ( n17090 , n16728 );
nand ( n17091 , n17089 , n17090 );
buf ( n17092 , n17091 );
not ( n17093 , n17092 );
nand ( n17094 , n17083 , n17084 , n17093 );
not ( n17095 , n17094 );
or ( n17096 , n17081 , n17095 );
not ( n17097 , n17075 );
buf ( n17098 , n17079 );
not ( n17099 , n17098 );
buf ( n17100 , n17099 );
nand ( n17101 , n17097 , n17100 );
nand ( n17102 , n17083 , n17084 , n17093 , n17101 );
nand ( n17103 , n17096 , n17102 );
not ( n17104 , n16905 );
nand ( n17105 , n17104 , n16854 );
nand ( n17106 , n16906 , n17103 , n17105 );
nand ( n17107 , n16847 , n17106 );
not ( n17108 , n17107 );
nand ( n17109 , n16538 , n17108 );
xor ( n17110 , n16878 , n16894 );
and ( n17111 , n17110 , n16899 );
and ( n17112 , n16878 , n16894 );
or ( n17113 , n17111 , n17112 );
or ( n17114 , n6939 , n9327 );
nand ( n17115 , n17114 , n548 );
not ( n17116 , n9575 );
not ( n17117 , n16868 );
or ( n17118 , n17116 , n17117 );
not ( n17119 , n6949 );
not ( n17120 , n15731 );
or ( n17121 , n17119 , n17120 );
nand ( n17122 , n15734 , n546 );
nand ( n17123 , n17121 , n17122 );
nand ( n17124 , n17123 , n7179 );
nand ( n17125 , n17118 , n17124 );
xor ( n17126 , n17115 , n17125 );
and ( n17127 , n544 , n16808 );
xor ( n17128 , n17126 , n17127 );
not ( n17129 , n16877 );
not ( n17130 , n9417 );
not ( n17131 , n16880 );
or ( n17132 , n17130 , n17131 );
xor ( n17133 , n544 , n15763 );
nand ( n17134 , n17133 , n9409 );
nand ( n17135 , n17132 , n17134 );
xor ( n17136 , n17129 , n17135 );
xor ( n17137 , n16862 , n16872 );
and ( n17138 , n17137 , n16877 );
and ( n17139 , n16862 , n16872 );
or ( n17140 , n17138 , n17139 );
xor ( n17141 , n17136 , n17140 );
xor ( n17142 , n17128 , n17141 );
xor ( n17143 , n16884 , n16888 );
and ( n17144 , n17143 , n16893 );
and ( n17145 , n16884 , n16888 );
or ( n17146 , n17144 , n17145 );
xor ( n17147 , n17142 , n17146 );
nor ( n17148 , n17113 , n17147 );
not ( n17149 , n17148 );
nand ( n17150 , n17113 , n17147 );
nand ( n17151 , n17149 , n17150 );
not ( n17152 , n17151 );
not ( n17153 , n16849 );
not ( n17154 , n16776 );
or ( n17155 , n17153 , n17154 );
nand ( n17156 , n17155 , n16853 );
nand ( n17157 , n16860 , n16901 );
nand ( n17158 , n17156 , n17157 );
buf ( n17159 , n16904 );
nand ( n17160 , n17158 , n17159 );
not ( n17161 , n17160 );
or ( n17162 , n17152 , n17161 );
not ( n17163 , n17159 );
nor ( n17164 , n17163 , n17151 );
nand ( n17165 , n17164 , n17158 );
nand ( n17166 , n17162 , n17165 );
not ( n17167 , n17166 );
buf ( n17168 , n16732 );
buf ( n17169 , n17079 );
nor ( n17170 , n17168 , n17169 );
buf ( n17171 , n17170 );
buf ( n17172 , n17171 );
not ( n17173 , n17172 );
buf ( n17174 , n16753 );
not ( n17175 , n17174 );
or ( n17176 , n17173 , n17175 );
buf ( n17177 , n17100 );
buf ( n17178 , n16725 );
and ( n17179 , n17177 , n17178 );
buf ( n17180 , n17075 );
nor ( n17181 , n17179 , n17180 );
buf ( n17182 , n17181 );
buf ( n17183 , n17182 );
nand ( n17184 , n17176 , n17183 );
buf ( n17185 , n17184 );
not ( n17186 , n17185 );
buf ( n17187 , n16742 );
buf ( n17188 , n17171 );
and ( n17189 , n17187 , n17188 );
buf ( n17190 , n17189 );
nand ( n17191 , n17190 , n16143 );
buf ( n17192 , n16129 );
buf ( n17193 , n16118 );
buf ( n17194 , n17193 );
buf ( n17195 , n17194 );
buf ( n17196 , n17195 );
buf ( n17197 , n17190 );
nand ( n17198 , n17192 , n17196 , n17197 );
buf ( n17199 , n17198 );
nand ( n17200 , n17186 , n17191 , n17199 );
xor ( n17201 , n16918 , n17063 );
and ( n17202 , n17201 , n17070 );
and ( n17203 , n16918 , n17063 );
or ( n17204 , n17202 , n17203 );
buf ( n17205 , n17204 );
buf ( n17206 , n17205 );
not ( n17207 , n17206 );
xor ( n17208 , n16951 , n16979 );
and ( n17209 , n17208 , n16986 );
and ( n17210 , n16951 , n16979 );
or ( n17211 , n17209 , n17210 );
buf ( n17212 , n17211 );
buf ( n17213 , n17212 );
xor ( n17214 , n17025 , n17042 );
and ( n17215 , n17214 , n17050 );
and ( n17216 , n17025 , n17042 );
or ( n17217 , n17215 , n17216 );
buf ( n17218 , n17217 );
buf ( n17219 , n17218 );
and ( n17220 , n16691 , n16692 );
buf ( n17221 , n17220 );
buf ( n17222 , n17221 );
buf ( n17223 , n17003 );
not ( n17224 , n17223 );
buf ( n17225 , n14616 );
not ( n17226 , n17225 );
or ( n17227 , n17224 , n17226 );
buf ( n17228 , n9952 );
buf ( n17229 , n545 );
buf ( n17230 , n576 );
xor ( n17231 , n17229 , n17230 );
buf ( n17232 , n17231 );
buf ( n17233 , n17232 );
nand ( n17234 , n17228 , n17233 );
buf ( n17235 , n17234 );
buf ( n17236 , n17235 );
nand ( n17237 , n17227 , n17236 );
buf ( n17238 , n17237 );
buf ( n17239 , n17238 );
xor ( n17240 , n17222 , n17239 );
buf ( n17241 , n17035 );
not ( n17242 , n17241 );
buf ( n17243 , n14637 );
not ( n17244 , n17243 );
or ( n17245 , n17242 , n17244 );
buf ( n17246 , n8294 );
buf ( n17247 , n578 );
nand ( n17248 , n17246 , n17247 );
buf ( n17249 , n17248 );
buf ( n17250 , n17249 );
nand ( n17251 , n17245 , n17250 );
buf ( n17252 , n17251 );
buf ( n17253 , n17252 );
not ( n17254 , n17253 );
buf ( n17255 , n17254 );
buf ( n17256 , n17255 );
xor ( n17257 , n17240 , n17256 );
buf ( n17258 , n17257 );
buf ( n17259 , n17258 );
xor ( n17260 , n17219 , n17259 );
not ( n17261 , n16655 );
not ( n17262 , n17012 );
or ( n17263 , n17261 , n17262 );
nand ( n17264 , n17263 , n16993 );
nand ( n17265 , n17009 , n16654 );
nand ( n17266 , n17264 , n17265 );
buf ( n17267 , n17266 );
xor ( n17268 , n17260 , n17267 );
buf ( n17269 , n17268 );
buf ( n17270 , n17269 );
xor ( n17271 , n16923 , n16940 );
and ( n17272 , n17271 , n16948 );
and ( n17273 , n16923 , n16940 );
or ( n17274 , n17272 , n17273 );
buf ( n17275 , n17274 );
buf ( n17276 , n17275 );
not ( n17277 , n16962 );
not ( n17278 , n10380 );
or ( n17279 , n17277 , n17278 );
buf ( n17280 , n6595 );
buf ( n17281 , n560 );
buf ( n17282 , n545 );
xor ( n17283 , n17281 , n17282 );
buf ( n17284 , n17283 );
buf ( n17285 , n17284 );
nand ( n17286 , n17280 , n17285 );
buf ( n17287 , n17286 );
nand ( n17288 , n17279 , n17287 );
nand ( n17289 , n560 , n547 );
not ( n17290 , n17289 );
and ( n17291 , n17288 , n17290 );
not ( n17292 , n17288 );
and ( n17293 , n17292 , n17289 );
nor ( n17294 , n17291 , n17293 );
not ( n17295 , n562 );
not ( n17296 , n5801 );
or ( n17297 , n17295 , n17296 );
nand ( n17298 , n9798 , n16933 );
nand ( n17299 , n17297 , n17298 );
and ( n17300 , n17294 , n17299 );
not ( n17301 , n17294 );
not ( n17302 , n17299 );
and ( n17303 , n17301 , n17302 );
or ( n17304 , n17300 , n17303 );
buf ( n17305 , n17304 );
xor ( n17306 , n17276 , n17305 );
xor ( n17307 , n16952 , n16969 );
and ( n17308 , n17307 , n16976 );
and ( n17309 , n16952 , n16969 );
or ( n17310 , n17308 , n17309 );
buf ( n17311 , n17310 );
buf ( n17312 , n17311 );
xor ( n17313 , n17306 , n17312 );
buf ( n17314 , n17313 );
buf ( n17315 , n17314 );
xor ( n17316 , n17270 , n17315 );
xor ( n17317 , n17015 , n17019 );
and ( n17318 , n17317 , n17052 );
and ( n17319 , n17015 , n17019 );
or ( n17320 , n17318 , n17319 );
buf ( n17321 , n17320 );
xor ( n17322 , n17316 , n17321 );
buf ( n17323 , n17322 );
buf ( n17324 , n17323 );
xor ( n17325 , n17213 , n17324 );
xor ( n17326 , n16989 , n17054 );
and ( n17327 , n17326 , n17060 );
and ( n17328 , n16989 , n17054 );
or ( n17329 , n17327 , n17328 );
buf ( n17330 , n17329 );
buf ( n17331 , n17330 );
xor ( n17332 , n17325 , n17331 );
buf ( n17333 , n17332 );
buf ( n17334 , n17333 );
not ( n17335 , n17334 );
buf ( n17336 , n17335 );
buf ( n17337 , n17336 );
nand ( n17338 , n17207 , n17337 );
buf ( n17339 , n17338 );
buf ( n17340 , n17336 );
not ( n17341 , n17340 );
buf ( n17342 , n17205 );
nand ( n17343 , n17341 , n17342 );
buf ( n17344 , n17343 );
nand ( n17345 , n17339 , n17344 );
xor ( n17346 , n17200 , n17345 );
not ( n17347 , n17346 );
or ( n17348 , n17167 , n17347 );
not ( n17349 , n17157 );
nor ( n17350 , n17349 , n17148 );
not ( n17351 , n17350 );
not ( n17352 , n16849 );
not ( n17353 , n16776 );
or ( n17354 , n17352 , n17353 );
not ( n17355 , n16835 );
nand ( n17356 , n17355 , n16781 );
nand ( n17357 , n17354 , n17356 );
not ( n17358 , n17357 );
or ( n17359 , n17351 , n17358 );
not ( n17360 , n17159 );
not ( n17361 , n17148 );
and ( n17362 , n17360 , n17361 );
and ( n17363 , n17113 , n17147 );
nor ( n17364 , n17362 , n17363 );
nand ( n17365 , n17359 , n17364 );
xor ( n17366 , n17115 , n17125 );
and ( n17367 , n17366 , n17127 );
and ( n17368 , n17115 , n17125 );
or ( n17369 , n17367 , n17368 );
not ( n17370 , n9417 );
not ( n17371 , n17133 );
or ( n17372 , n17370 , n17371 );
xor ( n17373 , n544 , n15269 );
nand ( n17374 , n17373 , n9409 );
nand ( n17375 , n17372 , n17374 );
and ( n17376 , n17123 , n9575 );
and ( n17377 , n6945 , n546 );
nor ( n17378 , n17376 , n17377 );
xor ( n17379 , n17375 , n17378 );
and ( n17380 , n544 , n16472 );
xor ( n17381 , n17379 , n17380 );
xor ( n17382 , n17369 , n17381 );
xor ( n17383 , n17129 , n17135 );
and ( n17384 , n17383 , n17140 );
and ( n17385 , n17129 , n17135 );
or ( n17386 , n17384 , n17385 );
xor ( n17387 , n17382 , n17386 );
not ( n17388 , n17387 );
xor ( n17389 , n17128 , n17141 );
and ( n17390 , n17389 , n17146 );
and ( n17391 , n17128 , n17141 );
or ( n17392 , n17390 , n17391 );
not ( n17393 , n17392 );
nand ( n17394 , n17388 , n17393 );
or ( n17395 , n17388 , n17393 );
and ( n17396 , n17394 , n17395 );
xor ( n17397 , n17365 , n17396 );
nand ( n17398 , n17190 , n17339 );
not ( n17399 , n17398 );
not ( n17400 , n17399 );
buf ( n17401 , n16143 );
not ( n17402 , n17401 );
or ( n17403 , n17400 , n17402 );
not ( n17404 , n16129 );
nor ( n17405 , n17404 , n17398 );
and ( n17406 , n17405 , n17195 );
not ( n17407 , n17339 );
not ( n17408 , n17185 );
or ( n17409 , n17407 , n17408 );
nand ( n17410 , n17409 , n17344 );
nor ( n17411 , n17406 , n17410 );
nand ( n17412 , n17403 , n17411 );
xor ( n17413 , n17213 , n17324 );
and ( n17414 , n17413 , n17331 );
and ( n17415 , n17213 , n17324 );
or ( n17416 , n17414 , n17415 );
buf ( n17417 , n17416 );
buf ( n17418 , n17417 );
not ( n17419 , n17418 );
xor ( n17420 , n17276 , n17305 );
and ( n17421 , n17420 , n17312 );
and ( n17422 , n17276 , n17305 );
or ( n17423 , n17421 , n17422 );
buf ( n17424 , n17423 );
buf ( n17425 , n17424 );
buf ( n17426 , n17299 );
not ( n17427 , n17290 );
not ( n17428 , n17288 );
or ( n17429 , n17427 , n17428 );
not ( n17430 , n17288 );
nand ( n17431 , n17430 , n17289 );
nand ( n17432 , n17302 , n17431 );
nand ( n17433 , n17429 , n17432 );
buf ( n17434 , n17433 );
xor ( n17435 , n17426 , n17434 );
and ( n17436 , n16959 , n16960 );
buf ( n17437 , n17436 );
buf ( n17438 , n17437 );
or ( n17439 , n5801 , n9798 );
nand ( n17440 , n17439 , n562 );
buf ( n17441 , n17440 );
xor ( n17442 , n17438 , n17441 );
buf ( n17443 , n17284 );
not ( n17444 , n17443 );
buf ( n17445 , n10380 );
not ( n17446 , n17445 );
or ( n17447 , n17444 , n17446 );
buf ( n17448 , n560 );
buf ( n17449 , n544 );
xnor ( n17450 , n17448 , n17449 );
buf ( n17451 , n17450 );
buf ( n17452 , n17451 );
not ( n17453 , n17452 );
buf ( n17454 , n6595 );
nand ( n17455 , n17453 , n17454 );
buf ( n17456 , n17455 );
buf ( n17457 , n17456 );
nand ( n17458 , n17447 , n17457 );
buf ( n17459 , n17458 );
buf ( n17460 , n17459 );
xor ( n17461 , n17442 , n17460 );
buf ( n17462 , n17461 );
buf ( n17463 , n17462 );
xor ( n17464 , n17435 , n17463 );
buf ( n17465 , n17464 );
buf ( n17466 , n17465 );
buf ( n17467 , n17252 );
xor ( n17468 , n17222 , n17239 );
and ( n17469 , n17468 , n17256 );
and ( n17470 , n17222 , n17239 );
or ( n17471 , n17469 , n17470 );
buf ( n17472 , n17471 );
buf ( n17473 , n17472 );
xor ( n17474 , n17467 , n17473 );
and ( n17475 , n17000 , n17001 );
buf ( n17476 , n17475 );
buf ( n17477 , n17476 );
buf ( n17478 , n17232 );
not ( n17479 , n17478 );
buf ( n17480 , n14616 );
not ( n17481 , n17480 );
or ( n17482 , n17479 , n17481 );
buf ( n17483 , n576 );
buf ( n17484 , n544 );
xnor ( n17485 , n17483 , n17484 );
buf ( n17486 , n17485 );
buf ( n17487 , n17486 );
not ( n17488 , n17487 );
buf ( n17489 , n9952 );
nand ( n17490 , n17488 , n17489 );
buf ( n17491 , n17490 );
buf ( n17492 , n17491 );
nand ( n17493 , n17482 , n17492 );
buf ( n17494 , n17493 );
buf ( n17495 , n17494 );
xor ( n17496 , n17477 , n17495 );
buf ( n17497 , n8294 );
buf ( n17498 , n14637 );
or ( n17499 , n17497 , n17498 );
buf ( n17500 , n578 );
nand ( n17501 , n17499 , n17500 );
buf ( n17502 , n17501 );
buf ( n17503 , n17502 );
xor ( n17504 , n17496 , n17503 );
buf ( n17505 , n17504 );
buf ( n17506 , n17505 );
xor ( n17507 , n17474 , n17506 );
buf ( n17508 , n17507 );
buf ( n17509 , n17508 );
xor ( n17510 , n17466 , n17509 );
xor ( n17511 , n17219 , n17259 );
and ( n17512 , n17511 , n17267 );
and ( n17513 , n17219 , n17259 );
or ( n17514 , n17512 , n17513 );
buf ( n17515 , n17514 );
buf ( n17516 , n17515 );
xor ( n17517 , n17510 , n17516 );
buf ( n17518 , n17517 );
buf ( n17519 , n17518 );
xor ( n17520 , n17425 , n17519 );
xor ( n17521 , n17270 , n17315 );
and ( n17522 , n17521 , n17321 );
and ( n17523 , n17270 , n17315 );
or ( n17524 , n17522 , n17523 );
buf ( n17525 , n17524 );
buf ( n17526 , n17525 );
xor ( n17527 , n17520 , n17526 );
buf ( n17528 , n17527 );
buf ( n17529 , n17528 );
not ( n17530 , n17529 );
buf ( n17531 , n17530 );
buf ( n17532 , n17531 );
nand ( n17533 , n17419 , n17532 );
buf ( n17534 , n17533 );
buf ( n17535 , n17534 );
buf ( n17536 , n17531 );
not ( n17537 , n17536 );
buf ( n17538 , n17417 );
nand ( n17539 , n17537 , n17538 );
buf ( n17540 , n17539 );
buf ( n17541 , n17540 );
and ( n17542 , n17535 , n17541 );
buf ( n17543 , n17542 );
xnor ( n17544 , n17412 , n17543 );
nand ( n17545 , n17397 , n17544 );
nand ( n17546 , n17348 , n17545 );
not ( n17547 , n17546 );
buf ( n17548 , n17339 );
buf ( n17549 , n17534 );
and ( n17550 , n17548 , n17549 );
buf ( n17551 , n17550 );
buf ( n17552 , n17551 );
not ( n17553 , n17552 );
buf ( n17554 , n17185 );
not ( n17555 , n17554 );
or ( n17556 , n17553 , n17555 );
buf ( n17557 , n17344 );
not ( n17558 , n17557 );
buf ( n17559 , n17534 );
not ( n17560 , n17559 );
buf ( n17561 , n17560 );
buf ( n17562 , n17561 );
not ( n17563 , n17562 );
and ( n17564 , n17558 , n17563 );
buf ( n17565 , n17540 );
not ( n17566 , n17565 );
buf ( n17567 , n17566 );
buf ( n17568 , n17567 );
nor ( n17569 , n17564 , n17568 );
buf ( n17570 , n17569 );
buf ( n17571 , n17570 );
nand ( n17572 , n17556 , n17571 );
buf ( n17573 , n17572 );
buf ( n17574 , n17573 );
not ( n17575 , n17574 );
buf ( n17576 , n17401 );
buf ( n17577 , n17190 );
buf ( n17578 , n17551 );
and ( n17579 , n17577 , n17578 );
buf ( n17580 , n17579 );
buf ( n17581 , n17580 );
nand ( n17582 , n17576 , n17581 );
buf ( n17583 , n17582 );
buf ( n17584 , n17583 );
buf ( n17585 , n16129 );
buf ( n17586 , n17195 );
buf ( n17587 , n17580 );
nand ( n17588 , n17585 , n17586 , n17587 );
buf ( n17589 , n17588 );
buf ( n17590 , n17589 );
nand ( n17591 , n17575 , n17584 , n17590 );
buf ( n17592 , n17591 );
xor ( n17593 , n17425 , n17519 );
and ( n17594 , n17593 , n17526 );
and ( n17595 , n17425 , n17519 );
or ( n17596 , n17594 , n17595 );
buf ( n17597 , n17596 );
buf ( n17598 , n17597 );
xor ( n17599 , n17426 , n17434 );
and ( n17600 , n17599 , n17463 );
and ( n17601 , n17426 , n17434 );
or ( n17602 , n17600 , n17601 );
buf ( n17603 , n17602 );
buf ( n17604 , n17603 );
buf ( n17605 , n545 );
buf ( n17606 , n560 );
nand ( n17607 , n17605 , n17606 );
buf ( n17608 , n17607 );
buf ( n17609 , n17608 );
buf ( n17610 , n10380 );
not ( n17611 , n17610 );
buf ( n17612 , n17611 );
buf ( n17613 , n17612 );
buf ( n17614 , n17451 );
or ( n17615 , n17613 , n17614 );
buf ( n17616 , n6595 );
not ( n17617 , n17616 );
buf ( n17618 , n17617 );
buf ( n17619 , n17618 );
buf ( n17620 , n7962 );
or ( n17621 , n17619 , n17620 );
nand ( n17622 , n17615 , n17621 );
buf ( n17623 , n17622 );
buf ( n17624 , n17623 );
xor ( n17625 , n17609 , n17624 );
xor ( n17626 , n17438 , n17441 );
and ( n17627 , n17626 , n17460 );
and ( n17628 , n17438 , n17441 );
or ( n17629 , n17627 , n17628 );
buf ( n17630 , n17629 );
buf ( n17631 , n17630 );
xor ( n17632 , n17625 , n17631 );
buf ( n17633 , n17632 );
buf ( n17634 , n17633 );
buf ( n17635 , n545 );
buf ( n17636 , n576 );
nand ( n17637 , n17635 , n17636 );
buf ( n17638 , n17637 );
buf ( n17639 , n17638 );
buf ( n17640 , n14616 );
not ( n17641 , n17640 );
buf ( n17642 , n17641 );
buf ( n17643 , n17642 );
buf ( n17644 , n17486 );
or ( n17645 , n17643 , n17644 );
buf ( n17646 , n9952 );
not ( n17647 , n17646 );
buf ( n17648 , n17647 );
buf ( n17649 , n17648 );
buf ( n17650 , n7809 );
or ( n17651 , n17649 , n17650 );
nand ( n17652 , n17645 , n17651 );
buf ( n17653 , n17652 );
buf ( n17654 , n17653 );
xor ( n17655 , n17639 , n17654 );
xor ( n17656 , n17477 , n17495 );
and ( n17657 , n17656 , n17503 );
and ( n17658 , n17477 , n17495 );
or ( n17659 , n17657 , n17658 );
buf ( n17660 , n17659 );
buf ( n17661 , n17660 );
xor ( n17662 , n17655 , n17661 );
buf ( n17663 , n17662 );
buf ( n17664 , n17663 );
xor ( n17665 , n17634 , n17664 );
xor ( n17666 , n17467 , n17473 );
and ( n17667 , n17666 , n17506 );
and ( n17668 , n17467 , n17473 );
or ( n17669 , n17667 , n17668 );
buf ( n17670 , n17669 );
buf ( n17671 , n17670 );
xor ( n17672 , n17665 , n17671 );
buf ( n17673 , n17672 );
buf ( n17674 , n17673 );
xor ( n17675 , n17604 , n17674 );
xor ( n17676 , n17466 , n17509 );
and ( n17677 , n17676 , n17516 );
and ( n17678 , n17466 , n17509 );
or ( n17679 , n17677 , n17678 );
buf ( n17680 , n17679 );
buf ( n17681 , n17680 );
xor ( n17682 , n17675 , n17681 );
buf ( n17683 , n17682 );
buf ( n17684 , n17683 );
and ( n17685 , n17598 , n17684 );
buf ( n17686 , n17685 );
buf ( n17687 , n17686 );
buf ( n17688 , n17597 );
buf ( n17689 , n17683 );
nor ( n17690 , n17688 , n17689 );
buf ( n17691 , n17690 );
buf ( n17692 , n17691 );
nor ( n17693 , n17687 , n17692 );
buf ( n17694 , n17693 );
not ( n17695 , n17694 );
and ( n17696 , n17592 , n17695 );
not ( n17697 , n17592 );
and ( n17698 , n17697 , n17694 );
or ( n17699 , n17696 , n17698 );
not ( n17700 , n17699 );
nand ( n17701 , n17365 , n17394 );
not ( n17702 , n17701 );
xor ( n17703 , n17369 , n17381 );
and ( n17704 , n17703 , n17386 );
and ( n17705 , n17369 , n17381 );
or ( n17706 , n17704 , n17705 );
not ( n17707 , n17706 );
and ( n17708 , n544 , n15763 );
xor ( n17709 , n17375 , n17378 );
and ( n17710 , n17709 , n17380 );
and ( n17711 , n17375 , n17378 );
or ( n17712 , n17710 , n17711 );
xor ( n17713 , n17708 , n17712 );
or ( n17714 , n9575 , n6945 );
nand ( n17715 , n17714 , n546 );
not ( n17716 , n17373 );
not ( n17717 , n9417 );
or ( n17718 , n17716 , n17717 );
and ( n17719 , n15734 , n544 );
and ( n17720 , n15731 , n8477 );
nor ( n17721 , n17719 , n17720 );
not ( n17722 , n9409 );
or ( n17723 , n17721 , n17722 );
nand ( n17724 , n17718 , n17723 );
xor ( n17725 , n17715 , n17724 );
not ( n17726 , n17378 );
xor ( n17727 , n17725 , n17726 );
xor ( n17728 , n17713 , n17727 );
not ( n17729 , n17728 );
nand ( n17730 , n17707 , n17729 );
not ( n17731 , n17730 );
nor ( n17732 , n17729 , n17707 );
nor ( n17733 , n17731 , n17732 );
and ( n17734 , n17733 , n17395 );
not ( n17735 , n17734 );
or ( n17736 , n17702 , n17735 );
not ( n17737 , n17395 );
not ( n17738 , n17701 );
or ( n17739 , n17737 , n17738 );
not ( n17740 , n17733 );
nand ( n17741 , n17739 , n17740 );
nand ( n17742 , n17736 , n17741 );
nand ( n17743 , n17700 , n17742 );
nand ( n17744 , n17547 , n17743 );
nor ( n17745 , n17109 , n17744 );
not ( n17746 , n17745 );
or ( n17747 , n15710 , n17746 );
not ( n17748 , n17744 );
nand ( n17749 , n16531 , n16536 );
not ( n17750 , n17749 );
not ( n17751 , n16451 );
not ( n17752 , n17751 );
or ( n17753 , n17750 , n17752 );
and ( n17754 , n15805 , n15791 );
not ( n17755 , n15805 );
and ( n17756 , n17755 , n15792 );
nor ( n17757 , n17754 , n17756 );
and ( n17758 , n16145 , n16151 );
not ( n17759 , n16145 );
and ( n17760 , n17759 , n16114 );
nor ( n17761 , n17758 , n17760 );
nand ( n17762 , n17757 , n17761 );
nand ( n17763 , n17753 , n17762 );
buf ( n17764 , n16537 );
nand ( n17765 , n17763 , n17108 , n17764 );
not ( n17766 , n17103 );
not ( n17767 , n17766 );
not ( n17768 , n17104 );
not ( n17769 , n16855 );
or ( n17770 , n17768 , n17769 );
nand ( n17771 , n16854 , n16905 );
nand ( n17772 , n17770 , n17771 );
nand ( n17773 , n17767 , n17772 );
not ( n17774 , n16761 );
nor ( n17775 , n17774 , n16845 );
and ( n17776 , n17773 , n17775 );
nor ( n17777 , n17772 , n17103 );
nor ( n17778 , n17776 , n17777 );
nand ( n17779 , n17765 , n17778 );
buf ( n17780 , n17779 );
and ( n17781 , n17748 , n17780 );
not ( n17782 , n17743 );
nor ( n17783 , n17346 , n17166 );
not ( n17784 , n17783 );
not ( n17785 , n17545 );
or ( n17786 , n17784 , n17785 );
or ( n17787 , n17397 , n17544 );
nand ( n17788 , n17786 , n17787 );
not ( n17789 , n17788 );
or ( n17790 , n17782 , n17789 );
not ( n17791 , n17742 );
nand ( n17792 , n17791 , n17699 );
nand ( n17793 , n17790 , n17792 );
nor ( n17794 , n17781 , n17793 );
nand ( n17795 , n17747 , n17794 );
nand ( n17796 , n17394 , n17730 );
nor ( n17797 , n17148 , n17796 );
not ( n17798 , n17797 );
not ( n17799 , n17160 );
or ( n17800 , n17798 , n17799 );
not ( n17801 , n17394 );
not ( n17802 , n17363 );
or ( n17803 , n17801 , n17802 );
nand ( n17804 , n17803 , n17395 );
and ( n17805 , n17804 , n17730 );
nor ( n17806 , n17805 , n17732 );
nand ( n17807 , n17800 , n17806 );
xor ( n17808 , n17708 , n17712 );
and ( n17809 , n17808 , n17727 );
and ( n17810 , n17708 , n17712 );
or ( n17811 , n17809 , n17810 );
not ( n17812 , n17811 );
and ( n17813 , n544 , n15269 );
not ( n17814 , n17721 );
and ( n17815 , n17814 , n9417 );
and ( n17816 , n9409 , n544 );
nor ( n17817 , n17815 , n17816 );
xor ( n17818 , n17813 , n17817 );
xor ( n17819 , n17715 , n17724 );
and ( n17820 , n17819 , n17726 );
and ( n17821 , n17715 , n17724 );
or ( n17822 , n17820 , n17821 );
xor ( n17823 , n17818 , n17822 );
not ( n17824 , n17823 );
and ( n17825 , n17812 , n17824 );
and ( n17826 , n17811 , n17823 );
nor ( n17827 , n17825 , n17826 );
and ( n17828 , n17807 , n17827 );
not ( n17829 , n17807 );
not ( n17830 , n17827 );
and ( n17831 , n17829 , n17830 );
nor ( n17832 , n17828 , n17831 );
buf ( n17833 , n17551 );
not ( n17834 , n17833 );
buf ( n17835 , n17691 );
nor ( n17836 , n17834 , n17835 );
buf ( n17837 , n17836 );
buf ( n17838 , n17837 );
not ( n17839 , n17838 );
buf ( n17840 , n17185 );
not ( n17841 , n17840 );
or ( n17842 , n17839 , n17841 );
buf ( n17843 , n17570 );
not ( n17844 , n17843 );
buf ( n17845 , n17691 );
not ( n17846 , n17845 );
and ( n17847 , n17844 , n17846 );
buf ( n17848 , n17686 );
nor ( n17849 , n17847 , n17848 );
buf ( n17850 , n17849 );
buf ( n17851 , n17850 );
nand ( n17852 , n17842 , n17851 );
buf ( n17853 , n17852 );
buf ( n17854 , n17853 );
not ( n17855 , n17854 );
buf ( n17856 , n17401 );
buf ( n17857 , n17190 );
buf ( n17858 , n17837 );
and ( n17859 , n17857 , n17858 );
buf ( n17860 , n17859 );
buf ( n17861 , n17860 );
nand ( n17862 , n17856 , n17861 );
buf ( n17863 , n17862 );
buf ( n17864 , n17863 );
buf ( n17865 , n16129 );
buf ( n17866 , n17195 );
buf ( n17867 , n17860 );
nand ( n17868 , n17865 , n17866 , n17867 );
buf ( n17869 , n17868 );
buf ( n17870 , n17869 );
nand ( n17871 , n17855 , n17864 , n17870 );
buf ( n17872 , n17871 );
buf ( n17873 , n544 );
buf ( n17874 , n576 );
nand ( n17875 , n17873 , n17874 );
buf ( n17876 , n17875 );
buf ( n17877 , n17876 );
not ( n17878 , n17877 );
buf ( n17879 , n14616 );
buf ( n17880 , n9952 );
or ( n17881 , n17879 , n17880 );
buf ( n17882 , n576 );
nand ( n17883 , n17881 , n17882 );
buf ( n17884 , n17883 );
buf ( n17885 , n17884 );
not ( n17886 , n17885 );
or ( n17887 , n17878 , n17886 );
buf ( n17888 , n17884 );
buf ( n17889 , n17876 );
or ( n17890 , n17888 , n17889 );
nand ( n17891 , n17887 , n17890 );
buf ( n17892 , n17891 );
buf ( n17893 , n17892 );
buf ( n17894 , n17638 );
xnor ( n17895 , n17893 , n17894 );
buf ( n17896 , n17895 );
buf ( n17897 , n17896 );
not ( n17898 , n17897 );
xor ( n17899 , n17639 , n17654 );
and ( n17900 , n17899 , n17661 );
and ( n17901 , n17639 , n17654 );
or ( n17902 , n17900 , n17901 );
buf ( n17903 , n17902 );
buf ( n17904 , n17903 );
buf ( n17905 , n544 );
buf ( n17906 , n560 );
nand ( n17907 , n17905 , n17906 );
buf ( n17908 , n17907 );
buf ( n17909 , n17908 );
not ( n17910 , n17909 );
buf ( n17911 , n10380 );
buf ( n17912 , n6595 );
or ( n17913 , n17911 , n17912 );
buf ( n17914 , n560 );
nand ( n17915 , n17913 , n17914 );
buf ( n17916 , n17915 );
buf ( n17917 , n17916 );
not ( n17918 , n17917 );
or ( n17919 , n17910 , n17918 );
buf ( n17920 , n17916 );
buf ( n17921 , n17908 );
or ( n17922 , n17920 , n17921 );
nand ( n17923 , n17919 , n17922 );
buf ( n17924 , n17923 );
buf ( n17925 , n17924 );
buf ( n17926 , n17608 );
xnor ( n17927 , n17925 , n17926 );
buf ( n17928 , n17927 );
buf ( n17929 , n17928 );
xnor ( n17930 , n17904 , n17929 );
buf ( n17931 , n17930 );
buf ( n17932 , n17931 );
not ( n17933 , n17932 );
or ( n17934 , n17898 , n17933 );
buf ( n17935 , n17931 );
buf ( n17936 , n17896 );
or ( n17937 , n17935 , n17936 );
nand ( n17938 , n17934 , n17937 );
buf ( n17939 , n17938 );
buf ( n17940 , n17939 );
xor ( n17941 , n17634 , n17664 );
and ( n17942 , n17941 , n17671 );
and ( n17943 , n17634 , n17664 );
or ( n17944 , n17942 , n17943 );
buf ( n17945 , n17944 );
buf ( n17946 , n17945 );
xor ( n17947 , n17609 , n17624 );
and ( n17948 , n17947 , n17631 );
and ( n17949 , n17609 , n17624 );
or ( n17950 , n17948 , n17949 );
buf ( n17951 , n17950 );
buf ( n17952 , n17951 );
xnor ( n17953 , n17946 , n17952 );
buf ( n17954 , n17953 );
buf ( n17955 , n17954 );
xnor ( n17956 , n17940 , n17955 );
buf ( n17957 , n17956 );
buf ( n17958 , n17957 );
not ( n17959 , n17958 );
xor ( n17960 , n17604 , n17674 );
and ( n17961 , n17960 , n17681 );
and ( n17962 , n17604 , n17674 );
or ( n17963 , n17961 , n17962 );
buf ( n17964 , n17963 );
buf ( n17965 , n17964 );
not ( n17966 , n17965 );
or ( n17967 , n17959 , n17966 );
buf ( n17968 , n17964 );
buf ( n17969 , n17957 );
or ( n17970 , n17968 , n17969 );
nand ( n17971 , n17967 , n17970 );
buf ( n17972 , n17971 );
xor ( n17973 , n17872 , n17972 );
nand ( n17974 , n17832 , n17973 );
or ( n17975 , n17832 , n17973 );
nand ( n17976 , n17974 , n17975 );
not ( n17977 , n17976 );
and ( n17978 , n17795 , n17977 );
not ( n17979 , n17795 );
and ( n17980 , n17979 , n17976 );
nor ( n17981 , n17978 , n17980 );
nor ( n17982 , n17109 , n17546 );
not ( n17983 , n17982 );
not ( n17984 , n15709 );
or ( n17985 , n17983 , n17984 );
and ( n17986 , n17779 , n17547 );
nor ( n17987 , n17986 , n17788 );
nand ( n17988 , n17985 , n17987 );
not ( n17989 , n17699 );
nand ( n17990 , n17989 , n17742 );
nand ( n17991 , n17792 , n17990 );
and ( n17992 , n17988 , n17991 );
not ( n17993 , n17988 );
not ( n17994 , n17991 );
and ( n17995 , n17993 , n17994 );
nor ( n17996 , n17992 , n17995 );
not ( n17997 , n17996 );
nand ( n17998 , n17787 , n17545 );
not ( n17999 , n17998 );
nand ( n18000 , n17765 , n17778 );
nand ( n18001 , n17166 , n17346 );
buf ( n18002 , n18001 );
nand ( n18003 , n18000 , n18002 );
buf ( n18004 , n9492 );
and ( n18005 , n15707 , n18004 );
nand ( n18006 , n16845 , n16762 );
and ( n18007 , n16538 , n18001 , n17773 , n18006 );
nand ( n18008 , n18005 , n18007 );
not ( n18009 , n15694 );
not ( n18010 , n15692 );
or ( n18011 , n18009 , n18010 );
not ( n18012 , n15704 );
nand ( n18013 , n18011 , n18012 );
and ( n18014 , n18007 , n18013 );
or ( n18015 , n17166 , n17346 );
not ( n18016 , n18015 );
nor ( n18017 , n18014 , n18016 );
nand ( n18018 , n18003 , n18008 , n18017 );
not ( n18019 , n18018 );
or ( n18020 , n17999 , n18019 );
not ( n18021 , n17998 );
nand ( n18022 , n18003 , n18008 , n18017 , n18021 );
nand ( n18023 , n18020 , n18022 );
and ( n18024 , n18002 , n18015 );
nand ( n18025 , n17765 , n17778 );
not ( n18026 , n18025 );
not ( n18027 , n15694 );
not ( n18028 , n15692 );
or ( n18029 , n18027 , n18028 );
nand ( n18030 , n18029 , n18012 );
not ( n18031 , n17109 );
nand ( n18032 , n18030 , n18031 );
not ( n18033 , n17109 );
nand ( n18034 , n18033 , n15707 , n18004 );
nand ( n18035 , n18026 , n18032 , n18034 );
xor ( n18036 , n18024 , n18035 );
nand ( n18037 , n18023 , n18036 );
not ( n18038 , n18037 );
nand ( n18039 , n15684 , n17981 , n17997 , n18038 );
and ( n18040 , n18006 , n16538 );
nand ( n18041 , n18040 , n18030 );
not ( n18042 , n15689 );
or ( n18043 , n17757 , n17761 );
nand ( n18044 , n18043 , n9492 );
nor ( n18045 , n18042 , n18044 );
not ( n18046 , n18045 );
not ( n18047 , n13699 );
nor ( n18048 , n18047 , n14748 );
not ( n18049 , n18048 );
or ( n18050 , n18046 , n18049 );
not ( n18051 , n17763 );
nand ( n18052 , n18050 , n18051 );
and ( n18053 , n17764 , n18006 );
and ( n18054 , n18052 , n18053 );
nor ( n18055 , n18054 , n17775 );
nand ( n18056 , n18041 , n18055 );
not ( n18057 , n18056 );
not ( n18058 , n17772 );
or ( n18059 , n17766 , n18058 );
not ( n18060 , n17777 );
nand ( n18061 , n18059 , n18060 );
not ( n18062 , n18061 );
not ( n18063 , n18062 );
or ( n18064 , n18057 , n18063 );
nand ( n18065 , n18041 , n18055 , n18061 );
nand ( n18066 , n18064 , n18065 );
not ( n18067 , n18066 );
not ( n18068 , n9492 );
not ( n18069 , n15707 );
or ( n18070 , n18068 , n18069 );
nand ( n18071 , n18070 , n15705 );
buf ( n18072 , n17762 );
buf ( n18073 , n16154 );
buf ( n18074 , n15810 );
nand ( n18075 , n18073 , n18074 );
nand ( n18076 , n18072 , n18075 );
not ( n18077 , n18076 );
and ( n18078 , n18071 , n18077 );
not ( n18079 , n18071 );
and ( n18080 , n18079 , n18076 );
nor ( n18081 , n18078 , n18080 );
buf ( n18082 , n18081 );
nand ( n18083 , n18042 , n15703 );
not ( n18084 , n18083 );
not ( n18085 , n14747 );
not ( n18086 , n13696 );
or ( n18087 , n18085 , n18086 );
nor ( n18088 , n15221 , n15702 );
nand ( n18089 , n18087 , n18088 );
not ( n18090 , n18089 );
or ( n18091 , n18084 , n18090 );
not ( n18092 , n15692 );
not ( n18093 , n18092 );
not ( n18094 , n13700 );
and ( n18095 , n18093 , n18094 );
nor ( n18096 , n18095 , n17763 );
nand ( n18097 , n18091 , n18096 );
not ( n18098 , n18075 );
and ( n18099 , n18051 , n18098 );
not ( n18100 , n17764 );
nor ( n18101 , n18099 , n18100 );
nand ( n18102 , n18097 , n18101 );
not ( n18103 , n17775 );
not ( n18104 , n18006 );
not ( n18105 , n18104 );
nand ( n18106 , n18103 , n18105 );
and ( n18107 , n18102 , n18106 );
not ( n18108 , n18102 );
not ( n18109 , n18106 );
and ( n18110 , n18108 , n18109 );
nor ( n18111 , n18107 , n18110 );
nand ( n18112 , n18089 , n18083 , n18075 );
not ( n18113 , n17751 );
not ( n18114 , n17749 );
or ( n18115 , n18113 , n18114 );
or ( n18116 , n17751 , n17749 );
nand ( n18117 , n18115 , n18116 );
not ( n18118 , n18117 );
nor ( n18119 , n18112 , n18118 );
not ( n18120 , n18119 );
not ( n18121 , n15707 );
nand ( n18122 , n18118 , n18072 );
not ( n18123 , n18122 );
nand ( n18124 , n18121 , n18112 , n18123 );
not ( n18125 , n18044 );
not ( n18126 , n18125 );
nand ( n18127 , n18112 , n18123 , n18126 );
not ( n18128 , n15706 );
nand ( n18129 , n18117 , n18125 );
not ( n18130 , n18129 );
and ( n18131 , n18128 , n18130 );
not ( n18132 , n18072 );
not ( n18133 , n18118 );
and ( n18134 , n18132 , n18133 );
nor ( n18135 , n18131 , n18134 );
nand ( n18136 , n18120 , n18124 , n18127 , n18135 );
buf ( n18137 , n18136 );
nand ( n18138 , n18067 , n18082 , n18111 , n18137 );
not ( n18139 , n18138 );
buf ( n18140 , n9517 );
nand ( n18141 , n18139 , n18140 );
nor ( n18142 , n18039 , n18141 );
not ( n18143 , n18000 );
and ( n18144 , n17990 , n17974 , n17547 );
not ( n18145 , n18144 );
or ( n18146 , n18143 , n18145 );
and ( n18147 , n17788 , n17974 , n17990 );
nand ( n18148 , n17832 , n17973 );
not ( n18149 , n18148 );
not ( n18150 , n17792 );
not ( n18151 , n18150 );
or ( n18152 , n18149 , n18151 );
nand ( n18153 , n18152 , n17975 );
nor ( n18154 , n18147 , n18153 );
nand ( n18155 , n18146 , n18154 );
not ( n18156 , n18155 );
not ( n18157 , n18004 );
not ( n18158 , n15707 );
or ( n18159 , n18157 , n18158 );
not ( n18160 , n18013 );
nand ( n18161 , n18159 , n18160 );
nand ( n18162 , n18144 , n18031 , n18161 );
nand ( n18163 , n18156 , n18162 );
not ( n18164 , n18163 );
buf ( n18165 , n18164 );
buf ( n18166 , n18165 );
buf ( n18167 , n18166 );
buf ( n18168 , n18167 );
not ( n18169 , n18168 );
buf ( n18170 , n18169 );
nor ( n18171 , n18142 , n18170 );
not ( n18172 , n18171 );
nand ( n18173 , n18170 , n18142 );
nand ( n18174 , n18172 , n18173 );
buf ( n18175 , n18174 );
not ( n18176 , n18171 );
not ( n18177 , n18176 );
nand ( n18178 , n15682 , n18082 , n18137 , n18140 );
not ( n18179 , n18109 );
nand ( n18180 , n18097 , n18101 );
not ( n18181 , n18180 );
or ( n18182 , n18179 , n18181 );
nand ( n18183 , n18097 , n18106 , n18101 );
nand ( n18184 , n18182 , n18183 );
buf ( n18185 , n18184 );
not ( n18186 , n18185 );
and ( n18187 , n18178 , n18186 );
not ( n18188 , n18178 );
and ( n18189 , n18188 , n18185 );
nor ( n18190 , n18187 , n18189 );
buf ( n18191 , n18190 );
not ( n18192 , n15681 );
nand ( n18193 , n18192 , n9521 );
not ( n18194 , n18193 );
buf ( n18195 , n18036 );
nand ( n18196 , n18139 , n18194 , n18195 );
not ( n18197 , n18196 );
not ( n18198 , n14256 );
and ( n18199 , n10819 , n13589 );
nand ( n18200 , n18198 , n18199 );
not ( n18201 , n18200 );
nand ( n18202 , n18201 , n9521 );
buf ( n18203 , n14254 );
buf ( n18204 , n18203 );
nand ( n18205 , n18201 , n18204 , n9521 );
buf ( n18206 , n15655 );
not ( n18207 , n15667 );
not ( n18208 , n18207 );
nand ( n18209 , n18206 , n18208 );
nand ( n18210 , n15680 , n18203 );
nor ( n18211 , n18209 , n18210 );
and ( n18212 , n18137 , n18211 );
nand ( n18213 , n15680 , n18203 );
buf ( n18214 , n17314 );
buf ( n18215 , n17212 );
nand ( n18216 , n6843 , n579 );
nand ( n18217 , n7578 , n580 );
nand ( n18218 , n18216 , n18217 );
buf ( n18219 , n18218 );
buf ( n18220 , n18219 );
not ( n18221 , n18220 );
buf ( n18222 , n578 );
not ( n18223 , n18222 );
buf ( n18224 , n10184 );
not ( n18225 , n18224 );
buf ( n18226 , n18225 );
buf ( n18227 , n18226 );
not ( n18228 , n18227 );
or ( n18229 , n18223 , n18228 );
buf ( n18230 , n10854 );
buf ( n18231 , n578 );
not ( n18232 , n18231 );
buf ( n18233 , n18232 );
buf ( n18234 , n18233 );
nand ( n18235 , n18230 , n18234 );
buf ( n18236 , n18235 );
buf ( n18237 , n18236 );
nand ( n18238 , n18229 , n18237 );
buf ( n18239 , n18238 );
buf ( n18240 , n18239 );
not ( n18241 , n18240 );
or ( n18242 , n18221 , n18241 );
buf ( n18243 , n578 );
not ( n18244 , n18243 );
buf ( n18245 , n9498 );
not ( n18246 , n18245 );
or ( n18247 , n18244 , n18246 );
buf ( n18248 , n9497 );
buf ( n18249 , n18233 );
nand ( n18250 , n18248 , n18249 );
buf ( n18251 , n18250 );
buf ( n18252 , n18251 );
nand ( n18253 , n18247 , n18252 );
buf ( n18254 , n18253 );
buf ( n18255 , n18254 );
buf ( n18256 , n578 );
buf ( n18257 , n579 );
nor ( n18258 , n18256 , n18257 );
buf ( n18259 , n18258 );
not ( n18260 , n18259 );
and ( n18261 , n578 , n579 );
nor ( n18262 , n18261 , n18219 );
nand ( n18263 , n18260 , n18262 );
not ( n18264 , n18263 );
buf ( n18265 , n18264 );
nand ( n18266 , n18255 , n18265 );
buf ( n18267 , n18266 );
buf ( n18268 , n18267 );
nand ( n18269 , n18242 , n18268 );
buf ( n18270 , n18269 );
buf ( n18271 , n18270 );
buf ( n18272 , n4783 );
buf ( n18273 , n584 );
or ( n18274 , n18272 , n18273 );
buf ( n18275 , n584 );
not ( n18276 , n18275 );
buf ( n18277 , n18276 );
buf ( n18278 , n18277 );
buf ( n18279 , n583 );
or ( n18280 , n18278 , n18279 );
nand ( n18281 , n18274 , n18280 );
buf ( n18282 , n18281 );
buf ( n18283 , n18282 );
buf ( n18284 , n18283 );
buf ( n18285 , n18284 );
buf ( n18286 , n18285 );
not ( n18287 , n18286 );
xor ( n18288 , n582 , n15680 );
buf ( n18289 , n18288 );
not ( n18290 , n18289 );
or ( n18291 , n18287 , n18290 );
buf ( n18292 , n582 );
not ( n18293 , n18292 );
buf ( n18294 , n18203 );
not ( n18295 , n18294 );
buf ( n18296 , n18295 );
buf ( n18297 , n18296 );
not ( n18298 , n18297 );
or ( n18299 , n18293 , n18298 );
buf ( n18300 , n18203 );
buf ( n18301 , n582 );
not ( n18302 , n18301 );
buf ( n18303 , n18302 );
buf ( n18304 , n18303 );
nand ( n18305 , n18300 , n18304 );
buf ( n18306 , n18305 );
buf ( n18307 , n18306 );
nand ( n18308 , n18299 , n18307 );
buf ( n18309 , n18308 );
buf ( n18310 , n18309 );
not ( n18311 , n18282 );
and ( n18312 , n582 , n583 );
and ( n18313 , n18303 , n4783 );
nor ( n18314 , n18312 , n18313 );
nand ( n18315 , n18311 , n18314 );
not ( n18316 , n18315 );
buf ( n18317 , n18316 );
nand ( n18318 , n18310 , n18317 );
buf ( n18319 , n18318 );
buf ( n18320 , n18319 );
nand ( n18321 , n18291 , n18320 );
buf ( n18322 , n18321 );
buf ( n18323 , n18322 );
xor ( n18324 , n18271 , n18323 );
buf ( n18325 , n576 );
nand ( n18326 , n7546 , n7549 );
buf ( n18327 , n18326 );
not ( n18328 , n18327 );
buf ( n18329 , n18328 );
buf ( n18330 , n18329 );
not ( n18331 , n18330 );
buf ( n18332 , n18331 );
buf ( n18333 , n18332 );
and ( n18334 , n18325 , n18333 );
buf ( n18335 , n18334 );
buf ( n18336 , n18335 );
buf ( n18337 , n577 );
buf ( n18338 , n578 );
xor ( n18339 , n18337 , n18338 );
buf ( n18340 , n18339 );
buf ( n18341 , n18340 );
not ( n18342 , n18341 );
buf ( n18343 , n576 );
buf ( n18344 , n8542 );
buf ( n18345 , n18344 );
xor ( n18346 , n18343 , n18345 );
buf ( n18347 , n18346 );
buf ( n18348 , n18347 );
not ( n18349 , n18348 );
or ( n18350 , n18342 , n18349 );
buf ( n18351 , n576 );
not ( n18352 , n7375 );
not ( n18353 , n7467 );
or ( n18354 , n18352 , n18353 );
nand ( n18355 , n18354 , n7471 );
not ( n18356 , n18355 );
not ( n18357 , n18356 );
buf ( n18358 , n18357 );
xor ( n18359 , n18351 , n18358 );
buf ( n18360 , n18359 );
buf ( n18361 , n18360 );
and ( n18362 , n576 , n577 );
nor ( n18363 , n18362 , n18340 );
or ( n18364 , n576 , n577 );
and ( n18365 , n18363 , n18364 );
buf ( n18366 , n18365 );
nand ( n18367 , n18361 , n18366 );
buf ( n18368 , n18367 );
buf ( n18369 , n18368 );
nand ( n18370 , n18350 , n18369 );
buf ( n18371 , n18370 );
buf ( n18372 , n18371 );
xor ( n18373 , n18336 , n18372 );
buf ( n18374 , n580 );
buf ( n18375 , n581 );
and ( n18376 , n18374 , n18375 );
and ( n18377 , n581 , n582 );
not ( n18378 , n581 );
and ( n18379 , n18378 , n18303 );
nor ( n18380 , n18377 , n18379 );
buf ( n18381 , n18380 );
buf ( n18382 , n580 );
buf ( n18383 , n581 );
nor ( n18384 , n18382 , n18383 );
buf ( n18385 , n18384 );
buf ( n18386 , n18385 );
nor ( n18387 , n18376 , n18381 , n18386 );
buf ( n18388 , n18387 );
buf ( n18389 , n18388 );
buf ( n18390 , n18389 );
buf ( n18391 , n18390 );
buf ( n18392 , n18391 );
not ( n18393 , n18392 );
not ( n18394 , n580 );
buf ( n18395 , n10819 );
not ( n18396 , n18395 );
buf ( n18397 , n18396 );
not ( n18398 , n18397 );
or ( n18399 , n18394 , n18398 );
buf ( n18400 , n580 );
not ( n18401 , n18400 );
buf ( n18402 , n18401 );
nand ( n18403 , n18402 , n10819 );
nand ( n18404 , n18399 , n18403 );
not ( n18405 , n18404 );
or ( n18406 , n18393 , n18405 );
buf ( n18407 , n13589 );
not ( n18408 , n18407 );
buf ( n18409 , n18408 );
nand ( n18410 , n18409 , n580 );
not ( n18411 , n18410 );
buf ( n18412 , n13592 );
buf ( n18413 , n18402 );
nand ( n18414 , n18412 , n18413 );
buf ( n18415 , n18414 );
not ( n18416 , n18415 );
or ( n18417 , n18411 , n18416 );
buf ( n18418 , n18380 );
nand ( n18419 , n18417 , n18418 );
nand ( n18420 , n18406 , n18419 );
buf ( n18421 , n18420 );
xor ( n18422 , n18373 , n18421 );
buf ( n18423 , n18422 );
buf ( n18424 , n18423 );
xor ( n18425 , n18324 , n18424 );
buf ( n18426 , n18425 );
buf ( n18427 , n18426 );
buf ( n18428 , n585 );
buf ( n18429 , n586 );
xor ( n18430 , n18428 , n18429 );
buf ( n18431 , n18430 );
buf ( n18432 , n18431 );
not ( n18433 , n18432 );
buf ( n18434 , n584 );
not ( n18435 , n18434 );
not ( n18436 , n15657 );
not ( n18437 , n15663 );
or ( n18438 , n18436 , n18437 );
nand ( n18439 , n18438 , n15666 );
buf ( n18440 , n18439 );
not ( n18441 , n18440 );
buf ( n18442 , n18441 );
buf ( n18443 , n18442 );
not ( n18444 , n18443 );
or ( n18445 , n18435 , n18444 );
nand ( n18446 , n15667 , n18277 );
buf ( n18447 , n18446 );
nand ( n18448 , n18445 , n18447 );
buf ( n18449 , n18448 );
buf ( n18450 , n18449 );
not ( n18451 , n18450 );
or ( n18452 , n18433 , n18451 );
buf ( n18453 , n584 );
not ( n18454 , n18453 );
buf ( n18455 , n15680 );
not ( n18456 , n18455 );
buf ( n18457 , n18456 );
buf ( n18458 , n18457 );
not ( n18459 , n18458 );
or ( n18460 , n18454 , n18459 );
buf ( n18461 , n15680 );
buf ( n18462 , n18277 );
nand ( n18463 , n18461 , n18462 );
buf ( n18464 , n18463 );
buf ( n18465 , n18464 );
nand ( n18466 , n18460 , n18465 );
buf ( n18467 , n18466 );
buf ( n18468 , n18467 );
buf ( n18469 , n584 );
buf ( n18470 , n585 );
and ( n18471 , n18469 , n18470 );
buf ( n18472 , n18431 );
buf ( n18473 , n584 );
buf ( n18474 , n585 );
nor ( n18475 , n18473 , n18474 );
buf ( n18476 , n18475 );
buf ( n18477 , n18476 );
nor ( n18478 , n18471 , n18472 , n18477 );
buf ( n18479 , n18478 );
buf ( n18480 , n18479 );
nand ( n18481 , n18468 , n18480 );
buf ( n18482 , n18481 );
buf ( n18483 , n18482 );
nand ( n18484 , n18452 , n18483 );
buf ( n18485 , n18484 );
buf ( n18486 , n18485 );
buf ( n18487 , n576 );
not ( n18488 , n18487 );
buf ( n18489 , n7541 );
buf ( n18490 , n18489 );
not ( n18491 , n18490 );
buf ( n18492 , n18491 );
buf ( n18493 , n18492 );
buf ( n18494 , n18493 );
nor ( n18495 , n18488 , n18494 );
buf ( n18496 , n18495 );
buf ( n18497 , n18496 );
buf ( n18498 , n18340 );
not ( n18499 , n18498 );
buf ( n18500 , n18360 );
not ( n18501 , n18500 );
or ( n18502 , n18499 , n18501 );
xor ( n18503 , n18325 , n18333 );
buf ( n18504 , n18503 );
buf ( n18505 , n18504 );
buf ( n18506 , n18365 );
nand ( n18507 , n18505 , n18506 );
buf ( n18508 , n18507 );
buf ( n18509 , n18508 );
nand ( n18510 , n18502 , n18509 );
buf ( n18511 , n18510 );
buf ( n18512 , n18511 );
xor ( n18513 , n18497 , n18512 );
buf ( n18514 , n18392 );
not ( n18515 , n18514 );
and ( n18516 , n10184 , n18402 );
not ( n18517 , n10184 );
and ( n18518 , n18517 , n580 );
or ( n18519 , n18516 , n18518 );
buf ( n18520 , n18519 );
not ( n18521 , n18520 );
or ( n18522 , n18515 , n18521 );
buf ( n18523 , n18380 );
not ( n18524 , n18523 );
buf ( n18525 , n18524 );
not ( n18526 , n18525 );
nand ( n18527 , n18526 , n18404 );
buf ( n18528 , n18527 );
nand ( n18529 , n18522 , n18528 );
buf ( n18530 , n18529 );
buf ( n18531 , n18530 );
xor ( n18532 , n18513 , n18531 );
buf ( n18533 , n18532 );
buf ( n18534 , n18533 );
xor ( n18535 , n18486 , n18534 );
buf ( n18536 , n13665 );
not ( n18537 , n18536 );
buf ( n18538 , n18537 );
buf ( n18539 , n18538 );
not ( n18540 , n18539 );
buf ( n18541 , n18540 );
buf ( n18542 , n18541 );
buf ( n18543 , n576 );
and ( n18544 , n18542 , n18543 );
buf ( n18545 , n18544 );
buf ( n18546 , n18545 );
buf ( n18547 , n18340 );
not ( n18548 , n18547 );
buf ( n18549 , n576 );
not ( n18550 , n18549 );
buf ( n18551 , n18492 );
not ( n18552 , n18551 );
or ( n18553 , n18550 , n18552 );
buf ( n18554 , n18489 );
buf ( n18555 , n7809 );
nand ( n18556 , n18554 , n18555 );
buf ( n18557 , n18556 );
buf ( n18558 , n18557 );
nand ( n18559 , n18553 , n18558 );
buf ( n18560 , n18559 );
buf ( n18561 , n18560 );
not ( n18562 , n18561 );
or ( n18563 , n18548 , n18562 );
buf ( n18564 , n576 );
not ( n18565 , n18564 );
buf ( n18566 , n5363 );
buf ( n18567 , n18566 );
not ( n18568 , n18567 );
buf ( n18569 , n18568 );
buf ( n18570 , n18569 );
not ( n18571 , n18570 );
or ( n18572 , n18565 , n18571 );
buf ( n18573 , n18566 );
buf ( n18574 , n7809 );
nand ( n18575 , n18573 , n18574 );
buf ( n18576 , n18575 );
buf ( n18577 , n18576 );
nand ( n18578 , n18572 , n18577 );
buf ( n18579 , n18578 );
buf ( n18580 , n18579 );
buf ( n18581 , n18365 );
nand ( n18582 , n18580 , n18581 );
buf ( n18583 , n18582 );
buf ( n18584 , n18583 );
nand ( n18585 , n18563 , n18584 );
buf ( n18586 , n18585 );
buf ( n18587 , n18586 );
xor ( n18588 , n18546 , n18587 );
buf ( n18589 , n18219 );
not ( n18590 , n18589 );
xor ( n18591 , n578 , n18355 );
buf ( n18592 , n18591 );
not ( n18593 , n18592 );
or ( n18594 , n18590 , n18593 );
buf ( n18595 , n578 );
not ( n18596 , n18595 );
buf ( n18597 , n18326 );
not ( n18598 , n18597 );
buf ( n18599 , n18598 );
buf ( n18600 , n18599 );
not ( n18601 , n18600 );
or ( n18602 , n18596 , n18601 );
buf ( n18603 , n18599 );
not ( n18604 , n18603 );
buf ( n18605 , n18604 );
buf ( n18606 , n18605 );
buf ( n18607 , n18233 );
nand ( n18608 , n18606 , n18607 );
buf ( n18609 , n18608 );
buf ( n18610 , n18609 );
nand ( n18611 , n18602 , n18610 );
buf ( n18612 , n18611 );
buf ( n18613 , n18612 );
buf ( n18614 , n18264 );
nand ( n18615 , n18613 , n18614 );
buf ( n18616 , n18615 );
buf ( n18617 , n18616 );
nand ( n18618 , n18594 , n18617 );
buf ( n18619 , n18618 );
buf ( n18620 , n18619 );
and ( n18621 , n18588 , n18620 );
and ( n18622 , n18546 , n18587 );
or ( n18623 , n18621 , n18622 );
buf ( n18624 , n18623 );
buf ( n18625 , n18624 );
buf ( n18626 , n18418 );
not ( n18627 , n18626 );
buf ( n18628 , n18519 );
not ( n18629 , n18628 );
or ( n18630 , n18627 , n18629 );
buf ( n18631 , n580 );
not ( n18632 , n18631 );
buf ( n18633 , n9497 );
not ( n18634 , n18633 );
buf ( n18635 , n18634 );
buf ( n18636 , n18635 );
not ( n18637 , n18636 );
or ( n18638 , n18632 , n18637 );
buf ( n18639 , n9497 );
buf ( n18640 , n18402 );
nand ( n18641 , n18639 , n18640 );
buf ( n18642 , n18641 );
buf ( n18643 , n18642 );
nand ( n18644 , n18638 , n18643 );
buf ( n18645 , n18644 );
buf ( n18646 , n18645 );
buf ( n18647 , n18392 );
nand ( n18648 , n18646 , n18647 );
buf ( n18649 , n18648 );
buf ( n18650 , n18649 );
nand ( n18651 , n18630 , n18650 );
buf ( n18652 , n18651 );
buf ( n18653 , n18652 );
xor ( n18654 , n18625 , n18653 );
buf ( n18655 , n18285 );
buf ( n18656 , n18655 );
buf ( n18657 , n18656 );
buf ( n18658 , n18657 );
not ( n18659 , n18658 );
buf ( n18660 , n582 );
not ( n18661 , n18660 );
buf ( n18662 , n13600 );
not ( n18663 , n18662 );
or ( n18664 , n18661 , n18663 );
buf ( n18665 , n18409 );
not ( n18666 , n18665 );
buf ( n18667 , n18666 );
buf ( n18668 , n18667 );
buf ( n18669 , n18303 );
nand ( n18670 , n18668 , n18669 );
buf ( n18671 , n18670 );
buf ( n18672 , n18671 );
nand ( n18673 , n18664 , n18672 );
buf ( n18674 , n18673 );
buf ( n18675 , n18674 );
not ( n18676 , n18675 );
or ( n18677 , n18659 , n18676 );
buf ( n18678 , n582 );
not ( n18679 , n18678 );
buf ( n18680 , n10819 );
not ( n18681 , n18680 );
buf ( n18682 , n18681 );
buf ( n18683 , n18682 );
not ( n18684 , n18683 );
or ( n18685 , n18679 , n18684 );
nand ( n18686 , n10819 , n18303 );
buf ( n18687 , n18686 );
nand ( n18688 , n18685 , n18687 );
buf ( n18689 , n18688 );
buf ( n18690 , n18689 );
buf ( n18691 , n18316 );
nand ( n18692 , n18690 , n18691 );
buf ( n18693 , n18692 );
buf ( n18694 , n18693 );
nand ( n18695 , n18677 , n18694 );
buf ( n18696 , n18695 );
buf ( n18697 , n18696 );
and ( n18698 , n18654 , n18697 );
and ( n18699 , n18625 , n18653 );
or ( n18700 , n18698 , n18699 );
buf ( n18701 , n18700 );
buf ( n18702 , n18701 );
and ( n18703 , n18535 , n18702 );
and ( n18704 , n18486 , n18534 );
or ( n18705 , n18703 , n18704 );
buf ( n18706 , n18705 );
buf ( n18707 , n18706 );
xor ( n18708 , n18427 , n18707 );
xor ( n18709 , n18497 , n18512 );
and ( n18710 , n18709 , n18531 );
and ( n18711 , n18497 , n18512 );
or ( n18712 , n18710 , n18711 );
buf ( n18713 , n18712 );
buf ( n18714 , n18713 );
buf ( n18715 , n18431 );
not ( n18716 , n18715 );
buf ( n18717 , n584 );
not ( n18718 , n18717 );
nand ( n18719 , n15209 , n15227 );
not ( n18720 , n15654 );
and ( n18721 , n18719 , n18720 );
not ( n18722 , n18719 );
and ( n18723 , n18722 , n15654 );
nor ( n18724 , n18721 , n18723 );
buf ( n18725 , n18724 );
not ( n18726 , n18725 );
buf ( n18727 , n18726 );
not ( n18728 , n18727 );
or ( n18729 , n18718 , n18728 );
buf ( n18730 , n18725 );
buf ( n18731 , n18277 );
nand ( n18732 , n18730 , n18731 );
buf ( n18733 , n18732 );
buf ( n18734 , n18733 );
nand ( n18735 , n18729 , n18734 );
buf ( n18736 , n18735 );
buf ( n18737 , n18736 );
not ( n18738 , n18737 );
or ( n18739 , n18716 , n18738 );
buf ( n18740 , n18449 );
buf ( n18741 , n18479 );
nand ( n18742 , n18740 , n18741 );
buf ( n18743 , n18742 );
buf ( n18744 , n18743 );
nand ( n18745 , n18739 , n18744 );
buf ( n18746 , n18745 );
buf ( n18747 , n18746 );
xor ( n18748 , n18714 , n18747 );
buf ( n18749 , n18219 );
not ( n18750 , n18749 );
buf ( n18751 , n18254 );
not ( n18752 , n18751 );
or ( n18753 , n18750 , n18752 );
buf ( n18754 , n578 );
not ( n18755 , n18754 );
buf ( n18756 , n8543 );
not ( n18757 , n18756 );
or ( n18758 , n18755 , n18757 );
not ( n18759 , n8543 );
buf ( n18760 , n18759 );
buf ( n18761 , n18233 );
nand ( n18762 , n18760 , n18761 );
buf ( n18763 , n18762 );
buf ( n18764 , n18763 );
nand ( n18765 , n18758 , n18764 );
buf ( n18766 , n18765 );
buf ( n18767 , n18766 );
buf ( n18768 , n18264 );
nand ( n18769 , n18767 , n18768 );
buf ( n18770 , n18769 );
buf ( n18771 , n18770 );
nand ( n18772 , n18753 , n18771 );
buf ( n18773 , n18772 );
buf ( n18774 , n18773 );
buf ( n18775 , n18285 );
not ( n18776 , n18775 );
buf ( n18777 , n18309 );
not ( n18778 , n18777 );
or ( n18779 , n18776 , n18778 );
buf ( n18780 , n18674 );
buf ( n18781 , n18316 );
nand ( n18782 , n18780 , n18781 );
buf ( n18783 , n18782 );
buf ( n18784 , n18783 );
nand ( n18785 , n18779 , n18784 );
buf ( n18786 , n18785 );
buf ( n18787 , n18786 );
xor ( n18788 , n18774 , n18787 );
buf ( n18789 , n18566 );
buf ( n18790 , n576 );
and ( n18791 , n18789 , n18790 );
buf ( n18792 , n18791 );
buf ( n18793 , n18792 );
buf ( n18794 , n18340 );
not ( n18795 , n18794 );
buf ( n18796 , n18504 );
not ( n18797 , n18796 );
or ( n18798 , n18795 , n18797 );
buf ( n18799 , n18560 );
buf ( n18800 , n18365 );
nand ( n18801 , n18799 , n18800 );
buf ( n18802 , n18801 );
buf ( n18803 , n18802 );
nand ( n18804 , n18798 , n18803 );
buf ( n18805 , n18804 );
buf ( n18806 , n18805 );
xor ( n18807 , n18793 , n18806 );
buf ( n18808 , n18219 );
not ( n18809 , n18808 );
buf ( n18810 , n18766 );
not ( n18811 , n18810 );
or ( n18812 , n18809 , n18811 );
buf ( n18813 , n18591 );
buf ( n18814 , n18264 );
nand ( n18815 , n18813 , n18814 );
buf ( n18816 , n18815 );
buf ( n18817 , n18816 );
nand ( n18818 , n18812 , n18817 );
buf ( n18819 , n18818 );
buf ( n18820 , n18819 );
and ( n18821 , n18807 , n18820 );
and ( n18822 , n18793 , n18806 );
or ( n18823 , n18821 , n18822 );
buf ( n18824 , n18823 );
buf ( n18825 , n18824 );
and ( n18826 , n18788 , n18825 );
and ( n18827 , n18774 , n18787 );
or ( n18828 , n18826 , n18827 );
buf ( n18829 , n18828 );
buf ( n18830 , n18829 );
xor ( n18831 , n18748 , n18830 );
buf ( n18832 , n18831 );
buf ( n18833 , n18832 );
xor ( n18834 , n18708 , n18833 );
buf ( n18835 , n18834 );
buf ( n18836 , n18835 );
buf ( n18837 , n18725 );
buf ( n18838 , n586 );
not ( n18839 , n18838 );
buf ( n18840 , n18839 );
buf ( n18841 , n18840 );
nand ( n18842 , n18837 , n18841 );
buf ( n18843 , n18842 );
not ( n18844 , n18843 );
not ( n18845 , n18725 );
nand ( n18846 , n18845 , n586 );
not ( n18847 , n18846 );
or ( n18848 , n18844 , n18847 );
not ( n18849 , n588 );
and ( n18850 , n587 , n18849 );
not ( n18851 , n587 );
and ( n18852 , n18851 , n588 );
or ( n18853 , n18850 , n18852 );
buf ( n18854 , n18853 );
not ( n18855 , n18854 );
buf ( n18856 , n18855 );
not ( n18857 , n18856 );
nand ( n18858 , n18848 , n18857 );
buf ( n18859 , n18442 );
not ( n18860 , n18859 );
buf ( n18861 , n18860 );
buf ( n18862 , n18861 );
buf ( n18863 , n18840 );
nand ( n18864 , n18862 , n18863 );
buf ( n18865 , n18864 );
buf ( n18866 , n18439 );
not ( n18867 , n18866 );
buf ( n18868 , n18867 );
nand ( n18869 , n18868 , n586 );
nand ( n18870 , n18865 , n18869 );
buf ( n18871 , n586 );
buf ( n18872 , n587 );
and ( n18873 , n18871 , n18872 );
buf ( n18874 , n18853 );
buf ( n18875 , n586 );
buf ( n18876 , n587 );
nor ( n18877 , n18875 , n18876 );
buf ( n18878 , n18877 );
buf ( n18879 , n18878 );
nor ( n18880 , n18873 , n18874 , n18879 );
buf ( n18881 , n18880 );
buf ( n18882 , n18881 );
nand ( n18883 , n18870 , n18882 );
nand ( n18884 , n18858 , n18883 );
buf ( n18885 , n18884 );
buf ( n18886 , n18657 );
not ( n18887 , n18886 );
buf ( n18888 , n18689 );
not ( n18889 , n18888 );
or ( n18890 , n18887 , n18889 );
not ( n18891 , n582 );
buf ( n18892 , n10184 );
not ( n18893 , n18892 );
buf ( n18894 , n18893 );
not ( n18895 , n18894 );
or ( n18896 , n18891 , n18895 );
buf ( n18897 , n10184 );
buf ( n18898 , n18303 );
nand ( n18899 , n18897 , n18898 );
buf ( n18900 , n18899 );
nand ( n18901 , n18896 , n18900 );
nand ( n18902 , n18901 , n18316 );
buf ( n18903 , n18902 );
nand ( n18904 , n18890 , n18903 );
buf ( n18905 , n18904 );
buf ( n18906 , n18905 );
buf ( n18907 , n18203 );
buf ( n18908 , n18907 );
buf ( n18909 , n18908 );
buf ( n18910 , n18431 );
not ( n18911 , n18910 );
buf ( n18912 , n18911 );
buf ( n18913 , n18912 );
buf ( n18914 , n18277 );
nor ( n18915 , n18913 , n18914 );
buf ( n18916 , n18915 );
not ( n18917 , n18916 );
nor ( n18918 , n18909 , n18917 );
not ( n18919 , n18918 );
buf ( n18920 , n584 );
not ( n18921 , n18920 );
buf ( n18922 , n18409 );
not ( n18923 , n18922 );
or ( n18924 , n18921 , n18923 );
buf ( n18925 , n13592 );
buf ( n18926 , n18277 );
nand ( n18927 , n18925 , n18926 );
buf ( n18928 , n18927 );
buf ( n18929 , n18928 );
nand ( n18930 , n18924 , n18929 );
buf ( n18931 , n18930 );
nand ( n18932 , n18931 , n18479 );
buf ( n18933 , n18912 );
buf ( n18934 , n584 );
nor ( n18935 , n18933 , n18934 );
buf ( n18936 , n18935 );
nand ( n18937 , n18909 , n18936 );
nand ( n18938 , n18919 , n18932 , n18937 );
buf ( n18939 , n18938 );
xor ( n18940 , n18906 , n18939 );
buf ( n18941 , n18418 );
not ( n18942 , n18941 );
buf ( n18943 , n580 );
not ( n18944 , n18943 );
buf ( n18945 , n8543 );
not ( n18946 , n18945 );
or ( n18947 , n18944 , n18946 );
buf ( n18948 , n8542 );
buf ( n18949 , n18402 );
nand ( n18950 , n18948 , n18949 );
buf ( n18951 , n18950 );
buf ( n18952 , n18951 );
nand ( n18953 , n18947 , n18952 );
buf ( n18954 , n18953 );
buf ( n18955 , n18954 );
not ( n18956 , n18955 );
or ( n18957 , n18942 , n18956 );
buf ( n18958 , n580 );
not ( n18959 , n18958 );
not ( n18960 , n18355 );
buf ( n18961 , n18960 );
not ( n18962 , n18961 );
or ( n18963 , n18959 , n18962 );
buf ( n18964 , n18357 );
buf ( n18965 , n18402 );
nand ( n18966 , n18964 , n18965 );
buf ( n18967 , n18966 );
buf ( n18968 , n18967 );
nand ( n18969 , n18963 , n18968 );
buf ( n18970 , n18969 );
buf ( n18971 , n18970 );
buf ( n18972 , n18391 );
nand ( n18973 , n18971 , n18972 );
buf ( n18974 , n18973 );
buf ( n18975 , n18974 );
nand ( n18976 , n18957 , n18975 );
buf ( n18977 , n18976 );
buf ( n18978 , n18977 );
buf ( n18979 , n13663 );
not ( n18980 , n18979 );
buf ( n18981 , n18980 );
buf ( n18982 , n18981 );
buf ( n18983 , n7809 );
nor ( n18984 , n18982 , n18983 );
buf ( n18985 , n18984 );
buf ( n18986 , n18985 );
buf ( n18987 , n18340 );
not ( n18988 , n18987 );
and ( n18989 , n18541 , n7809 );
not ( n18990 , n18541 );
and ( n18991 , n18990 , n576 );
or ( n18992 , n18989 , n18991 );
buf ( n18993 , n18992 );
not ( n18994 , n18993 );
or ( n18995 , n18988 , n18994 );
buf ( n18996 , n576 );
nand ( n18997 , n4775 , n4776 );
buf ( n18998 , n18997 );
not ( n18999 , n18998 );
buf ( n19000 , n18999 );
buf ( n19001 , n19000 );
not ( n19002 , n19001 );
buf ( n19003 , n19002 );
buf ( n19004 , n19003 );
xor ( n19005 , n18996 , n19004 );
buf ( n19006 , n19005 );
buf ( n19007 , n19006 );
buf ( n19008 , n18365 );
nand ( n19009 , n19007 , n19008 );
buf ( n19010 , n19009 );
buf ( n19011 , n19010 );
nand ( n19012 , n18995 , n19011 );
buf ( n19013 , n19012 );
buf ( n19014 , n19013 );
xor ( n19015 , n18986 , n19014 );
buf ( n19016 , n18219 );
not ( n19017 , n19016 );
buf ( n19018 , n578 );
not ( n19019 , n19018 );
buf ( n19020 , n18489 );
not ( n19021 , n19020 );
buf ( n19022 , n19021 );
buf ( n19023 , n19022 );
not ( n19024 , n19023 );
or ( n19025 , n19019 , n19024 );
buf ( n19026 , n18492 );
not ( n19027 , n19026 );
buf ( n19028 , n18233 );
nand ( n19029 , n19027 , n19028 );
buf ( n19030 , n19029 );
buf ( n19031 , n19030 );
nand ( n19032 , n19025 , n19031 );
buf ( n19033 , n19032 );
buf ( n19034 , n19033 );
not ( n19035 , n19034 );
or ( n19036 , n19017 , n19035 );
buf ( n19037 , n578 );
not ( n19038 , n19037 );
buf ( n19039 , n18569 );
not ( n19040 , n19039 );
or ( n19041 , n19038 , n19040 );
buf ( n19042 , n18566 );
buf ( n19043 , n18233 );
nand ( n19044 , n19042 , n19043 );
buf ( n19045 , n19044 );
buf ( n19046 , n19045 );
nand ( n19047 , n19041 , n19046 );
buf ( n19048 , n19047 );
buf ( n19049 , n19048 );
buf ( n19050 , n18264 );
nand ( n19051 , n19049 , n19050 );
buf ( n19052 , n19051 );
buf ( n19053 , n19052 );
nand ( n19054 , n19036 , n19053 );
buf ( n19055 , n19054 );
buf ( n19056 , n19055 );
and ( n19057 , n19015 , n19056 );
and ( n19058 , n18986 , n19014 );
or ( n19059 , n19057 , n19058 );
buf ( n19060 , n19059 );
buf ( n19061 , n19060 );
xor ( n19062 , n18978 , n19061 );
and ( n19063 , n18996 , n19004 );
buf ( n19064 , n19063 );
buf ( n19065 , n19064 );
buf ( n19066 , n18340 );
not ( n19067 , n19066 );
buf ( n19068 , n18579 );
not ( n19069 , n19068 );
or ( n19070 , n19067 , n19069 );
buf ( n19071 , n18992 );
buf ( n19072 , n18365 );
nand ( n19073 , n19071 , n19072 );
buf ( n19074 , n19073 );
buf ( n19075 , n19074 );
nand ( n19076 , n19070 , n19075 );
buf ( n19077 , n19076 );
buf ( n19078 , n19077 );
xor ( n19079 , n19065 , n19078 );
buf ( n19080 , n18219 );
not ( n19081 , n19080 );
buf ( n19082 , n18612 );
not ( n19083 , n19082 );
or ( n19084 , n19081 , n19083 );
buf ( n19085 , n19033 );
buf ( n19086 , n18264 );
nand ( n19087 , n19085 , n19086 );
buf ( n19088 , n19087 );
buf ( n19089 , n19088 );
nand ( n19090 , n19084 , n19089 );
buf ( n19091 , n19090 );
buf ( n19092 , n19091 );
xor ( n19093 , n19079 , n19092 );
buf ( n19094 , n19093 );
buf ( n19095 , n19094 );
and ( n19096 , n19062 , n19095 );
and ( n19097 , n18978 , n19061 );
or ( n19098 , n19096 , n19097 );
buf ( n19099 , n19098 );
buf ( n19100 , n19099 );
and ( n19101 , n18940 , n19100 );
and ( n19102 , n18906 , n18939 );
or ( n19103 , n19101 , n19102 );
buf ( n19104 , n19103 );
buf ( n19105 , n19104 );
xor ( n19106 , n18885 , n19105 );
xor ( n19107 , n18625 , n18653 );
xor ( n19108 , n19107 , n18697 );
buf ( n19109 , n19108 );
buf ( n19110 , n19109 );
and ( n19111 , n19106 , n19110 );
and ( n19112 , n18885 , n19105 );
or ( n19113 , n19111 , n19112 );
buf ( n19114 , n19113 );
buf ( n19115 , n19114 );
not ( n19116 , n18843 );
not ( n19117 , n18846 );
or ( n19118 , n19116 , n19117 );
nand ( n19119 , n19118 , n18881 );
buf ( n19120 , n18082 );
not ( n19121 , n19120 );
buf ( n19122 , n18856 );
buf ( n19123 , n18840 );
nor ( n19124 , n19122 , n19123 );
buf ( n19125 , n19124 );
buf ( n19126 , n19125 );
nand ( n19127 , n19121 , n19126 );
buf ( n19128 , n19127 );
buf ( n19129 , n18082 );
buf ( n19130 , n18856 );
buf ( n19131 , n586 );
nor ( n19132 , n19130 , n19131 );
buf ( n19133 , n19132 );
buf ( n19134 , n19133 );
nand ( n19135 , n19129 , n19134 );
buf ( n19136 , n19135 );
nand ( n19137 , n19119 , n19128 , n19136 );
buf ( n19138 , n19137 );
and ( n19139 , n589 , n1203 );
not ( n19140 , n589 );
and ( n19141 , n19140 , n590 );
or ( n19142 , n19139 , n19141 );
buf ( n19143 , n19142 );
not ( n19144 , n19143 );
and ( n19145 , n588 , n589 );
buf ( n19146 , n588 );
buf ( n19147 , n589 );
nor ( n19148 , n19146 , n19147 );
buf ( n19149 , n19148 );
nor ( n19150 , n19145 , n19149 );
nand ( n19151 , n19144 , n19150 );
not ( n19152 , n19151 );
buf ( n19153 , n19152 );
not ( n19154 , n19153 );
buf ( n19155 , n588 );
not ( n19156 , n19155 );
buf ( n19157 , n18137 );
not ( n19158 , n19157 );
buf ( n19159 , n19158 );
buf ( n19160 , n19159 );
not ( n19161 , n19160 );
or ( n19162 , n19156 , n19161 );
buf ( n19163 , n588 );
not ( n19164 , n19163 );
buf ( n19165 , n19159 );
not ( n19166 , n19165 );
buf ( n19167 , n19166 );
buf ( n19168 , n19167 );
nand ( n19169 , n19164 , n19168 );
buf ( n19170 , n19169 );
buf ( n19171 , n19170 );
nand ( n19172 , n19162 , n19171 );
buf ( n19173 , n19172 );
buf ( n19174 , n19173 );
not ( n19175 , n19174 );
or ( n19176 , n19154 , n19175 );
not ( n19177 , n18849 );
not ( n19178 , n18109 );
not ( n19179 , n18180 );
or ( n19180 , n19178 , n19179 );
nand ( n19181 , n19180 , n18183 );
not ( n19182 , n19181 );
or ( n19183 , n19177 , n19182 );
or ( n19184 , n18184 , n18849 );
nand ( n19185 , n19183 , n19184 );
buf ( n19186 , n19185 );
buf ( n19187 , n19143 );
nand ( n19188 , n19186 , n19187 );
buf ( n19189 , n19188 );
buf ( n19190 , n19189 );
nand ( n19191 , n19176 , n19190 );
buf ( n19192 , n19191 );
buf ( n19193 , n19192 );
xor ( n19194 , n19138 , n19193 );
xor ( n19195 , n18774 , n18787 );
xor ( n19196 , n19195 , n18825 );
buf ( n19197 , n19196 );
buf ( n19198 , n19197 );
xor ( n19199 , n19194 , n19198 );
buf ( n19200 , n19199 );
buf ( n19201 , n19200 );
xor ( n19202 , n19115 , n19201 );
buf ( n19203 , n591 );
not ( n19204 , n19203 );
not ( n19205 , n18062 );
not ( n19206 , n18056 );
or ( n19207 , n19205 , n19206 );
nand ( n19208 , n19207 , n18065 );
not ( n19209 , n19208 );
xor ( n19210 , n590 , n19209 );
buf ( n19211 , n19210 );
not ( n19212 , n19211 );
or ( n19213 , n19204 , n19212 );
buf ( n19214 , n590 );
not ( n19215 , n19214 );
buf ( n19216 , n18184 );
not ( n19217 , n19216 );
buf ( n19218 , n19217 );
buf ( n19219 , n19218 );
not ( n19220 , n19219 );
or ( n19221 , n19215 , n19220 );
buf ( n19222 , n590 );
not ( n19223 , n19222 );
buf ( n19224 , n19181 );
nand ( n19225 , n19223 , n19224 );
buf ( n19226 , n19225 );
buf ( n19227 , n19226 );
nand ( n19228 , n19221 , n19227 );
buf ( n19229 , n19228 );
buf ( n19230 , n19229 );
buf ( n19231 , n590 );
not ( n19232 , n19231 );
buf ( n19233 , n591 );
nor ( n19234 , n19232 , n19233 );
buf ( n19235 , n19234 );
buf ( n19236 , n19235 );
buf ( n19237 , n19236 );
buf ( n19238 , n19237 );
buf ( n19239 , n19238 );
buf ( n19240 , n19239 );
buf ( n19241 , n19240 );
buf ( n19242 , n19241 );
buf ( n19243 , n19242 );
buf ( n19244 , n19243 );
buf ( n19245 , n19244 );
nand ( n19246 , n19230 , n19245 );
buf ( n19247 , n19246 );
buf ( n19248 , n19247 );
nand ( n19249 , n19213 , n19248 );
buf ( n19250 , n19249 );
buf ( n19251 , n19250 );
buf ( n19252 , n19152 );
not ( n19253 , n19252 );
not ( n19254 , n18082 );
and ( n19255 , n588 , n19254 );
not ( n19256 , n588 );
and ( n19257 , n19256 , n18082 );
or ( n19258 , n19255 , n19257 );
buf ( n19259 , n19258 );
not ( n19260 , n19259 );
or ( n19261 , n19253 , n19260 );
buf ( n19262 , n19173 );
buf ( n19263 , n19143 );
nand ( n19264 , n19262 , n19263 );
buf ( n19265 , n19264 );
buf ( n19266 , n19265 );
nand ( n19267 , n19261 , n19266 );
buf ( n19268 , n19267 );
buf ( n19269 , n19268 );
xor ( n19270 , n19251 , n19269 );
xor ( n19271 , n18793 , n18806 );
xor ( n19272 , n19271 , n18820 );
buf ( n19273 , n19272 );
buf ( n19274 , n19273 );
buf ( n19275 , n18431 );
not ( n19276 , n19275 );
buf ( n19277 , n18467 );
not ( n19278 , n19277 );
or ( n19279 , n19276 , n19278 );
buf ( n19280 , n18909 );
not ( n19281 , n19280 );
buf ( n19282 , n19281 );
buf ( n19283 , n19282 );
buf ( n19284 , n584 );
nand ( n19285 , n19283 , n19284 );
buf ( n19286 , n19285 );
buf ( n19287 , n19286 );
not ( n19288 , n19287 );
buf ( n19289 , n18909 );
buf ( n19290 , n18277 );
nand ( n19291 , n19289 , n19290 );
buf ( n19292 , n19291 );
buf ( n19293 , n19292 );
not ( n19294 , n19293 );
or ( n19295 , n19288 , n19294 );
buf ( n19296 , n18479 );
nand ( n19297 , n19295 , n19296 );
buf ( n19298 , n19297 );
buf ( n19299 , n19298 );
nand ( n19300 , n19279 , n19299 );
buf ( n19301 , n19300 );
buf ( n19302 , n19301 );
xor ( n19303 , n19274 , n19302 );
xor ( n19304 , n19065 , n19078 );
and ( n19305 , n19304 , n19092 );
and ( n19306 , n19065 , n19078 );
or ( n19307 , n19305 , n19306 );
buf ( n19308 , n19307 );
buf ( n19309 , n19308 );
xor ( n19310 , n18546 , n18587 );
xor ( n19311 , n19310 , n18620 );
buf ( n19312 , n19311 );
buf ( n19313 , n19312 );
xor ( n19314 , n19309 , n19313 );
buf ( n19315 , n18418 );
not ( n19316 , n19315 );
buf ( n19317 , n18645 );
not ( n19318 , n19317 );
or ( n19319 , n19316 , n19318 );
buf ( n19320 , n18954 );
buf ( n19321 , n18392 );
nand ( n19322 , n19320 , n19321 );
buf ( n19323 , n19322 );
buf ( n19324 , n19323 );
nand ( n19325 , n19319 , n19324 );
buf ( n19326 , n19325 );
buf ( n19327 , n19326 );
and ( n19328 , n19314 , n19327 );
and ( n19329 , n19309 , n19313 );
or ( n19330 , n19328 , n19329 );
buf ( n19331 , n19330 );
buf ( n19332 , n19331 );
xor ( n19333 , n19303 , n19332 );
buf ( n19334 , n19333 );
buf ( n19335 , n19334 );
and ( n19336 , n19270 , n19335 );
and ( n19337 , n19251 , n19269 );
or ( n19338 , n19336 , n19337 );
buf ( n19339 , n19338 );
buf ( n19340 , n19339 );
and ( n19341 , n19202 , n19340 );
and ( n19342 , n19115 , n19201 );
or ( n19343 , n19341 , n19342 );
buf ( n19344 , n19343 );
buf ( n19345 , n19344 );
xor ( n19346 , n18836 , n19345 );
xor ( n19347 , n19138 , n19193 );
and ( n19348 , n19347 , n19198 );
and ( n19349 , n19138 , n19193 );
or ( n19350 , n19348 , n19349 );
buf ( n19351 , n19350 );
buf ( n19352 , n19351 );
buf ( n19353 , n18881 );
not ( n19354 , n19353 );
and ( n19355 , n18082 , n18840 );
not ( n19356 , n18082 );
and ( n19357 , n19356 , n586 );
or ( n19358 , n19355 , n19357 );
buf ( n19359 , n19358 );
not ( n19360 , n19359 );
or ( n19361 , n19354 , n19360 );
buf ( n19362 , n18840 );
not ( n19363 , n19362 );
buf ( n19364 , n18137 );
not ( n19365 , n19364 );
or ( n19366 , n19363 , n19365 );
buf ( n19367 , n19159 );
buf ( n19368 , n586 );
nand ( n19369 , n19367 , n19368 );
buf ( n19370 , n19369 );
buf ( n19371 , n19370 );
nand ( n19372 , n19366 , n19371 );
buf ( n19373 , n19372 );
buf ( n19374 , n19373 );
buf ( n19375 , n18857 );
nand ( n19376 , n19374 , n19375 );
buf ( n19377 , n19376 );
buf ( n19378 , n19377 );
nand ( n19379 , n19361 , n19378 );
buf ( n19380 , n19379 );
buf ( n19381 , n19380 );
not ( n19382 , n19143 );
not ( n19383 , n18066 );
not ( n19384 , n19383 );
and ( n19385 , n588 , n19384 );
not ( n19386 , n588 );
not ( n19387 , n19208 );
and ( n19388 , n19386 , n19387 );
or ( n19389 , n19385 , n19388 );
not ( n19390 , n19389 );
or ( n19391 , n19382 , n19390 );
nand ( n19392 , n19185 , n19152 );
nand ( n19393 , n19391 , n19392 );
buf ( n19394 , n19393 );
xor ( n19395 , n19381 , n19394 );
buf ( n19396 , n591 );
not ( n19397 , n19396 );
buf ( n19398 , n18023 );
xor ( n19399 , n590 , n19398 );
buf ( n19400 , n19399 );
not ( n19401 , n19400 );
or ( n19402 , n19397 , n19401 );
buf ( n19403 , n18036 );
and ( n19404 , n19403 , n590 );
not ( n19405 , n19403 );
and ( n19406 , n19405 , n2103 );
nor ( n19407 , n19404 , n19406 );
buf ( n19408 , n19407 );
buf ( n19409 , n19244 );
nand ( n19410 , n19408 , n19409 );
buf ( n19411 , n19410 );
buf ( n19412 , n19411 );
nand ( n19413 , n19402 , n19412 );
buf ( n19414 , n19413 );
buf ( n19415 , n19414 );
xor ( n19416 , n19395 , n19415 );
buf ( n19417 , n19416 );
buf ( n19418 , n19417 );
xor ( n19419 , n19352 , n19418 );
not ( n19420 , n591 );
not ( n19421 , n19407 );
or ( n19422 , n19420 , n19421 );
buf ( n19423 , n19210 );
buf ( n19424 , n19244 );
nand ( n19425 , n19423 , n19424 );
buf ( n19426 , n19425 );
nand ( n19427 , n19422 , n19426 );
buf ( n19428 , n19427 );
xor ( n19429 , n19274 , n19302 );
and ( n19430 , n19429 , n19332 );
and ( n19431 , n19274 , n19302 );
or ( n19432 , n19430 , n19431 );
buf ( n19433 , n19432 );
buf ( n19434 , n19433 );
xor ( n19435 , n19428 , n19434 );
xor ( n19436 , n18486 , n18534 );
xor ( n19437 , n19436 , n18702 );
buf ( n19438 , n19437 );
buf ( n19439 , n19438 );
and ( n19440 , n19435 , n19439 );
and ( n19441 , n19428 , n19434 );
or ( n19442 , n19440 , n19441 );
buf ( n19443 , n19442 );
buf ( n19444 , n19443 );
xor ( n19445 , n19419 , n19444 );
buf ( n19446 , n19445 );
buf ( n19447 , n19446 );
xor ( n19448 , n19346 , n19447 );
buf ( n19449 , n19448 );
buf ( n19450 , n19449 );
buf ( n19451 , n19450 );
buf ( n19452 , n19451 );
not ( n19453 , n19452 );
xor ( n19454 , n19428 , n19434 );
xor ( n19455 , n19454 , n19439 );
buf ( n19456 , n19455 );
buf ( n19457 , n19456 );
not ( n19458 , n18882 );
buf ( n19459 , n586 );
not ( n19460 , n19459 );
buf ( n19461 , n18457 );
not ( n19462 , n19461 );
or ( n19463 , n19460 , n19462 );
buf ( n19464 , n15680 );
buf ( n19465 , n18840 );
nand ( n19466 , n19464 , n19465 );
buf ( n19467 , n19466 );
buf ( n19468 , n19467 );
nand ( n19469 , n19463 , n19468 );
buf ( n19470 , n19469 );
not ( n19471 , n19470 );
or ( n19472 , n19458 , n19471 );
not ( n19473 , n18869 );
not ( n19474 , n18865 );
or ( n19475 , n19473 , n19474 );
nand ( n19476 , n19475 , n18857 );
nand ( n19477 , n19472 , n19476 );
buf ( n19478 , n19477 );
xor ( n19479 , n19309 , n19313 );
xor ( n19480 , n19479 , n19327 );
buf ( n19481 , n19480 );
buf ( n19482 , n19481 );
xor ( n19483 , n19478 , n19482 );
buf ( n19484 , n18479 );
not ( n19485 , n19484 );
buf ( n19486 , n584 );
not ( n19487 , n19486 );
buf ( n19488 , n18397 );
not ( n19489 , n19488 );
or ( n19490 , n19487 , n19489 );
buf ( n19491 , n10819 );
buf ( n19492 , n18277 );
nand ( n19493 , n19491 , n19492 );
buf ( n19494 , n19493 );
buf ( n19495 , n19494 );
nand ( n19496 , n19490 , n19495 );
buf ( n19497 , n19496 );
buf ( n19498 , n19497 );
not ( n19499 , n19498 );
or ( n19500 , n19485 , n19499 );
buf ( n19501 , n18931 );
buf ( n19502 , n18431 );
nand ( n19503 , n19501 , n19502 );
buf ( n19504 , n19503 );
buf ( n19505 , n19504 );
nand ( n19506 , n19500 , n19505 );
buf ( n19507 , n19506 );
buf ( n19508 , n19507 );
not ( n19509 , n18285 );
not ( n19510 , n18901 );
or ( n19511 , n19509 , n19510 );
buf ( n19512 , n582 );
not ( n19513 , n19512 );
buf ( n19514 , n18635 );
not ( n19515 , n19514 );
or ( n19516 , n19513 , n19515 );
buf ( n19517 , n9497 );
buf ( n19518 , n18303 );
nand ( n19519 , n19517 , n19518 );
buf ( n19520 , n19519 );
buf ( n19521 , n19520 );
nand ( n19522 , n19516 , n19521 );
buf ( n19523 , n19522 );
buf ( n19524 , n19523 );
buf ( n19525 , n18316 );
nand ( n19526 , n19524 , n19525 );
buf ( n19527 , n19526 );
nand ( n19528 , n19511 , n19527 );
buf ( n19529 , n19528 );
xor ( n19530 , n19508 , n19529 );
buf ( n19531 , n4750 );
buf ( n19532 , n19531 );
buf ( n19533 , n19532 );
buf ( n19534 , n19533 );
buf ( n19535 , n19534 );
buf ( n19536 , n576 );
and ( n19537 , n19535 , n19536 );
buf ( n19538 , n19537 );
buf ( n19539 , n19538 );
buf ( n19540 , n18340 );
not ( n19541 , n19540 );
buf ( n19542 , n19006 );
not ( n19543 , n19542 );
or ( n19544 , n19541 , n19543 );
buf ( n19545 , n576 );
not ( n19546 , n19545 );
buf ( n19547 , n13663 );
not ( n19548 , n19547 );
buf ( n19549 , n19548 );
buf ( n19550 , n19549 );
not ( n19551 , n19550 );
or ( n19552 , n19546 , n19551 );
buf ( n19553 , n19549 );
not ( n19554 , n19553 );
buf ( n19555 , n19554 );
buf ( n19556 , n19555 );
buf ( n19557 , n7809 );
nand ( n19558 , n19556 , n19557 );
buf ( n19559 , n19558 );
buf ( n19560 , n19559 );
nand ( n19561 , n19552 , n19560 );
buf ( n19562 , n19561 );
buf ( n19563 , n19562 );
buf ( n19564 , n18365 );
nand ( n19565 , n19563 , n19564 );
buf ( n19566 , n19565 );
buf ( n19567 , n19566 );
nand ( n19568 , n19544 , n19567 );
buf ( n19569 , n19568 );
buf ( n19570 , n19569 );
xor ( n19571 , n19539 , n19570 );
buf ( n19572 , n18219 );
not ( n19573 , n19572 );
buf ( n19574 , n19048 );
not ( n19575 , n19574 );
or ( n19576 , n19573 , n19575 );
buf ( n19577 , n578 );
not ( n19578 , n19577 );
buf ( n19579 , n18538 );
not ( n19580 , n19579 );
or ( n19581 , n19578 , n19580 );
buf ( n19582 , n13665 );
buf ( n19583 , n18233 );
nand ( n19584 , n19582 , n19583 );
buf ( n19585 , n19584 );
buf ( n19586 , n19585 );
nand ( n19587 , n19581 , n19586 );
buf ( n19588 , n19587 );
buf ( n19589 , n19588 );
buf ( n19590 , n18264 );
nand ( n19591 , n19589 , n19590 );
buf ( n19592 , n19591 );
buf ( n19593 , n19592 );
nand ( n19594 , n19576 , n19593 );
buf ( n19595 , n19594 );
buf ( n19596 , n19595 );
and ( n19597 , n19571 , n19596 );
and ( n19598 , n19539 , n19570 );
or ( n19599 , n19597 , n19598 );
buf ( n19600 , n19599 );
buf ( n19601 , n19600 );
buf ( n19602 , n18418 );
not ( n19603 , n19602 );
buf ( n19604 , n18970 );
not ( n19605 , n19604 );
or ( n19606 , n19603 , n19605 );
buf ( n19607 , n580 );
not ( n19608 , n19607 );
buf ( n19609 , n18599 );
not ( n19610 , n19609 );
or ( n19611 , n19608 , n19610 );
buf ( n19612 , n18326 );
buf ( n19613 , n18402 );
nand ( n19614 , n19612 , n19613 );
buf ( n19615 , n19614 );
buf ( n19616 , n19615 );
nand ( n19617 , n19611 , n19616 );
buf ( n19618 , n19617 );
buf ( n19619 , n19618 );
buf ( n19620 , n18391 );
nand ( n19621 , n19619 , n19620 );
buf ( n19622 , n19621 );
buf ( n19623 , n19622 );
nand ( n19624 , n19606 , n19623 );
buf ( n19625 , n19624 );
buf ( n19626 , n19625 );
xor ( n19627 , n19601 , n19626 );
buf ( n19628 , n13664 );
not ( n19629 , n19628 );
buf ( n19630 , n19629 );
buf ( n19631 , n19630 );
buf ( n19632 , n19631 );
buf ( n19633 , n19632 );
buf ( n19634 , n19633 );
not ( n19635 , n19634 );
buf ( n19636 , n19635 );
buf ( n19637 , n19636 );
buf ( n19638 , n576 );
and ( n19639 , n19637 , n19638 );
buf ( n19640 , n19639 );
buf ( n19641 , n19640 );
buf ( n19642 , n18340 );
not ( n19643 , n19642 );
buf ( n19644 , n19562 );
not ( n19645 , n19644 );
or ( n19646 , n19643 , n19645 );
buf ( n19647 , n576 );
not ( n19648 , n19647 );
buf ( n19649 , n19534 );
not ( n19650 , n19649 );
buf ( n19651 , n19650 );
buf ( n19652 , n19651 );
not ( n19653 , n19652 );
or ( n19654 , n19648 , n19653 );
buf ( n19655 , n19534 );
buf ( n19656 , n7809 );
nand ( n19657 , n19655 , n19656 );
buf ( n19658 , n19657 );
buf ( n19659 , n19658 );
nand ( n19660 , n19654 , n19659 );
buf ( n19661 , n19660 );
buf ( n19662 , n19661 );
buf ( n19663 , n18365 );
nand ( n19664 , n19662 , n19663 );
buf ( n19665 , n19664 );
buf ( n19666 , n19665 );
nand ( n19667 , n19646 , n19666 );
buf ( n19668 , n19667 );
buf ( n19669 , n19668 );
xor ( n19670 , n19641 , n19669 );
buf ( n19671 , n18219 );
not ( n19672 , n19671 );
buf ( n19673 , n19588 );
not ( n19674 , n19673 );
or ( n19675 , n19672 , n19674 );
buf ( n19676 , n578 );
not ( n19677 , n19676 );
buf ( n19678 , n19000 );
not ( n19679 , n19678 );
or ( n19680 , n19677 , n19679 );
buf ( n19681 , n18997 );
buf ( n19682 , n18233 );
nand ( n19683 , n19681 , n19682 );
buf ( n19684 , n19683 );
buf ( n19685 , n19684 );
nand ( n19686 , n19680 , n19685 );
buf ( n19687 , n19686 );
buf ( n19688 , n19687 );
buf ( n19689 , n18264 );
nand ( n19690 , n19688 , n19689 );
buf ( n19691 , n19690 );
buf ( n19692 , n19691 );
nand ( n19693 , n19675 , n19692 );
buf ( n19694 , n19693 );
buf ( n19695 , n19694 );
and ( n19696 , n19670 , n19695 );
and ( n19697 , n19641 , n19669 );
or ( n19698 , n19696 , n19697 );
buf ( n19699 , n19698 );
buf ( n19700 , n19699 );
buf ( n19701 , n18418 );
not ( n19702 , n19701 );
buf ( n19703 , n19618 );
not ( n19704 , n19703 );
or ( n19705 , n19702 , n19704 );
buf ( n19706 , n580 );
not ( n19707 , n19706 );
buf ( n19708 , n19022 );
not ( n19709 , n19708 );
or ( n19710 , n19707 , n19709 );
buf ( n19711 , n18489 );
buf ( n19712 , n18402 );
nand ( n19713 , n19711 , n19712 );
buf ( n19714 , n19713 );
buf ( n19715 , n19714 );
nand ( n19716 , n19710 , n19715 );
buf ( n19717 , n19716 );
buf ( n19718 , n19717 );
buf ( n19719 , n18391 );
nand ( n19720 , n19718 , n19719 );
buf ( n19721 , n19720 );
buf ( n19722 , n19721 );
nand ( n19723 , n19705 , n19722 );
buf ( n19724 , n19723 );
buf ( n19725 , n19724 );
xor ( n19726 , n19700 , n19725 );
xor ( n19727 , n19539 , n19570 );
xor ( n19728 , n19727 , n19596 );
buf ( n19729 , n19728 );
buf ( n19730 , n19729 );
and ( n19731 , n19726 , n19730 );
and ( n19732 , n19700 , n19725 );
or ( n19733 , n19731 , n19732 );
buf ( n19734 , n19733 );
buf ( n19735 , n19734 );
and ( n19736 , n19627 , n19735 );
and ( n19737 , n19601 , n19626 );
or ( n19738 , n19736 , n19737 );
buf ( n19739 , n19738 );
buf ( n19740 , n19739 );
and ( n19741 , n19530 , n19740 );
and ( n19742 , n19508 , n19529 );
or ( n19743 , n19741 , n19742 );
buf ( n19744 , n19743 );
buf ( n19745 , n19744 );
and ( n19746 , n19483 , n19745 );
and ( n19747 , n19478 , n19482 );
or ( n19748 , n19746 , n19747 );
buf ( n19749 , n19748 );
buf ( n19750 , n19749 );
xor ( n19751 , n18885 , n19105 );
xor ( n19752 , n19751 , n19110 );
buf ( n19753 , n19752 );
buf ( n19754 , n19753 );
xor ( n19755 , n19750 , n19754 );
buf ( n19756 , n19143 );
not ( n19757 , n19756 );
buf ( n19758 , n19258 );
not ( n19759 , n19758 );
or ( n19760 , n19757 , n19759 );
not ( n19761 , n18725 );
and ( n19762 , n588 , n19761 );
not ( n19763 , n588 );
and ( n19764 , n19763 , n18725 );
or ( n19765 , n19762 , n19764 );
buf ( n19766 , n19765 );
buf ( n19767 , n19152 );
nand ( n19768 , n19766 , n19767 );
buf ( n19769 , n19768 );
buf ( n19770 , n19769 );
nand ( n19771 , n19760 , n19770 );
buf ( n19772 , n19771 );
buf ( n19773 , n19772 );
xor ( n19774 , n18906 , n18939 );
xor ( n19775 , n19774 , n19100 );
buf ( n19776 , n19775 );
buf ( n19777 , n19776 );
xor ( n19778 , n19773 , n19777 );
buf ( n19779 , n19244 );
not ( n19780 , n19779 );
buf ( n19781 , n19159 );
not ( n19782 , n19781 );
buf ( n19783 , n19782 );
xor ( n19784 , n590 , n19783 );
buf ( n19785 , n19784 );
not ( n19786 , n19785 );
or ( n19787 , n19780 , n19786 );
buf ( n19788 , n19229 );
buf ( n19789 , n591 );
nand ( n19790 , n19788 , n19789 );
buf ( n19791 , n19790 );
buf ( n19792 , n19791 );
nand ( n19793 , n19787 , n19792 );
buf ( n19794 , n19793 );
buf ( n19795 , n19794 );
and ( n19796 , n19778 , n19795 );
and ( n19797 , n19773 , n19777 );
or ( n19798 , n19796 , n19797 );
buf ( n19799 , n19798 );
buf ( n19800 , n19799 );
and ( n19801 , n19755 , n19800 );
and ( n19802 , n19750 , n19754 );
or ( n19803 , n19801 , n19802 );
buf ( n19804 , n19803 );
buf ( n19805 , n19804 );
xor ( n19806 , n19457 , n19805 );
xor ( n19807 , n19115 , n19201 );
xor ( n19808 , n19807 , n19340 );
buf ( n19809 , n19808 );
buf ( n19810 , n19809 );
and ( n19811 , n19806 , n19810 );
and ( n19812 , n19457 , n19805 );
or ( n19813 , n19811 , n19812 );
buf ( n19814 , n19813 );
not ( n19815 , n19814 );
nand ( n19816 , n19453 , n19815 );
buf ( n19817 , n19452 );
buf ( n19818 , n19814 );
nand ( n19819 , n19817 , n19818 );
buf ( n19820 , n19819 );
nand ( n19821 , n19816 , n19820 );
not ( n19822 , n19821 );
not ( n19823 , n19822 );
xor ( n19824 , n19457 , n19805 );
xor ( n19825 , n19824 , n19810 );
buf ( n19826 , n19825 );
xor ( n19827 , n19251 , n19269 );
xor ( n19828 , n19827 , n19335 );
buf ( n19829 , n19828 );
buf ( n19830 , n19829 );
buf ( n19831 , n18857 );
not ( n19832 , n19831 );
buf ( n19833 , n19470 );
not ( n19834 , n19833 );
or ( n19835 , n19832 , n19834 );
and ( n19836 , n18203 , n18840 );
not ( n19837 , n18203 );
and ( n19838 , n19837 , n586 );
or ( n19839 , n19836 , n19838 );
buf ( n19840 , n19839 );
buf ( n19841 , n18881 );
nand ( n19842 , n19840 , n19841 );
buf ( n19843 , n19842 );
buf ( n19844 , n19843 );
nand ( n19845 , n19835 , n19844 );
buf ( n19846 , n19845 );
buf ( n19847 , n19846 );
xor ( n19848 , n18978 , n19061 );
xor ( n19849 , n19848 , n19095 );
buf ( n19850 , n19849 );
buf ( n19851 , n19850 );
xor ( n19852 , n19847 , n19851 );
xor ( n19853 , n18986 , n19014 );
xor ( n19854 , n19853 , n19056 );
buf ( n19855 , n19854 );
buf ( n19856 , n19855 );
buf ( n19857 , n18657 );
not ( n19858 , n19857 );
buf ( n19859 , n19523 );
not ( n19860 , n19859 );
or ( n19861 , n19858 , n19860 );
buf ( n19862 , n582 );
not ( n19863 , n19862 );
buf ( n19864 , n8543 );
not ( n19865 , n19864 );
or ( n19866 , n19863 , n19865 );
buf ( n19867 , n18759 );
buf ( n19868 , n18303 );
nand ( n19869 , n19867 , n19868 );
buf ( n19870 , n19869 );
buf ( n19871 , n19870 );
nand ( n19872 , n19866 , n19871 );
buf ( n19873 , n19872 );
buf ( n19874 , n19873 );
buf ( n19875 , n18316 );
nand ( n19876 , n19874 , n19875 );
buf ( n19877 , n19876 );
buf ( n19878 , n19877 );
nand ( n19879 , n19861 , n19878 );
buf ( n19880 , n19879 );
buf ( n19881 , n19880 );
xor ( n19882 , n19856 , n19881 );
buf ( n19883 , n18479 );
not ( n19884 , n19883 );
and ( n19885 , n10854 , n18277 );
not ( n19886 , n10854 );
and ( n19887 , n19886 , n584 );
or ( n19888 , n19885 , n19887 );
buf ( n19889 , n19888 );
not ( n19890 , n19889 );
or ( n19891 , n19884 , n19890 );
buf ( n19892 , n19497 );
buf ( n19893 , n18431 );
nand ( n19894 , n19892 , n19893 );
buf ( n19895 , n19894 );
buf ( n19896 , n19895 );
nand ( n19897 , n19891 , n19896 );
buf ( n19898 , n19897 );
buf ( n19899 , n19898 );
and ( n19900 , n19882 , n19899 );
and ( n19901 , n19856 , n19881 );
or ( n19902 , n19900 , n19901 );
buf ( n19903 , n19902 );
buf ( n19904 , n19903 );
and ( n19905 , n19852 , n19904 );
and ( n19906 , n19847 , n19851 );
or ( n19907 , n19905 , n19906 );
buf ( n19908 , n19907 );
buf ( n19909 , n19908 );
xor ( n19910 , n19478 , n19482 );
xor ( n19911 , n19910 , n19745 );
buf ( n19912 , n19911 );
buf ( n19913 , n19912 );
xor ( n19914 , n19909 , n19913 );
buf ( n19915 , n19143 );
not ( n19916 , n19915 );
buf ( n19917 , n19765 );
not ( n19918 , n19917 );
or ( n19919 , n19916 , n19918 );
and ( n19920 , n588 , n18868 );
not ( n19921 , n588 );
and ( n19922 , n19921 , n18861 );
or ( n19923 , n19920 , n19922 );
buf ( n19924 , n19923 );
buf ( n19925 , n19152 );
nand ( n19926 , n19924 , n19925 );
buf ( n19927 , n19926 );
buf ( n19928 , n19927 );
nand ( n19929 , n19919 , n19928 );
buf ( n19930 , n19929 );
buf ( n19931 , n19930 );
xor ( n19932 , n19508 , n19529 );
xor ( n19933 , n19932 , n19740 );
buf ( n19934 , n19933 );
buf ( n19935 , n19934 );
xor ( n19936 , n19931 , n19935 );
buf ( n19937 , n18857 );
not ( n19938 , n19937 );
buf ( n19939 , n19839 );
not ( n19940 , n19939 );
or ( n19941 , n19938 , n19940 );
buf ( n19942 , n586 );
not ( n19943 , n19942 );
buf ( n19944 , n18667 );
not ( n19945 , n19944 );
buf ( n19946 , n19945 );
buf ( n19947 , n19946 );
not ( n19948 , n19947 );
or ( n19949 , n19943 , n19948 );
buf ( n19950 , n13592 );
buf ( n19951 , n18840 );
nand ( n19952 , n19950 , n19951 );
buf ( n19953 , n19952 );
buf ( n19954 , n19953 );
nand ( n19955 , n19949 , n19954 );
buf ( n19956 , n19955 );
buf ( n19957 , n19956 );
buf ( n19958 , n18881 );
nand ( n19959 , n19957 , n19958 );
buf ( n19960 , n19959 );
buf ( n19961 , n19960 );
nand ( n19962 , n19941 , n19961 );
buf ( n19963 , n19962 );
buf ( n19964 , n19963 );
xor ( n19965 , n19601 , n19626 );
xor ( n19966 , n19965 , n19735 );
buf ( n19967 , n19966 );
buf ( n19968 , n19967 );
xor ( n19969 , n19964 , n19968 );
buf ( n19970 , n2337 );
not ( n19971 , n19970 );
buf ( n19972 , n19971 );
buf ( n19973 , n19972 );
not ( n19974 , n19973 );
buf ( n19975 , n19974 );
buf ( n19976 , n19975 );
buf ( n19977 , n576 );
and ( n19978 , n19976 , n19977 );
buf ( n19979 , n19978 );
buf ( n19980 , n19979 );
buf ( n19981 , n18340 );
not ( n19982 , n19981 );
buf ( n19983 , n19661 );
not ( n19984 , n19983 );
or ( n19985 , n19982 , n19984 );
buf ( n19986 , n576 );
not ( n19987 , n19986 );
buf ( n19988 , n19633 );
not ( n19989 , n19988 );
or ( n19990 , n19987 , n19989 );
buf ( n19991 , n19636 );
buf ( n19992 , n7809 );
nand ( n19993 , n19991 , n19992 );
buf ( n19994 , n19993 );
buf ( n19995 , n19994 );
nand ( n19996 , n19990 , n19995 );
buf ( n19997 , n19996 );
buf ( n19998 , n19997 );
buf ( n19999 , n18365 );
nand ( n20000 , n19998 , n19999 );
buf ( n20001 , n20000 );
buf ( n20002 , n20001 );
nand ( n20003 , n19985 , n20002 );
buf ( n20004 , n20003 );
buf ( n20005 , n20004 );
xor ( n20006 , n19980 , n20005 );
buf ( n20007 , n18219 );
not ( n20008 , n20007 );
buf ( n20009 , n19687 );
not ( n20010 , n20009 );
or ( n20011 , n20008 , n20010 );
buf ( n20012 , n578 );
not ( n20013 , n20012 );
buf ( n20014 , n19549 );
not ( n20015 , n20014 );
or ( n20016 , n20013 , n20015 );
buf ( n20017 , n18233 );
buf ( n20018 , n13663 );
nand ( n20019 , n20017 , n20018 );
buf ( n20020 , n20019 );
buf ( n20021 , n20020 );
nand ( n20022 , n20016 , n20021 );
buf ( n20023 , n20022 );
buf ( n20024 , n20023 );
buf ( n20025 , n18264 );
nand ( n20026 , n20024 , n20025 );
buf ( n20027 , n20026 );
buf ( n20028 , n20027 );
nand ( n20029 , n20011 , n20028 );
buf ( n20030 , n20029 );
buf ( n20031 , n20030 );
and ( n20032 , n20006 , n20031 );
and ( n20033 , n19980 , n20005 );
or ( n20034 , n20032 , n20033 );
buf ( n20035 , n20034 );
buf ( n20036 , n20035 );
xor ( n20037 , n19641 , n19669 );
xor ( n20038 , n20037 , n19695 );
buf ( n20039 , n20038 );
buf ( n20040 , n20039 );
xor ( n20041 , n20036 , n20040 );
buf ( n20042 , n18418 );
not ( n20043 , n20042 );
buf ( n20044 , n19717 );
not ( n20045 , n20044 );
or ( n20046 , n20043 , n20045 );
not ( n20047 , n580 );
not ( n20048 , n18569 );
or ( n20049 , n20047 , n20048 );
buf ( n20050 , n18566 );
buf ( n20051 , n18402 );
nand ( n20052 , n20050 , n20051 );
buf ( n20053 , n20052 );
nand ( n20054 , n20049 , n20053 );
nand ( n20055 , n20054 , n18391 );
buf ( n20056 , n20055 );
nand ( n20057 , n20046 , n20056 );
buf ( n20058 , n20057 );
buf ( n20059 , n20058 );
and ( n20060 , n20041 , n20059 );
and ( n20061 , n20036 , n20040 );
or ( n20062 , n20060 , n20061 );
buf ( n20063 , n20062 );
buf ( n20064 , n20063 );
buf ( n20065 , n18285 );
not ( n20066 , n20065 );
buf ( n20067 , n19873 );
not ( n20068 , n20067 );
or ( n20069 , n20066 , n20068 );
buf ( n20070 , n582 );
not ( n20071 , n20070 );
buf ( n20072 , n18960 );
not ( n20073 , n20072 );
or ( n20074 , n20071 , n20073 );
buf ( n20075 , n18357 );
buf ( n20076 , n18303 );
nand ( n20077 , n20075 , n20076 );
buf ( n20078 , n20077 );
buf ( n20079 , n20078 );
nand ( n20080 , n20074 , n20079 );
buf ( n20081 , n20080 );
buf ( n20082 , n20081 );
buf ( n20083 , n18316 );
nand ( n20084 , n20082 , n20083 );
buf ( n20085 , n20084 );
buf ( n20086 , n20085 );
nand ( n20087 , n20069 , n20086 );
buf ( n20088 , n20087 );
buf ( n20089 , n20088 );
xor ( n20090 , n20064 , n20089 );
xor ( n20091 , n19700 , n19725 );
xor ( n20092 , n20091 , n19730 );
buf ( n20093 , n20092 );
buf ( n20094 , n20093 );
and ( n20095 , n20090 , n20094 );
and ( n20096 , n20064 , n20089 );
or ( n20097 , n20095 , n20096 );
buf ( n20098 , n20097 );
buf ( n20099 , n20098 );
and ( n20100 , n19969 , n20099 );
and ( n20101 , n19964 , n19968 );
or ( n20102 , n20100 , n20101 );
buf ( n20103 , n20102 );
buf ( n20104 , n20103 );
and ( n20105 , n19936 , n20104 );
and ( n20106 , n19931 , n19935 );
or ( n20107 , n20105 , n20106 );
buf ( n20108 , n20107 );
buf ( n20109 , n20108 );
and ( n20110 , n19914 , n20109 );
and ( n20111 , n19909 , n19913 );
or ( n20112 , n20110 , n20111 );
buf ( n20113 , n20112 );
buf ( n20114 , n20113 );
xor ( n20115 , n19830 , n20114 );
xor ( n20116 , n19750 , n19754 );
xor ( n20117 , n20116 , n19800 );
buf ( n20118 , n20117 );
buf ( n20119 , n20118 );
and ( n20120 , n20115 , n20119 );
and ( n20121 , n19830 , n20114 );
or ( n20122 , n20120 , n20121 );
buf ( n20123 , n20122 );
nor ( n20124 , n19826 , n20123 );
xor ( n20125 , n19830 , n20114 );
xor ( n20126 , n20125 , n20119 );
buf ( n20127 , n20126 );
buf ( n20128 , n20127 );
xor ( n20129 , n19773 , n19777 );
xor ( n20130 , n20129 , n19795 );
buf ( n20131 , n20130 );
buf ( n20132 , n20131 );
buf ( n20133 , n19244 );
not ( n20134 , n20133 );
and ( n20135 , n590 , n19254 );
not ( n20136 , n590 );
not ( n20137 , n19254 );
and ( n20138 , n20136 , n20137 );
or ( n20139 , n20135 , n20138 );
buf ( n20140 , n20139 );
not ( n20141 , n20140 );
or ( n20142 , n20134 , n20141 );
buf ( n20143 , n19784 );
buf ( n20144 , n591 );
nand ( n20145 , n20143 , n20144 );
buf ( n20146 , n20145 );
buf ( n20147 , n20146 );
nand ( n20148 , n20142 , n20147 );
buf ( n20149 , n20148 );
buf ( n20150 , n20149 );
xor ( n20151 , n19847 , n19851 );
xor ( n20152 , n20151 , n19904 );
buf ( n20153 , n20152 );
buf ( n20154 , n20153 );
xor ( n20155 , n20150 , n20154 );
buf ( n20156 , n19152 );
not ( n20157 , n20156 );
buf ( n20158 , n15680 );
buf ( n20159 , n20158 );
buf ( n20160 , n20159 );
buf ( n20161 , n20160 );
not ( n20162 , n20161 );
buf ( n20163 , n20162 );
and ( n20164 , n588 , n20163 );
not ( n20165 , n588 );
and ( n20166 , n20165 , n20160 );
or ( n20167 , n20164 , n20166 );
buf ( n20168 , n20167 );
not ( n20169 , n20168 );
or ( n20170 , n20157 , n20169 );
buf ( n20171 , n19923 );
buf ( n20172 , n19143 );
nand ( n20173 , n20171 , n20172 );
buf ( n20174 , n20173 );
buf ( n20175 , n20174 );
nand ( n20176 , n20170 , n20175 );
buf ( n20177 , n20176 );
buf ( n20178 , n20177 );
xor ( n20179 , n19856 , n19881 );
xor ( n20180 , n20179 , n19899 );
buf ( n20181 , n20180 );
buf ( n20182 , n20181 );
xor ( n20183 , n20178 , n20182 );
buf ( n20184 , n18431 );
not ( n20185 , n20184 );
buf ( n20186 , n19888 );
not ( n20187 , n20186 );
or ( n20188 , n20185 , n20187 );
and ( n20189 , n584 , n9498 );
not ( n20190 , n584 );
and ( n20191 , n20190 , n9497 );
or ( n20192 , n20189 , n20191 );
buf ( n20193 , n20192 );
buf ( n20194 , n18479 );
nand ( n20195 , n20193 , n20194 );
buf ( n20196 , n20195 );
buf ( n20197 , n20196 );
nand ( n20198 , n20188 , n20197 );
buf ( n20199 , n20198 );
buf ( n20200 , n20199 );
buf ( n20201 , n18857 );
not ( n20202 , n20201 );
buf ( n20203 , n19956 );
not ( n20204 , n20203 );
or ( n20205 , n20202 , n20204 );
buf ( n20206 , n586 );
not ( n20207 , n20206 );
buf ( n20208 , n18682 );
not ( n20209 , n20208 );
or ( n20210 , n20207 , n20209 );
buf ( n20211 , n10822 );
buf ( n20212 , n18840 );
nand ( n20213 , n20211 , n20212 );
buf ( n20214 , n20213 );
buf ( n20215 , n20214 );
nand ( n20216 , n20210 , n20215 );
buf ( n20217 , n20216 );
buf ( n20218 , n20217 );
buf ( n20219 , n18881 );
nand ( n20220 , n20218 , n20219 );
buf ( n20221 , n20220 );
buf ( n20222 , n20221 );
nand ( n20223 , n20205 , n20222 );
buf ( n20224 , n20223 );
buf ( n20225 , n20224 );
xor ( n20226 , n20200 , n20225 );
buf ( n20227 , n18285 );
not ( n20228 , n20227 );
buf ( n20229 , n20081 );
not ( n20230 , n20229 );
or ( n20231 , n20228 , n20230 );
buf ( n20232 , n582 );
not ( n20233 , n20232 );
buf ( n20234 , n18329 );
not ( n20235 , n20234 );
or ( n20236 , n20233 , n20235 );
buf ( n20237 , n18605 );
buf ( n20238 , n18303 );
nand ( n20239 , n20237 , n20238 );
buf ( n20240 , n20239 );
buf ( n20241 , n20240 );
nand ( n20242 , n20236 , n20241 );
buf ( n20243 , n20242 );
buf ( n20244 , n20243 );
buf ( n20245 , n18316 );
nand ( n20246 , n20244 , n20245 );
buf ( n20247 , n20246 );
buf ( n20248 , n20247 );
nand ( n20249 , n20231 , n20248 );
buf ( n20250 , n20249 );
buf ( n20251 , n20250 );
not ( n20252 , n18380 );
not ( n20253 , n20054 );
or ( n20254 , n20252 , n20253 );
and ( n20255 , n18538 , n580 );
not ( n20256 , n18538 );
and ( n20257 , n20256 , n18402 );
or ( n20258 , n20255 , n20257 );
nand ( n20259 , n20258 , n18391 );
nand ( n20260 , n20254 , n20259 );
buf ( n20261 , n20260 );
buf ( n20262 , n576 );
buf ( n20263 , n13666 );
and ( n20264 , n20262 , n20263 );
buf ( n20265 , n20264 );
buf ( n20266 , n20265 );
buf ( n20267 , n18340 );
not ( n20268 , n20267 );
buf ( n20269 , n19997 );
not ( n20270 , n20269 );
or ( n20271 , n20268 , n20270 );
buf ( n20272 , n576 );
not ( n20273 , n20272 );
buf ( n20274 , n19972 );
not ( n20275 , n20274 );
or ( n20276 , n20273 , n20275 );
buf ( n20277 , n19975 );
buf ( n20278 , n7809 );
nand ( n20279 , n20277 , n20278 );
buf ( n20280 , n20279 );
buf ( n20281 , n20280 );
nand ( n20282 , n20276 , n20281 );
buf ( n20283 , n20282 );
buf ( n20284 , n20283 );
buf ( n20285 , n18365 );
nand ( n20286 , n20284 , n20285 );
buf ( n20287 , n20286 );
buf ( n20288 , n20287 );
nand ( n20289 , n20271 , n20288 );
buf ( n20290 , n20289 );
buf ( n20291 , n20290 );
xor ( n20292 , n20266 , n20291 );
buf ( n20293 , n18219 );
not ( n20294 , n20293 );
buf ( n20295 , n20023 );
not ( n20296 , n20295 );
or ( n20297 , n20294 , n20296 );
buf ( n20298 , n578 );
not ( n20299 , n20298 );
buf ( n20300 , n19651 );
not ( n20301 , n20300 );
or ( n20302 , n20299 , n20301 );
buf ( n20303 , n19534 );
buf ( n20304 , n18233 );
nand ( n20305 , n20303 , n20304 );
buf ( n20306 , n20305 );
buf ( n20307 , n20306 );
nand ( n20308 , n20302 , n20307 );
buf ( n20309 , n20308 );
buf ( n20310 , n20309 );
buf ( n20311 , n18264 );
nand ( n20312 , n20310 , n20311 );
buf ( n20313 , n20312 );
buf ( n20314 , n20313 );
nand ( n20315 , n20297 , n20314 );
buf ( n20316 , n20315 );
buf ( n20317 , n20316 );
and ( n20318 , n20292 , n20317 );
and ( n20319 , n20266 , n20291 );
or ( n20320 , n20318 , n20319 );
buf ( n20321 , n20320 );
buf ( n20322 , n20321 );
xor ( n20323 , n20261 , n20322 );
xor ( n20324 , n19980 , n20005 );
xor ( n20325 , n20324 , n20031 );
buf ( n20326 , n20325 );
buf ( n20327 , n20326 );
and ( n20328 , n20323 , n20327 );
and ( n20329 , n20261 , n20322 );
or ( n20330 , n20328 , n20329 );
buf ( n20331 , n20330 );
buf ( n20332 , n20331 );
xor ( n20333 , n20251 , n20332 );
xor ( n20334 , n20036 , n20040 );
xor ( n20335 , n20334 , n20059 );
buf ( n20336 , n20335 );
buf ( n20337 , n20336 );
and ( n20338 , n20333 , n20337 );
and ( n20339 , n20251 , n20332 );
or ( n20340 , n20338 , n20339 );
buf ( n20341 , n20340 );
buf ( n20342 , n20341 );
and ( n20343 , n20226 , n20342 );
and ( n20344 , n20200 , n20225 );
or ( n20345 , n20343 , n20344 );
buf ( n20346 , n20345 );
buf ( n20347 , n20346 );
and ( n20348 , n20183 , n20347 );
and ( n20349 , n20178 , n20182 );
or ( n20350 , n20348 , n20349 );
buf ( n20351 , n20350 );
buf ( n20352 , n20351 );
and ( n20353 , n20155 , n20352 );
and ( n20354 , n20150 , n20154 );
or ( n20355 , n20353 , n20354 );
buf ( n20356 , n20355 );
buf ( n20357 , n20356 );
xor ( n20358 , n20132 , n20357 );
xor ( n20359 , n19909 , n19913 );
xor ( n20360 , n20359 , n20109 );
buf ( n20361 , n20360 );
buf ( n20362 , n20361 );
and ( n20363 , n20358 , n20362 );
and ( n20364 , n20132 , n20357 );
or ( n20365 , n20363 , n20364 );
buf ( n20366 , n20365 );
buf ( n20367 , n20366 );
nor ( n20368 , n20128 , n20367 );
buf ( n20369 , n20368 );
nor ( n20370 , n20124 , n20369 );
buf ( n20371 , n20370 );
not ( n20372 , n20371 );
xor ( n20373 , n20132 , n20357 );
xor ( n20374 , n20373 , n20362 );
buf ( n20375 , n20374 );
xor ( n20376 , n19931 , n19935 );
xor ( n20377 , n20376 , n20104 );
buf ( n20378 , n20377 );
buf ( n20379 , n20378 );
xor ( n20380 , n19964 , n19968 );
xor ( n20381 , n20380 , n20099 );
buf ( n20382 , n20381 );
buf ( n20383 , n20382 );
buf ( n20384 , n591 );
not ( n20385 , n20384 );
buf ( n20386 , n20139 );
not ( n20387 , n20386 );
or ( n20388 , n20385 , n20387 );
not ( n20389 , n18726 );
and ( n20390 , n590 , n20389 );
not ( n20391 , n590 );
and ( n20392 , n20391 , n18726 );
nor ( n20393 , n20390 , n20392 );
buf ( n20394 , n20393 );
buf ( n20395 , n19244 );
nand ( n20396 , n20394 , n20395 );
buf ( n20397 , n20396 );
buf ( n20398 , n20397 );
nand ( n20399 , n20388 , n20398 );
buf ( n20400 , n20399 );
buf ( n20401 , n20400 );
xor ( n20402 , n20383 , n20401 );
xor ( n20403 , n20064 , n20089 );
xor ( n20404 , n20403 , n20094 );
buf ( n20405 , n20404 );
buf ( n20406 , n20405 );
buf ( n20407 , n19143 );
not ( n20408 , n20407 );
buf ( n20409 , n20167 );
not ( n20410 , n20409 );
or ( n20411 , n20408 , n20410 );
xor ( n20412 , n588 , n18909 );
buf ( n20413 , n20412 );
buf ( n20414 , n19152 );
nand ( n20415 , n20413 , n20414 );
buf ( n20416 , n20415 );
buf ( n20417 , n20416 );
nand ( n20418 , n20411 , n20417 );
buf ( n20419 , n20418 );
buf ( n20420 , n20419 );
xor ( n20421 , n20406 , n20420 );
buf ( n20422 , n18431 );
not ( n20423 , n20422 );
buf ( n20424 , n20192 );
not ( n20425 , n20424 );
or ( n20426 , n20423 , n20425 );
buf ( n20427 , n584 );
not ( n20428 , n20427 );
not ( n20429 , n18344 );
buf ( n20430 , n20429 );
not ( n20431 , n20430 );
or ( n20432 , n20428 , n20431 );
buf ( n20433 , n18759 );
buf ( n20434 , n18277 );
nand ( n20435 , n20433 , n20434 );
buf ( n20436 , n20435 );
buf ( n20437 , n20436 );
nand ( n20438 , n20432 , n20437 );
buf ( n20439 , n20438 );
buf ( n20440 , n20439 );
buf ( n20441 , n18479 );
nand ( n20442 , n20440 , n20441 );
buf ( n20443 , n20442 );
buf ( n20444 , n20443 );
nand ( n20445 , n20426 , n20444 );
buf ( n20446 , n20445 );
buf ( n20447 , n20446 );
buf ( n20448 , n576 );
buf ( n20449 , n2323 );
buf ( n20450 , n20449 );
not ( n20451 , n20450 );
buf ( n20452 , n20451 );
buf ( n20453 , n20452 );
not ( n20454 , n20453 );
buf ( n20455 , n20454 );
buf ( n20456 , n20455 );
and ( n20457 , n20448 , n20456 );
buf ( n20458 , n20457 );
buf ( n20459 , n20458 );
buf ( n20460 , n18340 );
not ( n20461 , n20460 );
buf ( n20462 , n20283 );
not ( n20463 , n20462 );
or ( n20464 , n20461 , n20463 );
xor ( n20465 , n20262 , n20263 );
buf ( n20466 , n20465 );
buf ( n20467 , n20466 );
buf ( n20468 , n18365 );
nand ( n20469 , n20467 , n20468 );
buf ( n20470 , n20469 );
buf ( n20471 , n20470 );
nand ( n20472 , n20464 , n20471 );
buf ( n20473 , n20472 );
buf ( n20474 , n20473 );
xor ( n20475 , n20459 , n20474 );
buf ( n20476 , n18219 );
not ( n20477 , n20476 );
buf ( n20478 , n20309 );
not ( n20479 , n20478 );
or ( n20480 , n20477 , n20479 );
buf ( n20481 , n13664 );
not ( n20482 , n20481 );
buf ( n20483 , n20482 );
nand ( n20484 , n20483 , n578 );
not ( n20485 , n20484 );
buf ( n20486 , n13664 );
buf ( n20487 , n20486 );
buf ( n20488 , n20487 );
buf ( n20489 , n20488 );
buf ( n20490 , n18233 );
nand ( n20491 , n20489 , n20490 );
buf ( n20492 , n20491 );
not ( n20493 , n20492 );
or ( n20494 , n20485 , n20493 );
nand ( n20495 , n20494 , n18264 );
buf ( n20496 , n20495 );
nand ( n20497 , n20480 , n20496 );
buf ( n20498 , n20497 );
buf ( n20499 , n20498 );
and ( n20500 , n20475 , n20499 );
and ( n20501 , n20459 , n20474 );
or ( n20502 , n20500 , n20501 );
buf ( n20503 , n20502 );
buf ( n20504 , n20503 );
buf ( n20505 , n18418 );
not ( n20506 , n20505 );
buf ( n20507 , n20258 );
not ( n20508 , n20507 );
or ( n20509 , n20506 , n20508 );
buf ( n20510 , n580 );
not ( n20511 , n20510 );
buf ( n20512 , n19000 );
not ( n20513 , n20512 );
or ( n20514 , n20511 , n20513 );
buf ( n20515 , n19003 );
buf ( n20516 , n18402 );
nand ( n20517 , n20515 , n20516 );
buf ( n20518 , n20517 );
buf ( n20519 , n20518 );
nand ( n20520 , n20514 , n20519 );
buf ( n20521 , n20520 );
buf ( n20522 , n20521 );
buf ( n20523 , n18391 );
nand ( n20524 , n20522 , n20523 );
buf ( n20525 , n20524 );
buf ( n20526 , n20525 );
nand ( n20527 , n20509 , n20526 );
buf ( n20528 , n20527 );
buf ( n20529 , n20528 );
xor ( n20530 , n20504 , n20529 );
xor ( n20531 , n20266 , n20291 );
xor ( n20532 , n20531 , n20317 );
buf ( n20533 , n20532 );
buf ( n20534 , n20533 );
and ( n20535 , n20530 , n20534 );
and ( n20536 , n20504 , n20529 );
or ( n20537 , n20535 , n20536 );
buf ( n20538 , n20537 );
buf ( n20539 , n20538 );
buf ( n20540 , n18285 );
not ( n20541 , n20540 );
buf ( n20542 , n20243 );
not ( n20543 , n20542 );
or ( n20544 , n20541 , n20543 );
buf ( n20545 , n582 );
not ( n20546 , n20545 );
buf ( n20547 , n19022 );
not ( n20548 , n20547 );
or ( n20549 , n20546 , n20548 );
buf ( n20550 , n18489 );
buf ( n20551 , n18303 );
nand ( n20552 , n20550 , n20551 );
buf ( n20553 , n20552 );
buf ( n20554 , n20553 );
nand ( n20555 , n20549 , n20554 );
buf ( n20556 , n20555 );
buf ( n20557 , n20556 );
buf ( n20558 , n18316 );
nand ( n20559 , n20557 , n20558 );
buf ( n20560 , n20559 );
buf ( n20561 , n20560 );
nand ( n20562 , n20544 , n20561 );
buf ( n20563 , n20562 );
buf ( n20564 , n20563 );
xor ( n20565 , n20539 , n20564 );
xor ( n20566 , n20261 , n20322 );
xor ( n20567 , n20566 , n20327 );
buf ( n20568 , n20567 );
buf ( n20569 , n20568 );
and ( n20570 , n20565 , n20569 );
and ( n20571 , n20539 , n20564 );
or ( n20572 , n20570 , n20571 );
buf ( n20573 , n20572 );
buf ( n20574 , n20573 );
xor ( n20575 , n20447 , n20574 );
buf ( n20576 , n18857 );
not ( n20577 , n20576 );
buf ( n20578 , n20217 );
not ( n20579 , n20578 );
or ( n20580 , n20577 , n20579 );
and ( n20581 , n18226 , n586 );
not ( n20582 , n18226 );
and ( n20583 , n20582 , n1766 );
or ( n20584 , n20581 , n20583 );
nand ( n20585 , n20584 , n18881 );
buf ( n20586 , n20585 );
nand ( n20587 , n20580 , n20586 );
buf ( n20588 , n20587 );
buf ( n20589 , n20588 );
and ( n20590 , n20575 , n20589 );
and ( n20591 , n20447 , n20574 );
or ( n20592 , n20590 , n20591 );
buf ( n20593 , n20592 );
buf ( n20594 , n20593 );
and ( n20595 , n20421 , n20594 );
and ( n20596 , n20406 , n20420 );
or ( n20597 , n20595 , n20596 );
buf ( n20598 , n20597 );
buf ( n20599 , n20598 );
and ( n20600 , n20402 , n20599 );
and ( n20601 , n20383 , n20401 );
or ( n20602 , n20600 , n20601 );
buf ( n20603 , n20602 );
buf ( n20604 , n20603 );
xor ( n20605 , n20379 , n20604 );
xor ( n20606 , n20150 , n20154 );
xor ( n20607 , n20606 , n20352 );
buf ( n20608 , n20607 );
buf ( n20609 , n20608 );
and ( n20610 , n20605 , n20609 );
and ( n20611 , n20379 , n20604 );
or ( n20612 , n20610 , n20611 );
buf ( n20613 , n20612 );
nor ( n20614 , n20375 , n20613 );
buf ( n20615 , n591 );
not ( n20616 , n20615 );
buf ( n20617 , n20393 );
not ( n20618 , n20617 );
or ( n20619 , n20616 , n20618 );
buf ( n20620 , n19244 );
not ( n20621 , n20620 );
buf ( n20622 , n20621 );
buf ( n20623 , n20622 );
not ( n20624 , n20623 );
and ( n20625 , n590 , n18442 );
not ( n20626 , n590 );
buf ( n20627 , n18868 );
not ( n20628 , n20627 );
buf ( n20629 , n20628 );
and ( n20630 , n20626 , n20629 );
or ( n20631 , n20625 , n20630 );
buf ( n20632 , n20631 );
nand ( n20633 , n20624 , n20632 );
buf ( n20634 , n20633 );
buf ( n20635 , n20634 );
nand ( n20636 , n20619 , n20635 );
buf ( n20637 , n20636 );
buf ( n20638 , n20637 );
xor ( n20639 , n20200 , n20225 );
xor ( n20640 , n20639 , n20342 );
buf ( n20641 , n20640 );
buf ( n20642 , n20641 );
xor ( n20643 , n20638 , n20642 );
xor ( n20644 , n20251 , n20332 );
xor ( n20645 , n20644 , n20337 );
buf ( n20646 , n20645 );
buf ( n20647 , n20646 );
buf ( n20648 , n19143 );
not ( n20649 , n20648 );
buf ( n20650 , n20412 );
not ( n20651 , n20650 );
or ( n20652 , n20649 , n20651 );
and ( n20653 , n588 , n19946 );
not ( n20654 , n588 );
and ( n20655 , n20654 , n13592 );
or ( n20656 , n20653 , n20655 );
buf ( n20657 , n20656 );
buf ( n20658 , n19152 );
nand ( n20659 , n20657 , n20658 );
buf ( n20660 , n20659 );
buf ( n20661 , n20660 );
nand ( n20662 , n20652 , n20661 );
buf ( n20663 , n20662 );
buf ( n20664 , n20663 );
xor ( n20665 , n20647 , n20664 );
buf ( n20666 , n19244 );
not ( n20667 , n20666 );
and ( n20668 , n590 , n20163 );
not ( n20669 , n590 );
and ( n20670 , n20669 , n20160 );
or ( n20671 , n20668 , n20670 );
buf ( n20672 , n20671 );
not ( n20673 , n20672 );
or ( n20674 , n20667 , n20673 );
buf ( n20675 , n20631 );
buf ( n20676 , n591 );
nand ( n20677 , n20675 , n20676 );
buf ( n20678 , n20677 );
buf ( n20679 , n20678 );
nand ( n20680 , n20674 , n20679 );
buf ( n20681 , n20680 );
buf ( n20682 , n20681 );
and ( n20683 , n20665 , n20682 );
and ( n20684 , n20647 , n20664 );
or ( n20685 , n20683 , n20684 );
buf ( n20686 , n20685 );
buf ( n20687 , n20686 );
and ( n20688 , n20643 , n20687 );
and ( n20689 , n20638 , n20642 );
or ( n20690 , n20688 , n20689 );
buf ( n20691 , n20690 );
buf ( n20692 , n20691 );
xor ( n20693 , n20178 , n20182 );
xor ( n20694 , n20693 , n20347 );
buf ( n20695 , n20694 );
buf ( n20696 , n20695 );
xor ( n20697 , n20692 , n20696 );
xor ( n20698 , n20383 , n20401 );
xor ( n20699 , n20698 , n20599 );
buf ( n20700 , n20699 );
buf ( n20701 , n20700 );
xor ( n20702 , n20697 , n20701 );
buf ( n20703 , n20702 );
xor ( n20704 , n20406 , n20420 );
xor ( n20705 , n20704 , n20594 );
buf ( n20706 , n20705 );
buf ( n20707 , n20706 );
xor ( n20708 , n20638 , n20642 );
xor ( n20709 , n20708 , n20687 );
buf ( n20710 , n20709 );
buf ( n20711 , n20710 );
xor ( n20712 , n20707 , n20711 );
buf ( n20713 , n18431 );
not ( n20714 , n20713 );
buf ( n20715 , n20439 );
not ( n20716 , n20715 );
or ( n20717 , n20714 , n20716 );
buf ( n20718 , n584 );
not ( n20719 , n20718 );
buf ( n20720 , n18960 );
not ( n20721 , n20720 );
or ( n20722 , n20719 , n20721 );
buf ( n20723 , n18357 );
buf ( n20724 , n18277 );
nand ( n20725 , n20723 , n20724 );
buf ( n20726 , n20725 );
buf ( n20727 , n20726 );
nand ( n20728 , n20722 , n20727 );
buf ( n20729 , n20728 );
buf ( n20730 , n20729 );
buf ( n20731 , n18479 );
nand ( n20732 , n20730 , n20731 );
buf ( n20733 , n20732 );
buf ( n20734 , n20733 );
nand ( n20735 , n20717 , n20734 );
buf ( n20736 , n20735 );
buf ( n20737 , n20736 );
buf ( n20738 , C0 );
buf ( n20739 , n20738 );
buf ( n20740 , n18340 );
not ( n20741 , n20740 );
buf ( n20742 , n20466 );
not ( n20743 , n20742 );
or ( n20744 , n20741 , n20743 );
xor ( n20745 , n20448 , n20456 );
buf ( n20746 , n20745 );
buf ( n20747 , n20746 );
buf ( n20748 , n18365 );
nand ( n20749 , n20747 , n20748 );
buf ( n20750 , n20749 );
buf ( n20751 , n20750 );
nand ( n20752 , n20744 , n20751 );
buf ( n20753 , n20752 );
buf ( n20754 , n20753 );
xor ( n20755 , n20739 , n20754 );
buf ( n20756 , C0 );
buf ( n20757 , n20756 );
buf ( n20758 , C0 );
buf ( n20759 , n20758 );
buf ( n20760 , n576 );
not ( n20761 , n20760 );
buf ( n20762 , C1 );
or ( n20763 , n20761 , C0 );
buf ( n20764 , C1 );
buf ( n20765 , n20764 );
nand ( n20766 , n20763 , n20765 );
buf ( n20767 , n20766 );
not ( n20768 , n20767 );
not ( n20769 , n18340 );
or ( n20770 , n20768 , n20769 );
buf ( n20771 , n576 );
not ( n20772 , n20771 );
buf ( n20773 , C1 );
or ( n20774 , n20772 , C0 );
buf ( n20775 , C1 );
buf ( n20776 , n20775 );
nand ( n20777 , n20774 , n20776 );
buf ( n20778 , n20777 );
buf ( n20779 , n20778 );
buf ( n20780 , n18365 );
nand ( n20781 , n20779 , n20780 );
buf ( n20782 , n20781 );
nand ( n20783 , n20770 , n20782 );
buf ( n20784 , n20783 );
xor ( n20785 , n20759 , n20784 );
buf ( n20786 , C1 );
buf ( n20787 , n20786 );
buf ( n20788 , n577 );
buf ( n20789 , n578 );
and ( n20790 , n20788 , n20789 );
buf ( n20791 , n7809 );
nor ( n20792 , n20790 , n20791 );
buf ( n20793 , n20792 );
buf ( n20794 , n20793 );
and ( n20795 , n20787 , n20794 );
buf ( n20796 , n20795 );
buf ( n20797 , n20796 );
not ( n20798 , n20778 );
not ( n20799 , n18340 );
or ( n20800 , n20798 , n20799 );
buf ( n20801 , n576 );
buf ( n20802 , C0 );
xor ( n20803 , n20801 , n20802 );
buf ( n20804 , n20803 );
buf ( n20805 , n20804 );
buf ( n20806 , n18365 );
nand ( n20807 , n20805 , n20806 );
buf ( n20808 , n20807 );
nand ( n20809 , n20800 , n20808 );
buf ( n20810 , n20809 );
and ( n20811 , n20797 , n20810 );
buf ( n20812 , n20811 );
buf ( n20813 , n20812 );
and ( n20814 , n20785 , n20813 );
or ( n20815 , n20814 , C0 );
buf ( n20816 , n20815 );
buf ( n20817 , n20816 );
xor ( n20818 , n20757 , n20817 );
buf ( n20819 , n18340 );
not ( n20820 , n20819 );
buf ( n20821 , n20746 );
not ( n20822 , n20821 );
or ( n20823 , n20820 , n20822 );
buf ( n20824 , n20767 );
buf ( n20825 , n18365 );
nand ( n20826 , n20824 , n20825 );
buf ( n20827 , n20826 );
buf ( n20828 , n20827 );
nand ( n20829 , n20823 , n20828 );
buf ( n20830 , n20829 );
buf ( n20831 , n20830 );
and ( n20832 , n20818 , n20831 );
or ( n20833 , n20832 , C0 );
buf ( n20834 , n20833 );
buf ( n20835 , n20834 );
and ( n20836 , n20755 , n20835 );
or ( n20837 , n20836 , C0 );
buf ( n20838 , n20837 );
buf ( n20839 , n20838 );
xor ( n20840 , n20459 , n20474 );
xor ( n20841 , n20840 , n20499 );
buf ( n20842 , n20841 );
buf ( n20843 , n20842 );
xor ( n20844 , n20839 , n20843 );
buf ( n20845 , n18418 );
not ( n20846 , n20845 );
buf ( n20847 , n20521 );
not ( n20848 , n20847 );
or ( n20849 , n20846 , n20848 );
not ( n20850 , n580 );
not ( n20851 , n18981 );
or ( n20852 , n20850 , n20851 );
buf ( n20853 , n19555 );
buf ( n20854 , n18402 );
nand ( n20855 , n20853 , n20854 );
buf ( n20856 , n20855 );
nand ( n20857 , n20852 , n20856 );
nand ( n20858 , n20857 , n18391 );
buf ( n20859 , n20858 );
nand ( n20860 , n20849 , n20859 );
buf ( n20861 , n20860 );
buf ( n20862 , n20861 );
and ( n20863 , n20844 , n20862 );
and ( n20864 , n20839 , n20843 );
or ( n20865 , n20863 , n20864 );
buf ( n20866 , n20865 );
buf ( n20867 , n20866 );
buf ( n20868 , n18285 );
not ( n20869 , n20868 );
buf ( n20870 , n20556 );
not ( n20871 , n20870 );
or ( n20872 , n20869 , n20871 );
buf ( n20873 , n582 );
not ( n20874 , n20873 );
buf ( n20875 , n18569 );
not ( n20876 , n20875 );
or ( n20877 , n20874 , n20876 );
buf ( n20878 , n18566 );
buf ( n20879 , n18303 );
nand ( n20880 , n20878 , n20879 );
buf ( n20881 , n20880 );
buf ( n20882 , n20881 );
nand ( n20883 , n20877 , n20882 );
buf ( n20884 , n20883 );
buf ( n20885 , n20884 );
buf ( n20886 , n18316 );
nand ( n20887 , n20885 , n20886 );
buf ( n20888 , n20887 );
buf ( n20889 , n20888 );
nand ( n20890 , n20872 , n20889 );
buf ( n20891 , n20890 );
buf ( n20892 , n20891 );
xor ( n20893 , n20867 , n20892 );
xor ( n20894 , n20504 , n20529 );
xor ( n20895 , n20894 , n20534 );
buf ( n20896 , n20895 );
buf ( n20897 , n20896 );
and ( n20898 , n20893 , n20897 );
and ( n20899 , n20867 , n20892 );
or ( n20900 , n20898 , n20899 );
buf ( n20901 , n20900 );
buf ( n20902 , n20901 );
xor ( n20903 , n20737 , n20902 );
xor ( n20904 , n20539 , n20564 );
xor ( n20905 , n20904 , n20569 );
buf ( n20906 , n20905 );
buf ( n20907 , n20906 );
and ( n20908 , n20903 , n20907 );
and ( n20909 , n20737 , n20902 );
or ( n20910 , n20908 , n20909 );
buf ( n20911 , n20910 );
buf ( n20912 , n20911 );
xor ( n20913 , n20447 , n20574 );
xor ( n20914 , n20913 , n20589 );
buf ( n20915 , n20914 );
buf ( n20916 , n20915 );
xor ( n20917 , n20912 , n20916 );
buf ( n20918 , n18857 );
not ( n20919 , n20918 );
buf ( n20920 , n20584 );
not ( n20921 , n20920 );
or ( n20922 , n20919 , n20921 );
buf ( n20923 , n586 );
not ( n20924 , n20923 );
buf ( n20925 , n9498 );
not ( n20926 , n20925 );
or ( n20927 , n20924 , n20926 );
buf ( n20928 , n9497 );
buf ( n20929 , n18840 );
nand ( n20930 , n20928 , n20929 );
buf ( n20931 , n20930 );
buf ( n20932 , n20931 );
nand ( n20933 , n20927 , n20932 );
buf ( n20934 , n20933 );
buf ( n20935 , n20934 );
buf ( n20936 , n18881 );
nand ( n20937 , n20935 , n20936 );
buf ( n20938 , n20937 );
buf ( n20939 , n20938 );
nand ( n20940 , n20922 , n20939 );
buf ( n20941 , n20940 );
buf ( n20942 , n20941 );
buf ( n20943 , n19152 );
not ( n20944 , n20943 );
xnor ( n20945 , n588 , n18682 );
buf ( n20946 , n20945 );
not ( n20947 , n20946 );
or ( n20948 , n20944 , n20947 );
buf ( n20949 , n20656 );
buf ( n20950 , n19143 );
nand ( n20951 , n20949 , n20950 );
buf ( n20952 , n20951 );
buf ( n20953 , n20952 );
nand ( n20954 , n20948 , n20953 );
buf ( n20955 , n20954 );
buf ( n20956 , n20955 );
xor ( n20957 , n20942 , n20956 );
buf ( n20958 , n18431 );
not ( n20959 , n20958 );
buf ( n20960 , n20729 );
not ( n20961 , n20960 );
or ( n20962 , n20959 , n20961 );
buf ( n20963 , n584 );
not ( n20964 , n20963 );
buf ( n20965 , n18329 );
not ( n20966 , n20965 );
or ( n20967 , n20964 , n20966 );
buf ( n20968 , n18599 );
not ( n20969 , n20968 );
buf ( n20970 , n18277 );
nand ( n20971 , n20969 , n20970 );
buf ( n20972 , n20971 );
buf ( n20973 , n20972 );
nand ( n20974 , n20967 , n20973 );
buf ( n20975 , n20974 );
buf ( n20976 , n20975 );
buf ( n20977 , n18479 );
nand ( n20978 , n20976 , n20977 );
buf ( n20979 , n20978 );
buf ( n20980 , n20979 );
nand ( n20981 , n20962 , n20980 );
buf ( n20982 , n20981 );
buf ( n20983 , n20982 );
buf ( n20984 , n18219 );
not ( n20985 , n20984 );
nand ( n20986 , n20492 , n20484 );
buf ( n20987 , n20986 );
not ( n20988 , n20987 );
or ( n20989 , n20985 , n20988 );
buf ( n20990 , n578 );
not ( n20991 , n20990 );
buf ( n20992 , n19972 );
not ( n20993 , n20992 );
or ( n20994 , n20991 , n20993 );
buf ( n20995 , n18233 );
buf ( n20996 , n2337 );
buf ( n20997 , n20996 );
buf ( n20998 , n20997 );
buf ( n20999 , n20998 );
nand ( n21000 , n20995 , n20999 );
buf ( n21001 , n21000 );
buf ( n21002 , n21001 );
nand ( n21003 , n20994 , n21002 );
buf ( n21004 , n21003 );
buf ( n21005 , n21004 );
buf ( n21006 , n18264 );
nand ( n21007 , n21005 , n21006 );
buf ( n21008 , n21007 );
buf ( n21009 , n21008 );
nand ( n21010 , n20989 , n21009 );
buf ( n21011 , n21010 );
buf ( n21012 , n21011 );
xor ( n21013 , n20739 , n20754 );
xor ( n21014 , n21013 , n20835 );
buf ( n21015 , n21014 );
buf ( n21016 , n21015 );
xor ( n21017 , n21012 , n21016 );
not ( n21018 , n18418 );
not ( n21019 , n20857 );
or ( n21020 , n21018 , n21019 );
buf ( n21021 , n580 );
not ( n21022 , n21021 );
buf ( n21023 , n19651 );
not ( n21024 , n21023 );
or ( n21025 , n21022 , n21024 );
buf ( n21026 , n19534 );
buf ( n21027 , n18402 );
nand ( n21028 , n21026 , n21027 );
buf ( n21029 , n21028 );
buf ( n21030 , n21029 );
nand ( n21031 , n21025 , n21030 );
buf ( n21032 , n21031 );
buf ( n21033 , n21032 );
buf ( n21034 , n18391 );
nand ( n21035 , n21033 , n21034 );
buf ( n21036 , n21035 );
nand ( n21037 , n21020 , n21036 );
buf ( n21038 , n21037 );
and ( n21039 , n21017 , n21038 );
and ( n21040 , n21012 , n21016 );
or ( n21041 , n21039 , n21040 );
buf ( n21042 , n21041 );
buf ( n21043 , n21042 );
buf ( n21044 , n18285 );
not ( n21045 , n21044 );
buf ( n21046 , n20884 );
not ( n21047 , n21046 );
or ( n21048 , n21045 , n21047 );
buf ( n21049 , n582 );
not ( n21050 , n21049 );
buf ( n21051 , n18538 );
not ( n21052 , n21051 );
or ( n21053 , n21050 , n21052 );
buf ( n21054 , n18541 );
buf ( n21055 , n18303 );
nand ( n21056 , n21054 , n21055 );
buf ( n21057 , n21056 );
buf ( n21058 , n21057 );
nand ( n21059 , n21053 , n21058 );
buf ( n21060 , n21059 );
buf ( n21061 , n21060 );
buf ( n21062 , n18316 );
nand ( n21063 , n21061 , n21062 );
buf ( n21064 , n21063 );
buf ( n21065 , n21064 );
nand ( n21066 , n21048 , n21065 );
buf ( n21067 , n21066 );
buf ( n21068 , n21067 );
xor ( n21069 , n21043 , n21068 );
xor ( n21070 , n20839 , n20843 );
xor ( n21071 , n21070 , n20862 );
buf ( n21072 , n21071 );
buf ( n21073 , n21072 );
and ( n21074 , n21069 , n21073 );
and ( n21075 , n21043 , n21068 );
or ( n21076 , n21074 , n21075 );
buf ( n21077 , n21076 );
buf ( n21078 , n21077 );
xor ( n21079 , n20983 , n21078 );
xor ( n21080 , n20867 , n20892 );
xor ( n21081 , n21080 , n20897 );
buf ( n21082 , n21081 );
buf ( n21083 , n21082 );
and ( n21084 , n21079 , n21083 );
and ( n21085 , n20983 , n21078 );
or ( n21086 , n21084 , n21085 );
buf ( n21087 , n21086 );
buf ( n21088 , n21087 );
and ( n21089 , n20957 , n21088 );
and ( n21090 , n20942 , n20956 );
or ( n21091 , n21089 , n21090 );
buf ( n21092 , n21091 );
buf ( n21093 , n21092 );
and ( n21094 , n20917 , n21093 );
and ( n21095 , n20912 , n20916 );
or ( n21096 , n21094 , n21095 );
buf ( n21097 , n21096 );
buf ( n21098 , n21097 );
and ( n21099 , n20712 , n21098 );
and ( n21100 , n20707 , n20711 );
or ( n21101 , n21099 , n21100 );
buf ( n21102 , n21101 );
nor ( n21103 , n20703 , n21102 );
xor ( n21104 , n20379 , n20604 );
xor ( n21105 , n21104 , n20609 );
buf ( n21106 , n21105 );
xor ( n21107 , n20692 , n20696 );
and ( n21108 , n21107 , n20701 );
and ( n21109 , n20692 , n20696 );
or ( n21110 , n21108 , n21109 );
buf ( n21111 , n21110 );
nor ( n21112 , n21106 , n21111 );
nor ( n21113 , n20614 , n21103 , n21112 );
not ( n21114 , n21113 );
xor ( n21115 , n20707 , n20711 );
xor ( n21116 , n21115 , n21098 );
buf ( n21117 , n21116 );
buf ( n21118 , n21117 );
not ( n21119 , n21118 );
buf ( n21120 , n21119 );
buf ( n21121 , n21120 );
xor ( n21122 , n20647 , n20664 );
xor ( n21123 , n21122 , n20682 );
buf ( n21124 , n21123 );
buf ( n21125 , n21124 );
buf ( n21126 , n591 );
not ( n21127 , n21126 );
buf ( n21128 , n20671 );
not ( n21129 , n21128 );
or ( n21130 , n21127 , n21129 );
buf ( n21131 , n590 );
not ( n21132 , n21131 );
buf ( n21133 , n19282 );
not ( n21134 , n21133 );
or ( n21135 , n21132 , n21134 );
buf ( n21136 , n590 );
not ( n21137 , n21136 );
buf ( n21138 , n18909 );
nand ( n21139 , n21137 , n21138 );
buf ( n21140 , n21139 );
buf ( n21141 , n21140 );
nand ( n21142 , n21135 , n21141 );
buf ( n21143 , n21142 );
buf ( n21144 , n21143 );
buf ( n21145 , n21144 );
buf ( n21146 , n21145 );
buf ( n21147 , n21146 );
buf ( n21148 , n19244 );
nand ( n21149 , n21147 , n21148 );
buf ( n21150 , n21149 );
buf ( n21151 , n21150 );
nand ( n21152 , n21130 , n21151 );
buf ( n21153 , n21152 );
buf ( n21154 , n21153 );
buf ( n21155 , n18857 );
not ( n21156 , n21155 );
buf ( n21157 , n20934 );
not ( n21158 , n21157 );
or ( n21159 , n21156 , n21158 );
buf ( n21160 , n586 );
not ( n21161 , n21160 );
buf ( n21162 , n20429 );
not ( n21163 , n21162 );
or ( n21164 , n21161 , n21163 );
buf ( n21165 , n18344 );
buf ( n21166 , n18840 );
nand ( n21167 , n21165 , n21166 );
buf ( n21168 , n21167 );
buf ( n21169 , n21168 );
nand ( n21170 , n21164 , n21169 );
buf ( n21171 , n21170 );
buf ( n21172 , n21171 );
buf ( n21173 , n18881 );
nand ( n21174 , n21172 , n21173 );
buf ( n21175 , n21174 );
buf ( n21176 , n21175 );
nand ( n21177 , n21159 , n21176 );
buf ( n21178 , n21177 );
buf ( n21179 , n21178 );
buf ( n21180 , n18431 );
not ( n21181 , n21180 );
buf ( n21182 , n20975 );
not ( n21183 , n21182 );
or ( n21184 , n21181 , n21183 );
buf ( n21185 , n584 );
not ( n21186 , n21185 );
buf ( n21187 , n19022 );
not ( n21188 , n21187 );
or ( n21189 , n21186 , n21188 );
buf ( n21190 , n18489 );
buf ( n21191 , n18277 );
nand ( n21192 , n21190 , n21191 );
buf ( n21193 , n21192 );
buf ( n21194 , n21193 );
nand ( n21195 , n21189 , n21194 );
buf ( n21196 , n21195 );
buf ( n21197 , n21196 );
buf ( n21198 , n18479 );
nand ( n21199 , n21197 , n21198 );
buf ( n21200 , n21199 );
buf ( n21201 , n21200 );
nand ( n21202 , n21184 , n21201 );
buf ( n21203 , n21202 );
buf ( n21204 , n21203 );
buf ( n21205 , n18219 );
not ( n21206 , n21205 );
buf ( n21207 , n21004 );
not ( n21208 , n21207 );
or ( n21209 , n21206 , n21208 );
buf ( n21210 , n578 );
not ( n21211 , n21210 );
buf ( n21212 , n13666 );
not ( n21213 , n21212 );
buf ( n21214 , n21213 );
buf ( n21215 , n21214 );
not ( n21216 , n21215 );
or ( n21217 , n21211 , n21216 );
buf ( n21218 , n13666 );
not ( n21219 , n21218 );
buf ( n21220 , n21219 );
buf ( n21221 , n21220 );
not ( n21222 , n21221 );
buf ( n21223 , n21222 );
buf ( n21224 , n21223 );
buf ( n21225 , n18233 );
nand ( n21226 , n21224 , n21225 );
buf ( n21227 , n21226 );
buf ( n21228 , n21227 );
nand ( n21229 , n21217 , n21228 );
buf ( n21230 , n21229 );
buf ( n21231 , n21230 );
buf ( n21232 , n18264 );
nand ( n21233 , n21231 , n21232 );
buf ( n21234 , n21233 );
buf ( n21235 , n21234 );
nand ( n21236 , n21209 , n21235 );
buf ( n21237 , n21236 );
buf ( n21238 , n21237 );
buf ( n21239 , C0 );
buf ( n21240 , n21239 );
xor ( n21241 , n21238 , n21240 );
buf ( n21242 , n18418 );
not ( n21243 , n21242 );
buf ( n21244 , n21032 );
not ( n21245 , n21244 );
or ( n21246 , n21243 , n21245 );
buf ( n21247 , n580 );
not ( n21248 , n21247 );
buf ( n21249 , n19633 );
not ( n21250 , n21249 );
or ( n21251 , n21248 , n21250 );
buf ( n21252 , n20488 );
buf ( n21253 , n18402 );
nand ( n21254 , n21252 , n21253 );
buf ( n21255 , n21254 );
buf ( n21256 , n21255 );
nand ( n21257 , n21251 , n21256 );
buf ( n21258 , n21257 );
buf ( n21259 , n21258 );
buf ( n21260 , n18391 );
nand ( n21261 , n21259 , n21260 );
buf ( n21262 , n21261 );
buf ( n21263 , n21262 );
nand ( n21264 , n21246 , n21263 );
buf ( n21265 , n21264 );
buf ( n21266 , n21265 );
and ( n21267 , n21241 , n21266 );
or ( n21268 , n21267 , C0 );
buf ( n21269 , n21268 );
buf ( n21270 , n21269 );
buf ( n21271 , n18285 );
not ( n21272 , n21271 );
buf ( n21273 , n21060 );
not ( n21274 , n21273 );
or ( n21275 , n21272 , n21274 );
buf ( n21276 , n582 );
not ( n21277 , n21276 );
buf ( n21278 , n19000 );
not ( n21279 , n21278 );
or ( n21280 , n21277 , n21279 );
buf ( n21281 , n18997 );
buf ( n21282 , n18303 );
nand ( n21283 , n21281 , n21282 );
buf ( n21284 , n21283 );
buf ( n21285 , n21284 );
nand ( n21286 , n21280 , n21285 );
buf ( n21287 , n21286 );
buf ( n21288 , n21287 );
buf ( n21289 , n18316 );
nand ( n21290 , n21288 , n21289 );
buf ( n21291 , n21290 );
buf ( n21292 , n21291 );
nand ( n21293 , n21275 , n21292 );
buf ( n21294 , n21293 );
buf ( n21295 , n21294 );
xor ( n21296 , n21270 , n21295 );
xor ( n21297 , n21012 , n21016 );
xor ( n21298 , n21297 , n21038 );
buf ( n21299 , n21298 );
buf ( n21300 , n21299 );
and ( n21301 , n21296 , n21300 );
and ( n21302 , n21270 , n21295 );
or ( n21303 , n21301 , n21302 );
buf ( n21304 , n21303 );
buf ( n21305 , n21304 );
xor ( n21306 , n21204 , n21305 );
xor ( n21307 , n21043 , n21068 );
xor ( n21308 , n21307 , n21073 );
buf ( n21309 , n21308 );
buf ( n21310 , n21309 );
and ( n21311 , n21306 , n21310 );
and ( n21312 , n21204 , n21305 );
or ( n21313 , n21311 , n21312 );
buf ( n21314 , n21313 );
buf ( n21315 , n21314 );
xor ( n21316 , n21179 , n21315 );
not ( n21317 , n19143 );
not ( n21318 , n20945 );
or ( n21319 , n21317 , n21318 );
buf ( n21320 , n588 );
not ( n21321 , n21320 );
buf ( n21322 , n18894 );
not ( n21323 , n21322 );
or ( n21324 , n21321 , n21323 );
buf ( n21325 , n18894 );
buf ( n21326 , n588 );
or ( n21327 , n21325 , n21326 );
buf ( n21328 , n21327 );
buf ( n21329 , n21328 );
nand ( n21330 , n21324 , n21329 );
buf ( n21331 , n21330 );
nand ( n21332 , n19152 , n21331 );
nand ( n21333 , n21319 , n21332 );
buf ( n21334 , n21333 );
and ( n21335 , n21316 , n21334 );
and ( n21336 , n21179 , n21315 );
or ( n21337 , n21335 , n21336 );
buf ( n21338 , n21337 );
buf ( n21339 , n21338 );
xor ( n21340 , n21154 , n21339 );
xor ( n21341 , n20737 , n20902 );
xor ( n21342 , n21341 , n20907 );
buf ( n21343 , n21342 );
buf ( n21344 , n21343 );
and ( n21345 , n21340 , n21344 );
and ( n21346 , n21154 , n21339 );
or ( n21347 , n21345 , n21346 );
buf ( n21348 , n21347 );
buf ( n21349 , n21348 );
xor ( n21350 , n21125 , n21349 );
xor ( n21351 , n20912 , n20916 );
xor ( n21352 , n21351 , n21093 );
buf ( n21353 , n21352 );
buf ( n21354 , n21353 );
and ( n21355 , n21350 , n21354 );
and ( n21356 , n21125 , n21349 );
or ( n21357 , n21355 , n21356 );
buf ( n21358 , n21357 );
buf ( n21359 , n21358 );
not ( n21360 , n21359 );
buf ( n21361 , n21360 );
buf ( n21362 , n21361 );
nand ( n21363 , n21121 , n21362 );
buf ( n21364 , n21363 );
not ( n21365 , n21364 );
xor ( n21366 , n21125 , n21349 );
xor ( n21367 , n21366 , n21354 );
buf ( n21368 , n21367 );
buf ( n21369 , n21368 );
xor ( n21370 , n20942 , n20956 );
xor ( n21371 , n21370 , n21088 );
buf ( n21372 , n21371 );
buf ( n21373 , n21372 );
buf ( n21374 , n591 );
not ( n21375 , n21374 );
buf ( n21376 , n21143 );
not ( n21377 , n21376 );
or ( n21378 , n21375 , n21377 );
and ( n21379 , n590 , n13600 );
not ( n21380 , n590 );
and ( n21381 , n21380 , n13592 );
or ( n21382 , n21379 , n21381 );
buf ( n21383 , n21382 );
buf ( n21384 , n19244 );
nand ( n21385 , n21383 , n21384 );
buf ( n21386 , n21385 );
buf ( n21387 , n21386 );
nand ( n21388 , n21378 , n21387 );
buf ( n21389 , n21388 );
buf ( n21390 , n21389 );
xor ( n21391 , n20983 , n21078 );
xor ( n21392 , n21391 , n21083 );
buf ( n21393 , n21392 );
buf ( n21394 , n21393 );
xor ( n21395 , n21390 , n21394 );
buf ( n21396 , C0 );
buf ( n21397 , n21396 );
buf ( n21398 , n18219 );
not ( n21399 , n21398 );
buf ( n21400 , n21230 );
not ( n21401 , n21400 );
or ( n21402 , n21399 , n21401 );
not ( n21403 , n578 );
buf ( n21404 , n20449 );
not ( n21405 , n21404 );
buf ( n21406 , n21405 );
not ( n21407 , n21406 );
or ( n21408 , n21403 , n21407 );
buf ( n21409 , n18233 );
buf ( n21410 , n20449 );
nand ( n21411 , n21409 , n21410 );
buf ( n21412 , n21411 );
nand ( n21413 , n21408 , n21412 );
buf ( n21414 , n21413 );
buf ( n21415 , n18264 );
nand ( n21416 , n21414 , n21415 );
buf ( n21417 , n21416 );
buf ( n21418 , n21417 );
nand ( n21419 , n21402 , n21418 );
buf ( n21420 , n21419 );
buf ( n21421 , n21420 );
xor ( n21422 , n21397 , n21421 );
buf ( n21423 , C0 );
buf ( n21424 , n21423 );
not ( n21425 , n18219 );
not ( n21426 , n21413 );
or ( n21427 , n21425 , n21426 );
buf ( n21428 , n578 );
not ( n21429 , n21428 );
or ( n21430 , n21429 , C0 );
buf ( n21431 , C1 );
buf ( n21432 , n21431 );
nand ( n21433 , n21430 , n21432 );
buf ( n21434 , n21433 );
nand ( n21435 , n21434 , n18264 );
nand ( n21436 , n21427 , n21435 );
buf ( n21437 , n21436 );
xor ( n21438 , n21424 , n21437 );
buf ( n21439 , C0 );
buf ( n21440 , n21439 );
buf ( n21441 , n18219 );
not ( n21442 , n21441 );
buf ( n21443 , n21434 );
not ( n21444 , n21443 );
or ( n21445 , n21442 , n21444 );
buf ( n21446 , n578 );
not ( n21447 , n21446 );
or ( n21448 , n21447 , C0 );
buf ( n21449 , C1 );
buf ( n21450 , n21449 );
nand ( n21451 , n21448 , n21450 );
buf ( n21452 , n21451 );
buf ( n21453 , n21452 );
buf ( n21454 , n18264 );
nand ( n21455 , n21453 , n21454 );
buf ( n21456 , n21455 );
buf ( n21457 , n21456 );
nand ( n21458 , n21445 , n21457 );
buf ( n21459 , n21458 );
buf ( n21460 , n21459 );
xor ( n21461 , n21440 , n21460 );
buf ( n21462 , C1 );
buf ( n21463 , n21462 );
buf ( n21464 , n579 );
buf ( n21465 , n580 );
and ( n21466 , n21464 , n21465 );
buf ( n21467 , n18233 );
nor ( n21468 , n21466 , n21467 );
buf ( n21469 , n21468 );
buf ( n21470 , n21469 );
and ( n21471 , n21463 , n21470 );
buf ( n21472 , n21471 );
buf ( n21473 , n21472 );
buf ( n21474 , n18219 );
not ( n21475 , n21474 );
buf ( n21476 , n21452 );
not ( n21477 , n21476 );
or ( n21478 , n21475 , n21477 );
buf ( n21479 , C0 );
buf ( n21480 , n18233 );
or ( n21481 , n21479 , n21480 );
nand ( n21482 , n21481 , C1 );
buf ( n21483 , n21482 );
buf ( n21484 , n21483 );
buf ( n21485 , n18264 );
nand ( n21486 , n21484 , n21485 );
buf ( n21487 , n21486 );
buf ( n21488 , n21487 );
nand ( n21489 , n21478 , n21488 );
buf ( n21490 , n21489 );
buf ( n21491 , n21490 );
and ( n21492 , n21473 , n21491 );
buf ( n21493 , n21492 );
buf ( n21494 , n21493 );
and ( n21495 , n21461 , n21494 );
or ( n21496 , n21495 , C0 );
buf ( n21497 , n21496 );
buf ( n21498 , n21497 );
and ( n21499 , n21438 , n21498 );
or ( n21500 , n21499 , C0 );
buf ( n21501 , n21500 );
buf ( n21502 , n21501 );
and ( n21503 , n21422 , n21502 );
or ( n21504 , n21503 , C0 );
buf ( n21505 , n21504 );
buf ( n21506 , n21505 );
xor ( n21507 , n21238 , n21240 );
xor ( n21508 , n21507 , n21266 );
buf ( n21509 , n21508 );
buf ( n21510 , n21509 );
xor ( n21511 , n21506 , n21510 );
buf ( n21512 , n18285 );
not ( n21513 , n21512 );
buf ( n21514 , n21287 );
not ( n21515 , n21514 );
or ( n21516 , n21513 , n21515 );
and ( n21517 , n13663 , n18303 );
not ( n21518 , n13663 );
and ( n21519 , n21518 , n582 );
or ( n21520 , n21517 , n21519 );
buf ( n21521 , n21520 );
buf ( n21522 , n18316 );
nand ( n21523 , n21521 , n21522 );
buf ( n21524 , n21523 );
buf ( n21525 , n21524 );
nand ( n21526 , n21516 , n21525 );
buf ( n21527 , n21526 );
buf ( n21528 , n21527 );
and ( n21529 , n21511 , n21528 );
and ( n21530 , n21506 , n21510 );
or ( n21531 , n21529 , n21530 );
buf ( n21532 , n21531 );
buf ( n21533 , n21532 );
buf ( n21534 , n18431 );
not ( n21535 , n21534 );
buf ( n21536 , n21196 );
not ( n21537 , n21536 );
or ( n21538 , n21535 , n21537 );
buf ( n21539 , n584 );
not ( n21540 , n21539 );
buf ( n21541 , n18569 );
not ( n21542 , n21541 );
or ( n21543 , n21540 , n21542 );
buf ( n21544 , n18566 );
buf ( n21545 , n18277 );
nand ( n21546 , n21544 , n21545 );
buf ( n21547 , n21546 );
buf ( n21548 , n21547 );
nand ( n21549 , n21543 , n21548 );
buf ( n21550 , n21549 );
buf ( n21551 , n21550 );
buf ( n21552 , n18479 );
nand ( n21553 , n21551 , n21552 );
buf ( n21554 , n21553 );
buf ( n21555 , n21554 );
nand ( n21556 , n21538 , n21555 );
buf ( n21557 , n21556 );
buf ( n21558 , n21557 );
xor ( n21559 , n21533 , n21558 );
xor ( n21560 , n21270 , n21295 );
xor ( n21561 , n21560 , n21300 );
buf ( n21562 , n21561 );
buf ( n21563 , n21562 );
and ( n21564 , n21559 , n21563 );
and ( n21565 , n21533 , n21558 );
or ( n21566 , n21564 , n21565 );
buf ( n21567 , n21566 );
buf ( n21568 , n21567 );
buf ( n21569 , n18857 );
not ( n21570 , n21569 );
buf ( n21571 , n21171 );
not ( n21572 , n21571 );
or ( n21573 , n21570 , n21572 );
and ( n21574 , n586 , n18960 );
not ( n21575 , n586 );
and ( n21576 , n21575 , n18357 );
or ( n21577 , n21574 , n21576 );
buf ( n21578 , n21577 );
buf ( n21579 , n18881 );
nand ( n21580 , n21578 , n21579 );
buf ( n21581 , n21580 );
buf ( n21582 , n21581 );
nand ( n21583 , n21573 , n21582 );
buf ( n21584 , n21583 );
buf ( n21585 , n21584 );
xor ( n21586 , n21568 , n21585 );
buf ( n21587 , n19143 );
not ( n21588 , n21587 );
buf ( n21589 , n21331 );
not ( n21590 , n21589 );
or ( n21591 , n21588 , n21590 );
buf ( n21592 , n18635 );
buf ( n21593 , n588 );
nand ( n21594 , n21592 , n21593 );
buf ( n21595 , n21594 );
buf ( n21596 , n21595 );
not ( n21597 , n21596 );
buf ( n21598 , n588 );
not ( n21599 , n21598 );
buf ( n21600 , n9497 );
nand ( n21601 , n21599 , n21600 );
buf ( n21602 , n21601 );
buf ( n21603 , n21602 );
not ( n21604 , n21603 );
or ( n21605 , n21597 , n21604 );
buf ( n21606 , n19152 );
nand ( n21607 , n21605 , n21606 );
buf ( n21608 , n21607 );
buf ( n21609 , n21608 );
nand ( n21610 , n21591 , n21609 );
buf ( n21611 , n21610 );
buf ( n21612 , n21611 );
and ( n21613 , n21586 , n21612 );
and ( n21614 , n21568 , n21585 );
or ( n21615 , n21613 , n21614 );
buf ( n21616 , n21615 );
buf ( n21617 , n21616 );
and ( n21618 , n21395 , n21617 );
and ( n21619 , n21390 , n21394 );
or ( n21620 , n21618 , n21619 );
buf ( n21621 , n21620 );
buf ( n21622 , n21621 );
xor ( n21623 , n21373 , n21622 );
xor ( n21624 , n21154 , n21339 );
xor ( n21625 , n21624 , n21344 );
buf ( n21626 , n21625 );
buf ( n21627 , n21626 );
and ( n21628 , n21623 , n21627 );
and ( n21629 , n21373 , n21622 );
or ( n21630 , n21628 , n21629 );
buf ( n21631 , n21630 );
buf ( n21632 , n21631 );
nor ( n21633 , n21369 , n21632 );
buf ( n21634 , n21633 );
buf ( n21635 , n21634 );
xor ( n21636 , n21373 , n21622 );
xor ( n21637 , n21636 , n21627 );
buf ( n21638 , n21637 );
xor ( n21639 , n21179 , n21315 );
xor ( n21640 , n21639 , n21334 );
buf ( n21641 , n21640 );
buf ( n21642 , n21641 );
xor ( n21643 , n21204 , n21305 );
xor ( n21644 , n21643 , n21310 );
buf ( n21645 , n21644 );
buf ( n21646 , n21645 );
buf ( n21647 , n19244 );
not ( n21648 , n21647 );
xor ( n21649 , n590 , n10822 );
buf ( n21650 , n21649 );
not ( n21651 , n21650 );
or ( n21652 , n21648 , n21651 );
buf ( n21653 , n21382 );
buf ( n21654 , n591 );
nand ( n21655 , n21653 , n21654 );
buf ( n21656 , n21655 );
buf ( n21657 , n21656 );
nand ( n21658 , n21652 , n21657 );
buf ( n21659 , n21658 );
buf ( n21660 , n21659 );
xor ( n21661 , n21646 , n21660 );
buf ( n21662 , n18857 );
not ( n21663 , n21662 );
buf ( n21664 , n21577 );
not ( n21665 , n21664 );
or ( n21666 , n21663 , n21665 );
buf ( n21667 , n586 );
not ( n21668 , n21667 );
buf ( n21669 , n18329 );
not ( n21670 , n21669 );
or ( n21671 , n21668 , n21670 );
buf ( n21672 , n18605 );
buf ( n21673 , n18840 );
nand ( n21674 , n21672 , n21673 );
buf ( n21675 , n21674 );
buf ( n21676 , n21675 );
nand ( n21677 , n21671 , n21676 );
buf ( n21678 , n21677 );
buf ( n21679 , n21678 );
buf ( n21680 , n18881 );
nand ( n21681 , n21679 , n21680 );
buf ( n21682 , n21681 );
buf ( n21683 , n21682 );
nand ( n21684 , n21666 , n21683 );
buf ( n21685 , n21684 );
buf ( n21686 , n21685 );
buf ( n21687 , n18418 );
not ( n21688 , n21687 );
buf ( n21689 , n21258 );
not ( n21690 , n21689 );
or ( n21691 , n21688 , n21690 );
buf ( n21692 , n580 );
not ( n21693 , n21692 );
buf ( n21694 , n19972 );
not ( n21695 , n21694 );
or ( n21696 , n21693 , n21695 );
buf ( n21697 , n18402 );
buf ( n21698 , n20998 );
nand ( n21699 , n21697 , n21698 );
buf ( n21700 , n21699 );
buf ( n21701 , n21700 );
nand ( n21702 , n21696 , n21701 );
buf ( n21703 , n21702 );
buf ( n21704 , n21703 );
buf ( n21705 , n18391 );
nand ( n21706 , n21704 , n21705 );
buf ( n21707 , n21706 );
buf ( n21708 , n21707 );
nand ( n21709 , n21691 , n21708 );
buf ( n21710 , n21709 );
buf ( n21711 , n21710 );
xor ( n21712 , n21397 , n21421 );
xor ( n21713 , n21712 , n21502 );
buf ( n21714 , n21713 );
buf ( n21715 , n21714 );
xor ( n21716 , n21711 , n21715 );
buf ( n21717 , n18285 );
not ( n21718 , n21717 );
buf ( n21719 , n21520 );
not ( n21720 , n21719 );
or ( n21721 , n21718 , n21720 );
buf ( n21722 , n582 );
not ( n21723 , n21722 );
buf ( n21724 , n19531 );
not ( n21725 , n21724 );
buf ( n21726 , n21725 );
buf ( n21727 , n21726 );
not ( n21728 , n21727 );
or ( n21729 , n21723 , n21728 );
nand ( n21730 , n18303 , n4754 );
buf ( n21731 , n21730 );
nand ( n21732 , n21729 , n21731 );
buf ( n21733 , n21732 );
buf ( n21734 , n21733 );
buf ( n21735 , n18316 );
nand ( n21736 , n21734 , n21735 );
buf ( n21737 , n21736 );
buf ( n21738 , n21737 );
nand ( n21739 , n21721 , n21738 );
buf ( n21740 , n21739 );
buf ( n21741 , n21740 );
and ( n21742 , n21716 , n21741 );
and ( n21743 , n21711 , n21715 );
or ( n21744 , n21742 , n21743 );
buf ( n21745 , n21744 );
buf ( n21746 , n21745 );
buf ( n21747 , n18431 );
not ( n21748 , n21747 );
buf ( n21749 , n21550 );
not ( n21750 , n21749 );
or ( n21751 , n21748 , n21750 );
and ( n21752 , n13665 , n18277 );
not ( n21753 , n13665 );
and ( n21754 , n21753 , n584 );
or ( n21755 , n21752 , n21754 );
buf ( n21756 , n21755 );
buf ( n21757 , n18479 );
nand ( n21758 , n21756 , n21757 );
buf ( n21759 , n21758 );
buf ( n21760 , n21759 );
nand ( n21761 , n21751 , n21760 );
buf ( n21762 , n21761 );
buf ( n21763 , n21762 );
xor ( n21764 , n21746 , n21763 );
xor ( n21765 , n21506 , n21510 );
xor ( n21766 , n21765 , n21528 );
buf ( n21767 , n21766 );
buf ( n21768 , n21767 );
and ( n21769 , n21764 , n21768 );
and ( n21770 , n21746 , n21763 );
or ( n21771 , n21769 , n21770 );
buf ( n21772 , n21771 );
buf ( n21773 , n21772 );
xor ( n21774 , n21686 , n21773 );
xor ( n21775 , n21533 , n21558 );
xor ( n21776 , n21775 , n21563 );
buf ( n21777 , n21776 );
buf ( n21778 , n21777 );
and ( n21779 , n21774 , n21778 );
and ( n21780 , n21686 , n21773 );
or ( n21781 , n21779 , n21780 );
buf ( n21782 , n21781 );
buf ( n21783 , n21782 );
and ( n21784 , n21661 , n21783 );
and ( n21785 , n21646 , n21660 );
or ( n21786 , n21784 , n21785 );
buf ( n21787 , n21786 );
buf ( n21788 , n21787 );
xor ( n21789 , n21642 , n21788 );
xor ( n21790 , n21390 , n21394 );
xor ( n21791 , n21790 , n21617 );
buf ( n21792 , n21791 );
buf ( n21793 , n21792 );
and ( n21794 , n21789 , n21793 );
and ( n21795 , n21642 , n21788 );
or ( n21796 , n21794 , n21795 );
buf ( n21797 , n21796 );
nor ( n21798 , n21638 , n21797 );
buf ( n21799 , n21798 );
nor ( n21800 , n21635 , n21799 );
buf ( n21801 , n21800 );
not ( n21802 , n21801 );
xor ( n21803 , n21642 , n21788 );
xor ( n21804 , n21803 , n21793 );
buf ( n21805 , n21804 );
buf ( n21806 , n21805 );
not ( n21807 , n21806 );
buf ( n21808 , n18635 );
buf ( n21809 , n588 );
not ( n21810 , n21809 );
buf ( n21811 , n19143 );
not ( n21812 , n21811 );
buf ( n21813 , n21812 );
buf ( n21814 , n21813 );
nor ( n21815 , n21810 , n21814 );
buf ( n21816 , n21815 );
buf ( n21817 , n21816 );
nand ( n21818 , n21808 , n21817 );
buf ( n21819 , n21818 );
buf ( n21820 , n21819 );
buf ( n21821 , n18635 );
not ( n21822 , n21821 );
buf ( n21823 , n21813 );
buf ( n21824 , n588 );
nor ( n21825 , n21823 , n21824 );
buf ( n21826 , n21825 );
buf ( n21827 , n21826 );
nand ( n21828 , n21822 , n21827 );
buf ( n21829 , n21828 );
buf ( n21830 , n21829 );
and ( n21831 , n588 , n20429 );
not ( n21832 , n588 );
and ( n21833 , n21832 , n18759 );
or ( n21834 , n21831 , n21833 );
buf ( n21835 , n21834 );
buf ( n21836 , n19152 );
nand ( n21837 , n21835 , n21836 );
buf ( n21838 , n21837 );
buf ( n21839 , n21838 );
nand ( n21840 , n21820 , n21830 , n21839 );
buf ( n21841 , n21840 );
buf ( n21842 , n21841 );
buf ( n21843 , n18857 );
not ( n21844 , n21843 );
buf ( n21845 , n21678 );
not ( n21846 , n21845 );
or ( n21847 , n21844 , n21846 );
buf ( n21848 , n586 );
not ( n21849 , n21848 );
buf ( n21850 , n19022 );
not ( n21851 , n21850 );
or ( n21852 , n21849 , n21851 );
buf ( n21853 , n18489 );
buf ( n21854 , n18840 );
nand ( n21855 , n21853 , n21854 );
buf ( n21856 , n21855 );
buf ( n21857 , n21856 );
nand ( n21858 , n21852 , n21857 );
buf ( n21859 , n21858 );
buf ( n21860 , n21859 );
buf ( n21861 , n18881 );
nand ( n21862 , n21860 , n21861 );
buf ( n21863 , n21862 );
buf ( n21864 , n21863 );
nand ( n21865 , n21847 , n21864 );
buf ( n21866 , n21865 );
buf ( n21867 , n21866 );
buf ( n21868 , n18418 );
not ( n21869 , n21868 );
buf ( n21870 , n21703 );
not ( n21871 , n21870 );
or ( n21872 , n21869 , n21871 );
buf ( n21873 , n580 );
not ( n21874 , n21873 );
buf ( n21875 , n21220 );
not ( n21876 , n21875 );
or ( n21877 , n21874 , n21876 );
buf ( n21878 , n18402 );
buf ( n21879 , n13666 );
nand ( n21880 , n21878 , n21879 );
buf ( n21881 , n21880 );
buf ( n21882 , n21881 );
nand ( n21883 , n21877 , n21882 );
buf ( n21884 , n21883 );
buf ( n21885 , n21884 );
buf ( n21886 , n18391 );
nand ( n21887 , n21885 , n21886 );
buf ( n21888 , n21887 );
buf ( n21889 , n21888 );
nand ( n21890 , n21872 , n21889 );
buf ( n21891 , n21890 );
buf ( n21892 , n21891 );
xor ( n21893 , n21424 , n21437 );
xor ( n21894 , n21893 , n21498 );
buf ( n21895 , n21894 );
buf ( n21896 , n21895 );
xor ( n21897 , n21892 , n21896 );
buf ( n21898 , n18285 );
not ( n21899 , n21898 );
buf ( n21900 , n21733 );
not ( n21901 , n21900 );
or ( n21902 , n21899 , n21901 );
buf ( n21903 , n582 );
not ( n21904 , n21903 );
buf ( n21905 , n13664 );
not ( n21906 , n21905 );
buf ( n21907 , n21906 );
buf ( n21908 , n21907 );
not ( n21909 , n21908 );
or ( n21910 , n21904 , n21909 );
buf ( n21911 , n13664 );
buf ( n21912 , n18303 );
nand ( n21913 , n21911 , n21912 );
buf ( n21914 , n21913 );
buf ( n21915 , n21914 );
nand ( n21916 , n21910 , n21915 );
buf ( n21917 , n21916 );
buf ( n21918 , n21917 );
buf ( n21919 , n18316 );
nand ( n21920 , n21918 , n21919 );
buf ( n21921 , n21920 );
buf ( n21922 , n21921 );
nand ( n21923 , n21902 , n21922 );
buf ( n21924 , n21923 );
buf ( n21925 , n21924 );
and ( n21926 , n21897 , n21925 );
and ( n21927 , n21892 , n21896 );
or ( n21928 , n21926 , n21927 );
buf ( n21929 , n21928 );
buf ( n21930 , n21929 );
nand ( n21931 , n18431 , n21755 );
and ( n21932 , n18997 , n18277 );
not ( n21933 , n18997 );
and ( n21934 , n21933 , n584 );
or ( n21935 , n21932 , n21934 );
buf ( n21936 , n21935 );
buf ( n21937 , n18479 );
nand ( n21938 , n21936 , n21937 );
buf ( n21939 , n21938 );
nand ( n21940 , n21931 , n21939 );
buf ( n21941 , n21940 );
xor ( n21942 , n21930 , n21941 );
xor ( n21943 , n21711 , n21715 );
xor ( n21944 , n21943 , n21741 );
buf ( n21945 , n21944 );
buf ( n21946 , n21945 );
and ( n21947 , n21942 , n21946 );
and ( n21948 , n21930 , n21941 );
or ( n21949 , n21947 , n21948 );
buf ( n21950 , n21949 );
buf ( n21951 , n21950 );
xor ( n21952 , n21867 , n21951 );
xor ( n21953 , n21746 , n21763 );
xor ( n21954 , n21953 , n21768 );
buf ( n21955 , n21954 );
buf ( n21956 , n21955 );
and ( n21957 , n21952 , n21956 );
and ( n21958 , n21867 , n21951 );
or ( n21959 , n21957 , n21958 );
buf ( n21960 , n21959 );
buf ( n21961 , n21960 );
xor ( n21962 , n21842 , n21961 );
buf ( n21963 , n19244 );
not ( n21964 , n21963 );
and ( n21965 , n590 , n18894 );
not ( n21966 , n590 );
and ( n21967 , n21966 , n10854 );
or ( n21968 , n21965 , n21967 );
buf ( n21969 , n21968 );
not ( n21970 , n21969 );
or ( n21971 , n21964 , n21970 );
buf ( n21972 , n21649 );
buf ( n21973 , n591 );
nand ( n21974 , n21972 , n21973 );
buf ( n21975 , n21974 );
buf ( n21976 , n21975 );
nand ( n21977 , n21971 , n21976 );
buf ( n21978 , n21977 );
buf ( n21979 , n21978 );
and ( n21980 , n21962 , n21979 );
and ( n21981 , n21842 , n21961 );
or ( n21982 , n21980 , n21981 );
buf ( n21983 , n21982 );
buf ( n21984 , n21983 );
xor ( n21985 , n21568 , n21585 );
xor ( n21986 , n21985 , n21612 );
buf ( n21987 , n21986 );
buf ( n21988 , n21987 );
xor ( n21989 , n21984 , n21988 );
xor ( n21990 , n21646 , n21660 );
xor ( n21991 , n21990 , n21783 );
buf ( n21992 , n21991 );
buf ( n21993 , n21992 );
and ( n21994 , n21989 , n21993 );
and ( n21995 , n21984 , n21988 );
or ( n21996 , n21994 , n21995 );
buf ( n21997 , n21996 );
buf ( n21998 , n21997 );
not ( n21999 , n21998 );
buf ( n22000 , n21999 );
buf ( n22001 , n22000 );
nand ( n22002 , n21807 , n22001 );
buf ( n22003 , n22002 );
xor ( n22004 , n21686 , n21773 );
xor ( n22005 , n22004 , n21778 );
buf ( n22006 , n22005 );
buf ( n22007 , n22006 );
buf ( n22008 , C0 );
buf ( n22009 , n22008 );
buf ( n22010 , n18418 );
not ( n22011 , n22010 );
buf ( n22012 , n21884 );
not ( n22013 , n22012 );
or ( n22014 , n22011 , n22013 );
and ( n22015 , n20449 , n18402 );
not ( n22016 , n20449 );
and ( n22017 , n22016 , n580 );
or ( n22018 , n22015 , n22017 );
buf ( n22019 , n22018 );
buf ( n22020 , n18391 );
nand ( n22021 , n22019 , n22020 );
buf ( n22022 , n22021 );
buf ( n22023 , n22022 );
nand ( n22024 , n22014 , n22023 );
buf ( n22025 , n22024 );
buf ( n22026 , n22025 );
xor ( n22027 , n22009 , n22026 );
buf ( n22028 , C0 );
buf ( n22029 , n22028 );
buf ( n22030 , n18380 );
not ( n22031 , n22030 );
buf ( n22032 , n22018 );
not ( n22033 , n22032 );
or ( n22034 , n22031 , n22033 );
buf ( n22035 , n580 );
not ( n22036 , n22035 );
or ( n22037 , n22036 , C0 );
buf ( n22038 , C1 );
buf ( n22039 , n22038 );
nand ( n22040 , n22037 , n22039 );
buf ( n22041 , n22040 );
buf ( n22042 , n22041 );
buf ( n22043 , n18391 );
nand ( n22044 , n22042 , n22043 );
buf ( n22045 , n22044 );
buf ( n22046 , n22045 );
nand ( n22047 , n22034 , n22046 );
buf ( n22048 , n22047 );
buf ( n22049 , n22048 );
xor ( n22050 , n22029 , n22049 );
buf ( n22051 , C0 );
buf ( n22052 , n22051 );
buf ( n22053 , n18380 );
not ( n22054 , n22053 );
buf ( n22055 , n22041 );
not ( n22056 , n22055 );
or ( n22057 , n22054 , n22056 );
buf ( n22058 , n580 );
not ( n22059 , n22058 );
or ( n22060 , n22059 , C0 );
buf ( n22061 , C1 );
buf ( n22062 , n22061 );
nand ( n22063 , n22060 , n22062 );
buf ( n22064 , n22063 );
buf ( n22065 , n22064 );
buf ( n22066 , n18391 );
nand ( n22067 , n22065 , n22066 );
buf ( n22068 , n22067 );
buf ( n22069 , n22068 );
nand ( n22070 , n22057 , n22069 );
buf ( n22071 , n22070 );
buf ( n22072 , n22071 );
xor ( n22073 , n22052 , n22072 );
buf ( n22074 , n18380 );
not ( n22075 , n22074 );
buf ( n22076 , n22064 );
not ( n22077 , n22076 );
or ( n22078 , n22075 , n22077 );
buf ( n22079 , C0 );
buf ( n22080 , n18402 );
or ( n22081 , n22079 , n22080 );
nand ( n22082 , n22081 , C1 );
buf ( n22083 , n22082 );
buf ( n22084 , n22083 );
buf ( n22085 , n18388 );
nand ( n22086 , n22084 , n22085 );
buf ( n22087 , n22086 );
buf ( n22088 , n22087 );
nand ( n22089 , n22078 , n22088 );
buf ( n22090 , n22089 );
buf ( n22091 , n22090 );
not ( n22092 , n22091 );
buf ( n22093 , C1 );
buf ( n22094 , n22093 );
buf ( n22095 , n581 );
buf ( n22096 , n582 );
nand ( n22097 , n22095 , n22096 );
buf ( n22098 , n22097 );
buf ( n22099 , n22098 );
buf ( n22100 , n580 );
nand ( n22101 , n22094 , n22099 , n22100 );
buf ( n22102 , n22101 );
buf ( n22103 , n22102 );
nor ( n22104 , n22092 , n22103 );
buf ( n22105 , n22104 );
buf ( n22106 , n22105 );
and ( n22107 , n22073 , n22106 );
or ( n22108 , n22107 , C0 );
buf ( n22109 , n22108 );
buf ( n22110 , n22109 );
and ( n22111 , n22050 , n22110 );
or ( n22112 , n22111 , C0 );
buf ( n22113 , n22112 );
buf ( n22114 , n22113 );
and ( n22115 , n22027 , n22114 );
or ( n22116 , n22115 , C0 );
buf ( n22117 , n22116 );
buf ( n22118 , n22117 );
xor ( n22119 , n21892 , n21896 );
xor ( n22120 , n22119 , n21925 );
buf ( n22121 , n22120 );
buf ( n22122 , n22121 );
xor ( n22123 , n22118 , n22122 );
buf ( n22124 , n18431 );
not ( n22125 , n22124 );
buf ( n22126 , n21935 );
not ( n22127 , n22126 );
or ( n22128 , n22125 , n22127 );
buf ( n22129 , n584 );
not ( n22130 , n22129 );
buf ( n22131 , n18981 );
not ( n22132 , n22131 );
or ( n22133 , n22130 , n22132 );
buf ( n22134 , n18277 );
buf ( n22135 , n13663 );
nand ( n22136 , n22134 , n22135 );
buf ( n22137 , n22136 );
buf ( n22138 , n22137 );
nand ( n22139 , n22133 , n22138 );
buf ( n22140 , n22139 );
buf ( n22141 , n22140 );
buf ( n22142 , n18479 );
nand ( n22143 , n22141 , n22142 );
buf ( n22144 , n22143 );
buf ( n22145 , n22144 );
nand ( n22146 , n22128 , n22145 );
buf ( n22147 , n22146 );
buf ( n22148 , n22147 );
and ( n22149 , n22123 , n22148 );
and ( n22150 , n22118 , n22122 );
or ( n22151 , n22149 , n22150 );
buf ( n22152 , n22151 );
buf ( n22153 , n22152 );
xor ( n22154 , n21930 , n21941 );
xor ( n22155 , n22154 , n21946 );
buf ( n22156 , n22155 );
buf ( n22157 , n22156 );
xor ( n22158 , n22153 , n22157 );
buf ( n22159 , n18857 );
not ( n22160 , n22159 );
buf ( n22161 , n21859 );
not ( n22162 , n22161 );
or ( n22163 , n22160 , n22162 );
buf ( n22164 , n586 );
buf ( n22165 , n18566 );
and ( n22166 , n22164 , n22165 );
not ( n22167 , n22164 );
buf ( n22168 , n18569 );
and ( n22169 , n22167 , n22168 );
nor ( n22170 , n22166 , n22169 );
buf ( n22171 , n22170 );
buf ( n22172 , n22171 );
buf ( n22173 , n18881 );
nand ( n22174 , n22172 , n22173 );
buf ( n22175 , n22174 );
buf ( n22176 , n22175 );
nand ( n22177 , n22163 , n22176 );
buf ( n22178 , n22177 );
buf ( n22179 , n22178 );
and ( n22180 , n22158 , n22179 );
and ( n22181 , n22153 , n22157 );
or ( n22182 , n22180 , n22181 );
buf ( n22183 , n22182 );
buf ( n22184 , n22183 );
buf ( n22185 , n19143 );
not ( n22186 , n22185 );
buf ( n22187 , n21834 );
not ( n22188 , n22187 );
or ( n22189 , n22186 , n22188 );
xnor ( n22190 , n588 , n18960 );
buf ( n22191 , n22190 );
buf ( n22192 , n19152 );
nand ( n22193 , n22191 , n22192 );
buf ( n22194 , n22193 );
buf ( n22195 , n22194 );
nand ( n22196 , n22189 , n22195 );
buf ( n22197 , n22196 );
buf ( n22198 , n22197 );
xor ( n22199 , n22184 , n22198 );
buf ( n22200 , n19244 );
not ( n22201 , n22200 );
and ( n22202 , n590 , n18635 );
not ( n22203 , n590 );
and ( n22204 , n22203 , n9497 );
or ( n22205 , n22202 , n22204 );
buf ( n22206 , n22205 );
not ( n22207 , n22206 );
or ( n22208 , n22201 , n22207 );
buf ( n22209 , n21968 );
buf ( n22210 , n591 );
nand ( n22211 , n22209 , n22210 );
buf ( n22212 , n22211 );
buf ( n22213 , n22212 );
nand ( n22214 , n22208 , n22213 );
buf ( n22215 , n22214 );
buf ( n22216 , n22215 );
and ( n22217 , n22199 , n22216 );
and ( n22218 , n22184 , n22198 );
or ( n22219 , n22217 , n22218 );
buf ( n22220 , n22219 );
buf ( n22221 , n22220 );
xor ( n22222 , n22007 , n22221 );
xor ( n22223 , n21842 , n21961 );
xor ( n22224 , n22223 , n21979 );
buf ( n22225 , n22224 );
buf ( n22226 , n22225 );
xor ( n22227 , n22222 , n22226 );
buf ( n22228 , n22227 );
not ( n22229 , n22228 );
xor ( n22230 , n21867 , n21951 );
xor ( n22231 , n22230 , n21956 );
buf ( n22232 , n22231 );
buf ( n22233 , n22232 );
buf ( n22234 , n19143 );
not ( n22235 , n22234 );
buf ( n22236 , n22190 );
not ( n22237 , n22236 );
or ( n22238 , n22235 , n22237 );
and ( n22239 , n588 , n18599 );
not ( n22240 , n588 );
and ( n22241 , n22240 , n18326 );
or ( n22242 , n22239 , n22241 );
buf ( n22243 , n22242 );
buf ( n22244 , n19152 );
nand ( n22245 , n22243 , n22244 );
buf ( n22246 , n22245 );
buf ( n22247 , n22246 );
nand ( n22248 , n22238 , n22247 );
buf ( n22249 , n22248 );
buf ( n22250 , n22249 );
buf ( n22251 , n18285 );
not ( n22252 , n22251 );
buf ( n22253 , n21917 );
not ( n22254 , n22253 );
or ( n22255 , n22252 , n22254 );
buf ( n22256 , n582 );
not ( n22257 , n22256 );
buf ( n22258 , n20998 );
not ( n22259 , n22258 );
buf ( n22260 , n22259 );
buf ( n22261 , n22260 );
not ( n22262 , n22261 );
or ( n22263 , n22257 , n22262 );
buf ( n22264 , n19975 );
buf ( n22265 , n18303 );
nand ( n22266 , n22264 , n22265 );
buf ( n22267 , n22266 );
buf ( n22268 , n22267 );
nand ( n22269 , n22263 , n22268 );
buf ( n22270 , n22269 );
buf ( n22271 , n22270 );
buf ( n22272 , n18316 );
nand ( n22273 , n22271 , n22272 );
buf ( n22274 , n22273 );
buf ( n22275 , n22274 );
nand ( n22276 , n22255 , n22275 );
buf ( n22277 , n22276 );
buf ( n22278 , n22277 );
xor ( n22279 , n22009 , n22026 );
xor ( n22280 , n22279 , n22114 );
buf ( n22281 , n22280 );
buf ( n22282 , n22281 );
xor ( n22283 , n22278 , n22282 );
buf ( n22284 , n18431 );
not ( n22285 , n22284 );
buf ( n22286 , n22140 );
not ( n22287 , n22286 );
or ( n22288 , n22285 , n22287 );
buf ( n22289 , n584 );
not ( n22290 , n22289 );
buf ( n22291 , n19651 );
not ( n22292 , n22291 );
or ( n22293 , n22290 , n22292 );
buf ( n22294 , n19534 );
buf ( n22295 , n18277 );
nand ( n22296 , n22294 , n22295 );
buf ( n22297 , n22296 );
buf ( n22298 , n22297 );
nand ( n22299 , n22293 , n22298 );
buf ( n22300 , n22299 );
buf ( n22301 , n22300 );
buf ( n22302 , n18479 );
nand ( n22303 , n22301 , n22302 );
buf ( n22304 , n22303 );
buf ( n22305 , n22304 );
nand ( n22306 , n22288 , n22305 );
buf ( n22307 , n22306 );
buf ( n22308 , n22307 );
and ( n22309 , n22283 , n22308 );
and ( n22310 , n22278 , n22282 );
or ( n22311 , n22309 , n22310 );
buf ( n22312 , n22311 );
buf ( n22313 , n22312 );
buf ( n22314 , n18857 );
not ( n22315 , n22314 );
buf ( n22316 , n22171 );
not ( n22317 , n22316 );
or ( n22318 , n22315 , n22317 );
and ( n22319 , n13665 , n18840 );
not ( n22320 , n13665 );
and ( n22321 , n22320 , n586 );
or ( n22322 , n22319 , n22321 );
buf ( n22323 , n22322 );
buf ( n22324 , n18881 );
nand ( n22325 , n22323 , n22324 );
buf ( n22326 , n22325 );
buf ( n22327 , n22326 );
nand ( n22328 , n22318 , n22327 );
buf ( n22329 , n22328 );
buf ( n22330 , n22329 );
xor ( n22331 , n22313 , n22330 );
xor ( n22332 , n22118 , n22122 );
xor ( n22333 , n22332 , n22148 );
buf ( n22334 , n22333 );
buf ( n22335 , n22334 );
and ( n22336 , n22331 , n22335 );
and ( n22337 , n22313 , n22330 );
or ( n22338 , n22336 , n22337 );
buf ( n22339 , n22338 );
buf ( n22340 , n22339 );
xor ( n22341 , n22250 , n22340 );
xor ( n22342 , n22153 , n22157 );
xor ( n22343 , n22342 , n22179 );
buf ( n22344 , n22343 );
buf ( n22345 , n22344 );
and ( n22346 , n22341 , n22345 );
and ( n22347 , n22250 , n22340 );
or ( n22348 , n22346 , n22347 );
buf ( n22349 , n22348 );
buf ( n22350 , n22349 );
xor ( n22351 , n22233 , n22350 );
xor ( n22352 , n22184 , n22198 );
xor ( n22353 , n22352 , n22216 );
buf ( n22354 , n22353 );
buf ( n22355 , n22354 );
and ( n22356 , n22351 , n22355 );
and ( n22357 , n22233 , n22350 );
or ( n22358 , n22356 , n22357 );
buf ( n22359 , n22358 );
not ( n22360 , n22359 );
and ( n22361 , n22229 , n22360 );
xor ( n22362 , n21984 , n21988 );
xor ( n22363 , n22362 , n21993 );
buf ( n22364 , n22363 );
buf ( n22365 , n22364 );
xor ( n22366 , n22007 , n22221 );
and ( n22367 , n22366 , n22226 );
and ( n22368 , n22007 , n22221 );
or ( n22369 , n22367 , n22368 );
buf ( n22370 , n22369 );
buf ( n22371 , n22370 );
nor ( n22372 , n22365 , n22371 );
buf ( n22373 , n22372 );
nor ( n22374 , n22361 , n22373 );
xor ( n22375 , n22233 , n22350 );
xor ( n22376 , n22375 , n22355 );
buf ( n22377 , n22376 );
buf ( n22378 , n22377 );
not ( n22379 , n22378 );
buf ( n22380 , n591 );
not ( n22381 , n22380 );
buf ( n22382 , n22205 );
not ( n22383 , n22382 );
or ( n22384 , n22381 , n22383 );
and ( n22385 , n590 , n20429 );
not ( n22386 , n590 );
and ( n22387 , n22386 , n18344 );
or ( n22388 , n22385 , n22387 );
buf ( n22389 , n22388 );
buf ( n22390 , n19244 );
nand ( n22391 , n22389 , n22390 );
buf ( n22392 , n22391 );
buf ( n22393 , n22392 );
nand ( n22394 , n22384 , n22393 );
buf ( n22395 , n22394 );
buf ( n22396 , n22395 );
buf ( n22397 , n19143 );
not ( n22398 , n22397 );
buf ( n22399 , n22242 );
not ( n22400 , n22399 );
or ( n22401 , n22398 , n22400 );
and ( n22402 , n588 , n18492 );
not ( n22403 , n588 );
and ( n22404 , n22403 , n18489 );
or ( n22405 , n22402 , n22404 );
buf ( n22406 , n22405 );
buf ( n22407 , n19152 );
nand ( n22408 , n22406 , n22407 );
buf ( n22409 , n22408 );
buf ( n22410 , n22409 );
nand ( n22411 , n22401 , n22410 );
buf ( n22412 , n22411 );
buf ( n22413 , n22412 );
buf ( n22414 , n18285 );
not ( n22415 , n22414 );
buf ( n22416 , n22270 );
not ( n22417 , n22416 );
or ( n22418 , n22415 , n22417 );
buf ( n22419 , n582 );
not ( n22420 , n22419 );
buf ( n22421 , n21214 );
not ( n22422 , n22421 );
or ( n22423 , n22420 , n22422 );
buf ( n22424 , n13666 );
buf ( n22425 , n18303 );
nand ( n22426 , n22424 , n22425 );
buf ( n22427 , n22426 );
buf ( n22428 , n22427 );
nand ( n22429 , n22423 , n22428 );
buf ( n22430 , n22429 );
buf ( n22431 , n22430 );
buf ( n22432 , n18316 );
nand ( n22433 , n22431 , n22432 );
buf ( n22434 , n22433 );
buf ( n22435 , n22434 );
nand ( n22436 , n22418 , n22435 );
buf ( n22437 , n22436 );
buf ( n22438 , n22437 );
xor ( n22439 , n22029 , n22049 );
xor ( n22440 , n22439 , n22110 );
buf ( n22441 , n22440 );
buf ( n22442 , n22441 );
xor ( n22443 , n22438 , n22442 );
buf ( n22444 , C0 );
buf ( n22445 , n22444 );
buf ( n22446 , n18285 );
not ( n22447 , n22446 );
buf ( n22448 , n22430 );
not ( n22449 , n22448 );
or ( n22450 , n22447 , n22449 );
and ( n22451 , n20449 , n18303 );
not ( n22452 , n20449 );
and ( n22453 , n22452 , n582 );
or ( n22454 , n22451 , n22453 );
buf ( n22455 , n22454 );
buf ( n22456 , n18316 );
nand ( n22457 , n22455 , n22456 );
buf ( n22458 , n22457 );
buf ( n22459 , n22458 );
nand ( n22460 , n22450 , n22459 );
buf ( n22461 , n22460 );
buf ( n22462 , n22461 );
xor ( n22463 , n22445 , n22462 );
buf ( n22464 , C0 );
buf ( n22465 , n22464 );
buf ( n22466 , n18285 );
not ( n22467 , n22466 );
buf ( n22468 , n22454 );
not ( n22469 , n22468 );
or ( n22470 , n22467 , n22469 );
buf ( n22471 , n582 );
not ( n22472 , n22471 );
or ( n22473 , n22472 , C0 );
buf ( n22474 , C1 );
buf ( n22475 , n22474 );
nand ( n22476 , n22473 , n22475 );
buf ( n22477 , n22476 );
buf ( n22478 , n22477 );
buf ( n22479 , n18316 );
nand ( n22480 , n22478 , n22479 );
buf ( n22481 , n22480 );
buf ( n22482 , n22481 );
nand ( n22483 , n22470 , n22482 );
buf ( n22484 , n22483 );
buf ( n22485 , n22484 );
xor ( n22486 , n22465 , n22485 );
buf ( n22487 , C0 );
buf ( n22488 , n22487 );
buf ( n22489 , n18285 );
not ( n22490 , n22489 );
buf ( n22491 , n22477 );
not ( n22492 , n22491 );
or ( n22493 , n22490 , n22492 );
buf ( n22494 , n582 );
not ( n22495 , n22494 );
or ( n22496 , n22495 , C0 );
buf ( n22497 , C1 );
buf ( n22498 , n22497 );
nand ( n22499 , n22496 , n22498 );
buf ( n22500 , n22499 );
buf ( n22501 , n22500 );
buf ( n22502 , n18316 );
nand ( n22503 , n22501 , n22502 );
buf ( n22504 , n22503 );
buf ( n22505 , n22504 );
nand ( n22506 , n22493 , n22505 );
buf ( n22507 , n22506 );
buf ( n22508 , n22507 );
xor ( n22509 , n22488 , n22508 );
buf ( n22510 , n18285 );
not ( n22511 , n22510 );
buf ( n22512 , n22500 );
not ( n22513 , n22512 );
or ( n22514 , n22511 , n22513 );
buf ( n22515 , C0 );
buf ( n22516 , n18303 );
or ( n22517 , n22515 , n22516 );
nand ( n22518 , n22517 , C1 );
buf ( n22519 , n22518 );
buf ( n22520 , n22519 );
buf ( n22521 , n18316 );
nand ( n22522 , n22520 , n22521 );
buf ( n22523 , n22522 );
buf ( n22524 , n22523 );
nand ( n22525 , n22514 , n22524 );
buf ( n22526 , n22525 );
buf ( n22527 , n22526 );
not ( n22528 , n22527 );
buf ( n22529 , C1 );
buf ( n22530 , n22529 );
buf ( n22531 , n583 );
buf ( n22532 , n584 );
and ( n22533 , n22531 , n22532 );
buf ( n22534 , n18303 );
nor ( n22535 , n22533 , n22534 );
buf ( n22536 , n22535 );
buf ( n22537 , n22536 );
and ( n22538 , n22530 , n22537 );
buf ( n22539 , n22538 );
buf ( n22540 , n22539 );
not ( n22541 , n22540 );
buf ( n22542 , n22541 );
buf ( n22543 , n22542 );
nor ( n22544 , n22528 , n22543 );
buf ( n22545 , n22544 );
buf ( n22546 , n22545 );
and ( n22547 , n22509 , n22546 );
or ( n22548 , n22547 , C0 );
buf ( n22549 , n22548 );
buf ( n22550 , n22549 );
and ( n22551 , n22486 , n22550 );
or ( n22552 , n22551 , C0 );
buf ( n22553 , n22552 );
buf ( n22554 , n22553 );
and ( n22555 , n22463 , n22554 );
or ( n22556 , n22555 , C0 );
buf ( n22557 , n22556 );
buf ( n22558 , n22557 );
and ( n22559 , n22443 , n22558 );
or ( n22560 , n22559 , C0 );
buf ( n22561 , n22560 );
buf ( n22562 , n22561 );
buf ( n22563 , n18857 );
not ( n22564 , n22563 );
buf ( n22565 , n22322 );
not ( n22566 , n22565 );
or ( n22567 , n22564 , n22566 );
buf ( n22568 , n586 );
not ( n22569 , n22568 );
buf ( n22570 , n19000 );
not ( n22571 , n22570 );
or ( n22572 , n22569 , n22571 );
buf ( n22573 , n18997 );
buf ( n22574 , n18840 );
nand ( n22575 , n22573 , n22574 );
buf ( n22576 , n22575 );
buf ( n22577 , n22576 );
nand ( n22578 , n22572 , n22577 );
buf ( n22579 , n22578 );
buf ( n22580 , n22579 );
buf ( n22581 , n18881 );
nand ( n22582 , n22580 , n22581 );
buf ( n22583 , n22582 );
buf ( n22584 , n22583 );
nand ( n22585 , n22567 , n22584 );
buf ( n22586 , n22585 );
buf ( n22587 , n22586 );
xor ( n22588 , n22562 , n22587 );
xor ( n22589 , n22278 , n22282 );
xor ( n22590 , n22589 , n22308 );
buf ( n22591 , n22590 );
buf ( n22592 , n22591 );
and ( n22593 , n22588 , n22592 );
and ( n22594 , n22562 , n22587 );
or ( n22595 , n22593 , n22594 );
buf ( n22596 , n22595 );
buf ( n22597 , n22596 );
xor ( n22598 , n22413 , n22597 );
xor ( n22599 , n22313 , n22330 );
xor ( n22600 , n22599 , n22335 );
buf ( n22601 , n22600 );
buf ( n22602 , n22601 );
and ( n22603 , n22598 , n22602 );
and ( n22604 , n22413 , n22597 );
or ( n22605 , n22603 , n22604 );
buf ( n22606 , n22605 );
buf ( n22607 , n22606 );
xor ( n22608 , n22396 , n22607 );
xor ( n22609 , n22250 , n22340 );
xor ( n22610 , n22609 , n22345 );
buf ( n22611 , n22610 );
buf ( n22612 , n22611 );
and ( n22613 , n22608 , n22612 );
and ( n22614 , n22396 , n22607 );
or ( n22615 , n22613 , n22614 );
buf ( n22616 , n22615 );
buf ( n22617 , n22616 );
not ( n22618 , n22617 );
buf ( n22619 , n22618 );
buf ( n22620 , n22619 );
nand ( n22621 , n22379 , n22620 );
buf ( n22622 , n22621 );
buf ( n22623 , n22622 );
not ( n22624 , n22623 );
buf ( n22625 , n591 );
not ( n22626 , n22625 );
and ( n22627 , n590 , n18960 );
not ( n22628 , n590 );
and ( n22629 , n22628 , n18357 );
or ( n22630 , n22627 , n22629 );
buf ( n22631 , n22630 );
not ( n22632 , n22631 );
or ( n22633 , n22626 , n22632 );
and ( n22634 , n590 , n18329 );
not ( n22635 , n590 );
and ( n22636 , n22635 , n18332 );
or ( n22637 , n22634 , n22636 );
buf ( n22638 , n22637 );
buf ( n22639 , n19244 );
nand ( n22640 , n22638 , n22639 );
buf ( n22641 , n22640 );
buf ( n22642 , n22641 );
nand ( n22643 , n22633 , n22642 );
buf ( n22644 , n22643 );
buf ( n22645 , n22644 );
buf ( n22646 , n18431 );
not ( n22647 , n22646 );
and ( n22648 , n20483 , n584 );
not ( n22649 , n20483 );
and ( n22650 , n22649 , n18277 );
or ( n22651 , n22648 , n22650 );
buf ( n22652 , n22651 );
not ( n22653 , n22652 );
or ( n22654 , n22647 , n22653 );
buf ( n22655 , n584 );
not ( n22656 , n22655 );
buf ( n22657 , n19972 );
not ( n22658 , n22657 );
or ( n22659 , n22656 , n22658 );
buf ( n22660 , n18277 );
buf ( n22661 , n20998 );
nand ( n22662 , n22660 , n22661 );
buf ( n22663 , n22662 );
buf ( n22664 , n22663 );
nand ( n22665 , n22659 , n22664 );
buf ( n22666 , n22665 );
buf ( n22667 , n22666 );
buf ( n22668 , n18479 );
nand ( n22669 , n22667 , n22668 );
buf ( n22670 , n22669 );
buf ( n22671 , n22670 );
nand ( n22672 , n22654 , n22671 );
buf ( n22673 , n22672 );
buf ( n22674 , n22673 );
xor ( n22675 , n22445 , n22462 );
xor ( n22676 , n22675 , n22554 );
buf ( n22677 , n22676 );
buf ( n22678 , n22677 );
xor ( n22679 , n22674 , n22678 );
buf ( n22680 , n18857 );
not ( n22681 , n22680 );
buf ( n22682 , n586 );
not ( n22683 , n22682 );
buf ( n22684 , n19549 );
not ( n22685 , n22684 );
or ( n22686 , n22683 , n22685 );
buf ( n22687 , n18840 );
buf ( n22688 , n13663 );
nand ( n22689 , n22687 , n22688 );
buf ( n22690 , n22689 );
buf ( n22691 , n22690 );
nand ( n22692 , n22686 , n22691 );
buf ( n22693 , n22692 );
buf ( n22694 , n22693 );
not ( n22695 , n22694 );
or ( n22696 , n22681 , n22695 );
buf ( n22697 , n586 );
not ( n22698 , n22697 );
buf ( n22699 , n21726 );
not ( n22700 , n22699 );
or ( n22701 , n22698 , n22700 );
buf ( n22702 , n21726 );
not ( n22703 , n22702 );
buf ( n22704 , n22703 );
buf ( n22705 , n22704 );
buf ( n22706 , n18840 );
nand ( n22707 , n22705 , n22706 );
buf ( n22708 , n22707 );
buf ( n22709 , n22708 );
nand ( n22710 , n22701 , n22709 );
buf ( n22711 , n22710 );
buf ( n22712 , n22711 );
buf ( n22713 , n18881 );
nand ( n22714 , n22712 , n22713 );
buf ( n22715 , n22714 );
buf ( n22716 , n22715 );
nand ( n22717 , n22696 , n22716 );
buf ( n22718 , n22717 );
buf ( n22719 , n22718 );
and ( n22720 , n22679 , n22719 );
and ( n22721 , n22674 , n22678 );
or ( n22722 , n22720 , n22721 );
buf ( n22723 , n22722 );
buf ( n22724 , n22723 );
buf ( n22725 , n19143 );
not ( n22726 , n22725 );
buf ( n22727 , n588 );
not ( n22728 , n22727 );
buf ( n22729 , n18569 );
not ( n22730 , n22729 );
or ( n22731 , n22728 , n22730 );
buf ( n22732 , n588 );
not ( n22733 , n22732 );
buf ( n22734 , n18566 );
nand ( n22735 , n22733 , n22734 );
buf ( n22736 , n22735 );
buf ( n22737 , n22736 );
nand ( n22738 , n22731 , n22737 );
buf ( n22739 , n22738 );
buf ( n22740 , n22739 );
not ( n22741 , n22740 );
or ( n22742 , n22726 , n22741 );
not ( n22743 , n18538 );
not ( n22744 , n588 );
or ( n22745 , n22743 , n22744 );
not ( n22746 , n588 );
nand ( n22747 , n22746 , n13665 );
nand ( n22748 , n22745 , n22747 );
nand ( n22749 , n22748 , n19152 );
buf ( n22750 , n22749 );
nand ( n22751 , n22742 , n22750 );
buf ( n22752 , n22751 );
buf ( n22753 , n22752 );
xor ( n22754 , n22724 , n22753 );
buf ( n22755 , n18431 );
not ( n22756 , n22755 );
buf ( n22757 , n22300 );
not ( n22758 , n22757 );
or ( n22759 , n22756 , n22758 );
buf ( n22760 , n22651 );
buf ( n22761 , n18479 );
nand ( n22762 , n22760 , n22761 );
buf ( n22763 , n22762 );
buf ( n22764 , n22763 );
nand ( n22765 , n22759 , n22764 );
buf ( n22766 , n22765 );
buf ( n22767 , n22766 );
xor ( n22768 , n22438 , n22442 );
xor ( n22769 , n22768 , n22558 );
buf ( n22770 , n22769 );
buf ( n22771 , n22770 );
xor ( n22772 , n22767 , n22771 );
buf ( n22773 , n18857 );
not ( n22774 , n22773 );
buf ( n22775 , n22579 );
not ( n22776 , n22775 );
or ( n22777 , n22774 , n22776 );
buf ( n22778 , n22693 );
buf ( n22779 , n18881 );
nand ( n22780 , n22778 , n22779 );
buf ( n22781 , n22780 );
buf ( n22782 , n22781 );
nand ( n22783 , n22777 , n22782 );
buf ( n22784 , n22783 );
buf ( n22785 , n22784 );
xor ( n22786 , n22772 , n22785 );
buf ( n22787 , n22786 );
buf ( n22788 , n22787 );
and ( n22789 , n22754 , n22788 );
and ( n22790 , n22724 , n22753 );
or ( n22791 , n22789 , n22790 );
buf ( n22792 , n22791 );
buf ( n22793 , n22792 );
xor ( n22794 , n22645 , n22793 );
xor ( n22795 , n22767 , n22771 );
and ( n22796 , n22795 , n22785 );
and ( n22797 , n22767 , n22771 );
or ( n22798 , n22796 , n22797 );
buf ( n22799 , n22798 );
buf ( n22800 , n22799 );
xor ( n22801 , n22562 , n22587 );
xor ( n22802 , n22801 , n22592 );
buf ( n22803 , n22802 );
buf ( n22804 , n22803 );
xor ( n22805 , n22800 , n22804 );
buf ( n22806 , n19143 );
not ( n22807 , n22806 );
buf ( n22808 , n22405 );
not ( n22809 , n22808 );
or ( n22810 , n22807 , n22809 );
buf ( n22811 , n22739 );
buf ( n22812 , n19152 );
nand ( n22813 , n22811 , n22812 );
buf ( n22814 , n22813 );
buf ( n22815 , n22814 );
nand ( n22816 , n22810 , n22815 );
buf ( n22817 , n22816 );
buf ( n22818 , n22817 );
xor ( n22819 , n22805 , n22818 );
buf ( n22820 , n22819 );
buf ( n22821 , n22820 );
and ( n22822 , n22794 , n22821 );
and ( n22823 , n22645 , n22793 );
or ( n22824 , n22822 , n22823 );
buf ( n22825 , n22824 );
not ( n22826 , n22825 );
xor ( n22827 , n22800 , n22804 );
and ( n22828 , n22827 , n22818 );
and ( n22829 , n22800 , n22804 );
or ( n22830 , n22828 , n22829 );
buf ( n22831 , n22830 );
buf ( n22832 , n22831 );
buf ( n22833 , n591 );
not ( n22834 , n22833 );
buf ( n22835 , n22388 );
not ( n22836 , n22835 );
or ( n22837 , n22834 , n22836 );
buf ( n22838 , n22630 );
buf ( n22839 , n19244 );
nand ( n22840 , n22838 , n22839 );
buf ( n22841 , n22840 );
buf ( n22842 , n22841 );
nand ( n22843 , n22837 , n22842 );
buf ( n22844 , n22843 );
buf ( n22845 , n22844 );
xor ( n22846 , n22832 , n22845 );
xor ( n22847 , n22413 , n22597 );
xor ( n22848 , n22847 , n22602 );
buf ( n22849 , n22848 );
buf ( n22850 , n22849 );
xor ( n22851 , n22846 , n22850 );
buf ( n22852 , n22851 );
not ( n22853 , n22852 );
and ( n22854 , n22826 , n22853 );
xor ( n22855 , n22645 , n22793 );
xor ( n22856 , n22855 , n22821 );
buf ( n22857 , n22856 );
buf ( n22858 , n22857 );
buf ( n22859 , n591 );
not ( n22860 , n22859 );
buf ( n22861 , n22637 );
not ( n22862 , n22861 );
or ( n22863 , n22860 , n22862 );
buf ( n22864 , n590 );
not ( n22865 , n22864 );
buf ( n22866 , n19022 );
not ( n22867 , n22866 );
or ( n22868 , n22865 , n22867 );
buf ( n22869 , n18489 );
buf ( n22870 , n590 );
not ( n22871 , n22870 );
buf ( n22872 , n22871 );
buf ( n22873 , n22872 );
nand ( n22874 , n22869 , n22873 );
buf ( n22875 , n22874 );
buf ( n22876 , n22875 );
nand ( n22877 , n22868 , n22876 );
buf ( n22878 , n22877 );
buf ( n22879 , n22878 );
buf ( n22880 , n19244 );
nand ( n22881 , n22879 , n22880 );
buf ( n22882 , n22881 );
buf ( n22883 , n22882 );
nand ( n22884 , n22863 , n22883 );
buf ( n22885 , n22884 );
buf ( n22886 , n22885 );
buf ( n22887 , n18431 );
not ( n22888 , n22887 );
buf ( n22889 , n22666 );
not ( n22890 , n22889 );
or ( n22891 , n22888 , n22890 );
buf ( n22892 , n584 );
not ( n22893 , n22892 );
buf ( n22894 , n21220 );
not ( n22895 , n22894 );
or ( n22896 , n22893 , n22895 );
buf ( n22897 , n21223 );
buf ( n22898 , n18277 );
nand ( n22899 , n22897 , n22898 );
buf ( n22900 , n22899 );
buf ( n22901 , n22900 );
nand ( n22902 , n22896 , n22901 );
buf ( n22903 , n22902 );
buf ( n22904 , n22903 );
buf ( n22905 , n18479 );
nand ( n22906 , n22904 , n22905 );
buf ( n22907 , n22906 );
buf ( n22908 , n22907 );
nand ( n22909 , n22891 , n22908 );
buf ( n22910 , n22909 );
buf ( n22911 , n22910 );
buf ( n22912 , C0 );
buf ( n22913 , n22912 );
xor ( n22914 , n22911 , n22913 );
buf ( n22915 , n18857 );
not ( n22916 , n22915 );
buf ( n22917 , n22711 );
not ( n22918 , n22917 );
or ( n22919 , n22916 , n22918 );
buf ( n22920 , n586 );
not ( n22921 , n22920 );
buf ( n22922 , n21907 );
not ( n22923 , n22922 );
or ( n22924 , n22921 , n22923 );
buf ( n22925 , n13664 );
buf ( n22926 , n18840 );
nand ( n22927 , n22925 , n22926 );
buf ( n22928 , n22927 );
buf ( n22929 , n22928 );
nand ( n22930 , n22924 , n22929 );
buf ( n22931 , n22930 );
buf ( n22932 , n22931 );
buf ( n22933 , n18881 );
nand ( n22934 , n22932 , n22933 );
buf ( n22935 , n22934 );
buf ( n22936 , n22935 );
nand ( n22937 , n22919 , n22936 );
buf ( n22938 , n22937 );
buf ( n22939 , n22938 );
and ( n22940 , n22914 , n22939 );
or ( n22941 , n22940 , C0 );
buf ( n22942 , n22941 );
buf ( n22943 , n22942 );
not ( n22944 , n19152 );
and ( n22945 , n588 , n19000 );
not ( n22946 , n588 );
and ( n22947 , n22946 , n18997 );
or ( n22948 , n22945 , n22947 );
not ( n22949 , n22948 );
or ( n22950 , n22944 , n22949 );
nand ( n22951 , n22748 , n19143 );
nand ( n22952 , n22950 , n22951 );
buf ( n22953 , n22952 );
xor ( n22954 , n22943 , n22953 );
xor ( n22955 , n22674 , n22678 );
xor ( n22956 , n22955 , n22719 );
buf ( n22957 , n22956 );
buf ( n22958 , n22957 );
and ( n22959 , n22954 , n22958 );
and ( n22960 , n22943 , n22953 );
or ( n22961 , n22959 , n22960 );
buf ( n22962 , n22961 );
buf ( n22963 , n22962 );
xor ( n22964 , n22886 , n22963 );
xor ( n22965 , n22724 , n22753 );
xor ( n22966 , n22965 , n22788 );
buf ( n22967 , n22966 );
buf ( n22968 , n22967 );
and ( n22969 , n22964 , n22968 );
and ( n22970 , n22886 , n22963 );
or ( n22971 , n22969 , n22970 );
buf ( n22972 , n22971 );
buf ( n22973 , n22972 );
nor ( n22974 , n22858 , n22973 );
buf ( n22975 , n22974 );
nor ( n22976 , n22854 , n22975 );
xor ( n22977 , n22886 , n22963 );
xor ( n22978 , n22977 , n22968 );
buf ( n22979 , n22978 );
buf ( n22980 , n22979 );
not ( n22981 , n22980 );
buf ( n22982 , C0 );
buf ( n22983 , n22982 );
buf ( n22984 , n18431 );
not ( n22985 , n22984 );
buf ( n22986 , n22903 );
not ( n22987 , n22986 );
or ( n22988 , n22985 , n22987 );
buf ( n22989 , n584 );
not ( n22990 , n22989 );
buf ( n22991 , n20452 );
not ( n22992 , n22991 );
or ( n22993 , n22990 , n22992 );
buf ( n22994 , n20455 );
buf ( n22995 , n18277 );
nand ( n22996 , n22994 , n22995 );
buf ( n22997 , n22996 );
buf ( n22998 , n22997 );
nand ( n22999 , n22993 , n22998 );
buf ( n23000 , n22999 );
buf ( n23001 , n23000 );
buf ( n23002 , n18479 );
nand ( n23003 , n23001 , n23002 );
buf ( n23004 , n23003 );
buf ( n23005 , n23004 );
nand ( n23006 , n22988 , n23005 );
buf ( n23007 , n23006 );
buf ( n23008 , n23007 );
xor ( n23009 , n22983 , n23008 );
buf ( n23010 , C0 );
buf ( n23011 , n23010 );
buf ( n23012 , C0 );
buf ( n23013 , n23012 );
buf ( n23014 , n584 );
not ( n23015 , n23014 );
or ( n23016 , n23015 , C0 );
buf ( n23017 , C1 );
buf ( n23018 , n23017 );
nand ( n23019 , n23016 , n23018 );
buf ( n23020 , n23019 );
not ( n23021 , n23020 );
not ( n23022 , n18431 );
or ( n23023 , n23021 , n23022 );
buf ( n23024 , n584 );
buf ( n23025 , n20773 );
and ( n23026 , n23024 , n23025 );
nor ( n23027 , n23026 , C0 );
buf ( n23028 , n23027 );
buf ( n23029 , n23028 );
not ( n23030 , n23029 );
buf ( n23031 , n18479 );
nand ( n23032 , n23030 , n23031 );
buf ( n23033 , n23032 );
nand ( n23034 , n23023 , n23033 );
buf ( n23035 , n23034 );
xor ( n23036 , n23013 , n23035 );
buf ( n23037 , C1 );
buf ( n23038 , n23037 );
buf ( n23039 , n585 );
buf ( n23040 , n586 );
and ( n23041 , n23039 , n23040 );
buf ( n23042 , n18277 );
nor ( n23043 , n23041 , n23042 );
buf ( n23044 , n23043 );
buf ( n23045 , n23044 );
and ( n23046 , n23038 , n23045 );
buf ( n23047 , n23046 );
buf ( n23048 , n23047 );
buf ( n23049 , n23028 );
buf ( n23050 , n18912 );
or ( n23051 , n23049 , n23050 );
buf ( n23052 , C1 );
buf ( n23053 , n23052 );
buf ( n23054 , n18479 );
not ( n23055 , n23054 );
buf ( n23056 , n23055 );
buf ( n23057 , n23056 );
buf ( n23058 , n18277 );
nor ( n23059 , n23057 , n23058 );
buf ( n23060 , n23059 );
buf ( n23061 , n23060 );
and ( n23062 , n23053 , n23061 );
nor ( n23063 , C0 , n23062 );
buf ( n23064 , n23063 );
buf ( n23065 , n23064 );
nand ( n23066 , n23051 , n23065 );
buf ( n23067 , n23066 );
buf ( n23068 , n23067 );
and ( n23069 , n23048 , n23068 );
buf ( n23070 , n23069 );
buf ( n23071 , n23070 );
and ( n23072 , n23036 , n23071 );
or ( n23073 , n23072 , C0 );
buf ( n23074 , n23073 );
buf ( n23075 , n23074 );
xor ( n23076 , n23011 , n23075 );
buf ( n23077 , n18431 );
not ( n23078 , n23077 );
buf ( n23079 , n23000 );
not ( n23080 , n23079 );
or ( n23081 , n23078 , n23080 );
buf ( n23082 , n23020 );
buf ( n23083 , n18479 );
nand ( n23084 , n23082 , n23083 );
buf ( n23085 , n23084 );
buf ( n23086 , n23085 );
nand ( n23087 , n23081 , n23086 );
buf ( n23088 , n23087 );
buf ( n23089 , n23088 );
and ( n23090 , n23076 , n23089 );
or ( n23091 , n23090 , C0 );
buf ( n23092 , n23091 );
buf ( n23093 , n23092 );
and ( n23094 , n23009 , n23093 );
or ( n23095 , n23094 , C0 );
buf ( n23096 , n23095 );
buf ( n23097 , n23096 );
xor ( n23098 , n22911 , n22913 );
xor ( n23099 , n23098 , n22939 );
buf ( n23100 , n23099 );
buf ( n23101 , n23100 );
xor ( n23102 , n23097 , n23101 );
buf ( n23103 , n19143 );
not ( n23104 , n23103 );
buf ( n23105 , n22948 );
not ( n23106 , n23105 );
or ( n23107 , n23104 , n23106 );
and ( n23108 , n588 , n19549 );
not ( n23109 , n588 );
and ( n23110 , n23109 , n13663 );
or ( n23111 , n23108 , n23110 );
buf ( n23112 , n23111 );
buf ( n23113 , n19152 );
nand ( n23114 , n23112 , n23113 );
buf ( n23115 , n23114 );
buf ( n23116 , n23115 );
nand ( n23117 , n23107 , n23116 );
buf ( n23118 , n23117 );
buf ( n23119 , n23118 );
and ( n23120 , n23102 , n23119 );
and ( n23121 , n23097 , n23101 );
or ( n23122 , n23120 , n23121 );
buf ( n23123 , n23122 );
buf ( n23124 , n23123 );
xor ( n23125 , n22943 , n22953 );
xor ( n23126 , n23125 , n22958 );
buf ( n23127 , n23126 );
buf ( n23128 , n23127 );
xor ( n23129 , n23124 , n23128 );
buf ( n23130 , n591 );
not ( n23131 , n23130 );
buf ( n23132 , n22878 );
not ( n23133 , n23132 );
or ( n23134 , n23131 , n23133 );
buf ( n23135 , n590 );
not ( n23136 , n23135 );
buf ( n23137 , n18569 );
not ( n23138 , n23137 );
or ( n23139 , n23136 , n23138 );
buf ( n23140 , n590 );
not ( n23141 , n23140 );
buf ( n23142 , n18566 );
nand ( n23143 , n23141 , n23142 );
buf ( n23144 , n23143 );
buf ( n23145 , n23144 );
nand ( n23146 , n23139 , n23145 );
buf ( n23147 , n23146 );
buf ( n23148 , n23147 );
buf ( n23149 , n19244 );
nand ( n23150 , n23148 , n23149 );
buf ( n23151 , n23150 );
buf ( n23152 , n23151 );
nand ( n23153 , n23134 , n23152 );
buf ( n23154 , n23153 );
buf ( n23155 , n23154 );
and ( n23156 , n23129 , n23155 );
and ( n23157 , n23124 , n23128 );
or ( n23158 , n23156 , n23157 );
buf ( n23159 , n23158 );
buf ( n23160 , n23159 );
not ( n23161 , n23160 );
buf ( n23162 , n23161 );
buf ( n23163 , n23162 );
nand ( n23164 , n22981 , n23163 );
buf ( n23165 , n23164 );
not ( n23166 , n23165 );
buf ( n23167 , C0 );
buf ( n23168 , n23167 );
buf ( n23169 , n18853 );
not ( n23170 , n23169 );
buf ( n23171 , n586 );
not ( n23172 , n23171 );
buf ( n23173 , n21214 );
not ( n23174 , n23173 );
or ( n23175 , n23172 , n23174 );
buf ( n23176 , n13666 );
buf ( n23177 , n18840 );
nand ( n23178 , n23176 , n23177 );
buf ( n23179 , n23178 );
buf ( n23180 , n23179 );
nand ( n23181 , n23175 , n23180 );
buf ( n23182 , n23181 );
buf ( n23183 , n23182 );
not ( n23184 , n23183 );
or ( n23185 , n23170 , n23184 );
buf ( n23186 , n586 );
not ( n23187 , n23186 );
buf ( n23188 , n21406 );
not ( n23189 , n23188 );
or ( n23190 , n23187 , n23189 );
buf ( n23191 , n20455 );
buf ( n23192 , n18840 );
nand ( n23193 , n23191 , n23192 );
buf ( n23194 , n23193 );
buf ( n23195 , n23194 );
nand ( n23196 , n23190 , n23195 );
buf ( n23197 , n23196 );
buf ( n23198 , n23197 );
buf ( n23199 , n18881 );
nand ( n23200 , n23198 , n23199 );
buf ( n23201 , n23200 );
buf ( n23202 , n23201 );
nand ( n23203 , n23185 , n23202 );
buf ( n23204 , n23203 );
buf ( n23205 , n23204 );
xor ( n23206 , n23168 , n23205 );
buf ( n23207 , C0 );
buf ( n23208 , n23207 );
buf ( n23209 , C0 );
buf ( n23210 , n23209 );
not ( n23211 , n18853 );
nor ( n23212 , n23211 , n18840 );
nand ( n23213 , C1 , n23212 );
buf ( n23214 , n586 );
not ( n23215 , n23214 );
or ( n23216 , n23215 , C0 );
buf ( n23217 , C1 );
buf ( n23218 , n23217 );
nand ( n23219 , n23216 , n23218 );
buf ( n23220 , n23219 );
nand ( n23221 , n23220 , n18881 );
nand ( n23222 , n23213 , C1 , n23221 );
buf ( n23223 , n23222 );
xor ( n23224 , n23210 , n23223 );
buf ( n23225 , C1 );
buf ( n23226 , n23225 );
buf ( n23227 , n587 );
buf ( n23228 , n588 );
and ( n23229 , n23227 , n23228 );
buf ( n23230 , n18840 );
nor ( n23231 , n23229 , n23230 );
buf ( n23232 , n23231 );
buf ( n23233 , n23232 );
and ( n23234 , n23226 , n23233 );
buf ( n23235 , n23234 );
buf ( n23236 , n23235 );
not ( n23237 , n23236 );
buf ( n23238 , n23220 );
buf ( n23239 , n18853 );
and ( n23240 , n23238 , n23239 );
buf ( n23241 , n23052 );
buf ( n23242 , n586 );
and ( n23243 , n23241 , n23242 );
nor ( n23244 , n23243 , C0 );
buf ( n23245 , n23244 );
buf ( n23246 , n23245 );
buf ( n23247 , n18881 );
not ( n23248 , n23247 );
buf ( n23249 , n23248 );
buf ( n23250 , n23249 );
nor ( n23251 , n23246 , n23250 );
buf ( n23252 , n23251 );
buf ( n23253 , n23252 );
nor ( n23254 , n23240 , n23253 );
buf ( n23255 , n23254 );
buf ( n23256 , n23255 );
nor ( n23257 , n23237 , n23256 );
buf ( n23258 , n23257 );
buf ( n23259 , n23258 );
and ( n23260 , n23224 , n23259 );
or ( n23261 , n23260 , C0 );
buf ( n23262 , n23261 );
buf ( n23263 , n23262 );
xor ( n23264 , n23208 , n23263 );
buf ( n23265 , n18853 );
not ( n23266 , n23265 );
buf ( n23267 , n23197 );
not ( n23268 , n23267 );
or ( n23269 , n23266 , n23268 );
and ( n23270 , n18840 , C1 );
nor ( n23271 , n23270 , C0 );
nand ( n23272 , n23271 , n18881 );
buf ( n23273 , n23272 );
nand ( n23274 , n23269 , n23273 );
buf ( n23275 , n23274 );
buf ( n23276 , n23275 );
and ( n23277 , n23264 , n23276 );
or ( n23278 , n23277 , C0 );
buf ( n23279 , n23278 );
buf ( n23280 , n23279 );
and ( n23281 , n23206 , n23280 );
or ( n23282 , n23281 , C0 );
buf ( n23283 , n23282 );
buf ( n23284 , n23283 );
buf ( n23285 , n18857 );
not ( n23286 , n23285 );
buf ( n23287 , n586 );
not ( n23288 , n23287 );
buf ( n23289 , n22260 );
not ( n23290 , n23289 );
or ( n23291 , n23288 , n23290 );
buf ( n23292 , n19975 );
buf ( n23293 , n18840 );
nand ( n23294 , n23292 , n23293 );
buf ( n23295 , n23294 );
buf ( n23296 , n23295 );
nand ( n23297 , n23291 , n23296 );
buf ( n23298 , n23297 );
buf ( n23299 , n23298 );
not ( n23300 , n23299 );
or ( n23301 , n23286 , n23300 );
buf ( n23302 , n23182 );
buf ( n23303 , n18881 );
nand ( n23304 , n23302 , n23303 );
buf ( n23305 , n23304 );
buf ( n23306 , n23305 );
nand ( n23307 , n23301 , n23306 );
buf ( n23308 , n23307 );
buf ( n23309 , n23308 );
buf ( n23310 , C0 );
buf ( n23311 , n23310 );
xor ( n23312 , n23309 , n23311 );
buf ( n23313 , n19143 );
not ( n23314 , n23313 );
xor ( n23315 , n588 , n19531 );
buf ( n23316 , n23315 );
not ( n23317 , n23316 );
or ( n23318 , n23314 , n23317 );
buf ( n23319 , n588 );
not ( n23320 , n23319 );
buf ( n23321 , n19630 );
not ( n23322 , n23321 );
or ( n23323 , n23320 , n23322 );
buf ( n23324 , n588 );
not ( n23325 , n23324 );
buf ( n23326 , n13664 );
nand ( n23327 , n23325 , n23326 );
buf ( n23328 , n23327 );
buf ( n23329 , n23328 );
nand ( n23330 , n23323 , n23329 );
buf ( n23331 , n23330 );
buf ( n23332 , n23331 );
buf ( n23333 , n19152 );
nand ( n23334 , n23332 , n23333 );
buf ( n23335 , n23334 );
buf ( n23336 , n23335 );
nand ( n23337 , n23318 , n23336 );
buf ( n23338 , n23337 );
buf ( n23339 , n23338 );
xor ( n23340 , n23312 , n23339 );
buf ( n23341 , n23340 );
buf ( n23342 , n23341 );
xor ( n23343 , n23284 , n23342 );
buf ( n23344 , n591 );
not ( n23345 , n23344 );
and ( n23346 , n590 , n19000 );
not ( n23347 , n590 );
and ( n23348 , n23347 , n18997 );
or ( n23349 , n23346 , n23348 );
buf ( n23350 , n23349 );
not ( n23351 , n23350 );
or ( n23352 , n23345 , n23351 );
buf ( n23353 , n590 );
not ( n23354 , n23353 );
buf ( n23355 , n18981 );
not ( n23356 , n23355 );
or ( n23357 , n23354 , n23356 );
buf ( n23358 , n590 );
not ( n23359 , n23358 );
buf ( n23360 , n13663 );
nand ( n23361 , n23359 , n23360 );
buf ( n23362 , n23361 );
buf ( n23363 , n23362 );
nand ( n23364 , n23357 , n23363 );
buf ( n23365 , n23364 );
buf ( n23366 , n23365 );
buf ( n23367 , n19241 );
nand ( n23368 , n23366 , n23367 );
buf ( n23369 , n23368 );
buf ( n23370 , n23369 );
nand ( n23371 , n23352 , n23370 );
buf ( n23372 , n23371 );
buf ( n23373 , n23372 );
xor ( n23374 , n23343 , n23373 );
buf ( n23375 , n23374 );
not ( n23376 , n23375 );
buf ( n23377 , n19143 );
not ( n23378 , n23377 );
buf ( n23379 , n23331 );
not ( n23380 , n23379 );
or ( n23381 , n23378 , n23380 );
and ( n23382 , n588 , n19972 );
not ( n23383 , n588 );
and ( n23384 , n23383 , n20998 );
or ( n23385 , n23382 , n23384 );
buf ( n23386 , n23385 );
buf ( n23387 , n19152 );
nand ( n23388 , n23386 , n23387 );
buf ( n23389 , n23388 );
buf ( n23390 , n23389 );
nand ( n23391 , n23381 , n23390 );
buf ( n23392 , n23391 );
buf ( n23393 , n23392 );
xor ( n23394 , n23168 , n23205 );
xor ( n23395 , n23394 , n23280 );
buf ( n23396 , n23395 );
buf ( n23397 , n23396 );
xor ( n23398 , n23393 , n23397 );
buf ( n23399 , n591 );
not ( n23400 , n23399 );
buf ( n23401 , n23365 );
not ( n23402 , n23401 );
or ( n23403 , n23400 , n23402 );
and ( n23404 , n19531 , n590 );
not ( n23405 , n19531 );
and ( n23406 , n23405 , n990 );
nor ( n23407 , n23404 , n23406 );
buf ( n23408 , n23407 );
buf ( n23409 , n19241 );
nand ( n23410 , n23408 , n23409 );
buf ( n23411 , n23410 );
buf ( n23412 , n23411 );
nand ( n23413 , n23403 , n23412 );
buf ( n23414 , n23413 );
buf ( n23415 , n23414 );
and ( n23416 , n23398 , n23415 );
and ( n23417 , n23393 , n23397 );
or ( n23418 , n23416 , n23417 );
buf ( n23419 , n23418 );
not ( n23420 , n23419 );
nand ( n23421 , n23376 , n23420 );
buf ( n23422 , n23421 );
not ( n23423 , n23422 );
buf ( n23424 , C0 );
buf ( n23425 , n19143 );
not ( n23426 , n23425 );
buf ( n23427 , n588 );
not ( n23428 , n23427 );
buf ( n23429 , n21406 );
and ( n23430 , n23428 , n23429 );
nor ( n23431 , C0 , n23430 );
buf ( n23432 , n23431 );
buf ( n23433 , n23432 );
not ( n23434 , n23433 );
or ( n23435 , n23426 , n23434 );
and ( n23436 , n588 , n20762 );
or ( n23437 , n23436 , C0 );
buf ( n23438 , n23437 );
buf ( n23439 , n19152 );
nand ( n23440 , n23438 , n23439 );
buf ( n23441 , n23440 );
buf ( n23442 , n23441 );
nand ( n23443 , n23435 , n23442 );
buf ( n23444 , n23443 );
buf ( n23445 , n23444 );
buf ( n23446 , C0 );
buf ( n23447 , n23446 );
not ( n23448 , n19152 );
buf ( n23449 , n588 );
not ( n23450 , n23449 );
buf ( n23451 , n23052 );
and ( n23452 , n23450 , n23451 );
nor ( n23453 , C0 , n23452 );
buf ( n23454 , n23453 );
not ( n23455 , n23454 );
or ( n23456 , n23448 , n23455 );
and ( n23457 , C1 , n18849 );
nor ( n23458 , C0 , n23457 );
nand ( n23459 , n23458 , n19143 );
nand ( n23460 , n23456 , n23459 );
buf ( n23461 , n23460 );
not ( n23462 , n23461 );
buf ( n23463 , C1 );
buf ( n23464 , n23463 );
buf ( n23465 , n589 );
buf ( n23466 , n590 );
nand ( n23467 , n23465 , n23466 );
buf ( n23468 , n23467 );
buf ( n23469 , n23468 );
buf ( n23470 , n588 );
nand ( n23471 , n23464 , n23469 , n23470 );
buf ( n23472 , n23471 );
buf ( n23473 , n23472 );
nor ( n23474 , n23462 , n23473 );
buf ( n23475 , n23474 );
buf ( n23476 , n23475 );
xor ( n23477 , n23447 , n23476 );
buf ( n23478 , n19143 );
not ( n23479 , n23478 );
buf ( n23480 , n23437 );
not ( n23481 , n23480 );
or ( n23482 , n23479 , n23481 );
buf ( n23483 , n23458 );
buf ( n23484 , n19152 );
nand ( n23485 , n23483 , n23484 );
buf ( n23486 , n23485 );
buf ( n23487 , n23486 );
nand ( n23488 , n23482 , n23487 );
buf ( n23489 , n23488 );
buf ( n23490 , n23489 );
and ( n23491 , n23477 , n23490 );
or ( n23492 , n23491 , C0 );
buf ( n23493 , n23492 );
buf ( n23494 , n23493 );
buf ( n23495 , C0 );
buf ( n23496 , n591 );
not ( n23497 , n23496 );
buf ( n23498 , n590 );
not ( n23499 , n23498 );
buf ( n23500 , n19972 );
not ( n23501 , n23500 );
or ( n23502 , n23499 , n23501 );
buf ( n23503 , n590 );
not ( n23504 , n23503 );
buf ( n23505 , n20998 );
nand ( n23506 , n23504 , n23505 );
buf ( n23507 , n23506 );
buf ( n23508 , n23507 );
nand ( n23509 , n23502 , n23508 );
buf ( n23510 , n23509 );
buf ( n23511 , n23510 );
not ( n23512 , n23511 );
or ( n23513 , n23497 , n23512 );
buf ( n23514 , n19238 );
buf ( n23515 , n590 );
not ( n23516 , n23515 );
buf ( n23517 , n13666 );
not ( n23518 , n23517 );
buf ( n23519 , n23518 );
buf ( n23520 , n23519 );
not ( n23521 , n23520 );
or ( n23522 , n23516 , n23521 );
buf ( n23523 , n590 );
not ( n23524 , n23523 );
buf ( n23525 , n13666 );
nand ( n23526 , n23524 , n23525 );
buf ( n23527 , n23526 );
buf ( n23528 , n23527 );
nand ( n23529 , n23522 , n23528 );
buf ( n23530 , n23529 );
buf ( n23531 , n23530 );
nand ( n23532 , n23514 , n23531 );
buf ( n23533 , n23532 );
buf ( n23534 , n23533 );
nand ( n23535 , n23513 , n23534 );
buf ( n23536 , n23535 );
buf ( n23537 , C1 );
buf ( n23538 , n23536 );
buf ( n23539 , n23495 );
nor ( n23540 , n23538 , n23539 );
buf ( n23541 , n23540 );
not ( n23542 , n23541 );
buf ( n23543 , n23530 );
buf ( n23544 , n591 );
and ( n23545 , n23543 , n23544 );
buf ( n23546 , n19238 );
not ( n23547 , n23546 );
buf ( n23548 , n20449 );
not ( n23549 , n23548 );
buf ( n23550 , n22872 );
not ( n23551 , n23550 );
and ( n23552 , n23549 , n23551 );
nor ( n23553 , n23552 , C0 );
buf ( n23554 , n23553 );
buf ( n23555 , n23554 );
nor ( n23556 , n23547 , n23555 );
buf ( n23557 , n23556 );
buf ( n23558 , n23557 );
nor ( n23559 , n23545 , n23558 );
buf ( n23560 , n23559 );
buf ( n23561 , C1 );
buf ( n23562 , n23560 );
buf ( n23563 , n23561 );
nand ( n23564 , n23562 , n23563 );
buf ( n23565 , n23564 );
buf ( n23566 , n591 );
not ( n23567 , n23566 );
buf ( n23568 , n23567 );
or ( n23569 , n23554 , n23568 );
buf ( n23570 , C0 );
buf ( n23571 , n590 );
xnor ( n23572 , n23570 , n23571 );
buf ( n23573 , n23572 );
buf ( n23574 , n23573 );
not ( n23575 , n23574 );
buf ( n23576 , n19238 );
nand ( n23577 , n23575 , n23576 );
buf ( n23578 , n23577 );
nand ( n23579 , n23569 , n23578 );
not ( n23580 , n23579 );
buf ( n23581 , C0 );
buf ( n23582 , n23581 );
xor ( n23583 , n590 , C0 );
buf ( n23584 , n23583 );
buf ( n23585 , n591 );
and ( n23586 , n23584 , n23585 );
buf ( n23587 , n19235 );
not ( n23588 , n23587 );
buf ( n23589 , C0 );
nor ( n23590 , n23588 , n23589 );
buf ( n23591 , n23590 );
buf ( n23592 , n23591 );
nor ( n23593 , n23586 , n23592 );
buf ( n23594 , n23593 );
buf ( n23595 , n23594 );
nand ( n23596 , C1 , n590 );
buf ( n23597 , n23596 );
nor ( n23598 , n23595 , n23597 );
buf ( n23599 , n23598 );
buf ( n23600 , n23599 );
xor ( n23601 , n23582 , n23600 );
not ( n23602 , n23583 );
not ( n23603 , n19238 );
or ( n23604 , n23602 , n23603 );
or ( n23605 , n23573 , n23568 );
nand ( n23606 , n23604 , n23605 );
buf ( n23607 , n23606 );
and ( n23608 , n23601 , n23607 );
or ( n23609 , n23608 , C0 );
buf ( n23610 , n23609 );
not ( n23611 , n23610 );
nand ( n23612 , n23611 , C1 );
not ( n23613 , n23612 );
or ( n23614 , n23580 , n23613 );
nand ( n23615 , n23614 , C1 );
nand ( n23616 , n23565 , n23615 );
buf ( n23617 , n23616 );
nand ( n23618 , C1 , n23617 );
buf ( n23619 , n23618 );
nand ( n23620 , n23542 , n23619 );
nand ( n23621 , n23537 , n23620 );
not ( n23622 , n23621 );
buf ( n23623 , C0 );
buf ( n23624 , n23623 );
buf ( n23625 , n19143 );
not ( n23626 , n23625 );
buf ( n23627 , n588 );
buf ( n23628 , n13666 );
and ( n23629 , n23627 , n23628 );
not ( n23630 , n23627 );
buf ( n23631 , n21214 );
and ( n23632 , n23630 , n23631 );
nor ( n23633 , n23629 , n23632 );
buf ( n23634 , n23633 );
buf ( n23635 , n23634 );
not ( n23636 , n23635 );
or ( n23637 , n23626 , n23636 );
buf ( n23638 , n19152 );
buf ( n23639 , n23432 );
nand ( n23640 , n23638 , n23639 );
buf ( n23641 , n23640 );
buf ( n23642 , n23641 );
nand ( n23643 , n23637 , n23642 );
buf ( n23644 , n23643 );
buf ( n23645 , n23644 );
xor ( n23646 , n23624 , n23645 );
xor ( n23647 , n23424 , n23445 );
and ( n23648 , n23647 , n23494 );
or ( n23649 , n23648 , C0 );
buf ( n23650 , n23649 );
buf ( n23651 , n23650 );
xor ( n23652 , n23646 , n23651 );
buf ( n23653 , n23652 );
buf ( n23654 , n591 );
not ( n23655 , n23654 );
xor ( n23656 , n13664 , n590 );
buf ( n23657 , n23656 );
not ( n23658 , n23657 );
or ( n23659 , n23655 , n23658 );
buf ( n23660 , n19241 );
buf ( n23661 , n23510 );
nand ( n23662 , n23660 , n23661 );
buf ( n23663 , n23662 );
buf ( n23664 , n23663 );
nand ( n23665 , n23659 , n23664 );
buf ( n23666 , n23665 );
nor ( n23667 , n23653 , n23666 );
not ( n23668 , n23667 );
not ( n23669 , n23668 );
or ( n23670 , n23622 , n23669 );
nand ( n23671 , n23653 , n23666 );
nand ( n23672 , n23670 , n23671 );
buf ( n23673 , n23672 );
not ( n23674 , n23673 );
buf ( n23675 , n23674 );
buf ( n23676 , n23675 );
buf ( n23677 , n19143 );
not ( n23678 , n23677 );
buf ( n23679 , n23385 );
not ( n23680 , n23679 );
or ( n23681 , n23678 , n23680 );
buf ( n23682 , n23634 );
buf ( n23683 , n19152 );
nand ( n23684 , n23682 , n23683 );
buf ( n23685 , n23684 );
buf ( n23686 , n23685 );
nand ( n23687 , n23681 , n23686 );
buf ( n23688 , n23687 );
buf ( n23689 , n23688 );
buf ( n23690 , C0 );
buf ( n23691 , n23690 );
xor ( n23692 , n23689 , n23691 );
buf ( n23693 , n591 );
not ( n23694 , n23693 );
buf ( n23695 , n23407 );
not ( n23696 , n23695 );
or ( n23697 , n23694 , n23696 );
buf ( n23698 , n23656 );
buf ( n23699 , n19238 );
nand ( n23700 , n23698 , n23699 );
buf ( n23701 , n23700 );
buf ( n23702 , n23701 );
nand ( n23703 , n23697 , n23702 );
buf ( n23704 , n23703 );
buf ( n23705 , n23704 );
xor ( n23706 , n23692 , n23705 );
buf ( n23707 , n23706 );
buf ( n23708 , n23707 );
buf ( n23709 , n23708 );
buf ( n23710 , n23709 );
buf ( n23711 , n23710 );
xor ( n23712 , n23624 , n23645 );
and ( n23713 , n23712 , n23651 );
or ( n23714 , n23713 , C0 );
buf ( n23715 , n23714 );
buf ( n23716 , n23715 );
nor ( n23717 , n23711 , n23716 );
buf ( n23718 , n23717 );
buf ( n23719 , n23718 );
or ( n23720 , n23676 , n23719 );
buf ( n23721 , n23710 );
buf ( n23722 , n23715 );
nand ( n23723 , n23721 , n23722 );
buf ( n23724 , n23723 );
buf ( n23725 , n23724 );
nand ( n23726 , n23720 , n23725 );
buf ( n23727 , n23726 );
buf ( n23728 , n23727 );
not ( n23729 , n23728 );
xor ( n23730 , n23393 , n23397 );
xor ( n23731 , n23730 , n23415 );
buf ( n23732 , n23731 );
not ( n23733 , n23732 );
xor ( n23734 , n23689 , n23691 );
and ( n23735 , n23734 , n23705 );
or ( n23736 , n23735 , C0 );
buf ( n23737 , n23736 );
buf ( n23738 , n23737 );
not ( n23739 , n23738 );
buf ( n23740 , n23739 );
nand ( n23741 , n23733 , n23740 );
buf ( n23742 , n23741 );
not ( n23743 , n23742 );
or ( n23744 , n23729 , n23743 );
buf ( n23745 , n23732 );
buf ( n23746 , n23737 );
nand ( n23747 , n23745 , n23746 );
buf ( n23748 , n23747 );
buf ( n23749 , n23748 );
nand ( n23750 , n23744 , n23749 );
buf ( n23751 , n23750 );
buf ( n23752 , n23751 );
not ( n23753 , n23752 );
or ( n23754 , n23423 , n23753 );
buf ( n23755 , n23375 );
buf ( n23756 , n23419 );
nand ( n23757 , n23755 , n23756 );
buf ( n23758 , n23757 );
buf ( n23759 , n23758 );
nand ( n23760 , n23754 , n23759 );
buf ( n23761 , n23760 );
buf ( n23762 , n23761 );
not ( n23763 , n23762 );
xor ( n23764 , n23309 , n23311 );
and ( n23765 , n23764 , n23339 );
or ( n23766 , n23765 , C0 );
buf ( n23767 , n23766 );
buf ( n23768 , n23767 );
buf ( n23769 , n591 );
not ( n23770 , n23769 );
and ( n23771 , n590 , n18538 );
not ( n23772 , n590 );
and ( n23773 , n23772 , n13665 );
or ( n23774 , n23771 , n23773 );
buf ( n23775 , n23774 );
not ( n23776 , n23775 );
or ( n23777 , n23770 , n23776 );
buf ( n23778 , n23349 );
buf ( n23779 , n19241 );
nand ( n23780 , n23778 , n23779 );
buf ( n23781 , n23780 );
buf ( n23782 , n23781 );
nand ( n23783 , n23777 , n23782 );
buf ( n23784 , n23783 );
buf ( n23785 , n23784 );
xor ( n23786 , n23768 , n23785 );
buf ( n23787 , n18857 );
not ( n23788 , n23787 );
buf ( n23789 , n22931 );
not ( n23790 , n23789 );
or ( n23791 , n23788 , n23790 );
buf ( n23792 , n23298 );
buf ( n23793 , n18881 );
nand ( n23794 , n23792 , n23793 );
buf ( n23795 , n23794 );
buf ( n23796 , n23795 );
nand ( n23797 , n23791 , n23796 );
buf ( n23798 , n23797 );
buf ( n23799 , n23798 );
xor ( n23800 , n22983 , n23008 );
xor ( n23801 , n23800 , n23093 );
buf ( n23802 , n23801 );
buf ( n23803 , n23802 );
xor ( n23804 , n23799 , n23803 );
buf ( n23805 , n19143 );
not ( n23806 , n23805 );
buf ( n23807 , n23111 );
not ( n23808 , n23807 );
or ( n23809 , n23806 , n23808 );
buf ( n23810 , n23315 );
buf ( n23811 , n19152 );
nand ( n23812 , n23810 , n23811 );
buf ( n23813 , n23812 );
buf ( n23814 , n23813 );
nand ( n23815 , n23809 , n23814 );
buf ( n23816 , n23815 );
buf ( n23817 , n23816 );
xor ( n23818 , n23804 , n23817 );
buf ( n23819 , n23818 );
buf ( n23820 , n23819 );
xor ( n23821 , n23786 , n23820 );
buf ( n23822 , n23821 );
xor ( n23823 , n23284 , n23342 );
and ( n23824 , n23823 , n23373 );
and ( n23825 , n23284 , n23342 );
or ( n23826 , n23824 , n23825 );
buf ( n23827 , n23826 );
or ( n23828 , n23822 , n23827 );
buf ( n23829 , n23828 );
not ( n23830 , n23829 );
or ( n23831 , n23763 , n23830 );
buf ( n23832 , n23822 );
buf ( n23833 , n23827 );
nand ( n23834 , n23832 , n23833 );
buf ( n23835 , n23834 );
buf ( n23836 , n23835 );
nand ( n23837 , n23831 , n23836 );
buf ( n23838 , n23837 );
not ( n23839 , n23838 );
buf ( n23840 , n591 );
not ( n23841 , n23840 );
buf ( n23842 , n23147 );
not ( n23843 , n23842 );
or ( n23844 , n23841 , n23843 );
buf ( n23845 , n23774 );
buf ( n23846 , n19244 );
nand ( n23847 , n23845 , n23846 );
buf ( n23848 , n23847 );
buf ( n23849 , n23848 );
nand ( n23850 , n23844 , n23849 );
buf ( n23851 , n23850 );
buf ( n23852 , n23851 );
xor ( n23853 , n23799 , n23803 );
and ( n23854 , n23853 , n23817 );
and ( n23855 , n23799 , n23803 );
or ( n23856 , n23854 , n23855 );
buf ( n23857 , n23856 );
buf ( n23858 , n23857 );
xor ( n23859 , n23852 , n23858 );
xor ( n23860 , n23097 , n23101 );
xor ( n23861 , n23860 , n23119 );
buf ( n23862 , n23861 );
buf ( n23863 , n23862 );
xor ( n23864 , n23859 , n23863 );
buf ( n23865 , n23864 );
buf ( n23866 , n23865 );
xor ( n23867 , n23768 , n23785 );
and ( n23868 , n23867 , n23820 );
and ( n23869 , n23768 , n23785 );
or ( n23870 , n23868 , n23869 );
buf ( n23871 , n23870 );
buf ( n23872 , n23871 );
or ( n23873 , n23866 , n23872 );
buf ( n23874 , n23873 );
not ( n23875 , n23874 );
or ( n23876 , n23839 , n23875 );
buf ( n23877 , n23865 );
buf ( n23878 , n23871 );
nand ( n23879 , n23877 , n23878 );
buf ( n23880 , n23879 );
nand ( n23881 , n23876 , n23880 );
buf ( n23882 , n23881 );
not ( n23883 , n23882 );
xor ( n23884 , n23124 , n23128 );
xor ( n23885 , n23884 , n23155 );
buf ( n23886 , n23885 );
not ( n23887 , n23886 );
buf ( n23888 , n23887 );
xor ( n23889 , n23852 , n23858 );
and ( n23890 , n23889 , n23863 );
and ( n23891 , n23852 , n23858 );
or ( n23892 , n23890 , n23891 );
buf ( n23893 , n23892 );
buf ( n23894 , n23893 );
not ( n23895 , n23894 );
buf ( n23896 , n23895 );
buf ( n23897 , n23896 );
nand ( n23898 , n23888 , n23897 );
buf ( n23899 , n23898 );
buf ( n23900 , n23899 );
not ( n23901 , n23900 );
or ( n23902 , n23883 , n23901 );
buf ( n23903 , n23886 );
buf ( n23904 , n23893 );
nand ( n23905 , n23903 , n23904 );
buf ( n23906 , n23905 );
buf ( n23907 , n23906 );
nand ( n23908 , n23902 , n23907 );
buf ( n23909 , n23908 );
not ( n23910 , n23909 );
or ( n23911 , n23166 , n23910 );
buf ( n23912 , n22979 );
buf ( n23913 , n23912 );
buf ( n23914 , n23913 );
buf ( n23915 , n23914 );
buf ( n23916 , n23159 );
nand ( n23917 , n23915 , n23916 );
buf ( n23918 , n23917 );
nand ( n23919 , n23911 , n23918 );
buf ( n23920 , n23919 );
and ( n23921 , n22976 , n23920 );
buf ( n23922 , n22857 );
not ( n23923 , n23922 );
buf ( n23924 , n22972 );
not ( n23925 , n23924 );
buf ( n23926 , n23925 );
buf ( n23927 , n23926 );
nor ( n23928 , n23923 , n23927 );
buf ( n23929 , n23928 );
not ( n23930 , n23929 );
buf ( n23931 , n22852 );
not ( n23932 , n23931 );
buf ( n23933 , n23932 );
buf ( n23934 , n23933 );
buf ( n23935 , n22825 );
not ( n23936 , n23935 );
buf ( n23937 , n23936 );
buf ( n23938 , n23937 );
nand ( n23939 , n23934 , n23938 );
buf ( n23940 , n23939 );
not ( n23941 , n23940 );
or ( n23942 , n23930 , n23941 );
buf ( n23943 , n22852 );
buf ( n23944 , n22825 );
nand ( n23945 , n23943 , n23944 );
buf ( n23946 , n23945 );
nand ( n23947 , n23942 , n23946 );
nor ( n23948 , n23921 , n23947 );
buf ( n23949 , n23948 );
xor ( n23950 , n22396 , n22607 );
xor ( n23951 , n23950 , n22612 );
buf ( n23952 , n23951 );
buf ( n23953 , n23952 );
xor ( n23954 , n22832 , n22845 );
and ( n23955 , n23954 , n22850 );
and ( n23956 , n22832 , n22845 );
or ( n23957 , n23955 , n23956 );
buf ( n23958 , n23957 );
buf ( n23959 , n23958 );
nor ( n23960 , n23953 , n23959 );
buf ( n23961 , n23960 );
buf ( n23962 , n23961 );
nor ( n23963 , n23949 , n23962 );
buf ( n23964 , n23963 );
buf ( n23965 , n23964 );
not ( n23966 , n23965 );
or ( n23967 , n22624 , n23966 );
buf ( n23968 , n22622 );
buf ( n23969 , n23952 );
buf ( n23970 , n23958 );
nand ( n23971 , n23969 , n23970 );
buf ( n23972 , n23971 );
buf ( n23973 , n23972 );
not ( n23974 , n23973 );
buf ( n23975 , n23974 );
buf ( n23976 , n23975 );
and ( n23977 , n23968 , n23976 );
buf ( n23978 , n22377 );
buf ( n23979 , n22616 );
nand ( n23980 , n23978 , n23979 );
buf ( n23981 , n23980 );
buf ( n23982 , n23981 );
not ( n23983 , n23982 );
buf ( n23984 , n23983 );
buf ( n23985 , n23984 );
nor ( n23986 , n23977 , n23985 );
buf ( n23987 , n23986 );
buf ( n23988 , n23987 );
nand ( n23989 , n23967 , n23988 );
buf ( n23990 , n23989 );
nand ( n23991 , n22003 , n22374 , n23990 );
buf ( n23992 , n21805 );
not ( n23993 , n23992 );
buf ( n23994 , n22000 );
nand ( n23995 , n23993 , n23994 );
buf ( n23996 , n23995 );
or ( n23997 , n22364 , n22370 );
buf ( n23998 , n22364 );
buf ( n23999 , n22370 );
nand ( n24000 , n23998 , n23999 );
buf ( n24001 , n24000 );
buf ( n24002 , n24001 );
buf ( n24003 , n22228 );
buf ( n24004 , n22359 );
nand ( n24005 , n24003 , n24004 );
buf ( n24006 , n24005 );
buf ( n24007 , n24006 );
nand ( n24008 , n24002 , n24007 );
buf ( n24009 , n24008 );
nand ( n24010 , n23996 , n23997 , n24009 );
buf ( n24011 , n21805 );
buf ( n24012 , n24011 );
buf ( n24013 , n24012 );
nand ( n24014 , n24013 , n21997 );
nand ( n24015 , n23991 , n24010 , n24014 );
not ( n24016 , n24015 );
or ( n24017 , n21802 , n24016 );
buf ( n24018 , n21368 );
not ( n24019 , n24018 );
buf ( n24020 , n24019 );
buf ( n24021 , n24020 );
buf ( n24022 , n21631 );
not ( n24023 , n24022 );
buf ( n24024 , n24023 );
buf ( n24025 , n24024 );
nand ( n24026 , n24021 , n24025 );
buf ( n24027 , n24026 );
buf ( n24028 , n24027 );
buf ( n24029 , n21638 );
not ( n24030 , n24029 );
buf ( n24031 , n21797 );
not ( n24032 , n24031 );
buf ( n24033 , n24032 );
buf ( n24034 , n24033 );
nor ( n24035 , n24030 , n24034 );
buf ( n24036 , n24035 );
buf ( n24037 , n24036 );
and ( n24038 , n24028 , n24037 );
buf ( n24039 , n21368 );
buf ( n24040 , n21631 );
and ( n24041 , n24039 , n24040 );
buf ( n24042 , n24041 );
buf ( n24043 , n24042 );
nor ( n24044 , n24038 , n24043 );
buf ( n24045 , n24044 );
nand ( n24046 , n24017 , n24045 );
not ( n24047 , n24046 );
or ( n24048 , n21365 , n24047 );
buf ( n24049 , n21117 );
buf ( n24050 , n21358 );
nand ( n24051 , n24049 , n24050 );
buf ( n24052 , n24051 );
buf ( n24053 , n24052 );
nand ( n24054 , n24048 , n24053 );
not ( n24055 , n24054 );
or ( n24056 , n21114 , n24055 );
not ( n24057 , n21106 );
not ( n24058 , n21111 );
and ( n24059 , n24057 , n24058 );
nor ( n24060 , n20375 , n20613 );
nor ( n24061 , n24059 , n24060 );
nand ( n24062 , n21102 , n20703 );
not ( n24063 , n24062 );
and ( n24064 , n24061 , n24063 );
nand ( n24065 , n21106 , n21111 );
or ( n24066 , n20614 , n24065 );
nand ( n24067 , n20375 , n20613 );
nand ( n24068 , n24066 , n24067 );
nor ( n24069 , n24064 , n24068 );
nand ( n24070 , n24056 , n24069 );
buf ( n24071 , n24070 );
not ( n24072 , n24071 );
or ( n24073 , n20372 , n24072 );
not ( n24074 , n19826 );
not ( n24075 , n20123 );
or ( n24076 , n24074 , n24075 );
nor ( n24077 , n20123 , n19826 );
nand ( n24078 , n20366 , n20127 );
or ( n24079 , n24077 , n24078 );
nand ( n24080 , n24076 , n24079 );
buf ( n24081 , n24080 );
not ( n24082 , n24081 );
buf ( n24083 , n24082 );
buf ( n24084 , n24083 );
nand ( n24085 , n24073 , n24084 );
buf ( n24086 , n24085 );
not ( n24087 , n24086 );
not ( n24088 , n24087 );
or ( n24089 , n19823 , n24088 );
nand ( n24090 , n24086 , n19821 );
nand ( n24091 , n24089 , n24090 );
buf ( n24092 , n24091 );
buf ( n24093 , n24092 );
xor ( n24094 , n18214 , n18215 );
xor ( n24095 , n24094 , n24093 );
buf ( n24096 , n24095 );
xor ( n24097 , n18214 , n18215 );
and ( n24098 , n24097 , n24093 );
and ( n24099 , n18214 , n18215 );
or ( n24100 , n24098 , n24099 );
buf ( n24101 , n24100 );
buf ( n24102 , n17633 );
buf ( n24103 , n17603 );
buf ( n24104 , n18418 );
not ( n24105 , n24104 );
xor ( n24106 , n580 , n15680 );
buf ( n24107 , n24106 );
not ( n24108 , n24107 );
or ( n24109 , n24105 , n24108 );
not ( n24110 , n580 );
not ( n24111 , n18296 );
or ( n24112 , n24110 , n24111 );
nand ( n24113 , n18909 , n18402 );
nand ( n24114 , n24112 , n24113 );
buf ( n24115 , n24114 );
buf ( n24116 , n18392 );
nand ( n24117 , n24115 , n24116 );
buf ( n24118 , n24117 );
buf ( n24119 , n24118 );
nand ( n24120 , n24109 , n24119 );
buf ( n24121 , n24120 );
buf ( n24122 , n24121 );
buf ( n24123 , n18725 );
not ( n24124 , n24123 );
buf ( n24125 , n18285 );
not ( n24126 , n24125 );
buf ( n24127 , n24126 );
buf ( n24128 , n24127 );
buf ( n24129 , n18303 );
nor ( n24130 , n24128 , n24129 );
buf ( n24131 , n24130 );
buf ( n24132 , n24131 );
nand ( n24133 , n24124 , n24132 );
buf ( n24134 , n24133 );
not ( n24135 , n18725 );
buf ( n24136 , n24135 );
not ( n24137 , n24136 );
buf ( n24138 , n18657 );
not ( n24139 , n24138 );
buf ( n24140 , n582 );
nor ( n24141 , n24139 , n24140 );
buf ( n24142 , n24141 );
buf ( n24143 , n24142 );
nand ( n24144 , n24137 , n24143 );
buf ( n24145 , n24144 );
buf ( n24146 , n582 );
not ( n24147 , n24146 );
buf ( n24148 , n18868 );
not ( n24149 , n24148 );
or ( n24150 , n24147 , n24149 );
buf ( n24151 , n18303 );
buf ( n24152 , n18439 );
nand ( n24153 , n24151 , n24152 );
buf ( n24154 , n24153 );
buf ( n24155 , n24154 );
nand ( n24156 , n24150 , n24155 );
buf ( n24157 , n24156 );
buf ( n24158 , n24157 );
buf ( n24159 , n18316 );
nand ( n24160 , n24158 , n24159 );
buf ( n24161 , n24160 );
nand ( n24162 , n24134 , n24145 , n24161 );
buf ( n24163 , n24162 );
xor ( n24164 , n24122 , n24163 );
and ( n24165 , n18351 , n18358 );
buf ( n24166 , n24165 );
buf ( n24167 , n24166 );
buf ( n24168 , n18264 );
not ( n24169 , n24168 );
buf ( n24170 , n18239 );
not ( n24171 , n24170 );
or ( n24172 , n24169 , n24171 );
and ( n24173 , n10819 , n18233 );
not ( n24174 , n10819 );
and ( n24175 , n24174 , n578 );
or ( n24176 , n24173 , n24175 );
buf ( n24177 , n24176 );
buf ( n24178 , n18219 );
nand ( n24179 , n24177 , n24178 );
buf ( n24180 , n24179 );
buf ( n24181 , n24180 );
nand ( n24182 , n24172 , n24181 );
buf ( n24183 , n24182 );
buf ( n24184 , n24183 );
xor ( n24185 , n24167 , n24184 );
buf ( n24186 , n18340 );
not ( n24187 , n24186 );
buf ( n24188 , n576 );
buf ( n24189 , n9497 );
xor ( n24190 , n24188 , n24189 );
buf ( n24191 , n24190 );
buf ( n24192 , n24191 );
not ( n24193 , n24192 );
or ( n24194 , n24187 , n24193 );
buf ( n24195 , n18347 );
buf ( n24196 , n18365 );
nand ( n24197 , n24195 , n24196 );
buf ( n24198 , n24197 );
buf ( n24199 , n24198 );
nand ( n24200 , n24194 , n24199 );
buf ( n24201 , n24200 );
buf ( n24202 , n24201 );
and ( n24203 , n24185 , n24202 );
and ( n24204 , n24167 , n24184 );
or ( n24205 , n24203 , n24204 );
buf ( n24206 , n24205 );
buf ( n24207 , n24206 );
xor ( n24208 , n24164 , n24207 );
buf ( n24209 , n24208 );
buf ( n24210 , n24209 );
xor ( n24211 , n24167 , n24184 );
xor ( n24212 , n24211 , n24202 );
buf ( n24213 , n24212 );
buf ( n24214 , n24213 );
buf ( n24215 , n18431 );
not ( n24216 , n24215 );
buf ( n24217 , n18277 );
not ( n24218 , n18082 );
buf ( n24219 , n24218 );
and ( n24220 , n24217 , n24219 );
not ( n24221 , n24217 );
buf ( n24222 , n18082 );
and ( n24223 , n24221 , n24222 );
nor ( n24224 , n24220 , n24223 );
buf ( n24225 , n24224 );
buf ( n24226 , n24225 );
not ( n24227 , n24226 );
or ( n24228 , n24216 , n24227 );
buf ( n24229 , n18736 );
buf ( n24230 , n18479 );
nand ( n24231 , n24229 , n24230 );
buf ( n24232 , n24231 );
buf ( n24233 , n24232 );
nand ( n24234 , n24228 , n24233 );
buf ( n24235 , n24234 );
buf ( n24236 , n24235 );
xor ( n24237 , n24214 , n24236 );
buf ( n24238 , n18857 );
not ( n24239 , n24238 );
buf ( n24240 , n19218 );
buf ( n24241 , n586 );
and ( n24242 , n24240 , n24241 );
not ( n24243 , n24240 );
buf ( n24244 , n18840 );
and ( n24245 , n24243 , n24244 );
or ( n24246 , n24242 , n24245 );
buf ( n24247 , n24246 );
buf ( n24248 , n24247 );
not ( n24249 , n24248 );
or ( n24250 , n24239 , n24249 );
buf ( n24251 , n18881 );
buf ( n24252 , n19373 );
nand ( n24253 , n24251 , n24252 );
buf ( n24254 , n24253 );
buf ( n24255 , n24254 );
nand ( n24256 , n24250 , n24255 );
buf ( n24257 , n24256 );
buf ( n24258 , n24257 );
and ( n24259 , n24237 , n24258 );
and ( n24260 , n24214 , n24236 );
or ( n24261 , n24259 , n24260 );
buf ( n24262 , n24261 );
buf ( n24263 , n24262 );
xor ( n24264 , n24210 , n24263 );
and ( n24265 , n18343 , n18345 );
buf ( n24266 , n24265 );
buf ( n24267 , n24266 );
buf ( n24268 , n18264 );
not ( n24269 , n24268 );
buf ( n24270 , n24176 );
not ( n24271 , n24270 );
or ( n24272 , n24269 , n24271 );
nand ( n24273 , n18409 , n578 );
not ( n24274 , n24273 );
buf ( n24275 , n13592 );
buf ( n24276 , n18233 );
nand ( n24277 , n24275 , n24276 );
buf ( n24278 , n24277 );
not ( n24279 , n24278 );
or ( n24280 , n24274 , n24279 );
nand ( n24281 , n24280 , n18219 );
buf ( n24282 , n24281 );
nand ( n24283 , n24272 , n24282 );
buf ( n24284 , n24283 );
buf ( n24285 , n24284 );
xor ( n24286 , n24267 , n24285 );
not ( n24287 , n18340 );
not ( n24288 , n576 );
not ( n24289 , n18894 );
or ( n24290 , n24288 , n24289 );
buf ( n24291 , n10184 );
buf ( n24292 , n7809 );
nand ( n24293 , n24291 , n24292 );
buf ( n24294 , n24293 );
nand ( n24295 , n24290 , n24294 );
not ( n24296 , n24295 );
or ( n24297 , n24287 , n24296 );
buf ( n24298 , n24191 );
buf ( n24299 , n18365 );
nand ( n24300 , n24298 , n24299 );
buf ( n24301 , n24300 );
nand ( n24302 , n24297 , n24301 );
buf ( n24303 , n24302 );
xor ( n24304 , n24286 , n24303 );
buf ( n24305 , n24304 );
buf ( n24306 , n24305 );
buf ( n24307 , n19254 );
not ( n24308 , n24307 );
buf ( n24309 , n23056 );
buf ( n24310 , n584 );
nor ( n24311 , n24309 , n24310 );
buf ( n24312 , n24311 );
buf ( n24313 , n24312 );
nand ( n24314 , n24308 , n24313 );
buf ( n24315 , n24314 );
buf ( n24316 , n24315 );
buf ( n24317 , n19167 );
not ( n24318 , n24317 );
buf ( n24319 , n18917 );
not ( n24320 , n24319 );
and ( n24321 , n24318 , n24320 );
buf ( n24322 , n18137 );
not ( n24323 , n24322 );
buf ( n24324 , n24323 );
buf ( n24325 , n24324 );
not ( n24326 , n24325 );
buf ( n24327 , n24326 );
buf ( n24328 , n24327 );
buf ( n24329 , n18936 );
and ( n24330 , n24328 , n24329 );
nor ( n24331 , n24321 , n24330 );
buf ( n24332 , n24331 );
buf ( n24333 , n24332 );
nand ( n24334 , n24218 , n23060 );
buf ( n24335 , n24334 );
nand ( n24336 , n24316 , n24333 , n24335 );
buf ( n24337 , n24336 );
buf ( n24338 , n24337 );
xor ( n24339 , n24306 , n24338 );
not ( n24340 , n24247 );
not ( n24341 , n18881 );
or ( n24342 , n24340 , n24341 );
not ( n24343 , n18856 );
buf ( n24344 , n586 );
not ( n24345 , n24344 );
not ( n24346 , n19209 );
buf ( n24347 , n24346 );
not ( n24348 , n24347 );
or ( n24349 , n24345 , n24348 );
buf ( n24350 , n19387 );
buf ( n24351 , n18840 );
nand ( n24352 , n24350 , n24351 );
buf ( n24353 , n24352 );
buf ( n24354 , n24353 );
nand ( n24355 , n24349 , n24354 );
buf ( n24356 , n24355 );
nand ( n24357 , n24343 , n24356 );
nand ( n24358 , n24342 , n24357 );
buf ( n24359 , n24358 );
xor ( n24360 , n24339 , n24359 );
buf ( n24361 , n24360 );
buf ( n24362 , n24361 );
xor ( n24363 , n24264 , n24362 );
buf ( n24364 , n24363 );
buf ( n24365 , n24364 );
xor ( n24366 , n19381 , n19394 );
and ( n24367 , n24366 , n19415 );
and ( n24368 , n19381 , n19394 );
or ( n24369 , n24367 , n24368 );
buf ( n24370 , n24369 );
buf ( n24371 , n24370 );
not ( n24372 , n19152 );
not ( n24373 , n19389 );
or ( n24374 , n24372 , n24373 );
and ( n24375 , n19403 , n21826 );
not ( n24376 , n19403 );
and ( n24377 , n24376 , n21816 );
nor ( n24378 , n24375 , n24377 );
nand ( n24379 , n24374 , n24378 );
buf ( n24380 , n24379 );
xor ( n24381 , n18271 , n18323 );
and ( n24382 , n24381 , n18424 );
and ( n24383 , n18271 , n18323 );
or ( n24384 , n24382 , n24383 );
buf ( n24385 , n24384 );
buf ( n24386 , n24385 );
xor ( n24387 , n24380 , n24386 );
not ( n24388 , n18418 );
not ( n24389 , n24114 );
or ( n24390 , n24388 , n24389 );
not ( n24391 , n18415 );
not ( n24392 , n18410 );
or ( n24393 , n24391 , n24392 );
nand ( n24394 , n24393 , n18392 );
nand ( n24395 , n24390 , n24394 );
buf ( n24396 , n24395 );
buf ( n24397 , n18316 );
not ( n24398 , n24397 );
buf ( n24399 , n18288 );
not ( n24400 , n24399 );
or ( n24401 , n24398 , n24400 );
buf ( n24402 , n24157 );
buf ( n24403 , n18657 );
nand ( n24404 , n24402 , n24403 );
buf ( n24405 , n24404 );
buf ( n24406 , n24405 );
nand ( n24407 , n24401 , n24406 );
buf ( n24408 , n24407 );
buf ( n24409 , n24408 );
xor ( n24410 , n24396 , n24409 );
xor ( n24411 , n18336 , n18372 );
and ( n24412 , n24411 , n18421 );
and ( n24413 , n18336 , n18372 );
or ( n24414 , n24412 , n24413 );
buf ( n24415 , n24414 );
buf ( n24416 , n24415 );
xor ( n24417 , n24410 , n24416 );
buf ( n24418 , n24417 );
buf ( n24419 , n24418 );
xor ( n24420 , n24387 , n24419 );
buf ( n24421 , n24420 );
buf ( n24422 , n24421 );
xor ( n24423 , n24371 , n24422 );
xor ( n24424 , n18427 , n18707 );
and ( n24425 , n24424 , n18833 );
and ( n24426 , n18427 , n18707 );
or ( n24427 , n24425 , n24426 );
buf ( n24428 , n24427 );
buf ( n24429 , n24428 );
and ( n24430 , n24423 , n24429 );
and ( n24431 , n24371 , n24422 );
or ( n24432 , n24430 , n24431 );
buf ( n24433 , n24432 );
buf ( n24434 , n24433 );
xor ( n24435 , n24365 , n24434 );
xor ( n24436 , n24380 , n24386 );
and ( n24437 , n24436 , n24419 );
and ( n24438 , n24380 , n24386 );
or ( n24439 , n24437 , n24438 );
buf ( n24440 , n24439 );
buf ( n24441 , n24440 );
buf ( n24442 , n19152 );
not ( n24443 , n24442 );
buf ( n24444 , n588 );
buf ( n24445 , n19403 );
and ( n24446 , n24444 , n24445 );
not ( n24447 , n24444 );
buf ( n24448 , n19403 );
not ( n24449 , n24448 );
buf ( n24450 , n24449 );
buf ( n24451 , n24450 );
and ( n24452 , n24447 , n24451 );
nor ( n24453 , n24446 , n24452 );
buf ( n24454 , n24453 );
buf ( n24455 , n24454 );
not ( n24456 , n24455 );
or ( n24457 , n24443 , n24456 );
buf ( n24458 , n588 );
not ( n24459 , n24458 );
buf ( n24460 , n19398 );
not ( n24461 , n24460 );
buf ( n24462 , n24461 );
buf ( n24463 , n24462 );
not ( n24464 , n24463 );
or ( n24465 , n24459 , n24464 );
buf ( n24466 , n588 );
not ( n24467 , n24466 );
buf ( n24468 , n19398 );
nand ( n24469 , n24467 , n24468 );
buf ( n24470 , n24469 );
buf ( n24471 , n24470 );
nand ( n24472 , n24465 , n24471 );
buf ( n24473 , n24472 );
buf ( n24474 , n24473 );
buf ( n24475 , n19143 );
nand ( n24476 , n24474 , n24475 );
buf ( n24477 , n24476 );
buf ( n24478 , n24477 );
nand ( n24479 , n24457 , n24478 );
buf ( n24480 , n24479 );
buf ( n24481 , n24480 );
xor ( n24482 , n24396 , n24409 );
and ( n24483 , n24482 , n24416 );
and ( n24484 , n24396 , n24409 );
or ( n24485 , n24483 , n24484 );
buf ( n24486 , n24485 );
buf ( n24487 , n24486 );
xor ( n24488 , n24481 , n24487 );
buf ( n24489 , n590 );
not ( n24490 , n24489 );
buf ( n24491 , n17795 );
nand ( n24492 , n17975 , n17974 );
not ( n24493 , n24492 );
and ( n24494 , n24491 , n24493 );
not ( n24495 , n24491 );
and ( n24496 , n24495 , n24492 );
nor ( n24497 , n24494 , n24496 );
not ( n24498 , n24497 );
buf ( n24499 , n24498 );
not ( n24500 , n24499 );
or ( n24501 , n24490 , n24500 );
not ( n24502 , n590 );
nand ( n24503 , n24502 , n24497 );
buf ( n24504 , n24503 );
nand ( n24505 , n24501 , n24504 );
buf ( n24506 , n24505 );
not ( n24507 , n24506 );
not ( n24508 , n591 );
or ( n24509 , n24507 , n24508 );
buf ( n24510 , n17997 );
not ( n24511 , n24510 );
buf ( n24512 , n24511 );
and ( n24513 , n590 , n24512 );
not ( n24514 , n590 );
and ( n24515 , n24514 , n17997 );
or ( n24516 , n24513 , n24515 );
buf ( n24517 , n24516 );
buf ( n24518 , n19244 );
nand ( n24519 , n24517 , n24518 );
buf ( n24520 , n24519 );
nand ( n24521 , n24509 , n24520 );
buf ( n24522 , n24521 );
xor ( n24523 , n24488 , n24522 );
buf ( n24524 , n24523 );
buf ( n24525 , n24524 );
xor ( n24526 , n24441 , n24525 );
buf ( n24527 , n591 );
not ( n24528 , n24527 );
buf ( n24529 , n24516 );
not ( n24530 , n24529 );
or ( n24531 , n24528 , n24530 );
buf ( n24532 , n19399 );
buf ( n24533 , n19244 );
nand ( n24534 , n24532 , n24533 );
buf ( n24535 , n24534 );
buf ( n24536 , n24535 );
nand ( n24537 , n24531 , n24536 );
buf ( n24538 , n24537 );
buf ( n24539 , n24538 );
xor ( n24540 , n18714 , n18747 );
and ( n24541 , n24540 , n18830 );
and ( n24542 , n18714 , n18747 );
or ( n24543 , n24541 , n24542 );
buf ( n24544 , n24543 );
buf ( n24545 , n24544 );
xor ( n24546 , n24539 , n24545 );
xor ( n24547 , n24214 , n24236 );
xor ( n24548 , n24547 , n24258 );
buf ( n24549 , n24548 );
buf ( n24550 , n24549 );
and ( n24551 , n24546 , n24550 );
and ( n24552 , n24539 , n24545 );
or ( n24553 , n24551 , n24552 );
buf ( n24554 , n24553 );
buf ( n24555 , n24554 );
xor ( n24556 , n24526 , n24555 );
buf ( n24557 , n24556 );
buf ( n24558 , n24557 );
xor ( n24559 , n24435 , n24558 );
buf ( n24560 , n24559 );
buf ( n24561 , n24560 );
xor ( n24562 , n24539 , n24545 );
xor ( n24563 , n24562 , n24550 );
buf ( n24564 , n24563 );
buf ( n24565 , n24564 );
xor ( n24566 , n19352 , n19418 );
and ( n24567 , n24566 , n19444 );
and ( n24568 , n19352 , n19418 );
or ( n24569 , n24567 , n24568 );
buf ( n24570 , n24569 );
buf ( n24571 , n24570 );
xor ( n24572 , n24565 , n24571 );
xor ( n24573 , n24371 , n24422 );
xor ( n24574 , n24573 , n24429 );
buf ( n24575 , n24574 );
buf ( n24576 , n24575 );
and ( n24577 , n24572 , n24576 );
and ( n24578 , n24565 , n24571 );
or ( n24579 , n24577 , n24578 );
buf ( n24580 , n24579 );
buf ( n24581 , n24580 );
or ( n24582 , n24561 , n24581 );
buf ( n24583 , n24582 );
buf ( n24584 , n24560 );
buf ( n24585 , n24580 );
nand ( n24586 , n24584 , n24585 );
buf ( n24587 , n24586 );
and ( n24588 , n24583 , n24587 );
buf ( n24589 , n24070 );
not ( n24590 , n24589 );
xor ( n24591 , n24565 , n24571 );
xor ( n24592 , n24591 , n24576 );
buf ( n24593 , n24592 );
not ( n24594 , n24593 );
xor ( n24595 , n18836 , n19345 );
and ( n24596 , n24595 , n19447 );
and ( n24597 , n18836 , n19345 );
or ( n24598 , n24596 , n24597 );
buf ( n24599 , n24598 );
not ( n24600 , n24599 );
and ( n24601 , n24594 , n24600 );
buf ( n24602 , n19449 );
buf ( n24603 , n19814 );
nor ( n24604 , n24602 , n24603 );
buf ( n24605 , n24604 );
nor ( n24606 , n24601 , n24605 );
and ( n24607 , n20370 , n24606 );
buf ( n24608 , n24607 );
not ( n24609 , n24608 );
or ( n24610 , n24590 , n24609 );
not ( n24611 , n24080 );
not ( n24612 , n24606 );
or ( n24613 , n24611 , n24612 );
buf ( n24614 , n24599 );
buf ( n24615 , n24593 );
nor ( n24616 , n24614 , n24615 );
buf ( n24617 , n24616 );
buf ( n24618 , n19449 );
buf ( n24619 , n19814 );
nand ( n24620 , n24618 , n24619 );
buf ( n24621 , n24620 );
nor ( n24622 , n24617 , n24621 );
buf ( n24623 , n24593 );
buf ( n24624 , n24599 );
and ( n24625 , n24623 , n24624 );
buf ( n24626 , n24625 );
nor ( n24627 , n24622 , n24626 );
nand ( n24628 , n24613 , n24627 );
buf ( n24629 , n24628 );
not ( n24630 , n24629 );
buf ( n24631 , n24630 );
buf ( n24632 , n24631 );
nand ( n24633 , n24610 , n24632 );
buf ( n24634 , n24633 );
buf ( n24635 , n24634 );
buf ( n24636 , n24635 );
buf ( n24637 , n24636 );
xor ( n24638 , n24588 , n24637 );
buf ( n24639 , n24638 );
xor ( n24640 , n24102 , n24103 );
xor ( n24641 , n24640 , n24639 );
buf ( n24642 , n24641 );
xor ( n24643 , n24102 , n24103 );
and ( n24644 , n24643 , n24639 );
and ( n24645 , n24102 , n24103 );
or ( n24646 , n24644 , n24645 );
buf ( n24647 , n24646 );
buf ( n24648 , n977 );
buf ( n24649 , n1235 );
not ( n24650 , n23619 );
not ( n24651 , n24650 );
buf ( n24652 , n23541 );
not ( n24653 , n24652 );
buf ( n24654 , n23537 );
nand ( n24655 , n24653 , n24654 );
buf ( n24656 , n24655 );
not ( n24657 , n24656 );
not ( n24658 , n24657 );
or ( n24659 , n24651 , n24658 );
nand ( n24660 , n23619 , n24656 );
nand ( n24661 , n24659 , n24660 );
buf ( n24662 , n24661 );
xor ( n24663 , n24648 , n24649 );
xor ( n24664 , n24663 , n24662 );
buf ( n24665 , n24664 );
xor ( n24666 , n24648 , n24649 );
and ( n24667 , n24666 , n24662 );
and ( n24668 , n24648 , n24649 );
or ( n24669 , n24667 , n24668 );
buf ( n24670 , n24669 );
buf ( n24671 , n1143 );
buf ( n24672 , n13678 );
buf ( n24673 , n23667 );
not ( n24674 , n24673 );
buf ( n24675 , n23671 );
nand ( n24676 , n24674 , n24675 );
buf ( n24677 , n24676 );
buf ( n24678 , n24677 );
not ( n24679 , n23621 );
buf ( n24680 , n24679 );
and ( n24681 , n24678 , n24680 );
not ( n24682 , n24678 );
buf ( n24683 , n24679 );
not ( n24684 , n24683 );
buf ( n24685 , n24684 );
buf ( n24686 , n24685 );
and ( n24687 , n24682 , n24686 );
nor ( n24688 , n24681 , n24687 );
buf ( n24689 , n24688 );
buf ( n24690 , n24689 );
xor ( n24691 , n24671 , n24672 );
xor ( n24692 , n24691 , n24690 );
buf ( n24693 , n24692 );
xor ( n24694 , n24671 , n24672 );
and ( n24695 , n24694 , n24690 );
and ( n24696 , n24671 , n24672 );
or ( n24697 , n24695 , n24696 );
buf ( n24698 , n24697 );
buf ( n24699 , n2057 );
buf ( n24700 , n13677 );
not ( n24701 , n23672 );
and ( n24702 , n23707 , n23715 );
not ( n24703 , n23707 );
buf ( n24704 , n23715 );
not ( n24705 , n24704 );
buf ( n24706 , n24705 );
and ( n24707 , n24703 , n24706 );
or ( n24708 , n24702 , n24707 );
not ( n24709 , n24708 );
not ( n24710 , n24709 );
or ( n24711 , n24701 , n24710 );
nand ( n24712 , n23675 , n24708 );
nand ( n24713 , n24711 , n24712 );
not ( n24714 , n24713 );
buf ( n24715 , n24714 );
xor ( n24716 , n24699 , n24700 );
xor ( n24717 , n24716 , n24715 );
buf ( n24718 , n24717 );
xor ( n24719 , n24699 , n24700 );
and ( n24720 , n24719 , n24715 );
and ( n24721 , n24699 , n24700 );
or ( n24722 , n24720 , n24721 );
buf ( n24723 , n24722 );
buf ( n24724 , n3534 );
buf ( n24725 , n13676 );
buf ( n24726 , n23727 );
not ( n24727 , n24726 );
buf ( n24728 , n23732 );
not ( n24729 , n24728 );
buf ( n24730 , n23740 );
nand ( n24731 , n24729 , n24730 );
buf ( n24732 , n24731 );
buf ( n24733 , n24732 );
buf ( n24734 , n23748 );
nand ( n24735 , n24733 , n24734 );
buf ( n24736 , n24735 );
buf ( n24737 , n24736 );
not ( n24738 , n24737 );
or ( n24739 , n24727 , n24738 );
buf ( n24740 , n23727 );
not ( n24741 , n24740 );
buf ( n24742 , n24736 );
not ( n24743 , n24742 );
buf ( n24744 , n24743 );
buf ( n24745 , n24744 );
nand ( n24746 , n24741 , n24745 );
buf ( n24747 , n24746 );
buf ( n24748 , n24747 );
nand ( n24749 , n24739 , n24748 );
buf ( n24750 , n24749 );
buf ( n24751 , n24750 );
xor ( n24752 , n24724 , n24725 );
xor ( n24753 , n24752 , n24751 );
buf ( n24754 , n24753 );
xor ( n24755 , n24724 , n24725 );
and ( n24756 , n24755 , n24751 );
and ( n24757 , n24724 , n24725 );
or ( n24758 , n24756 , n24757 );
buf ( n24759 , n24758 );
buf ( n24760 , n4151 );
buf ( n24761 , n24760 );
buf ( n24762 , n4138 );
buf ( n24763 , n23761 );
not ( n24764 , n24763 );
buf ( n24765 , n23828 );
buf ( n24766 , n23835 );
nand ( n24767 , n24765 , n24766 );
buf ( n24768 , n24767 );
buf ( n24769 , n24768 );
not ( n24770 , n24769 );
or ( n24771 , n24764 , n24770 );
buf ( n24772 , n24768 );
not ( n24773 , n24772 );
buf ( n24774 , n24773 );
buf ( n24775 , n24774 );
buf ( n24776 , n23761 );
not ( n24777 , n24776 );
buf ( n24778 , n24777 );
buf ( n24779 , n24778 );
nand ( n24780 , n24775 , n24779 );
buf ( n24781 , n24780 );
buf ( n24782 , n24781 );
nand ( n24783 , n24771 , n24782 );
buf ( n24784 , n24783 );
buf ( n24785 , n24784 );
xor ( n24786 , n24761 , n24762 );
xor ( n24787 , n24786 , n24785 );
buf ( n24788 , n24787 );
xor ( n24789 , n24761 , n24762 );
and ( n24790 , n24789 , n24785 );
and ( n24791 , n24761 , n24762 );
or ( n24792 , n24790 , n24791 );
buf ( n24793 , n24792 );
buf ( n24794 , n13684 );
buf ( n24795 , n4464 );
not ( n24796 , n23838 );
buf ( n24797 , n23874 );
buf ( n24798 , n23880 );
nand ( n24799 , n24797 , n24798 );
buf ( n24800 , n24799 );
not ( n24801 , n24800 );
or ( n24802 , n24796 , n24801 );
buf ( n24803 , n23838 );
not ( n24804 , n24803 );
buf ( n24805 , n24800 );
not ( n24806 , n24805 );
buf ( n24807 , n24806 );
buf ( n24808 , n24807 );
nand ( n24809 , n24804 , n24808 );
buf ( n24810 , n24809 );
nand ( n24811 , n24802 , n24810 );
buf ( n24812 , n24811 );
xor ( n24813 , n24794 , n24795 );
xor ( n24814 , n24813 , n24812 );
buf ( n24815 , n24814 );
xor ( n24816 , n24794 , n24795 );
and ( n24817 , n24816 , n24812 );
and ( n24818 , n24794 , n24795 );
or ( n24819 , n24817 , n24818 );
buf ( n24820 , n24819 );
buf ( n24821 , n5006 );
buf ( n24822 , n4993 );
buf ( n24823 , n23886 );
buf ( n24824 , n23893 );
nand ( n24825 , n24823 , n24824 );
buf ( n24826 , n24825 );
nand ( n24827 , n23899 , n24826 );
buf ( n24828 , n23881 );
not ( n24829 , n24828 );
and ( n24830 , n24827 , n24829 );
not ( n24831 , n24827 );
and ( n24832 , n24831 , n24828 );
nor ( n24833 , n24830 , n24832 );
not ( n24834 , n24833 );
not ( n24835 , n24834 );
buf ( n24836 , n24835 );
xor ( n24837 , n24821 , n24822 );
xor ( n24838 , n24837 , n24836 );
buf ( n24839 , n24838 );
xor ( n24840 , n24821 , n24822 );
and ( n24841 , n24840 , n24836 );
and ( n24842 , n24821 , n24822 );
or ( n24843 , n24841 , n24842 );
buf ( n24844 , n24843 );
buf ( n24845 , n15071 );
buf ( n24846 , n14910 );
buf ( n24847 , n24046 );
buf ( n24848 , n24847 );
buf ( n24849 , n24848 );
buf ( n24850 , n24849 );
buf ( n24851 , n24052 );
buf ( n24852 , n21364 );
nand ( n24853 , n24851 , n24852 );
buf ( n24854 , n24853 );
not ( n24855 , n24854 );
buf ( n24856 , n24855 );
and ( n24857 , n24850 , n24856 );
not ( n24858 , n24850 );
buf ( n24859 , n24854 );
and ( n24860 , n24858 , n24859 );
nor ( n24861 , n24857 , n24860 );
buf ( n24862 , n24861 );
buf ( n24863 , n24862 );
xor ( n24864 , n24845 , n24846 );
xor ( n24865 , n24864 , n24863 );
buf ( n24866 , n24865 );
xor ( n24867 , n24845 , n24846 );
and ( n24868 , n24867 , n24863 );
and ( n24869 , n24845 , n24846 );
or ( n24870 , n24868 , n24869 );
buf ( n24871 , n24870 );
buf ( n24872 , n8108 );
buf ( n24873 , n13673 );
buf ( n24874 , n23952 );
buf ( n24875 , n23958 );
or ( n24876 , n24874 , n24875 );
buf ( n24877 , n24876 );
buf ( n24878 , n24877 );
buf ( n24879 , n23972 );
nand ( n24880 , n24878 , n24879 );
buf ( n24881 , n24880 );
buf ( n24882 , n23948 );
xor ( n24883 , n24881 , n24882 );
not ( n24884 , n24883 );
not ( n24885 , n24884 );
buf ( n24886 , n24885 );
xor ( n24887 , n24872 , n24873 );
xor ( n24888 , n24887 , n24886 );
buf ( n24889 , n24888 );
xor ( n24890 , n24872 , n24873 );
and ( n24891 , n24890 , n24886 );
and ( n24892 , n24872 , n24873 );
or ( n24893 , n24891 , n24892 );
buf ( n24894 , n24893 );
buf ( n24895 , n13230 );
buf ( n24896 , n13217 );
not ( n24897 , n24013 );
not ( n24898 , n21997 );
or ( n24899 , n24897 , n24898 );
buf ( n24900 , n22003 );
buf ( n24901 , n24900 );
buf ( n24902 , n24901 );
nand ( n24903 , n24899 , n24902 );
not ( n24904 , n23997 );
buf ( n24905 , n23990 );
buf ( n24906 , n22228 );
buf ( n24907 , n22359 );
or ( n24908 , n24906 , n24907 );
buf ( n24909 , n24908 );
buf ( n24910 , n24909 );
nand ( n24911 , n24905 , n24910 );
buf ( n24912 , n24911 );
buf ( n24913 , n24912 );
not ( n24914 , n24913 );
buf ( n24915 , n24914 );
not ( n24916 , n24915 );
or ( n24917 , n24904 , n24916 );
buf ( n24918 , n23997 );
buf ( n24919 , n24009 );
nand ( n24920 , n24918 , n24919 );
buf ( n24921 , n24920 );
nand ( n24922 , n24917 , n24921 );
xor ( n24923 , n24903 , n24922 );
buf ( n24924 , n24923 );
not ( n24925 , n24924 );
buf ( n24926 , n24925 );
buf ( n24927 , n24926 );
xor ( n24928 , n24895 , n24896 );
xor ( n24929 , n24928 , n24927 );
buf ( n24930 , n24929 );
xor ( n24931 , n24895 , n24896 );
and ( n24932 , n24931 , n24927 );
and ( n24933 , n24895 , n24896 );
or ( n24934 , n24932 , n24933 );
buf ( n24935 , n24934 );
buf ( n24936 , n14021 );
buf ( n24937 , n14008 );
buf ( n24938 , n24015 );
not ( n24939 , n21638 );
not ( n24940 , n24939 );
not ( n24941 , n24033 );
and ( n24942 , n24940 , n24941 );
and ( n24943 , n24939 , n24033 );
nor ( n24944 , n24942 , n24943 );
and ( n24945 , n24938 , n24944 );
not ( n24946 , n24938 );
not ( n24947 , n24944 );
and ( n24948 , n24946 , n24947 );
nor ( n24949 , n24945 , n24948 );
not ( n24950 , n24949 );
not ( n24951 , n24950 );
buf ( n24952 , n24951 );
xor ( n24953 , n24936 , n24937 );
xor ( n24954 , n24953 , n24952 );
buf ( n24955 , n24954 );
xor ( n24956 , n24936 , n24937 );
and ( n24957 , n24956 , n24952 );
and ( n24958 , n24936 , n24937 );
or ( n24959 , n24957 , n24958 );
buf ( n24960 , n24959 );
buf ( n24961 , n13682 );
buf ( n24962 , n13674 );
buf ( n24963 , n22857 );
not ( n24964 , n24963 );
buf ( n24965 , n24964 );
buf ( n24966 , n24965 );
buf ( n24967 , n23926 );
nand ( n24968 , n24966 , n24967 );
buf ( n24969 , n24968 );
buf ( n24970 , n24969 );
buf ( n24971 , n22857 );
buf ( n24972 , n22972 );
nand ( n24973 , n24971 , n24972 );
buf ( n24974 , n24973 );
buf ( n24975 , n24974 );
nand ( n24976 , n24970 , n24975 );
buf ( n24977 , n24976 );
xnor ( n24978 , n23919 , n24977 );
buf ( n24979 , n24978 );
xor ( n24980 , n24961 , n24962 );
xor ( n24981 , n24980 , n24979 );
buf ( n24982 , n24981 );
xor ( n24983 , n24961 , n24962 );
and ( n24984 , n24983 , n24979 );
and ( n24985 , n24961 , n24962 );
or ( n24986 , n24984 , n24985 );
buf ( n24987 , n24986 );
buf ( n24988 , n14545 );
buf ( n24989 , n14701 );
buf ( n24990 , n24042 );
buf ( n24991 , n21634 );
nor ( n24992 , n24990 , n24991 );
buf ( n24993 , n24992 );
buf ( n24994 , n24993 );
not ( n24995 , n24994 );
nor ( n24996 , n24939 , n24033 );
not ( n24997 , n24996 );
nor ( n24998 , n21638 , n21797 );
not ( n24999 , n24998 );
nand ( n25000 , n24999 , n24938 );
nand ( n25001 , n24997 , n25000 );
buf ( n25002 , n25001 );
not ( n25003 , n25002 );
buf ( n25004 , n25003 );
not ( n25005 , n25004 );
or ( n25006 , n24995 , n25005 );
not ( n25007 , n24993 );
nand ( n25008 , n25007 , n25001 );
nand ( n25009 , n25006 , n25008 );
buf ( n25010 , n25009 );
buf ( n25011 , n25010 );
xor ( n25012 , n24988 , n24989 );
xor ( n25013 , n25012 , n25011 );
buf ( n25014 , n25013 );
xor ( n25015 , n24988 , n24989 );
and ( n25016 , n25015 , n25011 );
and ( n25017 , n24988 , n24989 );
or ( n25018 , n25016 , n25017 );
buf ( n25019 , n25018 );
buf ( n25020 , n15487 );
buf ( n25021 , n15623 );
buf ( n25022 , n24054 );
buf ( n25023 , n25022 );
or ( n25024 , n21102 , n20703 );
nand ( n25025 , n25024 , n24062 );
buf ( n25026 , n25025 );
xnor ( n25027 , n25023 , n25026 );
buf ( n25028 , n25027 );
buf ( n25029 , n25028 );
xor ( n25030 , n25020 , n25021 );
xor ( n25031 , n25030 , n25029 );
buf ( n25032 , n25031 );
xor ( n25033 , n25020 , n25021 );
and ( n25034 , n25033 , n25029 );
and ( n25035 , n25020 , n25021 );
or ( n25036 , n25034 , n25035 );
buf ( n25037 , n25036 );
buf ( n25038 , n16202 );
buf ( n25039 , n16415 );
buf ( n25040 , n24060 );
not ( n25041 , n25040 );
buf ( n25042 , n20375 );
buf ( n25043 , n20613 );
nand ( n25044 , n25042 , n25043 );
buf ( n25045 , n25044 );
buf ( n25046 , n25045 );
nand ( n25047 , n25041 , n25046 );
buf ( n25048 , n25047 );
not ( n25049 , n25048 );
not ( n25050 , n25049 );
nand ( n25051 , n24057 , n24058 );
buf ( n25052 , n25051 );
not ( n25053 , n25052 );
not ( n25054 , n21103 );
not ( n25055 , n25054 );
not ( n25056 , n24054 );
or ( n25057 , n25055 , n25056 );
buf ( n25058 , n24062 );
nand ( n25059 , n25057 , n25058 );
buf ( n25060 , n25059 );
not ( n25061 , n25060 );
or ( n25062 , n25053 , n25061 );
buf ( n25063 , n24065 );
nand ( n25064 , n25062 , n25063 );
buf ( n25065 , n25064 );
not ( n25066 , n25065 );
not ( n25067 , n25066 );
or ( n25068 , n25050 , n25067 );
nand ( n25069 , n25048 , n25065 );
nand ( n25070 , n25068 , n25069 );
buf ( n25071 , n25070 );
xor ( n25072 , n25038 , n25039 );
xor ( n25073 , n25072 , n25071 );
buf ( n25074 , n25073 );
xor ( n25075 , n25038 , n25039 );
and ( n25076 , n25075 , n25071 );
and ( n25077 , n25038 , n25039 );
or ( n25078 , n25076 , n25077 );
buf ( n25079 , n25078 );
buf ( n25080 , n16988 );
buf ( n25081 , n16917 );
or ( n25082 , n20366 , n20127 );
buf ( n25083 , n25082 );
not ( n25084 , n25083 );
buf ( n25085 , n24070 );
not ( n25086 , n25085 );
or ( n25087 , n25084 , n25086 );
buf ( n25088 , n24078 );
nand ( n25089 , n25087 , n25088 );
buf ( n25090 , n25089 );
not ( n25091 , n20123 );
xor ( n25092 , n19826 , n25091 );
and ( n25093 , n25090 , n25092 );
not ( n25094 , n25090 );
not ( n25095 , n25092 );
and ( n25096 , n25094 , n25095 );
nor ( n25097 , n25093 , n25096 );
not ( n25098 , n25097 );
buf ( n25099 , n25098 );
xor ( n25100 , n25080 , n25081 );
xor ( n25101 , n25100 , n25099 );
buf ( n25102 , n25101 );
xor ( n25103 , n25080 , n25081 );
and ( n25104 , n25103 , n25099 );
and ( n25105 , n25080 , n25081 );
or ( n25106 , n25104 , n25105 );
buf ( n25107 , n25106 );
buf ( n25108 , n1253 );
buf ( n25109 , n1336 );
buf ( n25110 , n1336 );
buf ( n25111 , n1253 );
or ( n25112 , n25110 , n25111 );
buf ( n25113 , n25112 );
buf ( n25114 , n25113 );
not ( n25115 , n25108 );
not ( n25116 , n25109 );
or ( n25117 , n25115 , n25116 );
nand ( n25118 , n25117 , n25114 );
buf ( n25119 , n25118 );
buf ( n25120 , n17951 );
buf ( n25121 , n17928 );
xor ( n25122 , n25120 , n25121 );
buf ( n25123 , n25122 );
xor ( n25124 , n17465 , n17424 );
buf ( n25125 , n24617 );
buf ( n25126 , n25125 );
buf ( n25127 , n24626 );
or ( n25128 , n25126 , n25127 );
buf ( n25129 , n25128 );
not ( n25130 , n25129 );
not ( n25131 , n19816 );
not ( n25132 , n24086 );
or ( n25133 , n25131 , n25132 );
nand ( n25134 , n25133 , n19820 );
not ( n25135 , n25134 );
not ( n25136 , n25135 );
or ( n25137 , n25130 , n25136 );
or ( n25138 , n25129 , n25135 );
nand ( n25139 , n25137 , n25138 );
not ( n25140 , n25139 );
xor ( n25141 , n25124 , n25140 );
buf ( n25142 , n25141 );
buf ( n25143 , n24101 );
xor ( n25144 , n25142 , n25143 );
buf ( n25145 , n25107 );
buf ( n25146 , n24096 );
xor ( n25147 , n25145 , n25146 );
buf ( n25148 , n25102 );
xor ( n25149 , n16543 , n16632 );
xor ( n25150 , n20366 , n20127 );
not ( n25151 , n25150 );
not ( n25152 , n25151 );
not ( n25153 , n24070 );
not ( n25154 , n25153 );
not ( n25155 , n25154 );
or ( n25156 , n25152 , n25155 );
nand ( n25157 , n25153 , n25150 );
nand ( n25158 , n25156 , n25157 );
buf ( n25159 , n25158 );
buf ( n25160 , n25159 );
and ( n25161 , n25149 , n25160 );
and ( n25162 , n16543 , n16632 );
or ( n25163 , n25161 , n25162 );
buf ( n25164 , n25163 );
xor ( n25165 , n25148 , n25164 );
buf ( n25166 , n25079 );
xor ( n25167 , n16543 , n16632 );
xor ( n25168 , n25167 , n25160 );
buf ( n25169 , n25168 );
xor ( n25170 , n25166 , n25169 );
buf ( n25171 , n16082 );
buf ( n25172 , n15815 );
xor ( n25173 , n25171 , n25172 );
and ( n25174 , n25051 , n24065 );
and ( n25175 , n25059 , n25174 );
not ( n25176 , n25059 );
not ( n25177 , n25174 );
and ( n25178 , n25176 , n25177 );
nor ( n25179 , n25175 , n25178 );
buf ( n25180 , n25179 );
not ( n25181 , n25180 );
not ( n25182 , n25181 );
not ( n25183 , n25182 );
not ( n25184 , n25183 );
buf ( n25185 , n25184 );
and ( n25186 , n25173 , n25185 );
and ( n25187 , n25171 , n25172 );
or ( n25188 , n25186 , n25187 );
buf ( n25189 , n25188 );
buf ( n25190 , n25189 );
buf ( n25191 , n25074 );
xor ( n25192 , n25190 , n25191 );
buf ( n25193 , n25037 );
xor ( n25194 , n25171 , n25172 );
xor ( n25195 , n25194 , n25185 );
buf ( n25196 , n25195 );
buf ( n25197 , n25196 );
xor ( n25198 , n25193 , n25197 );
buf ( n25199 , n24871 );
buf ( n25200 , n25032 );
xor ( n25201 , n25199 , n25200 );
buf ( n25202 , n25019 );
buf ( n25203 , n24866 );
xor ( n25204 , n25202 , n25203 );
buf ( n25205 , n25014 );
buf ( n25206 , n24960 );
xor ( n25207 , n25205 , n25206 );
buf ( n25208 , n24935 );
buf ( n25209 , n24955 );
xor ( n25210 , n25208 , n25209 );
buf ( n25211 , n10571 );
buf ( n25212 , n10554 );
xor ( n25213 , n25211 , n25212 );
buf ( n25214 , n24912 );
buf ( n25215 , n24006 );
nand ( n25216 , n25214 , n25215 );
buf ( n25217 , n25216 );
buf ( n25218 , n25217 );
buf ( n25219 , n23997 );
buf ( n25220 , n24001 );
and ( n25221 , n25219 , n25220 );
buf ( n25222 , n25221 );
buf ( n25223 , n25222 );
xor ( n25224 , n25218 , n25223 );
buf ( n25225 , n25224 );
buf ( n25226 , n25225 );
not ( n25227 , n25226 );
not ( n25228 , n25227 );
buf ( n25229 , n25228 );
and ( n25230 , n25213 , n25229 );
and ( n25231 , n25211 , n25212 );
or ( n25232 , n25230 , n25231 );
buf ( n25233 , n25232 );
buf ( n25234 , n25233 );
buf ( n25235 , n24930 );
xor ( n25236 , n25234 , n25235 );
buf ( n25237 , n9925 );
buf ( n25238 , n9894 );
xor ( n25239 , n25237 , n25238 );
buf ( n25240 , n23990 );
buf ( n25241 , n25240 );
buf ( n25242 , n25241 );
buf ( n25243 , n25242 );
buf ( n25244 , n24909 );
buf ( n25245 , n24006 );
nand ( n25246 , n25244 , n25245 );
buf ( n25247 , n25246 );
buf ( n25248 , n25247 );
not ( n25249 , n25248 );
buf ( n25250 , n25249 );
buf ( n25251 , n25250 );
and ( n25252 , n25243 , n25251 );
not ( n25253 , n25243 );
buf ( n25254 , n25247 );
and ( n25255 , n25253 , n25254 );
nor ( n25256 , n25252 , n25255 );
buf ( n25257 , n25256 );
buf ( n25258 , n25257 );
and ( n25259 , n25239 , n25258 );
and ( n25260 , n25237 , n25238 );
or ( n25261 , n25259 , n25260 );
buf ( n25262 , n25261 );
buf ( n25263 , n25262 );
xor ( n25264 , n25211 , n25212 );
xor ( n25265 , n25264 , n25229 );
buf ( n25266 , n25265 );
buf ( n25267 , n25266 );
xor ( n25268 , n25263 , n25267 );
xor ( n25269 , n25237 , n25238 );
xor ( n25270 , n25269 , n25258 );
buf ( n25271 , n25270 );
not ( n25272 , n9008 );
not ( n25273 , n9042 );
or ( n25274 , n25272 , n25273 );
buf ( n25275 , n23964 );
not ( n25276 , n25275 );
buf ( n25277 , n23972 );
nand ( n25278 , n25276 , n25277 );
buf ( n25279 , n25278 );
buf ( n25280 , n25279 );
buf ( n25281 , n22622 );
buf ( n25282 , n23981 );
and ( n25283 , n25281 , n25282 );
buf ( n25284 , n25283 );
buf ( n25285 , n25284 );
xor ( n25286 , n25280 , n25285 );
buf ( n25287 , n25286 );
buf ( n25288 , n25287 );
buf ( n25289 , n25288 );
buf ( n25290 , n25289 );
buf ( n25291 , n25290 );
not ( n25292 , n25291 );
buf ( n25293 , n25292 );
nor ( n25294 , n9008 , n9042 );
or ( n25295 , n25293 , n25294 );
nand ( n25296 , n25274 , n25295 );
or ( n25297 , n25271 , n25296 );
buf ( n25298 , n25297 );
not ( n25299 , n25298 );
xor ( n25300 , n9008 , n9042 );
buf ( n25301 , n25287 );
not ( n25302 , n25301 );
buf ( n25303 , n25302 );
buf ( n25304 , n25303 );
not ( n25305 , n25304 );
buf ( n25306 , n25305 );
and ( n25307 , n25300 , n25306 );
not ( n25308 , n25300 );
and ( n25309 , n25308 , n25293 );
nor ( n25310 , n25307 , n25309 );
buf ( n25311 , n25310 );
not ( n25312 , n25311 );
buf ( n25313 , n24894 );
not ( n25314 , n25313 );
buf ( n25315 , n25314 );
buf ( n25316 , n25315 );
nand ( n25317 , n25312 , n25316 );
buf ( n25318 , n25317 );
buf ( n25319 , n25318 );
not ( n25320 , n25319 );
buf ( n25321 , n24889 );
not ( n25322 , n25321 );
buf ( n25323 , n6674 );
xor ( n25324 , n6659 , n25323 );
not ( n25325 , n24969 );
not ( n25326 , n23919 );
or ( n25327 , n25325 , n25326 );
nand ( n25328 , n25327 , n24974 );
not ( n25329 , n25328 );
not ( n25330 , n25329 );
xnor ( n25331 , n22852 , n22825 );
not ( n25332 , n25331 );
not ( n25333 , n25332 );
or ( n25334 , n25330 , n25333 );
nand ( n25335 , n25331 , n25328 );
nand ( n25336 , n25334 , n25335 );
and ( n25337 , n25324 , n25336 );
and ( n25338 , n6659 , n25323 );
or ( n25339 , n25337 , n25338 );
buf ( n25340 , n25339 );
not ( n25341 , n25340 );
buf ( n25342 , n25341 );
buf ( n25343 , n25342 );
nand ( n25344 , n25322 , n25343 );
buf ( n25345 , n25344 );
buf ( n25346 , n25345 );
not ( n25347 , n25346 );
xor ( n25348 , n6659 , n25323 );
xor ( n25349 , n25348 , n25336 );
buf ( n25350 , n25349 );
buf ( n25351 , n24987 );
or ( n25352 , n25350 , n25351 );
buf ( n25353 , n25352 );
buf ( n25354 , n25353 );
not ( n25355 , n25354 );
buf ( n25356 , n24982 );
buf ( n25357 , n13683 );
buf ( n25358 , n6408 );
xor ( n25359 , n25357 , n25358 );
buf ( n25360 , n23914 );
not ( n25361 , n25360 );
buf ( n25362 , n25361 );
buf ( n25363 , n25362 );
buf ( n25364 , n23162 );
nand ( n25365 , n25363 , n25364 );
buf ( n25366 , n25365 );
nand ( n25367 , n25366 , n23918 );
not ( n25368 , n25367 );
not ( n25369 , n25368 );
buf ( n25370 , n23909 );
buf ( n25371 , n25370 );
buf ( n25372 , n25371 );
buf ( n25373 , n25372 );
not ( n25374 , n25373 );
buf ( n25375 , n25374 );
not ( n25376 , n25375 );
or ( n25377 , n25369 , n25376 );
nand ( n25378 , n25367 , n25372 );
nand ( n25379 , n25377 , n25378 );
buf ( n25380 , n25379 );
not ( n25381 , n25380 );
buf ( n25382 , n25381 );
buf ( n25383 , n25382 );
not ( n25384 , n25383 );
buf ( n25385 , n25384 );
buf ( n25386 , n25385 );
and ( n25387 , n25359 , n25386 );
and ( n25388 , n25357 , n25358 );
or ( n25389 , n25387 , n25388 );
buf ( n25390 , n25389 );
buf ( n25391 , n25390 );
or ( n25392 , n25356 , n25391 );
buf ( n25393 , n25392 );
buf ( n25394 , n25393 );
not ( n25395 , n25394 );
xor ( n25396 , n25357 , n25358 );
xor ( n25397 , n25396 , n25386 );
buf ( n25398 , n25397 );
not ( n25399 , n25398 );
not ( n25400 , n24844 );
nand ( n25401 , n25399 , n25400 );
not ( n25402 , n25401 );
not ( n25403 , n24820 );
not ( n25404 , n25403 );
not ( n25405 , n24839 );
not ( n25406 , n25405 );
or ( n25407 , n25404 , n25406 );
buf ( n25408 , n24815 );
buf ( n25409 , n24793 );
nor ( n25410 , n25408 , n25409 );
buf ( n25411 , n25410 );
buf ( n25412 , n25411 );
buf ( n25413 , n24788 );
buf ( n25414 , n3865 );
buf ( n25415 , n3842 );
xor ( n25416 , n25414 , n25415 );
buf ( n25417 , n23421 );
buf ( n25418 , n23758 );
nand ( n25419 , n25417 , n25418 );
buf ( n25420 , n25419 );
buf ( n25421 , n25420 );
buf ( n25422 , n23751 );
not ( n25423 , n25422 );
buf ( n25424 , n25423 );
buf ( n25425 , n25424 );
and ( n25426 , n25421 , n25425 );
not ( n25427 , n25421 );
buf ( n25428 , n23751 );
and ( n25429 , n25427 , n25428 );
nor ( n25430 , n25426 , n25429 );
buf ( n25431 , n25430 );
buf ( n25432 , n25431 );
and ( n25433 , n25416 , n25432 );
and ( n25434 , n25414 , n25415 );
or ( n25435 , n25433 , n25434 );
buf ( n25436 , n25435 );
buf ( n25437 , n25436 );
or ( n25438 , n25413 , n25437 );
buf ( n25439 , n25438 );
not ( n25440 , n25439 );
buf ( n25441 , n24759 );
xor ( n25442 , n25414 , n25415 );
xor ( n25443 , n25442 , n25432 );
buf ( n25444 , n25443 );
buf ( n25445 , n25444 );
xor ( n25446 , n25441 , n25445 );
xor ( n25447 , n24718 , n24698 );
xor ( n25448 , n24693 , n24670 );
buf ( n25449 , n24665 );
not ( n25450 , n25449 );
buf ( n25451 , n25450 );
buf ( n25452 , n25451 );
buf ( n25453 , n25113 );
not ( n25454 , n25453 );
buf ( n25455 , n25454 );
buf ( n25456 , n25455 );
nand ( n25457 , n25452 , n25456 );
buf ( n25458 , n25457 );
not ( n25459 , n1479 );
buf ( n25460 , n25459 );
buf ( n25461 , n1558 );
and ( n25462 , n25460 , n25461 );
buf ( n25463 , n25462 );
buf ( n25464 , n25463 );
buf ( n25465 , n1482 );
or ( n25466 , n25464 , n25465 );
xor ( n25467 , n1324 , n1407 );
buf ( n25468 , n25467 );
nand ( n25469 , n25466 , n25468 );
buf ( n25470 , n25469 );
buf ( n25471 , n25470 );
not ( n25472 , n25471 );
buf ( n25473 , n25472 );
buf ( n25474 , n25473 );
and ( n25475 , n1324 , n1407 );
buf ( n25476 , n25475 );
xor ( n25477 , n25474 , n25476 );
buf ( n25478 , n25119 );
and ( n25479 , n25477 , n25478 );
or ( n25480 , n25479 , C0 );
buf ( n25481 , n25480 );
and ( n25482 , n25458 , n25481 );
buf ( n25483 , n25451 );
buf ( n25484 , n25455 );
nor ( n25485 , n25483 , n25484 );
buf ( n25486 , n25485 );
nor ( n25487 , n25482 , n25486 );
not ( n25488 , n25487 );
and ( n25489 , n25448 , n25488 );
and ( n25490 , n24693 , n24670 );
or ( n25491 , n25489 , n25490 );
and ( n25492 , n25447 , n25491 );
and ( n25493 , n24718 , n24698 );
nor ( n25494 , n25492 , n25493 );
buf ( n25495 , n25494 );
buf ( n25496 , n24754 );
buf ( n25497 , n24723 );
nor ( n25498 , n25496 , n25497 );
buf ( n25499 , n25498 );
buf ( n25500 , n25499 );
or ( n25501 , n25495 , n25500 );
buf ( n25502 , n24754 );
buf ( n25503 , n24723 );
nand ( n25504 , n25502 , n25503 );
buf ( n25505 , n25504 );
buf ( n25506 , n25505 );
nand ( n25507 , n25501 , n25506 );
buf ( n25508 , n25507 );
buf ( n25509 , n25508 );
and ( n25510 , n25446 , n25509 );
and ( n25511 , n25441 , n25445 );
or ( n25512 , n25510 , n25511 );
buf ( n25513 , n25512 );
not ( n25514 , n25513 );
or ( n25515 , n25440 , n25514 );
nand ( n25516 , n24788 , n25436 );
nand ( n25517 , n25515 , n25516 );
not ( n25518 , n25517 );
buf ( n25519 , n25518 );
or ( n25520 , n25412 , n25519 );
buf ( n25521 , n24815 );
buf ( n25522 , n24793 );
nand ( n25523 , n25521 , n25522 );
buf ( n25524 , n25523 );
buf ( n25525 , n25524 );
nand ( n25526 , n25520 , n25525 );
buf ( n25527 , n25526 );
nand ( n25528 , n25407 , n25527 );
nand ( n25529 , n24839 , n24820 );
nand ( n25530 , n25528 , n25529 );
not ( n25531 , n25530 );
or ( n25532 , n25402 , n25531 );
nand ( n25533 , n25398 , n24844 );
nand ( n25534 , n25532 , n25533 );
buf ( n25535 , n25534 );
not ( n25536 , n25535 );
or ( n25537 , n25395 , n25536 );
buf ( n25538 , n24982 );
buf ( n25539 , n25390 );
nand ( n25540 , n25538 , n25539 );
buf ( n25541 , n25540 );
buf ( n25542 , n25541 );
nand ( n25543 , n25537 , n25542 );
buf ( n25544 , n25543 );
buf ( n25545 , n25544 );
not ( n25546 , n25545 );
or ( n25547 , n25355 , n25546 );
buf ( n25548 , n25349 );
buf ( n25549 , n24987 );
nand ( n25550 , n25548 , n25549 );
buf ( n25551 , n25550 );
buf ( n25552 , n25551 );
nand ( n25553 , n25547 , n25552 );
buf ( n25554 , n25553 );
buf ( n25555 , n25554 );
not ( n25556 , n25555 );
or ( n25557 , n25347 , n25556 );
buf ( n25558 , n24889 );
buf ( n25559 , n25339 );
nand ( n25560 , n25558 , n25559 );
buf ( n25561 , n25560 );
buf ( n25562 , n25561 );
nand ( n25563 , n25557 , n25562 );
buf ( n25564 , n25563 );
buf ( n25565 , n25564 );
not ( n25566 , n25565 );
or ( n25567 , n25320 , n25566 );
buf ( n25568 , n25310 );
buf ( n25569 , n24894 );
nand ( n25570 , n25568 , n25569 );
buf ( n25571 , n25570 );
buf ( n25572 , n25571 );
nand ( n25573 , n25567 , n25572 );
buf ( n25574 , n25573 );
buf ( n25575 , n25574 );
not ( n25576 , n25575 );
or ( n25577 , n25299 , n25576 );
buf ( n25578 , n25271 );
buf ( n25579 , n25296 );
nand ( n25580 , n25578 , n25579 );
buf ( n25581 , n25580 );
buf ( n25582 , n25581 );
nand ( n25583 , n25577 , n25582 );
buf ( n25584 , n25583 );
buf ( n25585 , n25584 );
and ( n25586 , n25268 , n25585 );
and ( n25587 , n25263 , n25267 );
or ( n25588 , n25586 , n25587 );
buf ( n25589 , n25588 );
buf ( n25590 , n25589 );
and ( n25591 , n25236 , n25590 );
and ( n25592 , n25234 , n25235 );
or ( n25593 , n25591 , n25592 );
buf ( n25594 , n25593 );
buf ( n25595 , n25594 );
and ( n25596 , n25210 , n25595 );
and ( n25597 , n25208 , n25209 );
or ( n25598 , n25596 , n25597 );
buf ( n25599 , n25598 );
buf ( n25600 , n25599 );
and ( n25601 , n25207 , n25600 );
and ( n25602 , n25205 , n25206 );
or ( n25603 , n25601 , n25602 );
buf ( n25604 , n25603 );
buf ( n25605 , n25604 );
and ( n25606 , n25204 , n25605 );
and ( n25607 , n25202 , n25203 );
or ( n25608 , n25606 , n25607 );
buf ( n25609 , n25608 );
buf ( n25610 , n25609 );
and ( n25611 , n25201 , n25610 );
and ( n25612 , n25199 , n25200 );
or ( n25613 , n25611 , n25612 );
buf ( n25614 , n25613 );
buf ( n25615 , n25614 );
and ( n25616 , n25198 , n25615 );
and ( n25617 , n25193 , n25197 );
or ( n25618 , n25616 , n25617 );
buf ( n25619 , n25618 );
buf ( n25620 , n25619 );
and ( n25621 , n25192 , n25620 );
and ( n25622 , n25190 , n25191 );
or ( n25623 , n25621 , n25622 );
buf ( n25624 , n25623 );
buf ( n25625 , n25624 );
and ( n25626 , n25170 , n25625 );
and ( n25627 , n25166 , n25169 );
or ( n25628 , n25626 , n25627 );
buf ( n25629 , n25628 );
buf ( n25630 , n25629 );
and ( n25631 , n25165 , n25630 );
and ( n25632 , n25148 , n25164 );
or ( n25633 , n25631 , n25632 );
buf ( n25634 , n25633 );
buf ( n25635 , n25634 );
and ( n25636 , n25147 , n25635 );
and ( n25637 , n25145 , n25146 );
or ( n25638 , n25636 , n25637 );
buf ( n25639 , n25638 );
buf ( n25640 , n25639 );
and ( n25641 , n25144 , n25640 );
and ( n25642 , n25142 , n25143 );
or ( n25643 , n25641 , n25642 );
buf ( n25644 , n25643 );
buf ( n25645 , n25644 );
buf ( n25646 , n24642 );
not ( n25647 , n25646 );
buf ( n25648 , n25647 );
buf ( n25649 , n25648 );
xor ( n25650 , n17465 , n17424 );
and ( n25651 , n25650 , n25140 );
and ( n25652 , n17465 , n17424 );
or ( n25653 , n25651 , n25652 );
buf ( n25654 , n25653 );
not ( n25655 , n25654 );
buf ( n25656 , n25655 );
buf ( n25657 , n25656 );
nand ( n25658 , n25649 , n25657 );
buf ( n25659 , n25658 );
buf ( n25660 , n25659 );
and ( n25661 , n25645 , n25660 );
buf ( n25662 , n25648 );
buf ( n25663 , n25656 );
nor ( n25664 , n25662 , n25663 );
buf ( n25665 , n25664 );
buf ( n25666 , n25665 );
nor ( n25667 , n25661 , n25666 );
buf ( n25668 , n25667 );
buf ( n25669 , n25668 );
buf ( n25670 , n25644 );
not ( n25671 , n25670 );
buf ( n25672 , n25665 );
not ( n25673 , n25672 );
and ( n25674 , n25671 , n25673 );
buf ( n25675 , n25659 );
not ( n25676 , n25675 );
buf ( n25677 , n25676 );
buf ( n25678 , n25677 );
nor ( n25679 , n25674 , n25678 );
buf ( n25680 , n25679 );
buf ( n25681 , n25680 );
buf ( n25682 , n24647 );
buf ( n25683 , n25123 );
xor ( n25684 , n25682 , n25683 );
buf ( n25685 , n25684 );
buf ( n25686 , n25685 );
and ( n25687 , n25686 , n25681 );
not ( n25688 , n25686 );
and ( n25689 , n25688 , n25669 );
nor ( n25690 , n25687 , n25689 );
buf ( n25691 , n25690 );
buf ( n25692 , n25656 );
buf ( n25693 , n24642 );
and ( n25694 , n25692 , n25693 );
not ( n25695 , n25692 );
buf ( n25696 , n25648 );
and ( n25697 , n25695 , n25696 );
nor ( n25698 , n25694 , n25697 );
buf ( n25699 , n25698 );
buf ( n25700 , n25699 );
buf ( n25701 , n25644 );
buf ( n25702 , n25699 );
buf ( n25703 , n25644 );
not ( n25704 , n25700 );
not ( n25705 , n25701 );
or ( n25706 , n25704 , n25705 );
or ( n25707 , n25702 , n25703 );
nand ( n25708 , n25706 , n25707 );
buf ( n25709 , n25708 );
xor ( n25710 , n25142 , n25143 );
xor ( n25711 , n25710 , n25640 );
buf ( n25712 , n25711 );
xor ( n25713 , n25145 , n25146 );
xor ( n25714 , n25713 , n25635 );
buf ( n25715 , n25714 );
xor ( n25716 , n25148 , n25164 );
xor ( n25717 , n25716 , n25630 );
buf ( n25718 , n25717 );
xor ( n25719 , n25166 , n25169 );
xor ( n25720 , n25719 , n25625 );
buf ( n25721 , n25720 );
xor ( n25722 , n25190 , n25191 );
xor ( n25723 , n25722 , n25620 );
buf ( n25724 , n25723 );
xor ( n25725 , n25193 , n25197 );
xor ( n25726 , n25725 , n25615 );
buf ( n25727 , n25726 );
xor ( n25728 , n25199 , n25200 );
xor ( n25729 , n25728 , n25610 );
buf ( n25730 , n25729 );
xor ( n25731 , n25202 , n25203 );
xor ( n25732 , n25731 , n25605 );
buf ( n25733 , n25732 );
xor ( n25734 , n25205 , n25206 );
xor ( n25735 , n25734 , n25600 );
buf ( n25736 , n25735 );
xor ( n25737 , n25208 , n25209 );
xor ( n25738 , n25737 , n25595 );
buf ( n25739 , n25738 );
xor ( n25740 , n25234 , n25235 );
xor ( n25741 , n25740 , n25590 );
buf ( n25742 , n25741 );
xor ( n25743 , n25263 , n25267 );
xor ( n25744 , n25743 , n25585 );
buf ( n25745 , n25744 );
buf ( n25746 , n25574 );
buf ( n25747 , n25271 );
buf ( n25748 , n25296 );
xnor ( n25749 , n25747 , n25748 );
buf ( n25750 , n25749 );
buf ( n25751 , n25750 );
buf ( n25752 , n25750 );
buf ( n25753 , n25574 );
not ( n25754 , n25746 );
not ( n25755 , n25751 );
or ( n25756 , n25754 , n25755 );
or ( n25757 , n25752 , n25753 );
nand ( n25758 , n25756 , n25757 );
buf ( n25759 , n25758 );
buf ( n25760 , n25564 );
and ( n25761 , n25310 , n25315 );
not ( n25762 , n25310 );
and ( n25763 , n25762 , n24894 );
nor ( n25764 , n25761 , n25763 );
buf ( n25765 , n25764 );
buf ( n25766 , n25764 );
buf ( n25767 , n25564 );
not ( n25768 , n25760 );
not ( n25769 , n25765 );
or ( n25770 , n25768 , n25769 );
or ( n25771 , n25766 , n25767 );
nand ( n25772 , n25770 , n25771 );
buf ( n25773 , n25772 );
buf ( n25774 , n25554 );
buf ( n25775 , n24889 );
buf ( n25776 , n25339 );
xnor ( n25777 , n25775 , n25776 );
buf ( n25778 , n25777 );
buf ( n25779 , n25778 );
buf ( n25780 , n25778 );
buf ( n25781 , n25554 );
not ( n25782 , n25774 );
not ( n25783 , n25779 );
or ( n25784 , n25782 , n25783 );
or ( n25785 , n25780 , n25781 );
nand ( n25786 , n25784 , n25785 );
buf ( n25787 , n25786 );
buf ( n25788 , n25544 );
buf ( n25789 , n25349 );
buf ( n25790 , n24987 );
xor ( n25791 , n25789 , n25790 );
buf ( n25792 , n25791 );
buf ( n25793 , n25792 );
xor ( n25794 , n25788 , n25793 );
buf ( n25795 , n25794 );
buf ( n25796 , n25534 );
buf ( n25797 , n24982 );
buf ( n25798 , n25390 );
xor ( n25799 , n25797 , n25798 );
buf ( n25800 , n25799 );
buf ( n25801 , n25800 );
xor ( n25802 , n25796 , n25801 );
buf ( n25803 , n25802 );
buf ( n25804 , n25518 );
buf ( n25805 , n25517 );
buf ( n25806 , n24815 );
buf ( n25807 , n24793 );
xor ( n25808 , n25806 , n25807 );
buf ( n25809 , n25808 );
buf ( n25810 , n25809 );
and ( n25811 , n25810 , n25805 );
not ( n25812 , n25810 );
and ( n25813 , n25812 , n25804 );
nor ( n25814 , n25811 , n25813 );
buf ( n25815 , n25814 );
buf ( n25816 , n25513 );
buf ( n25817 , n24788 );
buf ( n25818 , n25436 );
xor ( n25819 , n25817 , n25818 );
buf ( n25820 , n25819 );
buf ( n25821 , n25820 );
xor ( n25822 , n25816 , n25821 );
buf ( n25823 , n25822 );
xor ( n25824 , n25441 , n25445 );
xor ( n25825 , n25824 , n25509 );
buf ( n25826 , n25825 );
buf ( n25827 , n24665 );
buf ( n25828 , n25113 );
xor ( n25829 , n25827 , n25828 );
buf ( n25830 , n25829 );
buf ( n25831 , n25830 );
buf ( n25832 , n25481 );
xor ( n25833 , n25831 , n25832 );
buf ( n25834 , n25833 );
xor ( n25835 , n25474 , n25476 );
xor ( n25836 , n25835 , n25478 );
buf ( n25837 , n25836 );
buf ( n25838 , n25463 );
not ( n25839 , n1407 );
and ( n25840 , n1324 , n1482 );
not ( n25841 , n1324 );
and ( n25842 , n25841 , n25459 );
nor ( n25843 , n25840 , n25842 );
not ( n25844 , n25843 );
or ( n25845 , n25839 , n25844 );
or ( n25846 , n1407 , n25843 );
nand ( n25847 , n25845 , n25846 );
buf ( n25848 , n25847 );
buf ( n25849 , n25463 );
buf ( n25850 , n25847 );
not ( n25851 , n25838 );
not ( n25852 , n25848 );
or ( n25853 , n25851 , n25852 );
or ( n25854 , n25849 , n25850 );
nand ( n25855 , n25853 , n25854 );
buf ( n25856 , n25855 );
xor ( n25857 , n25460 , n25461 );
buf ( n25858 , n25857 );
buf ( n25859 , n24839 );
buf ( n25860 , n24820 );
xor ( n25861 , n25859 , n25860 );
buf ( n25862 , n25861 );
buf ( n25863 , n25398 );
buf ( n25864 , n24844 );
xor ( n25865 , n25863 , n25864 );
buf ( n25866 , n25865 );
buf ( n25867 , n24754 );
buf ( n25868 , n24723 );
xor ( n25869 , n25867 , n25868 );
buf ( n25870 , n25869 );
buf ( n25871 , n25494 );
buf ( n25872 , n25870 );
xnor ( n25873 , n25871 , n25872 );
buf ( n25874 , n25873 );
buf ( n25875 , n1021 );
buf ( n25876 , n13675 );
xor ( n25877 , n12423 , n12427 );
xor ( n25878 , n25877 , n12550 );
buf ( n25879 , n25878 );
buf ( n25880 , n25879 );
xor ( n25881 , n25875 , n25876 );
xor ( n25882 , n25881 , n25880 );
buf ( n25883 , n25882 );
xor ( n25884 , n25875 , n25876 );
and ( n25885 , n25884 , n25880 );
and ( n25886 , n25875 , n25876 );
or ( n25887 , n25885 , n25886 );
buf ( n25888 , n25887 );
buf ( n25889 , n1097 );
buf ( n25890 , n13680 );
nor ( n25891 , n12408 , n12378 );
not ( n25892 , n12554 );
nand ( n25893 , n25891 , n25892 );
not ( n25894 , n12409 );
nand ( n25895 , n25894 , n12554 );
not ( n25896 , n12378 );
nor ( n25897 , n25896 , n12407 );
nand ( n25898 , n25892 , n25897 );
nand ( n25899 , n12556 , n12554 );
nand ( n25900 , n25893 , n25895 , n25898 , n25899 );
buf ( n25901 , n25900 );
xor ( n25902 , n25889 , n25890 );
xor ( n25903 , n25902 , n25901 );
buf ( n25904 , n25903 );
xor ( n25905 , n25889 , n25890 );
and ( n25906 , n25905 , n25901 );
and ( n25907 , n25889 , n25890 );
or ( n25908 , n25906 , n25907 );
buf ( n25909 , n25908 );
buf ( n25910 , n2062 );
buf ( n25911 , n13667 );
buf ( n25912 , n12573 );
not ( n25913 , n25912 );
buf ( n25914 , n12579 );
nand ( n25915 , n25913 , n25914 );
buf ( n25916 , n25915 );
buf ( n25917 , n25916 );
buf ( n25918 , n12557 );
and ( n25919 , n25917 , n25918 );
not ( n25920 , n25917 );
not ( n25921 , n12557 );
buf ( n25922 , n25921 );
and ( n25923 , n25920 , n25922 );
nor ( n25924 , n25919 , n25923 );
buf ( n25925 , n25924 );
buf ( n25926 , n25925 );
xor ( n25927 , n25910 , n25911 );
xor ( n25928 , n25927 , n25926 );
buf ( n25929 , n25928 );
xor ( n25930 , n25910 , n25911 );
and ( n25931 , n25930 , n25926 );
and ( n25932 , n25910 , n25911 );
or ( n25933 , n25931 , n25932 );
buf ( n25934 , n25933 );
buf ( n25935 , n3550 );
buf ( n25936 , n13681 );
xor ( n25937 , n12371 , n12374 );
xor ( n25938 , n25937 , n12582 );
buf ( n25939 , n25938 );
xor ( n25940 , n25935 , n25936 );
xor ( n25941 , n25940 , n25939 );
buf ( n25942 , n25941 );
xor ( n25943 , n25935 , n25936 );
and ( n25944 , n25943 , n25939 );
and ( n25945 , n25935 , n25936 );
or ( n25946 , n25944 , n25945 );
buf ( n25947 , n25946 );
buf ( n25948 , n3871 );
buf ( n25949 , n13672 );
xor ( n25950 , n12191 , n12194 );
xor ( n25951 , n25950 , n12585 );
buf ( n25952 , n25951 );
xor ( n25953 , n25948 , n25949 );
xor ( n25954 , n25953 , n25952 );
buf ( n25955 , n25954 );
xor ( n25956 , n25948 , n25949 );
and ( n25957 , n25956 , n25952 );
and ( n25958 , n25948 , n25949 );
or ( n25959 , n25957 , n25958 );
buf ( n25960 , n25959 );
buf ( n25961 , n4157 );
buf ( n25962 , n13685 );
buf ( n25963 , n12146 );
buf ( n25964 , n12594 );
nand ( n25965 , n25963 , n25964 );
buf ( n25966 , n25965 );
buf ( n25967 , n25966 );
not ( n25968 , n25967 );
buf ( n25969 , n12588 );
not ( n25970 , n25969 );
or ( n25971 , n25968 , n25970 );
not ( n25972 , n25966 );
not ( n25973 , n12588 );
nand ( n25974 , n25972 , n25973 );
buf ( n25975 , n25974 );
nand ( n25976 , n25971 , n25975 );
buf ( n25977 , n25976 );
buf ( n25978 , n25977 );
xor ( n25979 , n25961 , n25962 );
xor ( n25980 , n25979 , n25978 );
buf ( n25981 , n25980 );
xor ( n25982 , n25961 , n25962 );
and ( n25983 , n25982 , n25978 );
and ( n25984 , n25961 , n25962 );
or ( n25985 , n25983 , n25984 );
buf ( n25986 , n25985 );
buf ( n25987 , n4483 );
buf ( n25988 , n13671 );
not ( n25989 , n12666 );
not ( n25990 , n12602 );
or ( n25991 , n25989 , n25990 );
nand ( n25992 , n25991 , n12670 );
not ( n25993 , n25992 );
not ( n25994 , n12595 );
or ( n25995 , n25993 , n25994 );
or ( n25996 , n12595 , n25992 );
nand ( n25997 , n25995 , n25996 );
buf ( n25998 , n25997 );
xor ( n25999 , n25987 , n25988 );
xor ( n26000 , n25999 , n25998 );
buf ( n26001 , n26000 );
xor ( n26002 , n25987 , n25988 );
and ( n26003 , n26002 , n25998 );
and ( n26004 , n25987 , n25988 );
or ( n26005 , n26003 , n26004 );
buf ( n26006 , n26005 );
buf ( n26007 , n5012 );
buf ( n26008 , n13670 );
buf ( n26009 , n12681 );
not ( n26010 , n26009 );
buf ( n26011 , n12709 );
buf ( n26012 , n12715 );
nor ( n26013 , n26011 , n26012 );
buf ( n26014 , n26013 );
buf ( n26015 , n26014 );
not ( n26016 , n26015 );
buf ( n26017 , n12728 );
nand ( n26018 , n26016 , n26017 );
buf ( n26019 , n26018 );
buf ( n26020 , n26019 );
not ( n26021 , n26020 );
or ( n26022 , n26010 , n26021 );
buf ( n26023 , n12681 );
not ( n26024 , n26023 );
buf ( n26025 , n26019 );
not ( n26026 , n26025 );
buf ( n26027 , n26026 );
buf ( n26028 , n26027 );
nand ( n26029 , n26024 , n26028 );
buf ( n26030 , n26029 );
buf ( n26031 , n26030 );
nand ( n26032 , n26022 , n26031 );
buf ( n26033 , n26032 );
buf ( n26034 , n26033 );
xor ( n26035 , n26007 , n26008 );
xor ( n26036 , n26035 , n26034 );
buf ( n26037 , n26036 );
xor ( n26038 , n26007 , n26008 );
and ( n26039 , n26038 , n26034 );
and ( n26040 , n26007 , n26008 );
or ( n26041 , n26039 , n26040 );
buf ( n26042 , n26041 );
buf ( n26043 , n16703 );
buf ( n26044 , n16710 );
buf ( n26045 , n10882 );
not ( n26046 , n26045 );
buf ( n26047 , n606 );
not ( n26048 , n26047 );
or ( n26049 , n18194 , n24218 );
not ( n26050 , n18193 );
nand ( n26051 , n26050 , n24218 );
nand ( n26052 , n26049 , n26051 );
buf ( n26053 , n26052 );
buf ( n26054 , n26053 );
not ( n26055 , n26054 );
buf ( n26056 , n26055 );
buf ( n26057 , n26056 );
not ( n26058 , n26057 );
or ( n26059 , n26048 , n26058 );
buf ( n26060 , n26053 );
not ( n26061 , n26060 );
buf ( n26062 , n26061 );
buf ( n26063 , n26062 );
not ( n26064 , n26063 );
buf ( n26065 , n26064 );
buf ( n26066 , n26065 );
buf ( n26067 , n10836 );
nand ( n26068 , n26066 , n26067 );
buf ( n26069 , n26068 );
buf ( n26070 , n26069 );
nand ( n26071 , n26059 , n26070 );
buf ( n26072 , n26071 );
buf ( n26073 , n26072 );
not ( n26074 , n26073 );
or ( n26075 , n26046 , n26074 );
buf ( n26076 , n606 );
not ( n26077 , n26076 );
not ( n26078 , n24327 );
nand ( n26079 , n15682 , n9517 , n18082 );
not ( n26080 , n26079 );
or ( n26081 , n26078 , n26080 );
not ( n26082 , n9517 );
nor ( n26083 , n18137 , n26082 );
nand ( n26084 , n15682 , n26083 , n18082 );
nand ( n26085 , n26081 , n26084 );
buf ( n26086 , n26085 );
not ( n26087 , n26086 );
buf ( n26088 , n26087 );
buf ( n26089 , n26088 );
not ( n26090 , n26089 );
or ( n26091 , n26077 , n26090 );
buf ( n26092 , n26088 );
not ( n26093 , n26092 );
buf ( n26094 , n26093 );
buf ( n26095 , n26094 );
buf ( n26096 , n10836 );
nand ( n26097 , n26095 , n26096 );
buf ( n26098 , n26097 );
buf ( n26099 , n26098 );
nand ( n26100 , n26091 , n26099 );
buf ( n26101 , n26100 );
buf ( n26102 , n26101 );
buf ( n26103 , n607 );
nand ( n26104 , n26102 , n26103 );
buf ( n26105 , n26104 );
buf ( n26106 , n26105 );
nand ( n26107 , n26075 , n26106 );
buf ( n26108 , n26107 );
buf ( n26109 , n26108 );
buf ( n26110 , n2361 );
buf ( n26111 , n592 );
and ( n26112 , n26110 , n26111 );
buf ( n26113 , n26112 );
buf ( n26114 , n26113 );
buf ( n26115 , n2452 );
not ( n26116 , n26115 );
buf ( n26117 , n592 );
not ( n26118 , n26117 );
buf ( n26119 , n7754 );
not ( n26120 , n26119 );
or ( n26121 , n26118 , n26120 );
buf ( n26122 , n2416 );
buf ( n26123 , n7751 );
nand ( n26124 , n26122 , n26123 );
buf ( n26125 , n26124 );
buf ( n26126 , n26125 );
nand ( n26127 , n26121 , n26126 );
buf ( n26128 , n26127 );
buf ( n26129 , n26128 );
not ( n26130 , n26129 );
or ( n26131 , n26116 , n26130 );
buf ( n26132 , n592 );
not ( n26133 , n26132 );
buf ( n26134 , n5458 );
not ( n26135 , n26134 );
or ( n26136 , n26133 , n26135 );
buf ( n26137 , n2416 );
buf ( n26138 , n5464 );
nand ( n26139 , n26137 , n26138 );
buf ( n26140 , n26139 );
buf ( n26141 , n26140 );
nand ( n26142 , n26136 , n26141 );
buf ( n26143 , n26142 );
buf ( n26144 , n26143 );
buf ( n26145 , n2460 );
nand ( n26146 , n26144 , n26145 );
buf ( n26147 , n26146 );
buf ( n26148 , n26147 );
nand ( n26149 , n26131 , n26148 );
buf ( n26150 , n26149 );
buf ( n26151 , n26150 );
xor ( n26152 , n26114 , n26151 );
buf ( n26153 , n2541 );
not ( n26154 , n26153 );
buf ( n26155 , n594 );
not ( n26156 , n26155 );
buf ( n26157 , n5407 );
not ( n26158 , n26157 );
or ( n26159 , n26156 , n26158 );
buf ( n26160 , n5411 );
buf ( n26161 , n2481 );
nand ( n26162 , n26160 , n26161 );
buf ( n26163 , n26162 );
buf ( n26164 , n26163 );
nand ( n26165 , n26159 , n26164 );
buf ( n26166 , n26165 );
buf ( n26167 , n26166 );
not ( n26168 , n26167 );
or ( n26169 , n26154 , n26168 );
buf ( n26170 , n594 );
not ( n26171 , n26170 );
buf ( n26172 , n8639 );
not ( n26173 , n26172 );
or ( n26174 , n26171 , n26173 );
not ( n26175 , n5572 );
buf ( n26176 , n26175 );
buf ( n26177 , n2481 );
nand ( n26178 , n26176 , n26177 );
buf ( n26179 , n26178 );
buf ( n26180 , n26179 );
nand ( n26181 , n26174 , n26180 );
buf ( n26182 , n26181 );
buf ( n26183 , n26182 );
buf ( n26184 , n2592 );
nand ( n26185 , n26183 , n26184 );
buf ( n26186 , n26185 );
buf ( n26187 , n26186 );
nand ( n26188 , n26169 , n26187 );
buf ( n26189 , n26188 );
buf ( n26190 , n26189 );
and ( n26191 , n26152 , n26190 );
and ( n26192 , n26114 , n26151 );
or ( n26193 , n26191 , n26192 );
buf ( n26194 , n26193 );
buf ( n26195 , n26194 );
buf ( n26196 , n592 );
not ( n26197 , n26196 );
buf ( n26198 , n8595 );
nor ( n26199 , n26197 , n26198 );
buf ( n26200 , n26199 );
buf ( n26201 , n26200 );
buf ( n26202 , n2452 );
not ( n26203 , n26202 );
buf ( n26204 , n592 );
not ( n26205 , n26204 );
buf ( n26206 , n8639 );
not ( n26207 , n26206 );
or ( n26208 , n26205 , n26207 );
buf ( n26209 , n26175 );
buf ( n26210 , n2416 );
nand ( n26211 , n26209 , n26210 );
buf ( n26212 , n26211 );
buf ( n26213 , n26212 );
nand ( n26214 , n26208 , n26213 );
buf ( n26215 , n26214 );
buf ( n26216 , n26215 );
not ( n26217 , n26216 );
or ( n26218 , n26203 , n26217 );
buf ( n26219 , n26128 );
buf ( n26220 , n2460 );
nand ( n26221 , n26219 , n26220 );
buf ( n26222 , n26221 );
buf ( n26223 , n26222 );
nand ( n26224 , n26218 , n26223 );
buf ( n26225 , n26224 );
buf ( n26226 , n26225 );
xor ( n26227 , n26201 , n26226 );
buf ( n26228 , n2541 );
not ( n26229 , n26228 );
and ( n26230 , n594 , n5376 );
not ( n26231 , n594 );
and ( n26232 , n26231 , n5373 );
or ( n26233 , n26230 , n26232 );
buf ( n26234 , n26233 );
not ( n26235 , n26234 );
or ( n26236 , n26229 , n26235 );
buf ( n26237 , n26166 );
buf ( n26238 , n2592 );
nand ( n26239 , n26237 , n26238 );
buf ( n26240 , n26239 );
buf ( n26241 , n26240 );
nand ( n26242 , n26236 , n26241 );
buf ( n26243 , n26242 );
buf ( n26244 , n26243 );
xor ( n26245 , n26227 , n26244 );
buf ( n26246 , n26245 );
buf ( n26247 , n26246 );
xor ( n26248 , n26195 , n26247 );
buf ( n26249 , n825 );
not ( n26250 , n26249 );
buf ( n26251 , n596 );
not ( n26252 , n26251 );
buf ( n26253 , n7593 );
not ( n26254 , n26253 );
or ( n26255 , n26252 , n26254 );
nand ( n26256 , n11008 , n2371 );
buf ( n26257 , n26256 );
nand ( n26258 , n26255 , n26257 );
buf ( n26259 , n26258 );
buf ( n26260 , n26259 );
not ( n26261 , n26260 );
or ( n26262 , n26250 , n26261 );
buf ( n26263 , n596 );
not ( n26264 , n26263 );
buf ( n26265 , n8684 );
not ( n26266 , n26265 );
or ( n26267 , n26264 , n26266 );
buf ( n26268 , n7648 );
buf ( n26269 , n2371 );
nand ( n26270 , n26268 , n26269 );
buf ( n26271 , n26270 );
buf ( n26272 , n26271 );
nand ( n26273 , n26267 , n26272 );
buf ( n26274 , n26273 );
buf ( n26275 , n26274 );
buf ( n26276 , n2404 );
buf ( n26277 , n26276 );
buf ( n26278 , n26277 );
buf ( n26279 , n26278 );
nand ( n26280 , n26275 , n26279 );
buf ( n26281 , n26280 );
buf ( n26282 , n26281 );
nand ( n26283 , n26262 , n26282 );
buf ( n26284 , n26283 );
buf ( n26285 , n26284 );
and ( n26286 , n26248 , n26285 );
and ( n26287 , n26195 , n26247 );
or ( n26288 , n26286 , n26287 );
buf ( n26289 , n26288 );
buf ( n26290 , n26289 );
not ( n26291 , n5550 );
not ( n26292 , n818 );
not ( n26293 , n9527 );
or ( n26294 , n26292 , n26293 );
nand ( n26295 , n598 , n9524 );
nand ( n26296 , n26294 , n26295 );
not ( n26297 , n26296 );
or ( n26298 , n26291 , n26297 );
buf ( n26299 , n598 );
not ( n26300 , n26299 );
not ( n26301 , n8553 );
buf ( n26302 , n26301 );
not ( n26303 , n26302 );
or ( n26304 , n26300 , n26303 );
buf ( n26305 , n8553 );
buf ( n26306 , n818 );
nand ( n26307 , n26305 , n26306 );
buf ( n26308 , n26307 );
buf ( n26309 , n26308 );
nand ( n26310 , n26304 , n26309 );
buf ( n26311 , n26310 );
buf ( n26312 , n26311 );
buf ( n26313 , n5631 );
nand ( n26314 , n26312 , n26313 );
buf ( n26315 , n26314 );
nand ( n26316 , n26298 , n26315 );
buf ( n26317 , n26316 );
xor ( n26318 , n26290 , n26317 );
xor ( n26319 , n26201 , n26226 );
and ( n26320 , n26319 , n26244 );
and ( n26321 , n26201 , n26226 );
or ( n26322 , n26320 , n26321 );
buf ( n26323 , n26322 );
buf ( n26324 , n26323 );
not ( n26325 , n26259 );
not ( n26326 , n26278 );
or ( n26327 , n26325 , n26326 );
buf ( n26328 , n11218 );
buf ( n26329 , n596 );
nor ( n26330 , n26328 , n26329 );
buf ( n26331 , n26330 );
and ( n26332 , n7559 , n26331 );
not ( n26333 , n7559 );
buf ( n26334 , n11218 );
buf ( n26335 , n2371 );
nor ( n26336 , n26334 , n26335 );
buf ( n26337 , n26336 );
and ( n26338 , n26333 , n26337 );
nor ( n26339 , n26332 , n26338 );
nand ( n26340 , n26327 , n26339 );
buf ( n26341 , n26340 );
xor ( n26342 , n26324 , n26341 );
buf ( n26343 , n5607 );
buf ( n26344 , n592 );
and ( n26345 , n26343 , n26344 );
buf ( n26346 , n26345 );
buf ( n26347 , n26346 );
buf ( n26348 , n2452 );
not ( n26349 , n26348 );
buf ( n26350 , n592 );
not ( n26351 , n26350 );
buf ( n26352 , n5407 );
not ( n26353 , n26352 );
or ( n26354 , n26351 , n26353 );
buf ( n26355 , n5411 );
buf ( n26356 , n2416 );
nand ( n26357 , n26355 , n26356 );
buf ( n26358 , n26357 );
buf ( n26359 , n26358 );
nand ( n26360 , n26354 , n26359 );
buf ( n26361 , n26360 );
buf ( n26362 , n26361 );
not ( n26363 , n26362 );
or ( n26364 , n26349 , n26363 );
buf ( n26365 , n26215 );
buf ( n26366 , n2460 );
nand ( n26367 , n26365 , n26366 );
buf ( n26368 , n26367 );
buf ( n26369 , n26368 );
nand ( n26370 , n26364 , n26369 );
buf ( n26371 , n26370 );
buf ( n26372 , n26371 );
xor ( n26373 , n26347 , n26372 );
buf ( n26374 , n2540 );
buf ( n26375 , n594 );
nor ( n26376 , n26374 , n26375 );
buf ( n26377 , n26376 );
nand ( n26378 , n26377 , n7648 );
buf ( n26379 , n26233 );
buf ( n26380 , n2592 );
nand ( n26381 , n26379 , n26380 );
buf ( n26382 , n26381 );
buf ( n26383 , n2540 );
buf ( n26384 , n2481 );
nor ( n26385 , n26383 , n26384 );
buf ( n26386 , n26385 );
nand ( n26387 , n11802 , n26386 );
nand ( n26388 , n26378 , n26382 , n26387 );
buf ( n26389 , n26388 );
xor ( n26390 , n26373 , n26389 );
buf ( n26391 , n26390 );
buf ( n26392 , n26391 );
xor ( n26393 , n26342 , n26392 );
buf ( n26394 , n26393 );
buf ( n26395 , n26394 );
and ( n26396 , n26318 , n26395 );
and ( n26397 , n26290 , n26317 );
or ( n26398 , n26396 , n26397 );
buf ( n26399 , n26398 );
buf ( n26400 , n26399 );
xor ( n26401 , n26109 , n26400 );
xor ( n26402 , n26324 , n26341 );
and ( n26403 , n26402 , n26392 );
and ( n26404 , n26324 , n26341 );
or ( n26405 , n26403 , n26404 );
buf ( n26406 , n26405 );
buf ( n26407 , n26406 );
not ( n26408 , n5631 );
not ( n26409 , n26296 );
or ( n26410 , n26408 , n26409 );
nand ( n26411 , n5550 , n598 );
buf ( n26412 , n26411 );
not ( n26413 , n26412 );
buf ( n26414 , n26413 );
or ( n26415 , n26414 , n10858 );
not ( n26416 , n10855 );
not ( n26417 , n10856 );
or ( n26418 , n26416 , n26417 );
nor ( n26419 , n5618 , n598 );
not ( n26420 , n26419 );
nand ( n26421 , n26418 , n26420 );
nand ( n26422 , n26415 , n26421 );
nand ( n26423 , n26410 , n26422 );
buf ( n26424 , n26423 );
xor ( n26425 , n26407 , n26424 );
and ( n26426 , n8553 , n26331 );
not ( n26427 , n8553 );
and ( n26428 , n26427 , n26337 );
nor ( n26429 , n26426 , n26428 );
buf ( n26430 , n596 );
not ( n26431 , n26430 );
buf ( n26432 , n7562 );
not ( n26433 , n26432 );
or ( n26434 , n26431 , n26433 );
buf ( n26435 , n7559 );
buf ( n26436 , n2371 );
nand ( n26437 , n26435 , n26436 );
buf ( n26438 , n26437 );
buf ( n26439 , n26438 );
nand ( n26440 , n26434 , n26439 );
buf ( n26441 , n26440 );
buf ( n26442 , n26441 );
buf ( n26443 , n26278 );
nand ( n26444 , n26442 , n26443 );
buf ( n26445 , n26444 );
nand ( n26446 , n26429 , n26445 );
buf ( n26447 , n26446 );
xor ( n26448 , n26347 , n26372 );
and ( n26449 , n26448 , n26389 );
and ( n26450 , n26347 , n26372 );
or ( n26451 , n26449 , n26450 );
buf ( n26452 , n26451 );
buf ( n26453 , n26452 );
xor ( n26454 , n26447 , n26453 );
buf ( n26455 , n26175 );
buf ( n26456 , n592 );
and ( n26457 , n26455 , n26456 );
buf ( n26458 , n26457 );
buf ( n26459 , n26458 );
buf ( n26460 , n2452 );
not ( n26461 , n26460 );
not ( n26462 , n5369 );
xor ( n26463 , n592 , n26462 );
buf ( n26464 , n26463 );
not ( n26465 , n26464 );
or ( n26466 , n26461 , n26465 );
buf ( n26467 , n26361 );
buf ( n26468 , n2460 );
nand ( n26469 , n26467 , n26468 );
buf ( n26470 , n26469 );
buf ( n26471 , n26470 );
nand ( n26472 , n26466 , n26471 );
buf ( n26473 , n26472 );
buf ( n26474 , n26473 );
xor ( n26475 , n26459 , n26474 );
buf ( n26476 , n2541 );
not ( n26477 , n26476 );
buf ( n26478 , n594 );
not ( n26479 , n26478 );
buf ( n26480 , n7593 );
not ( n26481 , n26480 );
or ( n26482 , n26479 , n26481 );
buf ( n26483 , n11008 );
buf ( n26484 , n2481 );
nand ( n26485 , n26483 , n26484 );
buf ( n26486 , n26485 );
buf ( n26487 , n26486 );
nand ( n26488 , n26482 , n26487 );
buf ( n26489 , n26488 );
buf ( n26490 , n26489 );
not ( n26491 , n26490 );
or ( n26492 , n26477 , n26491 );
buf ( n26493 , n7648 );
buf ( n26494 , n2659 );
and ( n26495 , n26493 , n26494 );
buf ( n26496 , n8684 );
buf ( n26497 , n2669 );
and ( n26498 , n26496 , n26497 );
nor ( n26499 , n26495 , n26498 );
buf ( n26500 , n26499 );
buf ( n26501 , n26500 );
nand ( n26502 , n26492 , n26501 );
buf ( n26503 , n26502 );
buf ( n26504 , n26503 );
xor ( n26505 , n26475 , n26504 );
buf ( n26506 , n26505 );
buf ( n26507 , n26506 );
xor ( n26508 , n26454 , n26507 );
buf ( n26509 , n26508 );
buf ( n26510 , n26509 );
xor ( n26511 , n26425 , n26510 );
buf ( n26512 , n26511 );
buf ( n26513 , n26512 );
and ( n26514 , n26401 , n26513 );
and ( n26515 , n26109 , n26400 );
or ( n26516 , n26514 , n26515 );
buf ( n26517 , n26516 );
buf ( n26518 , n26517 );
buf ( n26519 , n5430 );
not ( n26520 , n26519 );
and ( n26521 , n600 , n10861 );
not ( n26522 , n600 );
and ( n26523 , n26522 , n10858 );
or ( n26524 , n26521 , n26523 );
buf ( n26525 , n26524 );
not ( n26526 , n26525 );
or ( n26527 , n26520 , n26526 );
buf ( n26528 , n600 );
not ( n26529 , n26528 );
not ( n26530 , n10829 );
buf ( n26531 , n26530 );
not ( n26532 , n26531 );
or ( n26533 , n26529 , n26532 );
buf ( n26534 , n10829 );
buf ( n26535 , n7650 );
nand ( n26536 , n26534 , n26535 );
buf ( n26537 , n26536 );
buf ( n26538 , n26537 );
nand ( n26539 , n26533 , n26538 );
buf ( n26540 , n26539 );
buf ( n26541 , n26540 );
buf ( n26542 , n2915 );
nand ( n26543 , n26541 , n26542 );
buf ( n26544 , n26543 );
buf ( n26545 , n26544 );
nand ( n26546 , n26527 , n26545 );
buf ( n26547 , n26546 );
buf ( n26548 , n26547 );
and ( n26549 , n12936 , n12938 );
buf ( n26550 , n26549 );
buf ( n26551 , n26550 );
buf ( n26552 , n2452 );
not ( n26553 , n26552 );
buf ( n26554 , n26143 );
not ( n26555 , n26554 );
or ( n26556 , n26553 , n26555 );
buf ( n26557 , n592 );
not ( n26558 , n26557 );
buf ( n26559 , n2364 );
not ( n26560 , n26559 );
or ( n26561 , n26558 , n26560 );
buf ( n26562 , n2361 );
buf ( n26563 , n2416 );
nand ( n26564 , n26562 , n26563 );
buf ( n26565 , n26564 );
buf ( n26566 , n26565 );
nand ( n26567 , n26561 , n26566 );
buf ( n26568 , n26567 );
buf ( n26569 , n26568 );
buf ( n26570 , n2460 );
nand ( n26571 , n26569 , n26570 );
buf ( n26572 , n26571 );
buf ( n26573 , n26572 );
nand ( n26574 , n26556 , n26573 );
buf ( n26575 , n26574 );
buf ( n26576 , n26575 );
xor ( n26577 , n26551 , n26576 );
buf ( n26578 , n2541 );
not ( n26579 , n26578 );
buf ( n26580 , n26182 );
not ( n26581 , n26580 );
or ( n26582 , n26579 , n26581 );
buf ( n26583 , n594 );
not ( n26584 , n26583 );
buf ( n26585 , n7754 );
not ( n26586 , n26585 );
or ( n26587 , n26584 , n26586 );
buf ( n26588 , n2481 );
buf ( n26589 , n7751 );
nand ( n26590 , n26588 , n26589 );
buf ( n26591 , n26590 );
buf ( n26592 , n26591 );
nand ( n26593 , n26587 , n26592 );
buf ( n26594 , n26593 );
buf ( n26595 , n26594 );
buf ( n26596 , n2592 );
nand ( n26597 , n26595 , n26596 );
buf ( n26598 , n26597 );
buf ( n26599 , n26598 );
nand ( n26600 , n26582 , n26599 );
buf ( n26601 , n26600 );
buf ( n26602 , n26601 );
and ( n26603 , n26577 , n26602 );
and ( n26604 , n26551 , n26576 );
or ( n26605 , n26603 , n26604 );
buf ( n26606 , n26605 );
buf ( n26607 , n26606 );
xor ( n26608 , n26114 , n26151 );
xor ( n26609 , n26608 , n26190 );
buf ( n26610 , n26609 );
buf ( n26611 , n26610 );
xor ( n26612 , n26607 , n26611 );
buf ( n26613 , n825 );
not ( n26614 , n26613 );
buf ( n26615 , n26274 );
not ( n26616 , n26615 );
or ( n26617 , n26614 , n26616 );
and ( n26618 , n5373 , n2371 );
not ( n26619 , n5373 );
and ( n26620 , n26619 , n596 );
or ( n26621 , n26618 , n26620 );
buf ( n26622 , n26621 );
buf ( n26623 , n26278 );
nand ( n26624 , n26622 , n26623 );
buf ( n26625 , n26624 );
buf ( n26626 , n26625 );
nand ( n26627 , n26617 , n26626 );
buf ( n26628 , n26627 );
buf ( n26629 , n26628 );
and ( n26630 , n26612 , n26629 );
and ( n26631 , n26607 , n26611 );
or ( n26632 , n26630 , n26631 );
buf ( n26633 , n26632 );
buf ( n26634 , n26633 );
buf ( n26635 , n5550 );
not ( n26636 , n26635 );
buf ( n26637 , n26311 );
not ( n26638 , n26637 );
or ( n26639 , n26636 , n26638 );
buf ( n26640 , n598 );
not ( n26641 , n26640 );
buf ( n26642 , n7562 );
not ( n26643 , n26642 );
or ( n26644 , n26641 , n26643 );
buf ( n26645 , n7559 );
buf ( n26646 , n818 );
nand ( n26647 , n26645 , n26646 );
buf ( n26648 , n26647 );
buf ( n26649 , n26648 );
nand ( n26650 , n26644 , n26649 );
buf ( n26651 , n26650 );
buf ( n26652 , n26651 );
buf ( n26653 , n5631 );
nand ( n26654 , n26652 , n26653 );
buf ( n26655 , n26654 );
buf ( n26656 , n26655 );
nand ( n26657 , n26639 , n26656 );
buf ( n26658 , n26657 );
buf ( n26659 , n26658 );
xor ( n26660 , n26634 , n26659 );
xor ( n26661 , n26195 , n26247 );
xor ( n26662 , n26661 , n26285 );
buf ( n26663 , n26662 );
buf ( n26664 , n26663 );
and ( n26665 , n26660 , n26664 );
and ( n26666 , n26634 , n26659 );
or ( n26667 , n26665 , n26666 );
buf ( n26668 , n26667 );
buf ( n26669 , n26668 );
xor ( n26670 , n26548 , n26669 );
not ( n26671 , n18202 );
not ( n26672 , n18204 );
and ( n26673 , n26671 , n26672 );
and ( n26674 , n18204 , n18202 );
nor ( n26675 , n26673 , n26674 );
not ( n26676 , n26675 );
buf ( n26677 , n26676 );
not ( n26678 , n26677 );
buf ( n26679 , n5652 );
buf ( n26680 , n2912 );
nor ( n26681 , n26679 , n26680 );
buf ( n26682 , n26681 );
buf ( n26683 , n26682 );
not ( n26684 , n26683 );
buf ( n26685 , n26684 );
buf ( n26686 , n26685 );
not ( n26687 , n26686 );
and ( n26688 , n26678 , n26687 );
buf ( n26689 , n26676 );
buf ( n26690 , n5655 );
buf ( n26691 , n2912 );
and ( n26692 , n26690 , n26691 );
buf ( n26693 , n26692 );
buf ( n26694 , n26693 );
and ( n26695 , n26689 , n26694 );
nor ( n26696 , n26688 , n26695 );
buf ( n26697 , n26696 );
buf ( n26698 , n26697 );
buf ( n26699 , n602 );
not ( n26700 , n26699 );
buf ( n26701 , n13605 );
not ( n26702 , n26701 );
or ( n26703 , n26700 , n26702 );
buf ( n26704 , n13602 );
buf ( n26705 , n2912 );
nand ( n26706 , n26704 , n26705 );
buf ( n26707 , n26706 );
buf ( n26708 , n26707 );
nand ( n26709 , n26703 , n26708 );
buf ( n26710 , n26709 );
buf ( n26711 , n26710 );
buf ( n26712 , n7619 );
nand ( n26713 , n26711 , n26712 );
buf ( n26714 , n26713 );
buf ( n26715 , n26714 );
nand ( n26716 , n26698 , n26715 );
buf ( n26717 , n26716 );
buf ( n26718 , n26717 );
and ( n26719 , n26670 , n26718 );
and ( n26720 , n26548 , n26669 );
or ( n26721 , n26719 , n26720 );
buf ( n26722 , n26721 );
buf ( n26723 , n26722 );
buf ( n26724 , n26676 );
not ( n26725 , n26724 );
buf ( n26726 , n11930 );
nand ( n26727 , n26725 , n26726 );
buf ( n26728 , n26727 );
buf ( n26729 , n26676 );
buf ( n26730 , n11923 );
nand ( n26731 , n26729 , n26730 );
buf ( n26732 , n26731 );
and ( n26733 , n18205 , n20163 );
not ( n26734 , n18205 );
and ( n26735 , n26734 , n20160 );
nor ( n26736 , n26733 , n26735 );
buf ( n26737 , n26736 );
buf ( n26738 , n26737 );
not ( n26739 , n26738 );
buf ( n26740 , n26739 );
buf ( n26741 , n26740 );
buf ( n26742 , n26682 );
nand ( n26743 , n26741 , n26742 );
buf ( n26744 , n26743 );
buf ( n26745 , n26737 );
buf ( n26746 , n26693 );
nand ( n26747 , n26745 , n26746 );
buf ( n26748 , n26747 );
nand ( n26749 , n26728 , n26732 , n26744 , n26748 );
buf ( n26750 , n26749 );
not ( n26751 , n26540 );
not ( n26752 , n5430 );
or ( n26753 , n26751 , n26752 );
buf ( n26754 , n11547 );
buf ( n26755 , n600 );
nor ( n26756 , n26754 , n26755 );
buf ( n26757 , n26756 );
and ( n26758 , n13611 , n26757 );
not ( n26759 , n13611 );
buf ( n26760 , n11547 );
buf ( n26761 , n7650 );
nor ( n26762 , n26760 , n26761 );
buf ( n26763 , n26762 );
and ( n26764 , n26759 , n26763 );
nor ( n26765 , n26758 , n26764 );
nand ( n26766 , n26753 , n26765 );
buf ( n26767 , n26766 );
xor ( n26768 , n26750 , n26767 );
not ( n26769 , n8581 );
not ( n26770 , n604 );
buf ( n26771 , n26770 );
not ( n26772 , n26771 );
not ( n26773 , n14256 );
nand ( n26774 , n26773 , n18199 );
not ( n26775 , n26774 );
nor ( n26776 , n9520 , n18213 );
nand ( n26777 , n26775 , n26776 );
and ( n26778 , n26777 , n18207 );
not ( n26779 , n26777 );
and ( n26780 , n26779 , n18208 );
nor ( n26781 , n26778 , n26780 );
buf ( n26782 , n26781 );
buf ( n26783 , n26782 );
not ( n26784 , n26783 );
or ( n26785 , n26772 , n26784 );
not ( n26786 , n26781 );
buf ( n26787 , n26786 );
not ( n26788 , n26787 );
buf ( n26789 , n26788 );
buf ( n26790 , n26789 );
not ( n26791 , n26790 );
buf ( n26792 , n604 );
nand ( n26793 , n26791 , n26792 );
buf ( n26794 , n26793 );
buf ( n26795 , n26794 );
nand ( n26796 , n26785 , n26795 );
buf ( n26797 , n26796 );
not ( n26798 , n26797 );
or ( n26799 , n26769 , n26798 );
not ( n26800 , n12329 );
not ( n26801 , n18200 );
not ( n26802 , n18210 );
nand ( n26803 , n26801 , n26802 , n18208 , n9521 );
not ( n26804 , n18206 );
and ( n26805 , n26803 , n26804 );
not ( n26806 , n26803 );
buf ( n26807 , n18725 );
and ( n26808 , n26806 , n26807 );
nor ( n26809 , n26805 , n26808 );
buf ( n26810 , n26809 );
not ( n26811 , n26810 );
or ( n26812 , n26800 , n26811 );
not ( n26813 , n26810 );
not ( n26814 , n26813 );
or ( n26815 , n26814 , n12329 );
nand ( n26816 , n26812 , n26815 );
nand ( n26817 , n26816 , n7789 );
nand ( n26818 , n26799 , n26817 );
buf ( n26819 , n26818 );
xor ( n26820 , n26768 , n26819 );
buf ( n26821 , n26820 );
buf ( n26822 , n26821 );
xor ( n26823 , n26723 , n26822 );
buf ( n26824 , n8581 );
not ( n26825 , n26824 );
buf ( n26826 , n26737 );
not ( n26827 , n26826 );
buf ( n26828 , n26827 );
and ( n26829 , n604 , n26828 );
not ( n26830 , n604 );
and ( n26831 , n26830 , n26737 );
or ( n26832 , n26829 , n26831 );
buf ( n26833 , n26832 );
not ( n26834 , n26833 );
or ( n26835 , n26825 , n26834 );
buf ( n26836 , n26797 );
buf ( n26837 , n7790 );
nand ( n26838 , n26836 , n26837 );
buf ( n26839 , n26838 );
buf ( n26840 , n26839 );
nand ( n26841 , n26835 , n26840 );
buf ( n26842 , n26841 );
buf ( n26843 , n26842 );
buf ( n26844 , n607 );
not ( n26845 , n26844 );
buf ( n26846 , n26072 );
not ( n26847 , n26846 );
or ( n26848 , n26845 , n26847 );
buf ( n26849 , n606 );
not ( n26850 , n26849 );
not ( n26851 , n26810 );
buf ( n26852 , n26851 );
not ( n26853 , n26852 );
or ( n26854 , n26850 , n26853 );
buf ( n26855 , n26810 );
buf ( n26856 , n10836 );
nand ( n26857 , n26855 , n26856 );
buf ( n26858 , n26857 );
buf ( n26859 , n26858 );
nand ( n26860 , n26854 , n26859 );
buf ( n26861 , n26860 );
buf ( n26862 , n26861 );
buf ( n26863 , n10882 );
nand ( n26864 , n26862 , n26863 );
buf ( n26865 , n26864 );
buf ( n26866 , n26865 );
nand ( n26867 , n26848 , n26866 );
buf ( n26868 , n26867 );
buf ( n26869 , n26868 );
xor ( n26870 , n26843 , n26869 );
xor ( n26871 , n26290 , n26317 );
xor ( n26872 , n26871 , n26395 );
buf ( n26873 , n26872 );
buf ( n26874 , n26873 );
and ( n26875 , n26870 , n26874 );
and ( n26876 , n26843 , n26869 );
or ( n26877 , n26875 , n26876 );
buf ( n26878 , n26877 );
buf ( n26879 , n26878 );
and ( n26880 , n26823 , n26879 );
and ( n26881 , n26723 , n26822 );
or ( n26882 , n26880 , n26881 );
buf ( n26883 , n26882 );
buf ( n26884 , n26883 );
xor ( n26885 , n26518 , n26884 );
xor ( n26886 , n26447 , n26453 );
and ( n26887 , n26886 , n26507 );
and ( n26888 , n26447 , n26453 );
or ( n26889 , n26887 , n26888 );
buf ( n26890 , n26889 );
buf ( n26891 , n26890 );
not ( n26892 , n5550 );
not ( n26893 , n598 );
not ( n26894 , n10829 );
not ( n26895 , n26894 );
or ( n26896 , n26893 , n26895 );
buf ( n26897 , n10829 );
buf ( n26898 , n818 );
nand ( n26899 , n26897 , n26898 );
buf ( n26900 , n26899 );
nand ( n26901 , n26896 , n26900 );
not ( n26902 , n26901 );
or ( n26903 , n26892 , n26902 );
buf ( n26904 , n10858 );
not ( n26905 , n26904 );
buf ( n26906 , n11237 );
not ( n26907 , n26906 );
and ( n26908 , n26905 , n26907 );
buf ( n26909 , n10858 );
buf ( n26910 , n11248 );
and ( n26911 , n26909 , n26910 );
nor ( n26912 , n26908 , n26911 );
buf ( n26913 , n26912 );
nand ( n26914 , n26903 , n26913 );
buf ( n26915 , n26914 );
xor ( n26916 , n26891 , n26915 );
buf ( n26917 , n10945 );
not ( n26918 , n26917 );
buf ( n26919 , n600 );
not ( n26920 , n26919 );
buf ( n26921 , n26675 );
buf ( n26922 , n26921 );
not ( n26923 , n26922 );
or ( n26924 , n26920 , n26923 );
buf ( n26925 , n26676 );
buf ( n26926 , n7650 );
nand ( n26927 , n26925 , n26926 );
buf ( n26928 , n26927 );
buf ( n26929 , n26928 );
nand ( n26930 , n26924 , n26929 );
buf ( n26931 , n26930 );
buf ( n26932 , n26931 );
not ( n26933 , n26932 );
or ( n26934 , n26918 , n26933 );
buf ( n26935 , n13611 );
not ( n26936 , n26935 );
buf ( n26937 , n11568 );
not ( n26938 , n26937 );
and ( n26939 , n26936 , n26938 );
buf ( n26940 , n13611 );
buf ( n26941 , n11561 );
and ( n26942 , n26940 , n26941 );
nor ( n26943 , n26939 , n26942 );
buf ( n26944 , n26943 );
buf ( n26945 , n26944 );
nand ( n26946 , n26934 , n26945 );
buf ( n26947 , n26946 );
buf ( n26948 , n26947 );
xor ( n26949 , n26916 , n26948 );
buf ( n26950 , n26949 );
buf ( n26951 , n26950 );
buf ( n26952 , n5655 );
not ( n26953 , n26952 );
buf ( n26954 , n602 );
not ( n26955 , n26954 );
buf ( n26956 , n26786 );
not ( n26957 , n26956 );
or ( n26958 , n26955 , n26957 );
buf ( n26959 , n26782 );
buf ( n26960 , n2912 );
nand ( n26961 , n26959 , n26960 );
buf ( n26962 , n26961 );
buf ( n26963 , n26962 );
nand ( n26964 , n26958 , n26963 );
buf ( n26965 , n26964 );
buf ( n26966 , n26965 );
not ( n26967 , n26966 );
or ( n26968 , n26953 , n26967 );
buf ( n26969 , n11930 );
not ( n26970 , n26969 );
buf ( n26971 , n26970 );
not ( n26972 , n26971 );
not ( n26973 , n26737 );
not ( n26974 , n26973 );
or ( n26975 , n26972 , n26974 );
not ( n26976 , n26737 );
or ( n26977 , n26976 , n11923 );
nand ( n26978 , n26975 , n26977 );
buf ( n26979 , n26978 );
nand ( n26980 , n26968 , n26979 );
buf ( n26981 , n26980 );
buf ( n26982 , n26981 );
not ( n26983 , n7788 );
not ( n26984 , n604 );
not ( n26985 , n26062 );
or ( n26986 , n26984 , n26985 );
nand ( n26987 , n26053 , n26770 );
nand ( n26988 , n26986 , n26987 );
not ( n26989 , n26988 );
or ( n26990 , n26983 , n26989 );
nand ( n26991 , n26816 , n8581 );
nand ( n26992 , n26990 , n26991 );
buf ( n26993 , n26992 );
xor ( n26994 , n26982 , n26993 );
not ( n26995 , n607 );
buf ( n26996 , n606 );
not ( n26997 , n26996 );
buf ( n26998 , n18191 );
not ( n26999 , n26998 );
buf ( n27000 , n26999 );
buf ( n27001 , n27000 );
not ( n27002 , n27001 );
or ( n27003 , n26997 , n27002 );
buf ( n27004 , n18191 );
buf ( n27005 , n10836 );
nand ( n27006 , n27004 , n27005 );
buf ( n27007 , n27006 );
buf ( n27008 , n27007 );
nand ( n27009 , n27003 , n27008 );
buf ( n27010 , n27009 );
not ( n27011 , n27010 );
or ( n27012 , n26995 , n27011 );
nand ( n27013 , n26101 , n10882 );
nand ( n27014 , n27012 , n27013 );
buf ( n27015 , n27014 );
xor ( n27016 , n26994 , n27015 );
buf ( n27017 , n27016 );
buf ( n27018 , n27017 );
xor ( n27019 , n26951 , n27018 );
xor ( n27020 , n26459 , n26474 );
and ( n27021 , n27020 , n26504 );
and ( n27022 , n26459 , n26474 );
or ( n27023 , n27021 , n27022 );
buf ( n27024 , n27023 );
buf ( n27025 , n27024 );
buf ( n27026 , n5411 );
buf ( n27027 , n592 );
and ( n27028 , n27026 , n27027 );
buf ( n27029 , n27028 );
buf ( n27030 , n27029 );
buf ( n27031 , n2452 );
not ( n27032 , n27031 );
buf ( n27033 , n592 );
not ( n27034 , n27033 );
buf ( n27035 , n8684 );
not ( n27036 , n27035 );
or ( n27037 , n27034 , n27036 );
buf ( n27038 , n7648 );
buf ( n27039 , n2416 );
nand ( n27040 , n27038 , n27039 );
buf ( n27041 , n27040 );
buf ( n27042 , n27041 );
nand ( n27043 , n27037 , n27042 );
buf ( n27044 , n27043 );
buf ( n27045 , n27044 );
not ( n27046 , n27045 );
or ( n27047 , n27032 , n27046 );
buf ( n27048 , n26463 );
buf ( n27049 , n2460 );
nand ( n27050 , n27048 , n27049 );
buf ( n27051 , n27050 );
buf ( n27052 , n27051 );
nand ( n27053 , n27047 , n27052 );
buf ( n27054 , n27053 );
buf ( n27055 , n27054 );
xor ( n27056 , n27030 , n27055 );
buf ( n27057 , n2541 );
not ( n27058 , n27057 );
and ( n27059 , n594 , n7562 );
not ( n27060 , n594 );
and ( n27061 , n27060 , n7559 );
or ( n27062 , n27059 , n27061 );
buf ( n27063 , n27062 );
not ( n27064 , n27063 );
or ( n27065 , n27058 , n27064 );
buf ( n27066 , n26489 );
buf ( n27067 , n2592 );
nand ( n27068 , n27066 , n27067 );
buf ( n27069 , n27068 );
buf ( n27070 , n27069 );
nand ( n27071 , n27065 , n27070 );
buf ( n27072 , n27071 );
buf ( n27073 , n27072 );
xor ( n27074 , n27056 , n27073 );
buf ( n27075 , n27074 );
buf ( n27076 , n27075 );
xor ( n27077 , n27025 , n27076 );
not ( n27078 , n825 );
not ( n27079 , n596 );
not ( n27080 , n10902 );
or ( n27081 , n27079 , n27080 );
buf ( n27082 , n9527 );
buf ( n27083 , n2371 );
nand ( n27084 , n27082 , n27083 );
buf ( n27085 , n27084 );
nand ( n27086 , n27081 , n27085 );
not ( n27087 , n27086 );
or ( n27088 , n27078 , n27087 );
and ( n27089 , n8553 , n2845 );
not ( n27090 , n8553 );
and ( n27091 , n27090 , n2843 );
nor ( n27092 , n27089 , n27091 );
nand ( n27093 , n27088 , n27092 );
buf ( n27094 , n27093 );
xor ( n27095 , n27077 , n27094 );
buf ( n27096 , n27095 );
buf ( n27097 , n27096 );
xor ( n27098 , n26407 , n26424 );
and ( n27099 , n27098 , n26510 );
and ( n27100 , n26407 , n26424 );
or ( n27101 , n27099 , n27100 );
buf ( n27102 , n27101 );
buf ( n27103 , n27102 );
xor ( n27104 , n27097 , n27103 );
xor ( n27105 , n26750 , n26767 );
and ( n27106 , n27105 , n26819 );
and ( n27107 , n26750 , n26767 );
or ( n27108 , n27106 , n27107 );
buf ( n27109 , n27108 );
buf ( n27110 , n27109 );
xor ( n27111 , n27104 , n27110 );
buf ( n27112 , n27111 );
buf ( n27113 , n27112 );
xor ( n27114 , n27019 , n27113 );
buf ( n27115 , n27114 );
buf ( n27116 , n27115 );
xor ( n27117 , n26885 , n27116 );
buf ( n27118 , n27117 );
buf ( n27119 , n27118 );
not ( n27120 , n27119 );
buf ( n27121 , n27120 );
buf ( n27122 , n27121 );
buf ( n27123 , n825 );
not ( n27124 , n27123 );
and ( n27125 , n5373 , n2371 );
not ( n27126 , n5373 );
and ( n27127 , n27126 , n596 );
or ( n27128 , n27125 , n27127 );
buf ( n27129 , n27128 );
not ( n27130 , n27129 );
or ( n27131 , n27124 , n27130 );
buf ( n27132 , n596 );
not ( n27133 , n27132 );
buf ( n27134 , n5407 );
not ( n27135 , n27134 );
or ( n27136 , n27133 , n27135 );
buf ( n27137 , n5411 );
buf ( n27138 , n2371 );
nand ( n27139 , n27137 , n27138 );
buf ( n27140 , n27139 );
buf ( n27141 , n27140 );
nand ( n27142 , n27136 , n27141 );
buf ( n27143 , n27142 );
buf ( n27144 , n27143 );
buf ( n27145 , n2404 );
nand ( n27146 , n27144 , n27145 );
buf ( n27147 , n27146 );
buf ( n27148 , n27147 );
nand ( n27149 , n27131 , n27148 );
buf ( n27150 , n27149 );
buf ( n27151 , n27150 );
buf ( n27152 , n7719 );
not ( n27153 , n27152 );
buf ( n27154 , n2416 );
nor ( n27155 , n27153 , n27154 );
buf ( n27156 , n27155 );
buf ( n27157 , n27156 );
buf ( n27158 , n2452 );
not ( n27159 , n27158 );
buf ( n27160 , n26568 );
not ( n27161 , n27160 );
or ( n27162 , n27159 , n27161 );
buf ( n27163 , n12940 );
buf ( n27164 , n2460 );
nand ( n27165 , n27163 , n27164 );
buf ( n27166 , n27165 );
buf ( n27167 , n27166 );
nand ( n27168 , n27162 , n27167 );
buf ( n27169 , n27168 );
buf ( n27170 , n27169 );
xor ( n27171 , n27157 , n27170 );
not ( n27172 , n2541 );
not ( n27173 , n26594 );
or ( n27174 , n27172 , n27173 );
not ( n27175 , n2591 );
nand ( n27176 , n27175 , n12920 );
nand ( n27177 , n27174 , n27176 );
buf ( n27178 , n27177 );
and ( n27179 , n27171 , n27178 );
and ( n27180 , n27157 , n27170 );
or ( n27181 , n27179 , n27180 );
buf ( n27182 , n27181 );
buf ( n27183 , n27182 );
xor ( n27184 , n27151 , n27183 );
xor ( n27185 , n26551 , n26576 );
xor ( n27186 , n27185 , n26602 );
buf ( n27187 , n27186 );
buf ( n27188 , n27187 );
and ( n27189 , n27184 , n27188 );
and ( n27190 , n27151 , n27183 );
or ( n27191 , n27189 , n27190 );
buf ( n27192 , n27191 );
buf ( n27193 , n27192 );
buf ( n27194 , n5550 );
not ( n27195 , n27194 );
buf ( n27196 , n26651 );
not ( n27197 , n27196 );
or ( n27198 , n27195 , n27197 );
and ( n27199 , n598 , n7593 );
not ( n27200 , n598 );
and ( n27201 , n27200 , n11008 );
or ( n27202 , n27199 , n27201 );
buf ( n27203 , n27202 );
buf ( n27204 , n5631 );
nand ( n27205 , n27203 , n27204 );
buf ( n27206 , n27205 );
buf ( n27207 , n27206 );
nand ( n27208 , n27198 , n27207 );
buf ( n27209 , n27208 );
buf ( n27210 , n27209 );
xor ( n27211 , n27193 , n27210 );
xor ( n27212 , n26607 , n26611 );
xor ( n27213 , n27212 , n26629 );
buf ( n27214 , n27213 );
buf ( n27215 , n27214 );
and ( n27216 , n27211 , n27215 );
and ( n27217 , n27193 , n27210 );
or ( n27218 , n27216 , n27217 );
buf ( n27219 , n27218 );
buf ( n27220 , n27219 );
buf ( n27221 , n10945 );
not ( n27222 , n27221 );
buf ( n27223 , n26524 );
not ( n27224 , n27223 );
or ( n27225 , n27222 , n27224 );
not ( n27226 , n9527 );
not ( n27227 , n600 );
not ( n27228 , n27227 );
or ( n27229 , n27226 , n27228 );
nand ( n27230 , n9524 , n600 );
nand ( n27231 , n27229 , n27230 );
buf ( n27232 , n27231 );
buf ( n27233 , n5430 );
nand ( n27234 , n27232 , n27233 );
buf ( n27235 , n27234 );
buf ( n27236 , n27235 );
nand ( n27237 , n27225 , n27236 );
buf ( n27238 , n27237 );
buf ( n27239 , n27238 );
xor ( n27240 , n27220 , n27239 );
xor ( n27241 , n26634 , n26659 );
xor ( n27242 , n27241 , n26664 );
buf ( n27243 , n27242 );
buf ( n27244 , n27243 );
and ( n27245 , n27240 , n27244 );
and ( n27246 , n27220 , n27239 );
or ( n27247 , n27245 , n27246 );
buf ( n27248 , n27247 );
buf ( n27249 , n27248 );
xor ( n27250 , n26548 , n26669 );
xor ( n27251 , n27250 , n26718 );
buf ( n27252 , n27251 );
buf ( n27253 , n27252 );
xor ( n27254 , n27249 , n27253 );
buf ( n27255 , n7619 );
not ( n27256 , n27255 );
buf ( n27257 , n602 );
not ( n27258 , n27257 );
buf ( n27259 , n26894 );
not ( n27260 , n27259 );
or ( n27261 , n27258 , n27260 );
buf ( n27262 , n10829 );
buf ( n27263 , n2912 );
nand ( n27264 , n27262 , n27263 );
buf ( n27265 , n27264 );
buf ( n27266 , n27265 );
nand ( n27267 , n27261 , n27266 );
buf ( n27268 , n27267 );
buf ( n27269 , n27268 );
not ( n27270 , n27269 );
or ( n27271 , n27256 , n27270 );
buf ( n27272 , n26710 );
buf ( n27273 , n5655 );
nand ( n27274 , n27272 , n27273 );
buf ( n27275 , n27274 );
buf ( n27276 , n27275 );
nand ( n27277 , n27271 , n27276 );
buf ( n27278 , n27277 );
buf ( n27279 , n27278 );
buf ( n27280 , n10882 );
not ( n27281 , n27280 );
buf ( n27282 , n10836 );
not ( n27283 , n27282 );
buf ( n27284 , n26782 );
not ( n27285 , n27284 );
or ( n27286 , n27283 , n27285 );
buf ( n27287 , n26786 );
buf ( n27288 , n606 );
nand ( n27289 , n27287 , n27288 );
buf ( n27290 , n27289 );
buf ( n27291 , n27290 );
nand ( n27292 , n27286 , n27291 );
buf ( n27293 , n27292 );
buf ( n27294 , n27293 );
not ( n27295 , n27294 );
or ( n27296 , n27281 , n27295 );
buf ( n27297 , n26861 );
buf ( n27298 , n607 );
nand ( n27299 , n27297 , n27298 );
buf ( n27300 , n27299 );
buf ( n27301 , n27300 );
nand ( n27302 , n27296 , n27301 );
buf ( n27303 , n27302 );
buf ( n27304 , n27303 );
xor ( n27305 , n27279 , n27304 );
buf ( n27306 , n8581 );
not ( n27307 , n27306 );
and ( n27308 , n604 , n26921 );
not ( n27309 , n604 );
buf ( n27310 , n26921 );
not ( n27311 , n27310 );
buf ( n27312 , n27311 );
and ( n27313 , n27309 , n27312 );
or ( n27314 , n27308 , n27313 );
buf ( n27315 , n27314 );
not ( n27316 , n27315 );
or ( n27317 , n27307 , n27316 );
buf ( n27318 , n26832 );
buf ( n27319 , n7790 );
nand ( n27320 , n27318 , n27319 );
buf ( n27321 , n27320 );
buf ( n27322 , n27321 );
nand ( n27323 , n27317 , n27322 );
buf ( n27324 , n27323 );
buf ( n27325 , n27324 );
and ( n27326 , n27305 , n27325 );
and ( n27327 , n27279 , n27304 );
or ( n27328 , n27326 , n27327 );
buf ( n27329 , n27328 );
buf ( n27330 , n27329 );
and ( n27331 , n27254 , n27330 );
and ( n27332 , n27249 , n27253 );
or ( n27333 , n27331 , n27332 );
buf ( n27334 , n27333 );
buf ( n27335 , n27334 );
xor ( n27336 , n26109 , n26400 );
xor ( n27337 , n27336 , n26513 );
buf ( n27338 , n27337 );
buf ( n27339 , n27338 );
xor ( n27340 , n27335 , n27339 );
xor ( n27341 , n26723 , n26822 );
xor ( n27342 , n27341 , n26879 );
buf ( n27343 , n27342 );
buf ( n27344 , n27343 );
and ( n27345 , n27340 , n27344 );
and ( n27346 , n27335 , n27339 );
or ( n27347 , n27345 , n27346 );
buf ( n27348 , n27347 );
buf ( n27349 , n27348 );
not ( n27350 , n27349 );
buf ( n27351 , n27350 );
buf ( n27352 , n27351 );
nand ( n27353 , n27122 , n27352 );
buf ( n27354 , n27353 );
xor ( n27355 , n27335 , n27339 );
xor ( n27356 , n27355 , n27344 );
buf ( n27357 , n27356 );
not ( n27358 , n27357 );
xor ( n27359 , n26843 , n26869 );
xor ( n27360 , n27359 , n26874 );
buf ( n27361 , n27360 );
buf ( n27362 , n27361 );
xor ( n27363 , n12933 , n12951 );
and ( n27364 , n27363 , n12958 );
and ( n27365 , n12933 , n12951 );
or ( n27366 , n27364 , n27365 );
buf ( n27367 , n27366 );
buf ( n27368 , n27367 );
buf ( n27369 , n825 );
not ( n27370 , n27369 );
buf ( n27371 , n27143 );
not ( n27372 , n27371 );
or ( n27373 , n27370 , n27372 );
buf ( n27374 , n12976 );
buf ( n27375 , n2404 );
nand ( n27376 , n27374 , n27375 );
buf ( n27377 , n27376 );
buf ( n27378 , n27377 );
nand ( n27379 , n27373 , n27378 );
buf ( n27380 , n27379 );
buf ( n27381 , n27380 );
xor ( n27382 , n27368 , n27381 );
xor ( n27383 , n27157 , n27170 );
xor ( n27384 , n27383 , n27178 );
buf ( n27385 , n27384 );
buf ( n27386 , n27385 );
and ( n27387 , n27382 , n27386 );
and ( n27388 , n27368 , n27381 );
or ( n27389 , n27387 , n27388 );
buf ( n27390 , n27389 );
buf ( n27391 , n27390 );
buf ( n27392 , n5550 );
not ( n27393 , n27392 );
buf ( n27394 , n27202 );
not ( n27395 , n27394 );
or ( n27396 , n27393 , n27395 );
buf ( n27397 , n598 );
not ( n27398 , n27397 );
buf ( n27399 , n8684 );
not ( n27400 , n27399 );
or ( n27401 , n27398 , n27400 );
buf ( n27402 , n7648 );
buf ( n27403 , n818 );
nand ( n27404 , n27402 , n27403 );
buf ( n27405 , n27404 );
buf ( n27406 , n27405 );
nand ( n27407 , n27401 , n27406 );
buf ( n27408 , n27407 );
buf ( n27409 , n27408 );
buf ( n27410 , n5631 );
nand ( n27411 , n27409 , n27410 );
buf ( n27412 , n27411 );
buf ( n27413 , n27412 );
nand ( n27414 , n27396 , n27413 );
buf ( n27415 , n27414 );
buf ( n27416 , n27415 );
xor ( n27417 , n27391 , n27416 );
xor ( n27418 , n27151 , n27183 );
xor ( n27419 , n27418 , n27188 );
buf ( n27420 , n27419 );
buf ( n27421 , n27420 );
and ( n27422 , n27417 , n27421 );
and ( n27423 , n27391 , n27416 );
or ( n27424 , n27422 , n27423 );
buf ( n27425 , n27424 );
buf ( n27426 , n27425 );
not ( n27427 , n10945 );
not ( n27428 , n27231 );
or ( n27429 , n27427 , n27428 );
buf ( n27430 , n600 );
not ( n27431 , n27430 );
buf ( n27432 , n26301 );
not ( n27433 , n27432 );
or ( n27434 , n27431 , n27433 );
buf ( n27435 , n8553 );
buf ( n27436 , n5383 );
nand ( n27437 , n27435 , n27436 );
buf ( n27438 , n27437 );
buf ( n27439 , n27438 );
nand ( n27440 , n27434 , n27439 );
buf ( n27441 , n27440 );
nand ( n27442 , n27441 , n5430 );
nand ( n27443 , n27429 , n27442 );
buf ( n27444 , n27443 );
xor ( n27445 , n27426 , n27444 );
xor ( n27446 , n27193 , n27210 );
xor ( n27447 , n27446 , n27215 );
buf ( n27448 , n27447 );
buf ( n27449 , n27448 );
and ( n27450 , n27445 , n27449 );
and ( n27451 , n27426 , n27444 );
or ( n27452 , n27450 , n27451 );
buf ( n27453 , n27452 );
buf ( n27454 , n27453 );
xor ( n27455 , n27220 , n27239 );
xor ( n27456 , n27455 , n27244 );
buf ( n27457 , n27456 );
buf ( n27458 , n27457 );
xor ( n27459 , n27454 , n27458 );
buf ( n27460 , n7619 );
not ( n27461 , n27460 );
buf ( n27462 , n602 );
not ( n27463 , n27462 );
buf ( n27464 , n10861 );
not ( n27465 , n27464 );
or ( n27466 , n27463 , n27465 );
buf ( n27467 , n10858 );
buf ( n27468 , n2912 );
nand ( n27469 , n27467 , n27468 );
buf ( n27470 , n27469 );
buf ( n27471 , n27470 );
nand ( n27472 , n27466 , n27471 );
buf ( n27473 , n27472 );
buf ( n27474 , n27473 );
not ( n27475 , n27474 );
or ( n27476 , n27461 , n27475 );
buf ( n27477 , n27268 );
buf ( n27478 , n5655 );
nand ( n27479 , n27477 , n27478 );
buf ( n27480 , n27479 );
buf ( n27481 , n27480 );
nand ( n27482 , n27476 , n27481 );
buf ( n27483 , n27482 );
buf ( n27484 , n27483 );
buf ( n27485 , n2915 );
not ( n27486 , n27485 );
buf ( n27487 , n27441 );
not ( n27488 , n27487 );
or ( n27489 , n27486 , n27488 );
buf ( n27490 , n7559 );
buf ( n27491 , n600 );
and ( n27492 , n27490 , n27491 );
not ( n27493 , n27490 );
buf ( n27494 , n7650 );
and ( n27495 , n27493 , n27494 );
nor ( n27496 , n27492 , n27495 );
buf ( n27497 , n27496 );
buf ( n27498 , n27497 );
buf ( n27499 , n5430 );
nand ( n27500 , n27498 , n27499 );
buf ( n27501 , n27500 );
buf ( n27502 , n27501 );
nand ( n27503 , n27489 , n27502 );
buf ( n27504 , n27503 );
buf ( n27505 , n27504 );
xor ( n27506 , n12928 , n12961 );
and ( n27507 , n27506 , n12987 );
and ( n27508 , n12928 , n12961 );
or ( n27509 , n27507 , n27508 );
buf ( n27510 , n27509 );
buf ( n27511 , n27510 );
buf ( n27512 , n5550 );
not ( n27513 , n27512 );
buf ( n27514 , n27408 );
not ( n27515 , n27514 );
or ( n27516 , n27513 , n27515 );
buf ( n27517 , n12908 );
buf ( n27518 , n5631 );
nand ( n27519 , n27517 , n27518 );
buf ( n27520 , n27519 );
buf ( n27521 , n27520 );
nand ( n27522 , n27516 , n27521 );
buf ( n27523 , n27522 );
buf ( n27524 , n27523 );
xor ( n27525 , n27511 , n27524 );
xor ( n27526 , n27368 , n27381 );
xor ( n27527 , n27526 , n27386 );
buf ( n27528 , n27527 );
buf ( n27529 , n27528 );
and ( n27530 , n27525 , n27529 );
and ( n27531 , n27511 , n27524 );
or ( n27532 , n27530 , n27531 );
buf ( n27533 , n27532 );
buf ( n27534 , n27533 );
xor ( n27535 , n27505 , n27534 );
xor ( n27536 , n27391 , n27416 );
xor ( n27537 , n27536 , n27421 );
buf ( n27538 , n27537 );
buf ( n27539 , n27538 );
and ( n27540 , n27535 , n27539 );
and ( n27541 , n27505 , n27534 );
or ( n27542 , n27540 , n27541 );
buf ( n27543 , n27542 );
buf ( n27544 , n27543 );
xor ( n27545 , n27484 , n27544 );
buf ( n27546 , n26737 );
not ( n27547 , n27546 );
buf ( n27548 , n27547 );
and ( n27549 , n10836 , n27548 );
not ( n27550 , n10836 );
buf ( n27551 , n26737 );
buf ( n27552 , n27551 );
buf ( n27553 , n27552 );
and ( n27554 , n27550 , n27553 );
nor ( n27555 , n27549 , n27554 );
not ( n27556 , n27555 );
not ( n27557 , n10882 );
or ( n27558 , n27556 , n27557 );
buf ( n27559 , n27293 );
buf ( n27560 , n607 );
nand ( n27561 , n27559 , n27560 );
buf ( n27562 , n27561 );
nand ( n27563 , n27558 , n27562 );
buf ( n27564 , n27563 );
and ( n27565 , n27545 , n27564 );
and ( n27566 , n27484 , n27544 );
or ( n27567 , n27565 , n27566 );
buf ( n27568 , n27567 );
buf ( n27569 , n27568 );
and ( n27570 , n27459 , n27569 );
and ( n27571 , n27454 , n27458 );
or ( n27572 , n27570 , n27571 );
buf ( n27573 , n27572 );
buf ( n27574 , n27573 );
xor ( n27575 , n27362 , n27574 );
xor ( n27576 , n27249 , n27253 );
xor ( n27577 , n27576 , n27330 );
buf ( n27578 , n27577 );
buf ( n27579 , n27578 );
and ( n27580 , n27575 , n27579 );
and ( n27581 , n27362 , n27574 );
or ( n27582 , n27580 , n27581 );
buf ( n27583 , n27582 );
not ( n27584 , n27583 );
nand ( n27585 , n27358 , n27584 );
nand ( n27586 , n27354 , n27585 );
not ( n27587 , n27586 );
not ( n27588 , n27587 );
xor ( n27589 , n12870 , n12892 );
and ( n27590 , n27589 , n12993 );
and ( n27591 , n12870 , n12892 );
or ( n27592 , n27590 , n27591 );
buf ( n27593 , n27592 );
buf ( n27594 , n27593 );
buf ( n27595 , n5655 );
not ( n27596 , n27595 );
buf ( n27597 , n602 );
not ( n27598 , n27597 );
buf ( n27599 , n10902 );
not ( n27600 , n27599 );
or ( n27601 , n27598 , n27600 );
buf ( n27602 , n9527 );
buf ( n27603 , n2912 );
nand ( n27604 , n27602 , n27603 );
buf ( n27605 , n27604 );
buf ( n27606 , n27605 );
nand ( n27607 , n27601 , n27606 );
buf ( n27608 , n27607 );
buf ( n27609 , n27608 );
not ( n27610 , n27609 );
or ( n27611 , n27596 , n27610 );
buf ( n27612 , n7619 );
buf ( n27613 , n12852 );
nand ( n27614 , n27612 , n27613 );
buf ( n27615 , n27614 );
buf ( n27616 , n27615 );
nand ( n27617 , n27611 , n27616 );
buf ( n27618 , n27617 );
buf ( n27619 , n27618 );
xor ( n27620 , n27594 , n27619 );
xor ( n27621 , n12899 , n12913 );
and ( n27622 , n27621 , n12990 );
and ( n27623 , n12899 , n12913 );
or ( n27624 , n27622 , n27623 );
buf ( n27625 , n27624 );
buf ( n27626 , n27625 );
buf ( n27627 , n2915 );
not ( n27628 , n27627 );
buf ( n27629 , n27497 );
not ( n27630 , n27629 );
or ( n27631 , n27628 , n27630 );
buf ( n27632 , n12884 );
buf ( n27633 , n5430 );
nand ( n27634 , n27632 , n27633 );
buf ( n27635 , n27634 );
buf ( n27636 , n27635 );
nand ( n27637 , n27631 , n27636 );
buf ( n27638 , n27637 );
buf ( n27639 , n27638 );
xor ( n27640 , n27626 , n27639 );
xor ( n27641 , n27511 , n27524 );
xor ( n27642 , n27641 , n27529 );
buf ( n27643 , n27642 );
buf ( n27644 , n27643 );
xor ( n27645 , n27640 , n27644 );
buf ( n27646 , n27645 );
buf ( n27647 , n27646 );
xor ( n27648 , n27620 , n27647 );
buf ( n27649 , n27648 );
buf ( n27650 , n27649 );
xor ( n27651 , n13012 , n13029 );
and ( n27652 , n27651 , n13629 );
and ( n27653 , n13012 , n13029 );
or ( n27654 , n27652 , n27653 );
buf ( n27655 , n27654 );
buf ( n27656 , n27655 );
xor ( n27657 , n27650 , n27656 );
buf ( n27658 , n7790 );
not ( n27659 , n27658 );
buf ( n27660 , n604 );
not ( n27661 , n27660 );
buf ( n27662 , n10831 );
not ( n27663 , n27662 );
or ( n27664 , n27661 , n27663 );
buf ( n27665 , n604 );
not ( n27666 , n27665 );
buf ( n27667 , n10830 );
nand ( n27668 , n27666 , n27667 );
buf ( n27669 , n27668 );
buf ( n27670 , n27669 );
nand ( n27671 , n27664 , n27670 );
buf ( n27672 , n27671 );
buf ( n27673 , n27672 );
not ( n27674 , n27673 );
or ( n27675 , n27659 , n27674 );
buf ( n27676 , n13018 );
buf ( n27677 , n8581 );
nand ( n27678 , n27676 , n27677 );
buf ( n27679 , n27678 );
buf ( n27680 , n27679 );
nand ( n27681 , n27675 , n27680 );
buf ( n27682 , n27681 );
buf ( n27683 , n27682 );
xor ( n27684 , n12838 , n12863 );
and ( n27685 , n27684 , n12996 );
and ( n27686 , n12838 , n12863 );
or ( n27687 , n27685 , n27686 );
buf ( n27688 , n27687 );
buf ( n27689 , n27688 );
xor ( n27690 , n27683 , n27689 );
buf ( n27691 , n607 );
not ( n27692 , n27691 );
buf ( n27693 , n606 );
not ( n27694 , n27693 );
buf ( n27695 , n26921 );
not ( n27696 , n27695 );
or ( n27697 , n27694 , n27696 );
buf ( n27698 , n27312 );
buf ( n27699 , n10836 );
nand ( n27700 , n27698 , n27699 );
buf ( n27701 , n27700 );
buf ( n27702 , n27701 );
nand ( n27703 , n27697 , n27702 );
buf ( n27704 , n27703 );
buf ( n27705 , n27704 );
not ( n27706 , n27705 );
or ( n27707 , n27692 , n27706 );
buf ( n27708 , n13618 );
buf ( n27709 , n10882 );
nand ( n27710 , n27708 , n27709 );
buf ( n27711 , n27710 );
buf ( n27712 , n27711 );
nand ( n27713 , n27707 , n27712 );
buf ( n27714 , n27713 );
buf ( n27715 , n27714 );
xor ( n27716 , n27690 , n27715 );
buf ( n27717 , n27716 );
buf ( n27718 , n27717 );
xor ( n27719 , n27657 , n27718 );
buf ( n27720 , n27719 );
buf ( n27721 , n27720 );
xor ( n27722 , n12999 , n13005 );
and ( n27723 , n27722 , n13632 );
and ( n27724 , n12999 , n13005 );
or ( n27725 , n27723 , n27724 );
buf ( n27726 , n27725 );
buf ( n27727 , n27726 );
nor ( n27728 , n27721 , n27727 );
buf ( n27729 , n27728 );
buf ( n27730 , n27729 );
not ( n27731 , n27730 );
buf ( n27732 , n13640 );
buf ( n27733 , n11048 );
nand ( n27734 , n27731 , n27732 , n27733 );
buf ( n27735 , n27734 );
not ( n27736 , n12827 );
or ( n27737 , n27735 , n27736 );
buf ( n27738 , n27720 );
not ( n27739 , n27738 );
buf ( n27740 , n27739 );
buf ( n27741 , n27740 );
buf ( n27742 , n27726 );
not ( n27743 , n27742 );
buf ( n27744 , n27743 );
buf ( n27745 , n27744 );
nand ( n27746 , n27741 , n27745 );
buf ( n27747 , n27746 );
buf ( n27748 , n27747 );
buf ( n27749 , n13634 );
buf ( n27750 , n13639 );
nor ( n27751 , n27749 , n27750 );
buf ( n27752 , n27751 );
or ( n27753 , n27752 , n12830 );
nand ( n27754 , n27753 , n13645 );
buf ( n27755 , n27754 );
and ( n27756 , n27748 , n27755 );
buf ( n27757 , n27720 );
buf ( n27758 , n27726 );
nand ( n27759 , n27757 , n27758 );
buf ( n27760 , n27759 );
buf ( n27761 , n27760 );
not ( n27762 , n27761 );
buf ( n27763 , n27762 );
buf ( n27764 , n27763 );
nor ( n27765 , n27756 , n27764 );
buf ( n27766 , n27765 );
nand ( n27767 , n27737 , n27766 );
not ( n27768 , n27767 );
xor ( n27769 , n27362 , n27574 );
xor ( n27770 , n27769 , n27579 );
buf ( n27771 , n27770 );
buf ( n27772 , n27771 );
not ( n27773 , n27772 );
buf ( n27774 , n27773 );
buf ( n27775 , n27774 );
xor ( n27776 , n27279 , n27304 );
xor ( n27777 , n27776 , n27325 );
buf ( n27778 , n27777 );
buf ( n27779 , n27778 );
buf ( n27780 , n7790 );
not ( n27781 , n27780 );
buf ( n27782 , n27314 );
not ( n27783 , n27782 );
or ( n27784 , n27781 , n27783 );
buf ( n27785 , n13611 );
not ( n27786 , n27785 );
buf ( n27787 , n27786 );
and ( n27788 , n604 , n27787 );
not ( n27789 , n604 );
and ( n27790 , n27789 , n13611 );
or ( n27791 , n27788 , n27790 );
buf ( n27792 , n27791 );
buf ( n27793 , n8581 );
nand ( n27794 , n27792 , n27793 );
buf ( n27795 , n27794 );
buf ( n27796 , n27795 );
nand ( n27797 , n27784 , n27796 );
buf ( n27798 , n27797 );
buf ( n27799 , n27798 );
xor ( n27800 , n27426 , n27444 );
xor ( n27801 , n27800 , n27449 );
buf ( n27802 , n27801 );
buf ( n27803 , n27802 );
xor ( n27804 , n27799 , n27803 );
xor ( n27805 , n27626 , n27639 );
and ( n27806 , n27805 , n27644 );
and ( n27807 , n27626 , n27639 );
or ( n27808 , n27806 , n27807 );
buf ( n27809 , n27808 );
buf ( n27810 , n27809 );
buf ( n27811 , n5655 );
not ( n27812 , n27811 );
buf ( n27813 , n27473 );
not ( n27814 , n27813 );
or ( n27815 , n27812 , n27814 );
buf ( n27816 , n27608 );
buf ( n27817 , n7619 );
nand ( n27818 , n27816 , n27817 );
buf ( n27819 , n27818 );
buf ( n27820 , n27819 );
nand ( n27821 , n27815 , n27820 );
buf ( n27822 , n27821 );
buf ( n27823 , n27822 );
xor ( n27824 , n27810 , n27823 );
buf ( n27825 , n7790 );
not ( n27826 , n27825 );
buf ( n27827 , n27791 );
not ( n27828 , n27827 );
or ( n27829 , n27826 , n27828 );
buf ( n27830 , n27672 );
buf ( n27831 , n8581 );
nand ( n27832 , n27830 , n27831 );
buf ( n27833 , n27832 );
buf ( n27834 , n27833 );
nand ( n27835 , n27829 , n27834 );
buf ( n27836 , n27835 );
buf ( n27837 , n27836 );
and ( n27838 , n27824 , n27837 );
and ( n27839 , n27810 , n27823 );
or ( n27840 , n27838 , n27839 );
buf ( n27841 , n27840 );
buf ( n27842 , n27841 );
and ( n27843 , n27804 , n27842 );
and ( n27844 , n27799 , n27803 );
or ( n27845 , n27843 , n27844 );
buf ( n27846 , n27845 );
buf ( n27847 , n27846 );
xor ( n27848 , n27779 , n27847 );
xor ( n27849 , n27454 , n27458 );
xor ( n27850 , n27849 , n27569 );
buf ( n27851 , n27850 );
buf ( n27852 , n27851 );
and ( n27853 , n27848 , n27852 );
and ( n27854 , n27779 , n27847 );
or ( n27855 , n27853 , n27854 );
buf ( n27856 , n27855 );
buf ( n27857 , n27856 );
not ( n27858 , n27857 );
buf ( n27859 , n27858 );
buf ( n27860 , n27859 );
nand ( n27861 , n27775 , n27860 );
buf ( n27862 , n27861 );
buf ( n27863 , n27862 );
xor ( n27864 , n27779 , n27847 );
xor ( n27865 , n27864 , n27852 );
buf ( n27866 , n27865 );
buf ( n27867 , n27866 );
not ( n27868 , n27867 );
xor ( n27869 , n27484 , n27544 );
xor ( n27870 , n27869 , n27564 );
buf ( n27871 , n27870 );
buf ( n27872 , n27871 );
xor ( n27873 , n27505 , n27534 );
xor ( n27874 , n27873 , n27539 );
buf ( n27875 , n27874 );
buf ( n27876 , n27875 );
buf ( n27877 , n10882 );
not ( n27878 , n27877 );
buf ( n27879 , n27704 );
not ( n27880 , n27879 );
or ( n27881 , n27878 , n27880 );
buf ( n27882 , n10836 );
buf ( n27883 , n27548 );
and ( n27884 , n27882 , n27883 );
not ( n27885 , n27882 );
buf ( n27886 , n27553 );
and ( n27887 , n27885 , n27886 );
nor ( n27888 , n27884 , n27887 );
buf ( n27889 , n27888 );
buf ( n27890 , n27889 );
buf ( n27891 , n607 );
nand ( n27892 , n27890 , n27891 );
buf ( n27893 , n27892 );
buf ( n27894 , n27893 );
nand ( n27895 , n27881 , n27894 );
buf ( n27896 , n27895 );
buf ( n27897 , n27896 );
xor ( n27898 , n27876 , n27897 );
xor ( n27899 , n27594 , n27619 );
and ( n27900 , n27899 , n27647 );
and ( n27901 , n27594 , n27619 );
or ( n27902 , n27900 , n27901 );
buf ( n27903 , n27902 );
buf ( n27904 , n27903 );
and ( n27905 , n27898 , n27904 );
and ( n27906 , n27876 , n27897 );
or ( n27907 , n27905 , n27906 );
buf ( n27908 , n27907 );
buf ( n27909 , n27908 );
xor ( n27910 , n27872 , n27909 );
xor ( n27911 , n27799 , n27803 );
xor ( n27912 , n27911 , n27842 );
buf ( n27913 , n27912 );
buf ( n27914 , n27913 );
and ( n27915 , n27910 , n27914 );
and ( n27916 , n27872 , n27909 );
or ( n27917 , n27915 , n27916 );
buf ( n27918 , n27917 );
buf ( n27919 , n27918 );
not ( n27920 , n27919 );
buf ( n27921 , n27920 );
buf ( n27922 , n27921 );
nand ( n27923 , n27868 , n27922 );
buf ( n27924 , n27923 );
buf ( n27925 , n27924 );
nand ( n27926 , n27863 , n27925 );
buf ( n27927 , n27926 );
buf ( n27928 , n27927 );
xor ( n27929 , n27872 , n27909 );
xor ( n27930 , n27929 , n27914 );
buf ( n27931 , n27930 );
xor ( n27932 , n27683 , n27689 );
and ( n27933 , n27932 , n27715 );
and ( n27934 , n27683 , n27689 );
or ( n27935 , n27933 , n27934 );
buf ( n27936 , n27935 );
buf ( n27937 , n27936 );
xor ( n27938 , n27810 , n27823 );
xor ( n27939 , n27938 , n27837 );
buf ( n27940 , n27939 );
buf ( n27941 , n27940 );
xor ( n27942 , n27937 , n27941 );
xor ( n27943 , n27876 , n27897 );
xor ( n27944 , n27943 , n27904 );
buf ( n27945 , n27944 );
buf ( n27946 , n27945 );
and ( n27947 , n27942 , n27946 );
and ( n27948 , n27937 , n27941 );
or ( n27949 , n27947 , n27948 );
buf ( n27950 , n27949 );
or ( n27951 , n27931 , n27950 );
xor ( n27952 , n27937 , n27941 );
xor ( n27953 , n27952 , n27946 );
buf ( n27954 , n27953 );
buf ( n27955 , n27954 );
not ( n27956 , n27955 );
xor ( n27957 , n27650 , n27656 );
and ( n27958 , n27957 , n27718 );
and ( n27959 , n27650 , n27656 );
or ( n27960 , n27958 , n27959 );
buf ( n27961 , n27960 );
buf ( n27962 , n27961 );
not ( n27963 , n27962 );
buf ( n27964 , n27963 );
buf ( n27965 , n27964 );
nand ( n27966 , n27956 , n27965 );
buf ( n27967 , n27966 );
nand ( n27968 , n27951 , n27967 );
buf ( n27969 , n27968 );
nor ( n27970 , n27928 , n27969 );
buf ( n27971 , n27970 );
not ( n27972 , n27971 );
or ( n27973 , n27768 , n27972 );
buf ( n27974 , n27927 );
not ( n27975 , n27974 );
buf ( n27976 , n27975 );
buf ( n27977 , n27976 );
buf ( n27978 , n27931 );
buf ( n27979 , n27950 );
nor ( n27980 , n27978 , n27979 );
buf ( n27981 , n27980 );
buf ( n27982 , n27981 );
buf ( n27983 , n27954 );
buf ( n27984 , n27961 );
nand ( n27985 , n27983 , n27984 );
buf ( n27986 , n27985 );
buf ( n27987 , n27986 );
or ( n27988 , n27982 , n27987 );
buf ( n27989 , n27931 );
buf ( n27990 , n27950 );
nand ( n27991 , n27989 , n27990 );
buf ( n27992 , n27991 );
buf ( n27993 , n27992 );
nand ( n27994 , n27988 , n27993 );
buf ( n27995 , n27994 );
buf ( n27996 , n27995 );
and ( n27997 , n27977 , n27996 );
buf ( n27998 , n27866 );
not ( n27999 , n27998 );
buf ( n28000 , n27999 );
buf ( n28001 , n28000 );
buf ( n28002 , n27921 );
nor ( n28003 , n28001 , n28002 );
buf ( n28004 , n28003 );
buf ( n28005 , n28004 );
not ( n28006 , n28005 );
buf ( n28007 , n27774 );
buf ( n28008 , n27859 );
nand ( n28009 , n28007 , n28008 );
buf ( n28010 , n28009 );
buf ( n28011 , n28010 );
not ( n28012 , n28011 );
or ( n28013 , n28006 , n28012 );
not ( n28014 , n27774 );
nand ( n28015 , n28014 , n27856 );
buf ( n28016 , n28015 );
nand ( n28017 , n28013 , n28016 );
buf ( n28018 , n28017 );
buf ( n28019 , n28018 );
nor ( n28020 , n27997 , n28019 );
buf ( n28021 , n28020 );
nand ( n28022 , n27973 , n28021 );
not ( n28023 , n28022 );
or ( n28024 , n27588 , n28023 );
not ( n28025 , n27118 );
not ( n28026 , n27348 );
or ( n28027 , n28025 , n28026 );
buf ( n28028 , n27583 );
buf ( n28029 , n27357 );
nand ( n28030 , n28028 , n28029 );
buf ( n28031 , n28030 );
nand ( n28032 , n28027 , n28031 );
buf ( n28033 , n28032 );
buf ( n28034 , n27354 );
and ( n28035 , n28033 , n28034 );
buf ( n28036 , n28035 );
buf ( n28037 , n28036 );
not ( n28038 , n28037 );
buf ( n28039 , n28038 );
nand ( n28040 , n28024 , n28039 );
xor ( n28041 , n27030 , n27055 );
and ( n28042 , n28041 , n27073 );
and ( n28043 , n27030 , n27055 );
or ( n28044 , n28042 , n28043 );
buf ( n28045 , n28044 );
buf ( n28046 , n28045 );
and ( n28047 , n592 , n26462 );
buf ( n28048 , n28047 );
buf ( n28049 , n2452 );
not ( n28050 , n28049 );
buf ( n28051 , n592 );
not ( n28052 , n28051 );
buf ( n28053 , n11011 );
not ( n28054 , n28053 );
or ( n28055 , n28052 , n28054 );
buf ( n28056 , n7599 );
buf ( n28057 , n2416 );
nand ( n28058 , n28056 , n28057 );
buf ( n28059 , n28058 );
buf ( n28060 , n28059 );
nand ( n28061 , n28055 , n28060 );
buf ( n28062 , n28061 );
buf ( n28063 , n28062 );
not ( n28064 , n28063 );
or ( n28065 , n28050 , n28064 );
buf ( n28066 , n27044 );
buf ( n28067 , n2460 );
nand ( n28068 , n28066 , n28067 );
buf ( n28069 , n28068 );
buf ( n28070 , n28069 );
nand ( n28071 , n28065 , n28070 );
buf ( n28072 , n28071 );
buf ( n28073 , n28072 );
xor ( n28074 , n28048 , n28073 );
buf ( n28075 , n2541 );
not ( n28076 , n28075 );
xor ( n28077 , n594 , n8553 );
buf ( n28078 , n28077 );
not ( n28079 , n28078 );
or ( n28080 , n28076 , n28079 );
buf ( n28081 , n27062 );
buf ( n28082 , n2592 );
nand ( n28083 , n28081 , n28082 );
buf ( n28084 , n28083 );
buf ( n28085 , n28084 );
nand ( n28086 , n28080 , n28085 );
buf ( n28087 , n28086 );
buf ( n28088 , n28087 );
xor ( n28089 , n28074 , n28088 );
buf ( n28090 , n28089 );
buf ( n28091 , n28090 );
xor ( n28092 , n28046 , n28091 );
buf ( n28093 , n26278 );
not ( n28094 , n28093 );
buf ( n28095 , n27086 );
not ( n28096 , n28095 );
or ( n28097 , n28094 , n28096 );
buf ( n28098 , n596 );
not ( n28099 , n28098 );
buf ( n28100 , n10861 );
not ( n28101 , n28100 );
or ( n28102 , n28099 , n28101 );
buf ( n28103 , n10858 );
buf ( n28104 , n2371 );
nand ( n28105 , n28103 , n28104 );
buf ( n28106 , n28105 );
buf ( n28107 , n28106 );
nand ( n28108 , n28102 , n28107 );
buf ( n28109 , n28108 );
buf ( n28110 , n28109 );
buf ( n28111 , n825 );
nand ( n28112 , n28110 , n28111 );
buf ( n28113 , n28112 );
buf ( n28114 , n28113 );
nand ( n28115 , n28097 , n28114 );
buf ( n28116 , n28115 );
buf ( n28117 , n28116 );
xor ( n28118 , n28092 , n28117 );
buf ( n28119 , n28118 );
buf ( n28120 , n28119 );
xor ( n28121 , n26891 , n26915 );
and ( n28122 , n28121 , n26948 );
and ( n28123 , n26891 , n26915 );
or ( n28124 , n28122 , n28123 );
buf ( n28125 , n28124 );
buf ( n28126 , n28125 );
xor ( n28127 , n28120 , n28126 );
xor ( n28128 , n26982 , n26993 );
and ( n28129 , n28128 , n27015 );
and ( n28130 , n26982 , n26993 );
or ( n28131 , n28129 , n28130 );
buf ( n28132 , n28131 );
buf ( n28133 , n28132 );
xor ( n28134 , n28127 , n28133 );
buf ( n28135 , n28134 );
buf ( n28136 , n28135 );
buf ( n28137 , n7619 );
not ( n28138 , n28137 );
buf ( n28139 , n26965 );
not ( n28140 , n28139 );
or ( n28141 , n28138 , n28140 );
buf ( n28142 , n26810 );
not ( n28143 , n28142 );
buf ( n28144 , n26685 );
not ( n28145 , n28144 );
and ( n28146 , n28143 , n28145 );
buf ( n28147 , n26810 );
buf ( n28148 , n26693 );
and ( n28149 , n28147 , n28148 );
nor ( n28150 , n28146 , n28149 );
buf ( n28151 , n28150 );
buf ( n28152 , n28151 );
nand ( n28153 , n28141 , n28152 );
buf ( n28154 , n28153 );
buf ( n28155 , n28154 );
not ( n28156 , n5631 );
not ( n28157 , n26901 );
or ( n28158 , n28156 , n28157 );
not ( n28159 , n818 );
buf ( n28160 , n13605 );
not ( n28161 , n28160 );
buf ( n28162 , n28161 );
not ( n28163 , n28162 );
or ( n28164 , n28159 , n28163 );
buf ( n28165 , n13602 );
not ( n28166 , n28165 );
buf ( n28167 , n598 );
nand ( n28168 , n28166 , n28167 );
buf ( n28169 , n28168 );
nand ( n28170 , n28164 , n28169 );
nand ( n28171 , n28170 , n5550 );
nand ( n28172 , n28158 , n28171 );
buf ( n28173 , n28172 );
xor ( n28174 , n28155 , n28173 );
buf ( n28175 , n10945 );
not ( n28176 , n28175 );
buf ( n28177 , n600 );
buf ( n28178 , n26737 );
buf ( n28179 , n28178 );
buf ( n28180 , n28179 );
buf ( n28181 , n28180 );
and ( n28182 , n28177 , n28181 );
not ( n28183 , n28177 );
buf ( n28184 , n26828 );
and ( n28185 , n28183 , n28184 );
nor ( n28186 , n28182 , n28185 );
buf ( n28187 , n28186 );
buf ( n28188 , n28187 );
not ( n28189 , n28188 );
or ( n28190 , n28176 , n28189 );
buf ( n28191 , n26931 );
buf ( n28192 , n5430 );
nand ( n28193 , n28191 , n28192 );
buf ( n28194 , n28193 );
buf ( n28195 , n28194 );
nand ( n28196 , n28190 , n28195 );
buf ( n28197 , n28196 );
buf ( n28198 , n28197 );
xor ( n28199 , n28174 , n28198 );
buf ( n28200 , n28199 );
buf ( n28201 , n28200 );
buf ( n28202 , n8581 );
not ( n28203 , n28202 );
buf ( n28204 , n26988 );
not ( n28205 , n28204 );
or ( n28206 , n28203 , n28205 );
and ( n28207 , n604 , n26088 );
not ( n28208 , n604 );
buf ( n28209 , n26085 );
buf ( n28210 , n28209 );
buf ( n28211 , n28210 );
and ( n28212 , n28208 , n28211 );
or ( n28213 , n28207 , n28212 );
buf ( n28214 , n28213 );
buf ( n28215 , n7790 );
nand ( n28216 , n28214 , n28215 );
buf ( n28217 , n28216 );
buf ( n28218 , n28217 );
nand ( n28219 , n28206 , n28218 );
buf ( n28220 , n28219 );
buf ( n28221 , n28220 );
xor ( n28222 , n27025 , n27076 );
and ( n28223 , n28222 , n27094 );
and ( n28224 , n27025 , n27076 );
or ( n28225 , n28223 , n28224 );
buf ( n28226 , n28225 );
buf ( n28227 , n28226 );
xor ( n28228 , n28221 , n28227 );
buf ( n28229 , n10882 );
not ( n28230 , n28229 );
buf ( n28231 , n27010 );
not ( n28232 , n28231 );
or ( n28233 , n28230 , n28232 );
not ( n28234 , n606 );
nand ( n28235 , n18111 , n9517 );
not ( n28236 , n28235 );
nand ( n28237 , n28236 , n15682 , n18082 , n18137 );
buf ( n28238 , n19384 );
and ( n28239 , n28237 , n28238 );
not ( n28240 , n28237 );
not ( n28241 , n24346 );
and ( n28242 , n28240 , n28241 );
nor ( n28243 , n28239 , n28242 );
not ( n28244 , n28243 );
not ( n28245 , n28244 );
or ( n28246 , n28234 , n28245 );
buf ( n28247 , n28243 );
nand ( n28248 , n28247 , n10836 );
nand ( n28249 , n28246 , n28248 );
buf ( n28250 , n28249 );
buf ( n28251 , n607 );
nand ( n28252 , n28250 , n28251 );
buf ( n28253 , n28252 );
buf ( n28254 , n28253 );
nand ( n28255 , n28233 , n28254 );
buf ( n28256 , n28255 );
buf ( n28257 , n28256 );
xor ( n28258 , n28228 , n28257 );
buf ( n28259 , n28258 );
buf ( n28260 , n28259 );
xor ( n28261 , n28201 , n28260 );
xor ( n28262 , n27097 , n27103 );
and ( n28263 , n28262 , n27110 );
and ( n28264 , n27097 , n27103 );
or ( n28265 , n28263 , n28264 );
buf ( n28266 , n28265 );
buf ( n28267 , n28266 );
xor ( n28268 , n28261 , n28267 );
buf ( n28269 , n28268 );
buf ( n28270 , n28269 );
xor ( n28271 , n28136 , n28270 );
xor ( n28272 , n26951 , n27018 );
and ( n28273 , n28272 , n27113 );
and ( n28274 , n26951 , n27018 );
or ( n28275 , n28273 , n28274 );
buf ( n28276 , n28275 );
buf ( n28277 , n28276 );
xor ( n28278 , n28271 , n28277 );
buf ( n28279 , n28278 );
buf ( n28280 , n28279 );
not ( n28281 , n28280 );
buf ( n28282 , n28281 );
buf ( n28283 , n28282 );
xor ( n28284 , n26518 , n26884 );
and ( n28285 , n28284 , n27116 );
and ( n28286 , n26518 , n26884 );
or ( n28287 , n28285 , n28286 );
buf ( n28288 , n28287 );
buf ( n28289 , n28288 );
not ( n28290 , n28289 );
buf ( n28291 , n28290 );
buf ( n28292 , n28291 );
nand ( n28293 , n28283 , n28292 );
buf ( n28294 , n28293 );
buf ( n28295 , n28294 );
buf ( n28296 , n28282 );
not ( n28297 , n28296 );
buf ( n28298 , n28288 );
nand ( n28299 , n28297 , n28298 );
buf ( n28300 , n28299 );
buf ( n28301 , n28300 );
nand ( n28302 , n28295 , n28301 );
buf ( n28303 , n28302 );
xnor ( n28304 , n28040 , n28303 );
buf ( n28305 , n28304 );
buf ( n28306 , n28305 );
buf ( n28307 , n28306 );
xor ( n28308 , n26043 , n26044 );
xor ( n28309 , n28308 , n28307 );
buf ( n28310 , n28309 );
xor ( n28311 , n26043 , n26044 );
and ( n28312 , n28311 , n28307 );
and ( n28313 , n26043 , n26044 );
or ( n28314 , n28312 , n28313 );
buf ( n28315 , n28314 );
buf ( n28316 , n9025 );
buf ( n28317 , n9234 );
buf ( n28318 , n13661 );
xor ( n28319 , n28316 , n28317 );
xor ( n28320 , n28319 , n28318 );
buf ( n28321 , n28320 );
xor ( n28322 , n28316 , n28317 );
and ( n28323 , n28322 , n28318 );
and ( n28324 , n28316 , n28317 );
or ( n28325 , n28323 , n28324 );
buf ( n28326 , n28325 );
buf ( n28327 , n9931 );
buf ( n28328 , n10153 );
not ( n28329 , n27736 );
not ( n28330 , n11045 );
not ( n28331 , n10894 );
not ( n28332 , n28331 );
or ( n28333 , n28330 , n28332 );
nand ( n28334 , n28333 , n12830 );
buf ( n28335 , n28334 );
not ( n28336 , n28335 );
buf ( n28337 , n28336 );
not ( n28338 , n28337 );
or ( n28339 , n28329 , n28338 );
buf ( n28340 , n28334 );
buf ( n28341 , n12827 );
nand ( n28342 , n28340 , n28341 );
buf ( n28343 , n28342 );
nand ( n28344 , n28339 , n28343 );
buf ( n28345 , n28344 );
xor ( n28346 , n28327 , n28328 );
xor ( n28347 , n28346 , n28345 );
buf ( n28348 , n28347 );
xor ( n28349 , n28327 , n28328 );
and ( n28350 , n28349 , n28345 );
and ( n28351 , n28327 , n28328 );
or ( n28352 , n28350 , n28351 );
buf ( n28353 , n28352 );
buf ( n28354 , n14179 );
buf ( n28355 , n14027 );
not ( n28356 , n27767 );
buf ( n28357 , n27967 );
buf ( n28358 , n27986 );
nand ( n28359 , n28357 , n28358 );
buf ( n28360 , n28359 );
and ( n28361 , n28356 , n28360 );
not ( n28362 , n28356 );
buf ( n28363 , n28360 );
not ( n28364 , n28363 );
buf ( n28365 , n28364 );
and ( n28366 , n28362 , n28365 );
nor ( n28367 , n28361 , n28366 );
buf ( n28368 , n28367 );
buf ( n28369 , n28368 );
xor ( n28370 , n28354 , n28355 );
xor ( n28371 , n28370 , n28369 );
buf ( n28372 , n28371 );
xor ( n28373 , n28354 , n28355 );
and ( n28374 , n28373 , n28369 );
and ( n28375 , n28354 , n28355 );
or ( n28376 , n28374 , n28375 );
buf ( n28377 , n28376 );
buf ( n28378 , n14920 );
buf ( n28379 , n15065 );
not ( n28380 , n27767 );
buf ( n28381 , n27968 );
not ( n28382 , n28381 );
buf ( n28383 , n28382 );
not ( n28384 , n28383 );
or ( n28385 , n28380 , n28384 );
buf ( n28386 , n27995 );
not ( n28387 , n28386 );
buf ( n28388 , n28387 );
nand ( n28389 , n28385 , n28388 );
not ( n28390 , n28389 );
buf ( n28391 , n28000 );
buf ( n28392 , n27921 );
nand ( n28393 , n28391 , n28392 );
buf ( n28394 , n28393 );
buf ( n28395 , n28394 );
buf ( n28396 , n28000 );
not ( n28397 , n28396 );
buf ( n28398 , n27918 );
nand ( n28399 , n28397 , n28398 );
buf ( n28400 , n28399 );
buf ( n28401 , n28400 );
nand ( n28402 , n28395 , n28401 );
buf ( n28403 , n28402 );
and ( n28404 , n28390 , n28403 );
not ( n28405 , n28390 );
buf ( n28406 , n28403 );
not ( n28407 , n28406 );
buf ( n28408 , n28407 );
and ( n28409 , n28405 , n28408 );
nor ( n28410 , n28404 , n28409 );
buf ( n28411 , n28410 );
buf ( n28412 , n28411 );
xor ( n28413 , n28378 , n28379 );
xor ( n28414 , n28413 , n28412 );
buf ( n28415 , n28414 );
xor ( n28416 , n28378 , n28379 );
and ( n28417 , n28416 , n28412 );
and ( n28418 , n28378 , n28379 );
or ( n28419 , n28417 , n28418 );
buf ( n28420 , n28419 );
buf ( n28421 , n6679 );
buf ( n28422 , n6866 );
and ( n28423 , n11721 , n12765 );
buf ( n28424 , n12759 );
and ( n28425 , n28423 , n28424 );
not ( n28426 , n28423 );
not ( n28427 , n28424 );
and ( n28428 , n28426 , n28427 );
nor ( n28429 , n28425 , n28428 );
buf ( n28430 , n28429 );
buf ( n28431 , n28430 );
xor ( n28432 , n28421 , n28422 );
xor ( n28433 , n28432 , n28431 );
buf ( n28434 , n28433 );
xor ( n28435 , n28421 , n28422 );
and ( n28436 , n28435 , n28431 );
and ( n28437 , n28421 , n28422 );
or ( n28438 , n28436 , n28437 );
buf ( n28439 , n28438 );
buf ( n28440 , n17053 );
buf ( n28441 , n17059 );
not ( n28442 , n28294 );
not ( n28443 , n28040 );
or ( n28444 , n28442 , n28443 );
nand ( n28445 , n28444 , n28300 );
xor ( n28446 , n28136 , n28270 );
and ( n28447 , n28446 , n28277 );
and ( n28448 , n28136 , n28270 );
or ( n28449 , n28447 , n28448 );
buf ( n28450 , n28449 );
buf ( n28451 , n28450 );
not ( n28452 , n28451 );
buf ( n28453 , n28452 );
buf ( n28454 , n28453 );
not ( n28455 , n28454 );
buf ( n28456 , n28455 );
buf ( n28457 , n28456 );
xor ( n28458 , n28155 , n28173 );
and ( n28459 , n28458 , n28198 );
and ( n28460 , n28155 , n28173 );
or ( n28461 , n28459 , n28460 );
buf ( n28462 , n28461 );
buf ( n28463 , n28462 );
xor ( n28464 , n28048 , n28073 );
and ( n28465 , n28464 , n28088 );
and ( n28466 , n28048 , n28073 );
or ( n28467 , n28465 , n28466 );
buf ( n28468 , n28467 );
buf ( n28469 , n28468 );
buf ( n28470 , n26278 );
not ( n28471 , n28470 );
buf ( n28472 , n28109 );
not ( n28473 , n28472 );
or ( n28474 , n28471 , n28473 );
and ( n28475 , n10829 , n2371 );
not ( n28476 , n10829 );
and ( n28477 , n28476 , n596 );
or ( n28478 , n28475 , n28477 );
buf ( n28479 , n28478 );
buf ( n28480 , n825 );
nand ( n28481 , n28479 , n28480 );
buf ( n28482 , n28481 );
buf ( n28483 , n28482 );
nand ( n28484 , n28474 , n28483 );
buf ( n28485 , n28484 );
buf ( n28486 , n28485 );
xor ( n28487 , n28469 , n28486 );
not ( n28488 , n5631 );
not ( n28489 , n28170 );
or ( n28490 , n28488 , n28489 );
buf ( n28491 , n27312 );
not ( n28492 , n28491 );
buf ( n28493 , n26411 );
not ( n28494 , n28493 );
and ( n28495 , n28492 , n28494 );
buf ( n28496 , n26676 );
buf ( n28497 , n26419 );
and ( n28498 , n28496 , n28497 );
nor ( n28499 , n28495 , n28498 );
buf ( n28500 , n28499 );
nand ( n28501 , n28490 , n28500 );
buf ( n28502 , n28501 );
xor ( n28503 , n28487 , n28502 );
buf ( n28504 , n28503 );
buf ( n28505 , n28504 );
xor ( n28506 , n28463 , n28505 );
not ( n28507 , n10945 );
buf ( n28508 , n600 );
not ( n28509 , n28508 );
buf ( n28510 , n26786 );
not ( n28511 , n28510 );
or ( n28512 , n28509 , n28511 );
buf ( n28513 , n26782 );
buf ( n28514 , n7650 );
nand ( n28515 , n28513 , n28514 );
buf ( n28516 , n28515 );
buf ( n28517 , n28516 );
nand ( n28518 , n28512 , n28517 );
buf ( n28519 , n28518 );
not ( n28520 , n28519 );
or ( n28521 , n28507 , n28520 );
or ( n28522 , n26976 , n11561 );
nand ( n28523 , n26976 , n11568 );
nand ( n28524 , n28522 , n28523 );
nand ( n28525 , n28521 , n28524 );
buf ( n28526 , n28525 );
buf ( n28527 , n7648 );
buf ( n28528 , n592 );
and ( n28529 , n28527 , n28528 );
buf ( n28530 , n28529 );
buf ( n28531 , n28530 );
buf ( n28532 , n2452 );
not ( n28533 , n28532 );
buf ( n28534 , n592 );
buf ( n28535 , n7559 );
xor ( n28536 , n28534 , n28535 );
buf ( n28537 , n28536 );
buf ( n28538 , n28537 );
not ( n28539 , n28538 );
or ( n28540 , n28533 , n28539 );
buf ( n28541 , n28062 );
buf ( n28542 , n2460 );
buf ( n28543 , n28542 );
buf ( n28544 , n28543 );
buf ( n28545 , n28544 );
nand ( n28546 , n28541 , n28545 );
buf ( n28547 , n28546 );
buf ( n28548 , n28547 );
nand ( n28549 , n28540 , n28548 );
buf ( n28550 , n28549 );
buf ( n28551 , n28550 );
xor ( n28552 , n28531 , n28551 );
and ( n28553 , n9527 , n26377 );
not ( n28554 , n9527 );
and ( n28555 , n28554 , n26386 );
nor ( n28556 , n28553 , n28555 );
buf ( n28557 , n28077 );
buf ( n28558 , n2592 );
nand ( n28559 , n28557 , n28558 );
buf ( n28560 , n28559 );
nand ( n28561 , n28556 , n28560 );
buf ( n28562 , n28561 );
xor ( n28563 , n28552 , n28562 );
buf ( n28564 , n28563 );
buf ( n28565 , n28564 );
xor ( n28566 , n28526 , n28565 );
buf ( n28567 , n7790 );
not ( n28568 , n28567 );
not ( n28569 , n604 );
not ( n28570 , n27000 );
or ( n28571 , n28569 , n28570 );
not ( n28572 , n604 );
nand ( n28573 , n28572 , n18191 );
nand ( n28574 , n28571 , n28573 );
buf ( n28575 , n28574 );
not ( n28576 , n28575 );
or ( n28577 , n28568 , n28576 );
buf ( n28578 , n28213 );
buf ( n28579 , n8581 );
nand ( n28580 , n28578 , n28579 );
buf ( n28581 , n28580 );
buf ( n28582 , n28581 );
nand ( n28583 , n28577 , n28582 );
buf ( n28584 , n28583 );
buf ( n28585 , n28584 );
xor ( n28586 , n28566 , n28585 );
buf ( n28587 , n28586 );
buf ( n28588 , n28587 );
xor ( n28589 , n28506 , n28588 );
buf ( n28590 , n28589 );
buf ( n28591 , n28590 );
xor ( n28592 , n28201 , n28260 );
and ( n28593 , n28592 , n28267 );
and ( n28594 , n28201 , n28260 );
or ( n28595 , n28593 , n28594 );
buf ( n28596 , n28595 );
buf ( n28597 , n28596 );
xor ( n28598 , n28591 , n28597 );
xor ( n28599 , n28221 , n28227 );
and ( n28600 , n28599 , n28257 );
and ( n28601 , n28221 , n28227 );
or ( n28602 , n28600 , n28601 );
buf ( n28603 , n28602 );
buf ( n28604 , n28603 );
buf ( n28605 , n5655 );
not ( n28606 , n28605 );
buf ( n28607 , n602 );
not ( n28608 , n28607 );
buf ( n28609 , n26053 );
not ( n28610 , n28609 );
buf ( n28611 , n28610 );
buf ( n28612 , n28611 );
not ( n28613 , n28612 );
or ( n28614 , n28608 , n28613 );
buf ( n28615 , n26053 );
buf ( n28616 , n2912 );
nand ( n28617 , n28615 , n28616 );
buf ( n28618 , n28617 );
buf ( n28619 , n28618 );
nand ( n28620 , n28614 , n28619 );
buf ( n28621 , n28620 );
buf ( n28622 , n28621 );
not ( n28623 , n28622 );
or ( n28624 , n28606 , n28623 );
not ( n28625 , n26810 );
not ( n28626 , n28625 );
buf ( n28627 , n28626 );
buf ( n28628 , n11923 );
and ( n28629 , n28627 , n28628 );
buf ( n28630 , n28625 );
buf ( n28631 , n11930 );
and ( n28632 , n28630 , n28631 );
nor ( n28633 , n28629 , n28632 );
buf ( n28634 , n28633 );
buf ( n28635 , n28634 );
nand ( n28636 , n28624 , n28635 );
buf ( n28637 , n28636 );
buf ( n28638 , n28637 );
xor ( n28639 , n28046 , n28091 );
and ( n28640 , n28639 , n28117 );
and ( n28641 , n28046 , n28091 );
or ( n28642 , n28640 , n28641 );
buf ( n28643 , n28642 );
buf ( n28644 , n28643 );
xor ( n28645 , n28638 , n28644 );
buf ( n28646 , n10882 );
not ( n28647 , n28646 );
buf ( n28648 , n28249 );
not ( n28649 , n28648 );
or ( n28650 , n28647 , n28649 );
buf ( n28651 , n606 );
not ( n28652 , n28651 );
not ( n28653 , n18195 );
and ( n28654 , n18082 , n19383 );
and ( n28655 , n18184 , n18201 , n18140 );
nand ( n28656 , n28654 , n18212 , n28655 );
not ( n28657 , n28656 );
or ( n28658 , n28653 , n28657 );
buf ( n28659 , n18195 );
not ( n28660 , n28659 );
buf ( n28661 , n28660 );
nand ( n28662 , n28654 , n18212 , n28655 , n28661 );
nand ( n28663 , n28658 , n28662 );
buf ( n28664 , n28663 );
buf ( n28665 , n28664 );
not ( n28666 , n28665 );
buf ( n28667 , n28666 );
buf ( n28668 , n28667 );
not ( n28669 , n28668 );
or ( n28670 , n28652 , n28669 );
buf ( n28671 , n28664 );
buf ( n28672 , n10836 );
nand ( n28673 , n28671 , n28672 );
buf ( n28674 , n28673 );
buf ( n28675 , n28674 );
nand ( n28676 , n28670 , n28675 );
buf ( n28677 , n28676 );
buf ( n28678 , n28677 );
buf ( n28679 , n607 );
nand ( n28680 , n28678 , n28679 );
buf ( n28681 , n28680 );
buf ( n28682 , n28681 );
nand ( n28683 , n28650 , n28682 );
buf ( n28684 , n28683 );
buf ( n28685 , n28684 );
xor ( n28686 , n28645 , n28685 );
buf ( n28687 , n28686 );
buf ( n28688 , n28687 );
xor ( n28689 , n28604 , n28688 );
xor ( n28690 , n28120 , n28126 );
and ( n28691 , n28690 , n28133 );
and ( n28692 , n28120 , n28126 );
or ( n28693 , n28691 , n28692 );
buf ( n28694 , n28693 );
buf ( n28695 , n28694 );
xor ( n28696 , n28689 , n28695 );
buf ( n28697 , n28696 );
buf ( n28698 , n28697 );
xor ( n28699 , n28598 , n28698 );
buf ( n28700 , n28699 );
buf ( n28701 , n28700 );
not ( n28702 , n28701 );
buf ( n28703 , n28702 );
buf ( n28704 , n28703 );
not ( n28705 , n28704 );
buf ( n28706 , n28705 );
buf ( n28707 , n28706 );
nand ( n28708 , n28457 , n28707 );
buf ( n28709 , n28708 );
buf ( n28710 , n28703 );
buf ( n28711 , n28453 );
nand ( n28712 , n28710 , n28711 );
buf ( n28713 , n28712 );
buf ( n28714 , n28713 );
nand ( n28715 , n28709 , n28714 );
not ( n28716 , n28715 );
and ( n28717 , n28445 , n28716 );
not ( n28718 , n28445 );
and ( n28719 , n28718 , n28715 );
nor ( n28720 , n28717 , n28719 );
buf ( n28721 , n28720 );
not ( n28722 , n28721 );
not ( n28723 , n28722 );
buf ( n28724 , n28723 );
xor ( n28725 , n28440 , n28441 );
xor ( n28726 , n28725 , n28724 );
buf ( n28727 , n28726 );
xor ( n28728 , n28440 , n28441 );
and ( n28729 , n28728 , n28724 );
and ( n28730 , n28440 , n28441 );
or ( n28731 , n28729 , n28730 );
buf ( n28732 , n28731 );
buf ( n28733 , n1274 );
buf ( n28734 , n1277 );
xor ( n28735 , n28733 , n28734 );
buf ( n28736 , n28735 );
and ( n28737 , n28733 , n28734 );
buf ( n28738 , n28737 );
buf ( n28739 , n17903 );
buf ( n28740 , n17896 );
xor ( n28741 , n28739 , n28740 );
buf ( n28742 , n28741 );
buf ( n28743 , n17508 );
buf ( n28744 , n17515 );
xor ( n28745 , n28743 , n28744 );
and ( n28746 , n10829 , n2371 );
not ( n28747 , n10829 );
and ( n28748 , n28747 , n596 );
or ( n28749 , n28746 , n28748 );
not ( n28750 , n28749 );
not ( n28751 , n26278 );
or ( n28752 , n28750 , n28751 );
and ( n28753 , n13602 , n26331 );
not ( n28754 , n13602 );
and ( n28755 , n28754 , n26337 );
nor ( n28756 , n28753 , n28755 );
nand ( n28757 , n28752 , n28756 );
buf ( n28758 , n28757 );
buf ( n28759 , n26676 );
buf ( n28760 , n11237 );
or ( n28761 , n28759 , n28760 );
buf ( n28762 , n28761 );
buf ( n28763 , n28762 );
buf ( n28764 , n26737 );
not ( n28765 , n28764 );
buf ( n28766 , n26414 );
nand ( n28767 , n28765 , n28766 );
buf ( n28768 , n28767 );
buf ( n28769 , n28768 );
buf ( n28770 , n26737 );
buf ( n28771 , n26419 );
nand ( n28772 , n28770 , n28771 );
buf ( n28773 , n28772 );
buf ( n28774 , n28773 );
buf ( n28775 , n26676 );
buf ( n28776 , n11248 );
nand ( n28777 , n28775 , n28776 );
buf ( n28778 , n28777 );
buf ( n28779 , n28778 );
nand ( n28780 , n28763 , n28769 , n28774 , n28779 );
buf ( n28781 , n28780 );
buf ( n28782 , n28781 );
xor ( n28783 , n28758 , n28782 );
not ( n28784 , n2915 );
and ( n28785 , n26810 , n7650 );
not ( n28786 , n26810 );
and ( n28787 , n28786 , n600 );
or ( n28788 , n28785 , n28787 );
not ( n28789 , n28788 );
or ( n28790 , n28784 , n28789 );
nand ( n28791 , n28519 , n5430 );
nand ( n28792 , n28790 , n28791 );
buf ( n28793 , n28792 );
xor ( n28794 , n28783 , n28793 );
buf ( n28795 , n28794 );
buf ( n28796 , n28795 );
xor ( n28797 , n28526 , n28565 );
and ( n28798 , n28797 , n28585 );
and ( n28799 , n28526 , n28565 );
or ( n28800 , n28798 , n28799 );
buf ( n28801 , n28800 );
buf ( n28802 , n28801 );
xor ( n28803 , n28796 , n28802 );
buf ( n28804 , n28211 );
not ( n28805 , n28804 );
buf ( n28806 , n26685 );
not ( n28807 , n28806 );
and ( n28808 , n28805 , n28807 );
buf ( n28809 , n26094 );
buf ( n28810 , n26693 );
and ( n28811 , n28809 , n28810 );
nor ( n28812 , n28808 , n28811 );
buf ( n28813 , n28812 );
buf ( n28814 , n26062 );
buf ( n28815 , n11930 );
nand ( n28816 , n28814 , n28815 );
buf ( n28817 , n28816 );
nand ( n28818 , n26053 , n11923 );
nand ( n28819 , n28813 , n28817 , n28818 );
buf ( n28820 , n28819 );
xor ( n28821 , n28531 , n28551 );
and ( n28822 , n28821 , n28562 );
and ( n28823 , n28531 , n28551 );
or ( n28824 , n28822 , n28823 );
buf ( n28825 , n28824 );
buf ( n28826 , n28825 );
xor ( n28827 , n28820 , n28826 );
buf ( n28828 , n11008 );
buf ( n28829 , n592 );
and ( n28830 , n28828 , n28829 );
buf ( n28831 , n28830 );
buf ( n28832 , n28831 );
buf ( n28833 , n2452 );
not ( n28834 , n28833 );
buf ( n28835 , n592 );
not ( n28836 , n28835 );
buf ( n28837 , n8554 );
not ( n28838 , n28837 );
or ( n28839 , n28836 , n28838 );
buf ( n28840 , n8553 );
buf ( n28841 , n2416 );
nand ( n28842 , n28840 , n28841 );
buf ( n28843 , n28842 );
buf ( n28844 , n28843 );
nand ( n28845 , n28839 , n28844 );
buf ( n28846 , n28845 );
buf ( n28847 , n28846 );
not ( n28848 , n28847 );
or ( n28849 , n28834 , n28848 );
buf ( n28850 , n28537 );
buf ( n28851 , n28544 );
nand ( n28852 , n28850 , n28851 );
buf ( n28853 , n28852 );
buf ( n28854 , n28853 );
nand ( n28855 , n28849 , n28854 );
buf ( n28856 , n28855 );
buf ( n28857 , n28856 );
xor ( n28858 , n28832 , n28857 );
buf ( n28859 , n2541 );
not ( n28860 , n28859 );
and ( n28861 , n594 , n10861 );
not ( n28862 , n594 );
and ( n28863 , n28862 , n10858 );
or ( n28864 , n28861 , n28863 );
buf ( n28865 , n28864 );
not ( n28866 , n28865 );
or ( n28867 , n28860 , n28866 );
not ( n28868 , n9524 );
buf ( n28869 , n28868 );
buf ( n28870 , n2659 );
and ( n28871 , n28869 , n28870 );
buf ( n28872 , n28868 );
buf ( n28873 , n2666 );
nor ( n28874 , n28872 , n28873 );
buf ( n28875 , n28874 );
buf ( n28876 , n28875 );
nor ( n28877 , n28871 , n28876 );
buf ( n28878 , n28877 );
buf ( n28879 , n28878 );
nand ( n28880 , n28867 , n28879 );
buf ( n28881 , n28880 );
buf ( n28882 , n28881 );
xor ( n28883 , n28858 , n28882 );
buf ( n28884 , n28883 );
buf ( n28885 , n28884 );
xor ( n28886 , n28827 , n28885 );
buf ( n28887 , n28886 );
buf ( n28888 , n28887 );
xor ( n28889 , n28803 , n28888 );
buf ( n28890 , n28889 );
buf ( n28891 , n28890 );
xor ( n28892 , n28604 , n28688 );
and ( n28893 , n28892 , n28695 );
and ( n28894 , n28604 , n28688 );
or ( n28895 , n28893 , n28894 );
buf ( n28896 , n28895 );
buf ( n28897 , n28896 );
xor ( n28898 , n28891 , n28897 );
xor ( n28899 , n28638 , n28644 );
and ( n28900 , n28899 , n28685 );
and ( n28901 , n28638 , n28644 );
or ( n28902 , n28900 , n28901 );
buf ( n28903 , n28902 );
buf ( n28904 , n28903 );
buf ( n28905 , n604 );
not ( n28906 , n28905 );
not ( n28907 , n28243 );
buf ( n28908 , n28907 );
not ( n28909 , n28908 );
or ( n28910 , n28906 , n28909 );
not ( n28911 , n604 );
nand ( n28912 , n28911 , n28243 );
buf ( n28913 , n28912 );
nand ( n28914 , n28910 , n28913 );
buf ( n28915 , n28914 );
not ( n28916 , n28915 );
not ( n28917 , n7790 );
or ( n28918 , n28916 , n28917 );
nand ( n28919 , n28574 , n8581 );
nand ( n28920 , n28918 , n28919 );
buf ( n28921 , n28920 );
xor ( n28922 , n28469 , n28486 );
and ( n28923 , n28922 , n28502 );
and ( n28924 , n28469 , n28486 );
or ( n28925 , n28923 , n28924 );
buf ( n28926 , n28925 );
buf ( n28927 , n28926 );
xor ( n28928 , n28921 , n28927 );
buf ( n28929 , n607 );
not ( n28930 , n28929 );
buf ( n28931 , n606 );
not ( n28932 , n28931 );
buf ( n28933 , n19398 );
not ( n28934 , n28933 );
not ( n28935 , n18196 );
or ( n28936 , n28934 , n28935 );
nand ( n28937 , n18197 , n24462 );
nand ( n28938 , n28936 , n28937 );
buf ( n28939 , n28938 );
not ( n28940 , n28939 );
buf ( n28941 , n28940 );
buf ( n28942 , n28941 );
not ( n28943 , n28942 );
or ( n28944 , n28932 , n28943 );
buf ( n28945 , n28941 );
not ( n28946 , n28945 );
buf ( n28947 , n28946 );
buf ( n28948 , n28947 );
buf ( n28949 , n10836 );
nand ( n28950 , n28948 , n28949 );
buf ( n28951 , n28950 );
buf ( n28952 , n28951 );
nand ( n28953 , n28944 , n28952 );
buf ( n28954 , n28953 );
buf ( n28955 , n28954 );
not ( n28956 , n28955 );
or ( n28957 , n28930 , n28956 );
buf ( n28958 , n28677 );
buf ( n28959 , n10882 );
nand ( n28960 , n28958 , n28959 );
buf ( n28961 , n28960 );
buf ( n28962 , n28961 );
nand ( n28963 , n28957 , n28962 );
buf ( n28964 , n28963 );
buf ( n28965 , n28964 );
xor ( n28966 , n28928 , n28965 );
buf ( n28967 , n28966 );
buf ( n28968 , n28967 );
xor ( n28969 , n28904 , n28968 );
xor ( n28970 , n28463 , n28505 );
and ( n28971 , n28970 , n28588 );
and ( n28972 , n28463 , n28505 );
or ( n28973 , n28971 , n28972 );
buf ( n28974 , n28973 );
buf ( n28975 , n28974 );
xor ( n28976 , n28969 , n28975 );
buf ( n28977 , n28976 );
buf ( n28978 , n28977 );
xor ( n28979 , n28898 , n28978 );
buf ( n28980 , n28979 );
xor ( n28981 , n28591 , n28597 );
and ( n28982 , n28981 , n28698 );
and ( n28983 , n28591 , n28597 );
or ( n28984 , n28982 , n28983 );
buf ( n28985 , n28984 );
or ( n28986 , n28980 , n28985 );
not ( n28987 , n28986 );
not ( n28988 , n28022 );
not ( n28989 , n28282 );
not ( n28990 , n28291 );
or ( n28991 , n28989 , n28990 );
not ( n28992 , n28700 );
nand ( n28993 , n28992 , n28453 );
nand ( n28994 , n28991 , n28993 );
nor ( n28995 , n28994 , n27586 );
not ( n28996 , n28995 );
or ( n28997 , n28988 , n28996 );
not ( n28998 , n28994 );
and ( n28999 , n28998 , n28036 );
buf ( n29000 , n28282 );
buf ( n29001 , n28291 );
nor ( n29002 , n29000 , n29001 );
buf ( n29003 , n29002 );
buf ( n29004 , n29003 );
not ( n29005 , n29004 );
buf ( n29006 , n28713 );
not ( n29007 , n29006 );
or ( n29008 , n29005 , n29007 );
buf ( n29009 , n28709 );
nand ( n29010 , n29008 , n29009 );
buf ( n29011 , n29010 );
nor ( n29012 , n28999 , n29011 );
nand ( n29013 , n28997 , n29012 );
not ( n29014 , n29013 );
or ( n29015 , n28987 , n29014 );
nand ( n29016 , n28980 , n28985 );
buf ( n29017 , n29016 );
nand ( n29018 , n29015 , n29017 );
not ( n29019 , n825 );
or ( n29020 , n2371 , n26676 );
nand ( n29021 , n26676 , n2371 );
nand ( n29022 , n29020 , n29021 );
not ( n29023 , n29022 );
or ( n29024 , n29019 , n29023 );
buf ( n29025 , n13611 );
buf ( n29026 , n2845 );
and ( n29027 , n29025 , n29026 );
buf ( n29028 , n27787 );
buf ( n29029 , n2843 );
and ( n29030 , n29028 , n29029 );
nor ( n29031 , n29027 , n29030 );
buf ( n29032 , n29031 );
nand ( n29033 , n29024 , n29032 );
buf ( n29034 , n29033 );
buf ( n29035 , n28180 );
buf ( n29036 , n11237 );
nor ( n29037 , n29035 , n29036 );
buf ( n29038 , n29037 );
buf ( n29039 , n29038 );
buf ( n29040 , n26737 );
buf ( n29041 , n11248 );
and ( n29042 , n29040 , n29041 );
buf ( n29043 , n29042 );
buf ( n29044 , n29043 );
nor ( n29045 , n29039 , n29044 );
buf ( n29046 , n29045 );
buf ( n29047 , n29046 );
not ( n29048 , n598 );
not ( n29049 , n26786 );
or ( n29050 , n29048 , n29049 );
buf ( n29051 , n26782 );
buf ( n29052 , n818 );
nand ( n29053 , n29051 , n29052 );
buf ( n29054 , n29053 );
nand ( n29055 , n29050 , n29054 );
buf ( n29056 , n29055 );
buf ( n29057 , n5550 );
nand ( n29058 , n29056 , n29057 );
buf ( n29059 , n29058 );
buf ( n29060 , n29059 );
nand ( n29061 , n29047 , n29060 );
buf ( n29062 , n29061 );
buf ( n29063 , n29062 );
xor ( n29064 , n29034 , n29063 );
not ( n29065 , n2915 );
not ( n29066 , n600 );
not ( n29067 , n26062 );
or ( n29068 , n29066 , n29067 );
nand ( n29069 , n26053 , n27227 );
nand ( n29070 , n29068 , n29069 );
not ( n29071 , n29070 );
or ( n29072 , n29065 , n29071 );
nand ( n29073 , n28788 , n5430 );
nand ( n29074 , n29072 , n29073 );
buf ( n29075 , n29074 );
xor ( n29076 , n29064 , n29075 );
buf ( n29077 , n29076 );
buf ( n29078 , n29077 );
xor ( n29079 , n28820 , n28826 );
and ( n29080 , n29079 , n28885 );
and ( n29081 , n28820 , n28826 );
or ( n29082 , n29080 , n29081 );
buf ( n29083 , n29082 );
buf ( n29084 , n29083 );
xor ( n29085 , n29078 , n29084 );
buf ( n29086 , n602 );
not ( n29087 , n29086 );
buf ( n29088 , n26088 );
not ( n29089 , n29088 );
or ( n29090 , n29087 , n29089 );
buf ( n29091 , n28211 );
buf ( n29092 , n2912 );
nand ( n29093 , n29091 , n29092 );
buf ( n29094 , n29093 );
buf ( n29095 , n29094 );
nand ( n29096 , n29090 , n29095 );
buf ( n29097 , n29096 );
not ( n29098 , n29097 );
not ( n29099 , n7619 );
or ( n29100 , n29098 , n29099 );
and ( n29101 , n18191 , n26693 );
not ( n29102 , n18191 );
and ( n29103 , n29102 , n26682 );
nor ( n29104 , n29101 , n29103 );
nand ( n29105 , n29100 , n29104 );
buf ( n29106 , n29105 );
and ( n29107 , n28534 , n28535 );
buf ( n29108 , n29107 );
buf ( n29109 , n29108 );
buf ( n29110 , n2452 );
not ( n29111 , n29110 );
and ( n29112 , n592 , n9524 );
not ( n29113 , n592 );
and ( n29114 , n29113 , n9527 );
or ( n29115 , n29112 , n29114 );
buf ( n29116 , n29115 );
not ( n29117 , n29116 );
or ( n29118 , n29111 , n29117 );
buf ( n29119 , n28846 );
buf ( n29120 , n28544 );
nand ( n29121 , n29119 , n29120 );
buf ( n29122 , n29121 );
buf ( n29123 , n29122 );
nand ( n29124 , n29118 , n29123 );
buf ( n29125 , n29124 );
buf ( n29126 , n29125 );
xor ( n29127 , n29109 , n29126 );
buf ( n29128 , n2592 );
not ( n29129 , n29128 );
buf ( n29130 , n28864 );
not ( n29131 , n29130 );
or ( n29132 , n29129 , n29131 );
buf ( n29133 , n10829 );
buf ( n29134 , n26377 );
and ( n29135 , n29133 , n29134 );
not ( n29136 , n29133 );
buf ( n29137 , n26386 );
and ( n29138 , n29136 , n29137 );
nor ( n29139 , n29135 , n29138 );
buf ( n29140 , n29139 );
buf ( n29141 , n29140 );
nand ( n29142 , n29132 , n29141 );
buf ( n29143 , n29142 );
buf ( n29144 , n29143 );
xor ( n29145 , n29127 , n29144 );
buf ( n29146 , n29145 );
buf ( n29147 , n29146 );
xor ( n29148 , n29106 , n29147 );
buf ( n29149 , n8581 );
not ( n29150 , n29149 );
buf ( n29151 , n28915 );
not ( n29152 , n29151 );
or ( n29153 , n29150 , n29152 );
xor ( n29154 , n604 , n28664 );
buf ( n29155 , n29154 );
buf ( n29156 , n7790 );
nand ( n29157 , n29155 , n29156 );
buf ( n29158 , n29157 );
buf ( n29159 , n29158 );
nand ( n29160 , n29153 , n29159 );
buf ( n29161 , n29160 );
buf ( n29162 , n29161 );
xor ( n29163 , n29148 , n29162 );
buf ( n29164 , n29163 );
buf ( n29165 , n29164 );
xor ( n29166 , n29085 , n29165 );
buf ( n29167 , n29166 );
buf ( n29168 , n29167 );
xor ( n29169 , n28921 , n28927 );
and ( n29170 , n29169 , n28965 );
and ( n29171 , n28921 , n28927 );
or ( n29172 , n29170 , n29171 );
buf ( n29173 , n29172 );
buf ( n29174 , n29173 );
xor ( n29175 , n28832 , n28857 );
and ( n29176 , n29175 , n28882 );
and ( n29177 , n28832 , n28857 );
or ( n29178 , n29176 , n29177 );
buf ( n29179 , n29178 );
buf ( n29180 , n29179 );
xor ( n29181 , n28758 , n28782 );
and ( n29182 , n29181 , n28793 );
and ( n29183 , n28758 , n28782 );
or ( n29184 , n29182 , n29183 );
buf ( n29185 , n29184 );
buf ( n29186 , n29185 );
xor ( n29187 , n29180 , n29186 );
buf ( n29188 , n10882 );
not ( n29189 , n29188 );
buf ( n29190 , n28954 );
not ( n29191 , n29190 );
or ( n29192 , n29189 , n29191 );
buf ( n29193 , n607 );
buf ( n29194 , n606 );
not ( n29195 , n29194 );
not ( n29196 , n17997 );
nand ( n29197 , n18139 , n18038 , n26050 );
not ( n29198 , n29197 );
or ( n29199 , n29196 , n29198 );
nand ( n29200 , n24512 , n18038 , n18139 , n26050 );
nand ( n29201 , n29199 , n29200 );
buf ( n29202 , n29201 );
not ( n29203 , n29202 );
buf ( n29204 , n29203 );
not ( n29205 , n29204 );
or ( n29206 , n29195 , n29205 );
buf ( n29207 , n29202 );
buf ( n29208 , n10836 );
nand ( n29209 , n29207 , n29208 );
buf ( n29210 , n29209 );
buf ( n29211 , n29210 );
nand ( n29212 , n29206 , n29211 );
buf ( n29213 , n29212 );
buf ( n29214 , n29213 );
nand ( n29215 , n29193 , n29214 );
buf ( n29216 , n29215 );
buf ( n29217 , n29216 );
nand ( n29218 , n29192 , n29217 );
buf ( n29219 , n29218 );
buf ( n29220 , n29219 );
xor ( n29221 , n29187 , n29220 );
buf ( n29222 , n29221 );
buf ( n29223 , n29222 );
xor ( n29224 , n29174 , n29223 );
xor ( n29225 , n28796 , n28802 );
and ( n29226 , n29225 , n28888 );
and ( n29227 , n28796 , n28802 );
or ( n29228 , n29226 , n29227 );
buf ( n29229 , n29228 );
buf ( n29230 , n29229 );
xor ( n29231 , n29224 , n29230 );
buf ( n29232 , n29231 );
buf ( n29233 , n29232 );
xor ( n29234 , n29168 , n29233 );
xor ( n29235 , n28904 , n28968 );
and ( n29236 , n29235 , n28975 );
and ( n29237 , n28904 , n28968 );
or ( n29238 , n29236 , n29237 );
buf ( n29239 , n29238 );
buf ( n29240 , n29239 );
xor ( n29241 , n29234 , n29240 );
buf ( n29242 , n29241 );
buf ( n29243 , n29242 );
xor ( n29244 , n28891 , n28897 );
and ( n29245 , n29244 , n28978 );
and ( n29246 , n28891 , n28897 );
or ( n29247 , n29245 , n29246 );
buf ( n29248 , n29247 );
buf ( n29249 , n29248 );
nor ( n29250 , n29243 , n29249 );
buf ( n29251 , n29250 );
buf ( n29252 , n29251 );
buf ( n29253 , n29252 );
buf ( n29254 , n29253 );
not ( n29255 , n29254 );
buf ( n29256 , n29242 );
buf ( n29257 , n29256 );
buf ( n29258 , n29257 );
buf ( n29259 , n29258 );
buf ( n29260 , n29248 );
nand ( n29261 , n29259 , n29260 );
buf ( n29262 , n29261 );
and ( n29263 , n29255 , n29262 );
and ( n29264 , n29018 , n29263 );
not ( n29265 , n29018 );
nand ( n29266 , n29255 , n29262 );
and ( n29267 , n29265 , n29266 );
nor ( n29268 , n29264 , n29267 );
buf ( n29269 , n29268 );
buf ( n29270 , n29269 );
buf ( n29271 , n29270 );
xor ( n29272 , n28745 , n29271 );
buf ( n29273 , n29272 );
buf ( n29274 , n29273 );
buf ( n29275 , n17269 );
buf ( n29276 , n17320 );
xor ( n29277 , n29275 , n29276 );
not ( n29278 , n29013 );
nand ( n29279 , n29016 , n28986 );
and ( n29280 , n29278 , n29279 );
not ( n29281 , n29278 );
not ( n29282 , n29279 );
and ( n29283 , n29281 , n29282 );
nor ( n29284 , n29280 , n29283 );
buf ( n29285 , n29284 );
buf ( n29286 , n29285 );
buf ( n29287 , n29286 );
buf ( n29288 , n29287 );
buf ( n29289 , n29288 );
buf ( n29290 , n29289 );
buf ( n29291 , n29290 );
buf ( n29292 , n29291 );
and ( n29293 , n29277 , n29292 );
and ( n29294 , n29275 , n29276 );
or ( n29295 , n29293 , n29294 );
buf ( n29296 , n29295 );
buf ( n29297 , n29296 );
xor ( n29298 , n29274 , n29297 );
buf ( n29299 , n28732 );
xor ( n29300 , n29275 , n29276 );
xor ( n29301 , n29300 , n29292 );
buf ( n29302 , n29301 );
buf ( n29303 , n29302 );
xor ( n29304 , n29299 , n29303 );
buf ( n29305 , n28727 );
buf ( n29306 , n28315 );
xor ( n29307 , n29305 , n29306 );
xor ( n29308 , n16319 , n16313 );
buf ( n29309 , n27121 );
buf ( n29310 , n27351 );
or ( n29311 , n29309 , n29310 );
buf ( n29312 , n29311 );
nand ( n29313 , n29312 , n27354 );
not ( n29314 , n29313 );
not ( n29315 , n27585 );
not ( n29316 , n28022 );
or ( n29317 , n29315 , n29316 );
nand ( n29318 , n27357 , n27583 );
nand ( n29319 , n29317 , n29318 );
not ( n29320 , n29319 );
not ( n29321 , n29320 );
or ( n29322 , n29314 , n29321 );
not ( n29323 , n29313 );
nand ( n29324 , n29319 , n29323 );
nand ( n29325 , n29322 , n29324 );
buf ( n29326 , n29325 );
not ( n29327 , n29326 );
buf ( n29328 , n29327 );
and ( n29329 , n29308 , n29328 );
and ( n29330 , n16319 , n16313 );
or ( n29331 , n29329 , n29330 );
buf ( n29332 , n29331 );
buf ( n29333 , n28310 );
xor ( n29334 , n29332 , n29333 );
buf ( n29335 , n15922 );
buf ( n29336 , n15937 );
xor ( n29337 , n29335 , n29336 );
buf ( n29338 , n27585 );
buf ( n29339 , n29318 );
nand ( n29340 , n29338 , n29339 );
buf ( n29341 , n29340 );
buf ( n29342 , n29341 );
not ( n29343 , n29342 );
buf ( n29344 , n29343 );
not ( n29345 , n29344 );
buf ( n29346 , n28022 );
buf ( n29347 , n29346 );
buf ( n29348 , n29347 );
buf ( n29349 , n29348 );
not ( n29350 , n29349 );
buf ( n29351 , n29350 );
not ( n29352 , n29351 );
or ( n29353 , n29345 , n29352 );
buf ( n29354 , n29348 );
buf ( n29355 , n29341 );
nand ( n29356 , n29354 , n29355 );
buf ( n29357 , n29356 );
nand ( n29358 , n29353 , n29357 );
not ( n29359 , n29358 );
not ( n29360 , n29359 );
buf ( n29361 , n29360 );
and ( n29362 , n29337 , n29361 );
and ( n29363 , n29335 , n29336 );
or ( n29364 , n29362 , n29363 );
buf ( n29365 , n29364 );
buf ( n29366 , n29365 );
xor ( n29367 , n15615 , n15499 );
not ( n29368 , n28394 );
not ( n29369 , n28389 );
or ( n29370 , n29368 , n29369 );
nand ( n29371 , n29370 , n28400 );
buf ( n29372 , n28015 );
buf ( n29373 , n29372 );
buf ( n29374 , n29373 );
nand ( n29375 , n29374 , n28010 );
not ( n29376 , n29375 );
and ( n29377 , n29371 , n29376 );
not ( n29378 , n29371 );
and ( n29379 , n29378 , n29375 );
nor ( n29380 , n29377 , n29379 );
and ( n29381 , n29367 , n29380 );
and ( n29382 , n15615 , n15499 );
or ( n29383 , n29381 , n29382 );
buf ( n29384 , n29383 );
xor ( n29385 , n29335 , n29336 );
xor ( n29386 , n29385 , n29361 );
buf ( n29387 , n29386 );
buf ( n29388 , n29387 );
xor ( n29389 , n29384 , n29388 );
buf ( n29390 , n28415 );
not ( n29391 , n29390 );
xor ( n29392 , n14707 , n14696 );
not ( n29393 , n27981 );
and ( n29394 , n29393 , n27992 );
not ( n29395 , n29394 );
not ( n29396 , n27967 );
not ( n29397 , n27767 );
or ( n29398 , n29396 , n29397 );
nand ( n29399 , n29398 , n27986 );
not ( n29400 , n29399 );
not ( n29401 , n29400 );
or ( n29402 , n29395 , n29401 );
not ( n29403 , n29394 );
nand ( n29404 , n29403 , n29399 );
nand ( n29405 , n29402 , n29404 );
not ( n29406 , n29405 );
not ( n29407 , n29406 );
and ( n29408 , n29392 , n29407 );
and ( n29409 , n14707 , n14696 );
or ( n29410 , n29408 , n29409 );
buf ( n29411 , n29410 );
not ( n29412 , n29411 );
buf ( n29413 , n29412 );
buf ( n29414 , n29413 );
nand ( n29415 , n29391 , n29414 );
buf ( n29416 , n29415 );
buf ( n29417 , n29416 );
not ( n29418 , n29417 );
xor ( n29419 , n14707 , n14696 );
xor ( n29420 , n29419 , n29407 );
buf ( n29421 , n29420 );
not ( n29422 , n29421 );
buf ( n29423 , n28377 );
not ( n29424 , n29423 );
buf ( n29425 , n29424 );
buf ( n29426 , n29425 );
nand ( n29427 , n29422 , n29426 );
buf ( n29428 , n29427 );
buf ( n29429 , n29428 );
not ( n29430 , n29429 );
buf ( n29431 , n28348 );
not ( n29432 , n29431 );
buf ( n29433 , n28326 );
not ( n29434 , n29433 );
buf ( n29435 , n29434 );
buf ( n29436 , n29435 );
nand ( n29437 , n29432 , n29436 );
buf ( n29438 , n29437 );
xor ( n29439 , n13686 , n10577 );
xor ( n29440 , n29439 , n13652 );
not ( n29441 , n29440 );
not ( n29442 , n28353 );
nand ( n29443 , n29441 , n29442 );
and ( n29444 , n29438 , n29443 );
not ( n29445 , n29444 );
buf ( n29446 , n13679 );
buf ( n29447 , n8325 );
buf ( n29448 , n29447 );
buf ( n29449 , n29448 );
xor ( n29450 , n29446 , n29449 );
not ( n29451 , n12794 );
not ( n29452 , n29451 );
not ( n29453 , n12788 );
not ( n29454 , n29453 );
or ( n29455 , n29452 , n29454 );
nand ( n29456 , n29455 , n12802 );
not ( n29457 , n29456 );
buf ( n29458 , n12766 );
not ( n29459 , n29458 );
or ( n29460 , n29457 , n29459 );
or ( n29461 , n29458 , n29456 );
nand ( n29462 , n29460 , n29461 );
buf ( n29463 , n29462 );
buf ( n29464 , n29463 );
xor ( n29465 , n29450 , n29464 );
buf ( n29466 , n29465 );
buf ( n29467 , n29466 );
not ( n29468 , n29467 );
buf ( n29469 , n28439 );
not ( n29470 , n29469 );
buf ( n29471 , n29470 );
buf ( n29472 , n29471 );
nand ( n29473 , n29468 , n29472 );
buf ( n29474 , n29473 );
buf ( n29475 , n29474 );
not ( n29476 , n29475 );
buf ( n29477 , n28434 );
buf ( n29478 , n6186 );
buf ( n29479 , n13668 );
xor ( n29480 , n29478 , n29479 );
buf ( n29481 , n11819 );
not ( n29482 , n29481 );
buf ( n29483 , n12758 );
nand ( n29484 , n29482 , n29483 );
buf ( n29485 , n29484 );
buf ( n29486 , n29485 );
buf ( n29487 , n12755 );
buf ( n29488 , n29487 );
buf ( n29489 , n29488 );
buf ( n29490 , n29489 );
not ( n29491 , n29490 );
buf ( n29492 , n29491 );
buf ( n29493 , n29492 );
and ( n29494 , n29486 , n29493 );
not ( n29495 , n29486 );
buf ( n29496 , n29489 );
and ( n29497 , n29495 , n29496 );
nor ( n29498 , n29494 , n29497 );
buf ( n29499 , n29498 );
buf ( n29500 , n29499 );
buf ( n29501 , n29500 );
and ( n29502 , n29480 , n29501 );
and ( n29503 , n29478 , n29479 );
or ( n29504 , n29502 , n29503 );
buf ( n29505 , n29504 );
buf ( n29506 , n29505 );
or ( n29507 , n29477 , n29506 );
xor ( n29508 , n29478 , n29479 );
xor ( n29509 , n29508 , n29501 );
buf ( n29510 , n29509 );
not ( n29511 , n29510 );
buf ( n29512 , n5951 );
buf ( n29513 , n13669 );
xor ( n29514 , n29512 , n29513 );
buf ( n29515 , n12745 );
not ( n29516 , n29515 );
buf ( n29517 , n12735 );
not ( n29518 , n29517 );
buf ( n29519 , n29518 );
buf ( n29520 , n29519 );
not ( n29521 , n29520 );
or ( n29522 , n29516 , n29521 );
buf ( n29523 , n12754 );
nand ( n29524 , n29522 , n29523 );
buf ( n29525 , n29524 );
buf ( n29526 , n29525 );
buf ( n29527 , n12731 );
not ( n29528 , n29527 );
buf ( n29529 , n29528 );
and ( n29530 , n29526 , n29529 );
not ( n29531 , n29526 );
buf ( n29532 , n29527 );
and ( n29533 , n29531 , n29532 );
nor ( n29534 , n29530 , n29533 );
buf ( n29535 , n29534 );
buf ( n29536 , n29535 );
xor ( n29537 , n29514 , n29536 );
buf ( n29538 , n29537 );
buf ( n29539 , n29538 );
buf ( n29540 , n26042 );
or ( n29541 , n29539 , n29540 );
buf ( n29542 , n29541 );
buf ( n29543 , n29542 );
not ( n29544 , n29543 );
buf ( n29545 , n25986 );
buf ( n29546 , n26001 );
xor ( n29547 , n29545 , n29546 );
buf ( n29548 , n25960 );
not ( n29549 , n29548 );
buf ( n29550 , n25981 );
not ( n29551 , n29550 );
or ( n29552 , n29549 , n29551 );
buf ( n29553 , n25960 );
buf ( n29554 , n25981 );
or ( n29555 , n29553 , n29554 );
buf ( n29556 , n25955 );
buf ( n29557 , n25947 );
or ( n29558 , n29556 , n29557 );
buf ( n29559 , n25942 );
buf ( n29560 , n25934 );
or ( n29561 , n29559 , n29560 );
buf ( n29562 , n25888 );
buf ( n29563 , n28738 );
buf ( n29564 , n1319 );
buf ( n29565 , n1412 );
not ( n29566 , n29565 );
buf ( n29567 , n29566 );
buf ( n29568 , n29567 );
xor ( n29569 , n29564 , n29568 );
buf ( n29570 , n1467 );
buf ( n29571 , n1539 );
xor ( n29572 , n29570 , n29571 );
buf ( n29573 , n1502 );
and ( n29574 , n29572 , n29573 );
or ( n29575 , n29574 , C0 );
buf ( n29576 , n29575 );
buf ( n29577 , n29576 );
and ( n29578 , n29569 , n29577 );
and ( n29579 , n29564 , n29568 );
or ( n29580 , n29578 , n29579 );
buf ( n29581 , n29580 );
buf ( n29582 , n29581 );
buf ( n29583 , n1412 );
xor ( n29584 , n29582 , n29583 );
buf ( n29585 , n28736 );
and ( n29586 , n29584 , n29585 );
and ( n29587 , n29582 , n29583 );
or ( n29588 , n29586 , n29587 );
buf ( n29589 , n29588 );
buf ( n29590 , n29589 );
xor ( n29591 , n29563 , n29590 );
buf ( n29592 , n25883 );
and ( n29593 , n29591 , n29592 );
and ( n29594 , n29563 , n29590 );
or ( n29595 , n29593 , n29594 );
buf ( n29596 , n29595 );
buf ( n29597 , n29596 );
xor ( n29598 , n29562 , n29597 );
buf ( n29599 , n25904 );
and ( n29600 , n29598 , n29599 );
and ( n29601 , n29562 , n29597 );
or ( n29602 , n29600 , n29601 );
buf ( n29603 , n29602 );
buf ( n29604 , n29603 );
not ( n29605 , n29604 );
buf ( n29606 , n29605 );
buf ( n29607 , n29606 );
buf ( n29608 , n25929 );
buf ( n29609 , n25909 );
nor ( n29610 , n29608 , n29609 );
buf ( n29611 , n29610 );
buf ( n29612 , n29611 );
or ( n29613 , n29607 , n29612 );
buf ( n29614 , n25929 );
buf ( n29615 , n25909 );
nand ( n29616 , n29614 , n29615 );
buf ( n29617 , n29616 );
buf ( n29618 , n29617 );
nand ( n29619 , n29613 , n29618 );
buf ( n29620 , n29619 );
buf ( n29621 , n29620 );
nand ( n29622 , n29561 , n29621 );
buf ( n29623 , n29622 );
buf ( n29624 , n29623 );
buf ( n29625 , n25942 );
buf ( n29626 , n25934 );
nand ( n29627 , n29625 , n29626 );
buf ( n29628 , n29627 );
buf ( n29629 , n29628 );
nand ( n29630 , n29624 , n29629 );
buf ( n29631 , n29630 );
buf ( n29632 , n29631 );
nand ( n29633 , n29558 , n29632 );
buf ( n29634 , n29633 );
buf ( n29635 , n29634 );
buf ( n29636 , n25947 );
buf ( n29637 , n25955 );
nand ( n29638 , n29636 , n29637 );
buf ( n29639 , n29638 );
buf ( n29640 , n29639 );
nand ( n29641 , n29635 , n29640 );
buf ( n29642 , n29641 );
buf ( n29643 , n29642 );
nand ( n29644 , n29555 , n29643 );
buf ( n29645 , n29644 );
buf ( n29646 , n29645 );
nand ( n29647 , n29552 , n29646 );
buf ( n29648 , n29647 );
buf ( n29649 , n29648 );
and ( n29650 , n29547 , n29649 );
and ( n29651 , n29545 , n29546 );
or ( n29652 , n29650 , n29651 );
buf ( n29653 , n29652 );
buf ( n29654 , n29653 );
not ( n29655 , n29654 );
buf ( n29656 , n29655 );
buf ( n29657 , n26037 );
buf ( n29658 , n26006 );
nor ( n29659 , n29657 , n29658 );
buf ( n29660 , n29659 );
or ( n29661 , n29656 , n29660 );
buf ( n29662 , n26037 );
buf ( n29663 , n26006 );
nand ( n29664 , n29662 , n29663 );
buf ( n29665 , n29664 );
nand ( n29666 , n29661 , n29665 );
buf ( n29667 , n29666 );
not ( n29668 , n29667 );
or ( n29669 , n29544 , n29668 );
buf ( n29670 , n29538 );
buf ( n29671 , n26042 );
nand ( n29672 , n29670 , n29671 );
buf ( n29673 , n29672 );
buf ( n29674 , n29673 );
nand ( n29675 , n29669 , n29674 );
buf ( n29676 , n29675 );
xor ( n29677 , n29512 , n29513 );
and ( n29678 , n29677 , n29536 );
and ( n29679 , n29512 , n29513 );
or ( n29680 , n29678 , n29679 );
buf ( n29681 , n29680 );
or ( n29682 , n29676 , n29681 );
not ( n29683 , n29682 );
or ( n29684 , n29511 , n29683 );
nand ( n29685 , n29676 , n29681 );
nand ( n29686 , n29684 , n29685 );
buf ( n29687 , n29686 );
nand ( n29688 , n29507 , n29687 );
buf ( n29689 , n29688 );
buf ( n29690 , n29689 );
buf ( n29691 , n28434 );
buf ( n29692 , n29505 );
nand ( n29693 , n29691 , n29692 );
buf ( n29694 , n29693 );
buf ( n29695 , n29694 );
nand ( n29696 , n29690 , n29695 );
buf ( n29697 , n29696 );
buf ( n29698 , n29697 );
not ( n29699 , n29698 );
or ( n29700 , n29476 , n29699 );
buf ( n29701 , n29466 );
buf ( n29702 , n28439 );
nand ( n29703 , n29701 , n29702 );
buf ( n29704 , n29703 );
buf ( n29705 , n29704 );
nand ( n29706 , n29700 , n29705 );
buf ( n29707 , n29706 );
buf ( n29708 , n29707 );
not ( n29709 , n29708 );
buf ( n29710 , n29709 );
buf ( n29711 , n29710 );
buf ( n29712 , n28321 );
xor ( n29713 , n29446 , n29449 );
and ( n29714 , n29713 , n29464 );
and ( n29715 , n29446 , n29449 );
or ( n29716 , n29714 , n29715 );
buf ( n29717 , n29716 );
buf ( n29718 , n29717 );
nor ( n29719 , n29712 , n29718 );
buf ( n29720 , n29719 );
buf ( n29721 , n29720 );
or ( n29722 , n29711 , n29721 );
buf ( n29723 , n28321 );
buf ( n29724 , n29717 );
nand ( n29725 , n29723 , n29724 );
buf ( n29726 , n29725 );
buf ( n29727 , n29726 );
nand ( n29728 , n29722 , n29727 );
buf ( n29729 , n29728 );
not ( n29730 , n29729 );
or ( n29731 , n29445 , n29730 );
buf ( n29732 , n28348 );
buf ( n29733 , n28326 );
nand ( n29734 , n29732 , n29733 );
buf ( n29735 , n29734 );
not ( n29736 , n29735 );
and ( n29737 , n29443 , n29736 );
and ( n29738 , n29440 , n28353 );
nor ( n29739 , n29737 , n29738 );
nand ( n29740 , n29731 , n29739 );
not ( n29741 , n29740 );
xor ( n29742 , n13415 , n13236 );
not ( n29743 , n13640 );
not ( n29744 , n12832 );
or ( n29745 , n29743 , n29744 );
buf ( n29746 , n13648 );
nand ( n29747 , n29745 , n29746 );
nand ( n29748 , n27747 , n27760 );
not ( n29749 , n29748 );
and ( n29750 , n29747 , n29749 );
not ( n29751 , n29747 );
and ( n29752 , n29751 , n29748 );
nor ( n29753 , n29750 , n29752 );
buf ( n29754 , n29753 );
and ( n29755 , n29742 , n29754 );
and ( n29756 , n13415 , n13236 );
or ( n29757 , n29755 , n29756 );
buf ( n29758 , n29757 );
not ( n29759 , n29758 );
buf ( n29760 , n29759 );
buf ( n29761 , n28372 );
not ( n29762 , n29761 );
buf ( n29763 , n29762 );
nand ( n29764 , n29760 , n29763 );
xor ( n29765 , n13686 , n10577 );
and ( n29766 , n29765 , n13652 );
and ( n29767 , n13686 , n10577 );
or ( n29768 , n29766 , n29767 );
not ( n29769 , n29768 );
xor ( n29770 , n13415 , n13236 );
xor ( n29771 , n29770 , n29754 );
buf ( n29772 , n29771 );
not ( n29773 , n29772 );
buf ( n29774 , n29773 );
nand ( n29775 , n29769 , n29774 );
and ( n29776 , n29764 , n29775 );
not ( n29777 , n29776 );
or ( n29778 , n29741 , n29777 );
nand ( n29779 , n29771 , n29768 );
not ( n29780 , n29779 );
and ( n29781 , n29764 , n29780 );
buf ( n29782 , n29763 );
not ( n29783 , n29782 );
buf ( n29784 , n29783 );
and ( n29785 , n29757 , n29784 );
nor ( n29786 , n29781 , n29785 );
nand ( n29787 , n29778 , n29786 );
buf ( n29788 , n29787 );
not ( n29789 , n29788 );
or ( n29790 , n29430 , n29789 );
buf ( n29791 , n29420 );
buf ( n29792 , n29425 );
not ( n29793 , n29792 );
buf ( n29794 , n29793 );
buf ( n29795 , n29794 );
nand ( n29796 , n29791 , n29795 );
buf ( n29797 , n29796 );
buf ( n29798 , n29797 );
nand ( n29799 , n29790 , n29798 );
buf ( n29800 , n29799 );
buf ( n29801 , n29800 );
not ( n29802 , n29801 );
or ( n29803 , n29418 , n29802 );
buf ( n29804 , n28415 );
buf ( n29805 , n29410 );
nand ( n29806 , n29804 , n29805 );
buf ( n29807 , n29806 );
buf ( n29808 , n29807 );
nand ( n29809 , n29803 , n29808 );
buf ( n29810 , n29809 );
buf ( n29811 , n29810 );
not ( n29812 , n29811 );
xor ( n29813 , n15615 , n15499 );
xor ( n29814 , n29813 , n29380 );
buf ( n29815 , n29814 );
not ( n29816 , n29815 );
buf ( n29817 , n28420 );
not ( n29818 , n29817 );
buf ( n29819 , n29818 );
buf ( n29820 , n29819 );
nand ( n29821 , n29816 , n29820 );
buf ( n29822 , n29821 );
buf ( n29823 , n29822 );
not ( n29824 , n29823 );
or ( n29825 , n29812 , n29824 );
buf ( n29826 , n28420 );
buf ( n29827 , n29814 );
nand ( n29828 , n29826 , n29827 );
buf ( n29829 , n29828 );
buf ( n29830 , n29829 );
nand ( n29831 , n29825 , n29830 );
buf ( n29832 , n29831 );
buf ( n29833 , n29832 );
and ( n29834 , n29389 , n29833 );
and ( n29835 , n29384 , n29388 );
or ( n29836 , n29834 , n29835 );
buf ( n29837 , n29836 );
buf ( n29838 , n29837 );
xor ( n29839 , n29366 , n29838 );
xor ( n29840 , n16319 , n16313 );
xor ( n29841 , n29840 , n29328 );
buf ( n29842 , n29841 );
and ( n29843 , n29839 , n29842 );
and ( n29844 , n29366 , n29838 );
or ( n29845 , n29843 , n29844 );
buf ( n29846 , n29845 );
buf ( n29847 , n29846 );
and ( n29848 , n29334 , n29847 );
and ( n29849 , n29332 , n29333 );
or ( n29850 , n29848 , n29849 );
buf ( n29851 , n29850 );
buf ( n29852 , n29851 );
and ( n29853 , n29307 , n29852 );
and ( n29854 , n29305 , n29306 );
or ( n29855 , n29853 , n29854 );
buf ( n29856 , n29855 );
buf ( n29857 , n29856 );
and ( n29858 , n29304 , n29857 );
and ( n29859 , n29299 , n29303 );
or ( n29860 , n29858 , n29859 );
buf ( n29861 , n29860 );
buf ( n29862 , n29861 );
and ( n29863 , n29298 , n29862 );
and ( n29864 , n29274 , n29297 );
or ( n29865 , n29863 , n29864 );
buf ( n29866 , n29865 );
buf ( n29867 , n29866 );
buf ( n29868 , n17663 );
buf ( n29869 , n17670 );
xor ( n29870 , n29868 , n29869 );
buf ( n29871 , n29251 );
buf ( n29872 , n28980 );
buf ( n29873 , n28985 );
nor ( n29874 , n29872 , n29873 );
buf ( n29875 , n29874 );
buf ( n29876 , n29875 );
nor ( n29877 , n29871 , n29876 );
buf ( n29878 , n29877 );
buf ( n29879 , n29878 );
buf ( n29880 , n29879 );
buf ( n29881 , n29880 );
not ( n29882 , n29881 );
not ( n29883 , n29013 );
or ( n29884 , n29882 , n29883 );
buf ( n29885 , n29254 );
not ( n29886 , n29885 );
buf ( n29887 , n29016 );
not ( n29888 , n29887 );
and ( n29889 , n29886 , n29888 );
buf ( n29890 , n29262 );
not ( n29891 , n29890 );
buf ( n29892 , n29891 );
buf ( n29893 , n29892 );
nor ( n29894 , n29889 , n29893 );
buf ( n29895 , n29894 );
nand ( n29896 , n29884 , n29895 );
not ( n29897 , n5550 );
not ( n29898 , n598 );
not ( n29899 , n26851 );
or ( n29900 , n29898 , n29899 );
nand ( n29901 , n26810 , n818 );
nand ( n29902 , n29900 , n29901 );
not ( n29903 , n29902 );
or ( n29904 , n29897 , n29903 );
nand ( n29905 , n29055 , n5631 );
nand ( n29906 , n29904 , n29905 );
buf ( n29907 , n29906 );
buf ( n29908 , n2541 );
not ( n29909 , n29908 );
buf ( n29910 , n594 );
not ( n29911 , n29910 );
buf ( n29912 , n13605 );
not ( n29913 , n29912 );
or ( n29914 , n29911 , n29913 );
buf ( n29915 , n13602 );
buf ( n29916 , n2481 );
nand ( n29917 , n29915 , n29916 );
buf ( n29918 , n29917 );
buf ( n29919 , n29918 );
nand ( n29920 , n29914 , n29919 );
buf ( n29921 , n29920 );
buf ( n29922 , n29921 );
not ( n29923 , n29922 );
or ( n29924 , n29909 , n29923 );
and ( n29925 , n10830 , n2659 );
buf ( n29926 , n10830 );
buf ( n29927 , n2666 );
nor ( n29928 , n29926 , n29927 );
buf ( n29929 , n29928 );
nor ( n29930 , n29925 , n29929 );
buf ( n29931 , n29930 );
nand ( n29932 , n29924 , n29931 );
buf ( n29933 , n29932 );
buf ( n29934 , n29933 );
xor ( n29935 , n29907 , n29934 );
buf ( n29936 , n5430 );
not ( n29937 , n29936 );
buf ( n29938 , n29070 );
not ( n29939 , n29938 );
or ( n29940 , n29937 , n29939 );
buf ( n29941 , n600 );
not ( n29942 , n29941 );
buf ( n29943 , n26088 );
not ( n29944 , n29943 );
or ( n29945 , n29942 , n29944 );
buf ( n29946 , n28211 );
buf ( n29947 , n7650 );
nand ( n29948 , n29946 , n29947 );
buf ( n29949 , n29948 );
buf ( n29950 , n29949 );
nand ( n29951 , n29945 , n29950 );
buf ( n29952 , n29951 );
buf ( n29953 , n29952 );
buf ( n29954 , n2915 );
nand ( n29955 , n29953 , n29954 );
buf ( n29956 , n29955 );
buf ( n29957 , n29956 );
nand ( n29958 , n29940 , n29957 );
buf ( n29959 , n29958 );
buf ( n29960 , n29959 );
xor ( n29961 , n29935 , n29960 );
buf ( n29962 , n29961 );
buf ( n29963 , n29962 );
xor ( n29964 , n29106 , n29147 );
and ( n29965 , n29964 , n29162 );
and ( n29966 , n29106 , n29147 );
or ( n29967 , n29965 , n29966 );
buf ( n29968 , n29967 );
buf ( n29969 , n29968 );
xor ( n29970 , n29963 , n29969 );
buf ( n29971 , n7619 );
not ( n29972 , n29971 );
buf ( n29973 , n602 );
buf ( n29974 , n18191 );
and ( n29975 , n29973 , n29974 );
not ( n29976 , n29973 );
buf ( n29977 , n27000 );
and ( n29978 , n29976 , n29977 );
nor ( n29979 , n29975 , n29978 );
buf ( n29980 , n29979 );
buf ( n29981 , n29980 );
not ( n29982 , n29981 );
or ( n29983 , n29972 , n29982 );
buf ( n29984 , n28247 );
buf ( n29985 , n26693 );
and ( n29986 , n29984 , n29985 );
buf ( n29987 , n28244 );
buf ( n29988 , n26682 );
and ( n29989 , n29987 , n29988 );
nor ( n29990 , n29986 , n29989 );
buf ( n29991 , n29990 );
buf ( n29992 , n29991 );
nand ( n29993 , n29983 , n29992 );
buf ( n29994 , n29993 );
buf ( n29995 , n29994 );
xor ( n29996 , n29109 , n29126 );
and ( n29997 , n29996 , n29144 );
and ( n29998 , n29109 , n29126 );
or ( n29999 , n29997 , n29998 );
buf ( n30000 , n29999 );
buf ( n30001 , n30000 );
xor ( n30002 , n29995 , n30001 );
buf ( n30003 , n607 );
not ( n30004 , n30003 );
buf ( n30005 , n606 );
not ( n30006 , n15683 );
not ( n30007 , n17996 );
not ( n30008 , n18037 );
and ( n30009 , n30006 , n30007 , n30008 );
nand ( n30010 , n18139 , n18140 );
not ( n30011 , n30010 );
and ( n30012 , n24491 , n24493 );
not ( n30013 , n24491 );
and ( n30014 , n30013 , n24492 );
nor ( n30015 , n30012 , n30014 );
not ( n30016 , n30015 );
nand ( n30017 , n30009 , n30011 , n30016 );
or ( n30018 , n15683 , n18037 );
not ( n30019 , n30007 );
or ( n30020 , n30018 , n30019 );
nand ( n30021 , n30020 , n30015 );
nand ( n30022 , n30010 , n30015 );
nand ( n30023 , n30017 , n30021 , n30022 );
buf ( n30024 , n30023 );
buf ( n30025 , n30024 );
buf ( n30026 , n30025 );
buf ( n30027 , n30026 );
and ( n30028 , n30005 , n30027 );
not ( n30029 , n30005 );
buf ( n30030 , n30026 );
not ( n30031 , n30030 );
buf ( n30032 , n30031 );
buf ( n30033 , n30032 );
and ( n30034 , n30029 , n30033 );
nor ( n30035 , n30028 , n30034 );
buf ( n30036 , n30035 );
buf ( n30037 , n30036 );
not ( n30038 , n30037 );
or ( n30039 , n30004 , n30038 );
buf ( n30040 , n29213 );
buf ( n30041 , n10882 );
nand ( n30042 , n30040 , n30041 );
buf ( n30043 , n30042 );
buf ( n30044 , n30043 );
nand ( n30045 , n30039 , n30044 );
buf ( n30046 , n30045 );
buf ( n30047 , n30046 );
xor ( n30048 , n30002 , n30047 );
buf ( n30049 , n30048 );
buf ( n30050 , n30049 );
xor ( n30051 , n29970 , n30050 );
buf ( n30052 , n30051 );
buf ( n30053 , n30052 );
xor ( n30054 , n29174 , n29223 );
and ( n30055 , n30054 , n29230 );
and ( n30056 , n29174 , n29223 );
or ( n30057 , n30055 , n30056 );
buf ( n30058 , n30057 );
buf ( n30059 , n30058 );
xor ( n30060 , n30053 , n30059 );
xor ( n30061 , n29180 , n29186 );
and ( n30062 , n30061 , n29220 );
and ( n30063 , n29180 , n29186 );
or ( n30064 , n30062 , n30063 );
buf ( n30065 , n30064 );
buf ( n30066 , n30065 );
buf ( n30067 , n7790 );
not ( n30068 , n30067 );
and ( n30069 , n604 , n28941 );
not ( n30070 , n604 );
buf ( n30071 , n28938 );
buf ( n30072 , n30071 );
buf ( n30073 , n30072 );
and ( n30074 , n30070 , n30073 );
or ( n30075 , n30069 , n30074 );
buf ( n30076 , n30075 );
not ( n30077 , n30076 );
or ( n30078 , n30068 , n30077 );
buf ( n30079 , n29154 );
buf ( n30080 , n8581 );
nand ( n30081 , n30079 , n30080 );
buf ( n30082 , n30081 );
buf ( n30083 , n30082 );
nand ( n30084 , n30078 , n30083 );
buf ( n30085 , n30084 );
buf ( n30086 , n30085 );
buf ( n30087 , n8553 );
buf ( n30088 , n592 );
and ( n30089 , n30087 , n30088 );
buf ( n30090 , n30089 );
buf ( n30091 , n30090 );
buf ( n30092 , n2452 );
not ( n30093 , n30092 );
buf ( n30094 , n592 );
not ( n30095 , n30094 );
buf ( n30096 , n10861 );
not ( n30097 , n30096 );
or ( n30098 , n30095 , n30097 );
buf ( n30099 , n10858 );
buf ( n30100 , n2416 );
nand ( n30101 , n30099 , n30100 );
buf ( n30102 , n30101 );
buf ( n30103 , n30102 );
nand ( n30104 , n30098 , n30103 );
buf ( n30105 , n30104 );
buf ( n30106 , n30105 );
not ( n30107 , n30106 );
or ( n30108 , n30093 , n30107 );
buf ( n30109 , n28544 );
buf ( n30110 , n29115 );
nand ( n30111 , n30109 , n30110 );
buf ( n30112 , n30111 );
buf ( n30113 , n30112 );
nand ( n30114 , n30108 , n30113 );
buf ( n30115 , n30114 );
buf ( n30116 , n30115 );
xor ( n30117 , n30091 , n30116 );
buf ( n30118 , n825 );
not ( n30119 , n30118 );
not ( n30120 , n596 );
not ( n30121 , n26973 );
or ( n30122 , n30120 , n30121 );
buf ( n30123 , n26737 );
buf ( n30124 , n2371 );
nand ( n30125 , n30123 , n30124 );
buf ( n30126 , n30125 );
nand ( n30127 , n30122 , n30126 );
buf ( n30128 , n30127 );
not ( n30129 , n30128 );
or ( n30130 , n30119 , n30129 );
nand ( n30131 , n29022 , n26278 );
buf ( n30132 , n30131 );
nand ( n30133 , n30130 , n30132 );
buf ( n30134 , n30133 );
buf ( n30135 , n30134 );
xor ( n30136 , n30117 , n30135 );
buf ( n30137 , n30136 );
buf ( n30138 , n30137 );
xor ( n30139 , n30086 , n30138 );
xor ( n30140 , n29034 , n29063 );
and ( n30141 , n30140 , n29075 );
and ( n30142 , n29034 , n29063 );
or ( n30143 , n30141 , n30142 );
buf ( n30144 , n30143 );
buf ( n30145 , n30144 );
xor ( n30146 , n30139 , n30145 );
buf ( n30147 , n30146 );
buf ( n30148 , n30147 );
xor ( n30149 , n30066 , n30148 );
xor ( n30150 , n29078 , n29084 );
and ( n30151 , n30150 , n29165 );
and ( n30152 , n29078 , n29084 );
or ( n30153 , n30151 , n30152 );
buf ( n30154 , n30153 );
buf ( n30155 , n30154 );
xor ( n30156 , n30149 , n30155 );
buf ( n30157 , n30156 );
buf ( n30158 , n30157 );
xor ( n30159 , n30060 , n30158 );
buf ( n30160 , n30159 );
buf ( n30161 , n30160 );
not ( n30162 , n30161 );
xor ( n30163 , n29168 , n29233 );
and ( n30164 , n30163 , n29240 );
and ( n30165 , n29168 , n29233 );
or ( n30166 , n30164 , n30165 );
buf ( n30167 , n30166 );
buf ( n30168 , n30167 );
not ( n30169 , n30168 );
buf ( n30170 , n30169 );
buf ( n30171 , n30170 );
nand ( n30172 , n30162 , n30171 );
buf ( n30173 , n30172 );
buf ( n30174 , n30173 );
buf ( n30175 , n30174 );
buf ( n30176 , n30175 );
buf ( n30177 , n30160 );
buf ( n30178 , n30167 );
nand ( n30179 , n30177 , n30178 );
buf ( n30180 , n30179 );
nand ( n30181 , n30176 , n30180 );
not ( n30182 , n30181 );
and ( n30183 , n29896 , n30182 );
not ( n30184 , n29896 );
and ( n30185 , n30184 , n30181 );
nor ( n30186 , n30183 , n30185 );
buf ( n30187 , n30186 );
buf ( n30188 , n30187 );
buf ( n30189 , n30188 );
xor ( n30190 , n29870 , n30189 );
buf ( n30191 , n30190 );
buf ( n30192 , n30191 );
not ( n30193 , n30192 );
buf ( n30194 , n30193 );
buf ( n30195 , n30194 );
xor ( n30196 , n28743 , n28744 );
and ( n30197 , n30196 , n29271 );
and ( n30198 , n28743 , n28744 );
or ( n30199 , n30197 , n30198 );
buf ( n30200 , n30199 );
buf ( n30201 , n30200 );
not ( n30202 , n30201 );
buf ( n30203 , n30202 );
buf ( n30204 , n30203 );
nand ( n30205 , n30195 , n30204 );
buf ( n30206 , n30205 );
buf ( n30207 , n30206 );
and ( n30208 , n29867 , n30207 );
buf ( n30209 , n30194 );
buf ( n30210 , n30203 );
nor ( n30211 , n30209 , n30210 );
buf ( n30212 , n30211 );
buf ( n30213 , n30212 );
nor ( n30214 , n30208 , n30213 );
buf ( n30215 , n30214 );
buf ( n30216 , n30215 );
buf ( n30217 , n29866 );
buf ( n30218 , n30212 );
or ( n30219 , n30217 , n30218 );
buf ( n30220 , n30206 );
nand ( n30221 , n30219 , n30220 );
buf ( n30222 , n30221 );
buf ( n30223 , n30222 );
not ( n30224 , n30223 );
buf ( n30225 , n30224 );
buf ( n30226 , n30225 );
xor ( n30227 , n29868 , n29869 );
and ( n30228 , n30227 , n30189 );
and ( n30229 , n29868 , n29869 );
or ( n30230 , n30228 , n30229 );
buf ( n30231 , n30230 );
buf ( n30232 , n30231 );
buf ( n30233 , n28742 );
xor ( n30234 , n30232 , n30233 );
buf ( n30235 , n30234 );
buf ( n30236 , n30235 );
and ( n30237 , n30236 , n30226 );
not ( n30238 , n30236 );
and ( n30239 , n30238 , n30216 );
nor ( n30240 , n30237 , n30239 );
buf ( n30241 , n30240 );
buf ( n30242 , n30203 );
buf ( n30243 , n30191 );
and ( n30244 , n30242 , n30243 );
not ( n30245 , n30242 );
buf ( n30246 , n30194 );
and ( n30247 , n30245 , n30246 );
nor ( n30248 , n30244 , n30247 );
buf ( n30249 , n30248 );
buf ( n30250 , n30249 );
buf ( n30251 , n29866 );
buf ( n30252 , n30249 );
buf ( n30253 , n29866 );
not ( n30254 , n30250 );
not ( n30255 , n30251 );
or ( n30256 , n30254 , n30255 );
or ( n30257 , n30252 , n30253 );
nand ( n30258 , n30256 , n30257 );
buf ( n30259 , n30258 );
xor ( n30260 , n29274 , n29297 );
xor ( n30261 , n30260 , n29862 );
buf ( n30262 , n30261 );
xor ( n30263 , n29299 , n29303 );
xor ( n30264 , n30263 , n29857 );
buf ( n30265 , n30264 );
xor ( n30266 , n29305 , n29306 );
xor ( n30267 , n30266 , n29852 );
buf ( n30268 , n30267 );
xor ( n30269 , n29332 , n29333 );
xor ( n30270 , n30269 , n29847 );
buf ( n30271 , n30270 );
buf ( n30272 , n29729 );
buf ( n30273 , n28348 );
buf ( n30274 , n29435 );
and ( n30275 , n30273 , n30274 );
not ( n30276 , n30273 );
buf ( n30277 , n28326 );
and ( n30278 , n30276 , n30277 );
nor ( n30279 , n30275 , n30278 );
buf ( n30280 , n30279 );
buf ( n30281 , n30280 );
buf ( n30282 , n30280 );
buf ( n30283 , n29729 );
not ( n30284 , n30272 );
not ( n30285 , n30281 );
or ( n30286 , n30284 , n30285 );
or ( n30287 , n30282 , n30283 );
nand ( n30288 , n30286 , n30287 );
buf ( n30289 , n30288 );
buf ( n30290 , n29710 );
buf ( n30291 , n29707 );
buf ( n30292 , n28321 );
buf ( n30293 , n29717 );
xor ( n30294 , n30292 , n30293 );
buf ( n30295 , n30294 );
buf ( n30296 , n30295 );
and ( n30297 , n30296 , n30291 );
not ( n30298 , n30296 );
and ( n30299 , n30298 , n30290 );
nor ( n30300 , n30297 , n30299 );
buf ( n30301 , n30300 );
buf ( n30302 , n29466 );
buf ( n30303 , n29471 );
and ( n30304 , n30302 , n30303 );
not ( n30305 , n30302 );
buf ( n30306 , n28439 );
and ( n30307 , n30305 , n30306 );
nor ( n30308 , n30304 , n30307 );
buf ( n30309 , n30308 );
buf ( n30310 , n30309 );
buf ( n30311 , n29697 );
buf ( n30312 , n30309 );
buf ( n30313 , n29697 );
not ( n30314 , n30310 );
not ( n30315 , n30311 );
or ( n30316 , n30314 , n30315 );
or ( n30317 , n30312 , n30313 );
nand ( n30318 , n30316 , n30317 );
buf ( n30319 , n30318 );
buf ( n30320 , n29686 );
buf ( n30321 , n28434 );
buf ( n30322 , n29505 );
xnor ( n30323 , n30321 , n30322 );
buf ( n30324 , n30323 );
buf ( n30325 , n30324 );
buf ( n30326 , n30324 );
buf ( n30327 , n29686 );
not ( n30328 , n30320 );
not ( n30329 , n30325 );
or ( n30330 , n30328 , n30329 );
or ( n30331 , n30326 , n30327 );
nand ( n30332 , n30330 , n30331 );
buf ( n30333 , n30332 );
buf ( n30334 , n29510 );
buf ( n30335 , n29681 );
xnor ( n30336 , n30334 , n30335 );
buf ( n30337 , n30336 );
buf ( n30338 , n30337 );
buf ( n30339 , n29676 );
buf ( n30340 , n29676 );
buf ( n30341 , n30337 );
not ( n30342 , n30338 );
not ( n30343 , n30339 );
or ( n30344 , n30342 , n30343 );
or ( n30345 , n30340 , n30341 );
nand ( n30346 , n30344 , n30345 );
buf ( n30347 , n30346 );
buf ( n30348 , n29656 );
buf ( n30349 , n29653 );
buf ( n30350 , n26037 );
buf ( n30351 , n26006 );
xor ( n30352 , n30350 , n30351 );
buf ( n30353 , n30352 );
buf ( n30354 , n30353 );
and ( n30355 , n30354 , n30349 );
not ( n30356 , n30354 );
and ( n30357 , n30356 , n30348 );
nor ( n30358 , n30355 , n30357 );
buf ( n30359 , n30358 );
xor ( n30360 , n29545 , n29546 );
xor ( n30361 , n30360 , n29649 );
buf ( n30362 , n30361 );
buf ( n30363 , n25981 );
buf ( n30364 , n25960 );
xor ( n30365 , n30363 , n30364 );
buf ( n30366 , n30365 );
buf ( n30367 , n30366 );
buf ( n30368 , n29642 );
xor ( n30369 , n30367 , n30368 );
buf ( n30370 , n30369 );
buf ( n30371 , n25955 );
buf ( n30372 , n25947 );
xor ( n30373 , n30371 , n30372 );
buf ( n30374 , n30373 );
buf ( n30375 , n30374 );
buf ( n30376 , n29631 );
xor ( n30377 , n30375 , n30376 );
buf ( n30378 , n30377 );
buf ( n30379 , n25942 );
buf ( n30380 , n25934 );
xor ( n30381 , n30379 , n30380 );
buf ( n30382 , n30381 );
buf ( n30383 , n30382 );
buf ( n30384 , n29620 );
xor ( n30385 , n30383 , n30384 );
buf ( n30386 , n30385 );
buf ( n30387 , n29606 );
buf ( n30388 , n29603 );
buf ( n30389 , n25929 );
buf ( n30390 , n25909 );
xor ( n30391 , n30389 , n30390 );
buf ( n30392 , n30391 );
buf ( n30393 , n30392 );
and ( n30394 , n30393 , n30388 );
not ( n30395 , n30393 );
and ( n30396 , n30395 , n30387 );
nor ( n30397 , n30394 , n30396 );
buf ( n30398 , n30397 );
xor ( n30399 , n29562 , n29597 );
xor ( n30400 , n30399 , n29599 );
buf ( n30401 , n30400 );
xor ( n30402 , n29563 , n29590 );
xor ( n30403 , n30402 , n29592 );
buf ( n30404 , n30403 );
xor ( n30405 , n29582 , n29583 );
xor ( n30406 , n30405 , n29585 );
buf ( n30407 , n30406 );
xor ( n30408 , n29564 , n29568 );
xor ( n30409 , n30408 , n29577 );
buf ( n30410 , n30409 );
buf ( n30411 , n29442 );
buf ( n30412 , n28353 );
buf ( n30413 , n29440 );
and ( n30414 , n30413 , n30412 );
not ( n30415 , n30413 );
and ( n30416 , n30415 , n30411 );
nor ( n30417 , n30414 , n30416 );
buf ( n30418 , n30417 );
buf ( n30419 , n29774 );
buf ( n30420 , n29771 );
buf ( n30421 , n29768 );
and ( n30422 , n30421 , n30420 );
not ( n30423 , n30421 );
and ( n30424 , n30423 , n30419 );
nor ( n30425 , n30422 , n30424 );
buf ( n30426 , n30425 );
buf ( n30427 , n29819 );
buf ( n30428 , n28420 );
buf ( n30429 , n29814 );
and ( n30430 , n30429 , n30428 );
not ( n30431 , n30429 );
and ( n30432 , n30431 , n30427 );
nor ( n30433 , n30430 , n30432 );
buf ( n30434 , n30433 );
buf ( n30435 , n29413 );
buf ( n30436 , n29410 );
buf ( n30437 , n28415 );
and ( n30438 , n30437 , n30436 );
not ( n30439 , n30437 );
and ( n30440 , n30439 , n30435 );
nor ( n30441 , n30438 , n30440 );
buf ( n30442 , n30441 );
buf ( n30443 , n29425 );
buf ( n30444 , n29794 );
buf ( n30445 , n29420 );
and ( n30446 , n30445 , n30444 );
not ( n30447 , n30445 );
and ( n30448 , n30447 , n30443 );
nor ( n30449 , n30446 , n30448 );
buf ( n30450 , n30449 );
buf ( n30451 , n29760 );
buf ( n30452 , n29757 );
buf ( n30453 , n29784 );
and ( n30454 , n30453 , n30452 );
not ( n30455 , n30453 );
and ( n30456 , n30455 , n30451 );
nor ( n30457 , n30454 , n30456 );
buf ( n30458 , n30457 );
not ( n30459 , n29438 );
not ( n30460 , n29729 );
or ( n30461 , n30459 , n30460 );
nand ( n30462 , n30461 , n29735 );
buf ( n30463 , n30462 );
buf ( n30464 , n30418 );
xor ( n30465 , n30463 , n30464 );
buf ( n30466 , n30465 );
buf ( n30467 , n29740 );
buf ( n30468 , n30426 );
xor ( n30469 , n30467 , n30468 );
buf ( n30470 , n30469 );
not ( n30471 , n29775 );
not ( n30472 , n29740 );
or ( n30473 , n30471 , n30472 );
nand ( n30474 , n30473 , n29779 );
buf ( n30475 , n30474 );
buf ( n30476 , n30458 );
xor ( n30477 , n30475 , n30476 );
buf ( n30478 , n30477 );
buf ( n30479 , n29787 );
buf ( n30480 , n30450 );
xor ( n30481 , n30479 , n30480 );
buf ( n30482 , n30481 );
buf ( n30483 , n29800 );
buf ( n30484 , n30442 );
xor ( n30485 , n30483 , n30484 );
buf ( n30486 , n30485 );
buf ( n30487 , n29810 );
buf ( n30488 , n30434 );
xor ( n30489 , n30487 , n30488 );
buf ( n30490 , n30489 );
buf ( n30491 , n18340 );
not ( n30492 , n30491 );
buf ( n30493 , n576 );
not ( n30494 , n30493 );
buf ( n30495 , n19403 );
buf ( n30496 , n30495 );
buf ( n30497 , n30496 );
buf ( n30498 , n30497 );
not ( n30499 , n30498 );
buf ( n30500 , n30499 );
buf ( n30501 , n30500 );
not ( n30502 , n30501 );
or ( n30503 , n30494 , n30502 );
buf ( n30504 , n30497 );
buf ( n30505 , n7809 );
nand ( n30506 , n30504 , n30505 );
buf ( n30507 , n30506 );
buf ( n30508 , n30507 );
nand ( n30509 , n30503 , n30508 );
buf ( n30510 , n30509 );
buf ( n30511 , n30510 );
not ( n30512 , n30511 );
or ( n30513 , n30492 , n30512 );
buf ( n30514 , n576 );
not ( n30515 , n30514 );
buf ( n30516 , n28238 );
not ( n30517 , n30516 );
or ( n30518 , n30515 , n30517 );
buf ( n30519 , n19209 );
buf ( n30520 , n7809 );
nand ( n30521 , n30519 , n30520 );
buf ( n30522 , n30521 );
buf ( n30523 , n30522 );
nand ( n30524 , n30518 , n30523 );
buf ( n30525 , n30524 );
buf ( n30526 , n30525 );
buf ( n30527 , n18365 );
buf ( n30528 , n30527 );
buf ( n30529 , n30528 );
buf ( n30530 , n30529 );
nand ( n30531 , n30526 , n30530 );
buf ( n30532 , n30531 );
buf ( n30533 , n30532 );
nand ( n30534 , n30513 , n30533 );
buf ( n30535 , n30534 );
buf ( n30536 , n30535 );
buf ( n30537 , n18264 );
buf ( n30538 , n578 );
not ( n30539 , n30538 );
buf ( n30540 , n19398 );
not ( n30541 , n30540 );
buf ( n30542 , n30541 );
buf ( n30543 , n30542 );
not ( n30544 , n30543 );
or ( n30545 , n30539 , n30544 );
buf ( n30546 , n30542 );
not ( n30547 , n30546 );
buf ( n30548 , n30547 );
buf ( n30549 , n30548 );
buf ( n30550 , n18233 );
nand ( n30551 , n30549 , n30550 );
buf ( n30552 , n30551 );
buf ( n30553 , n30552 );
nand ( n30554 , n30545 , n30553 );
buf ( n30555 , n30554 );
buf ( n30556 , n30555 );
nand ( n30557 , n30537 , n30556 );
buf ( n30558 , n30557 );
not ( n30559 , n578 );
buf ( n30560 , n17997 );
buf ( n30561 , n30560 );
buf ( n30562 , n30561 );
buf ( n30563 , n30562 );
not ( n30564 , n30563 );
buf ( n30565 , n30564 );
not ( n30566 , n30565 );
or ( n30567 , n30559 , n30566 );
buf ( n30568 , n30562 );
buf ( n30569 , n18233 );
nand ( n30570 , n30568 , n30569 );
buf ( n30571 , n30570 );
nand ( n30572 , n30567 , n30571 );
nand ( n30573 , n30572 , n18219 );
nand ( n30574 , n30558 , n30573 );
buf ( n30575 , n30574 );
xor ( n30576 , n30536 , n30575 );
buf ( n30577 , n19181 );
buf ( n30578 , n30577 );
buf ( n30579 , n30578 );
buf ( n30580 , n30579 );
not ( n30581 , n30580 );
buf ( n30582 , n30581 );
buf ( n30583 , n30582 );
not ( n30584 , n30583 );
buf ( n30585 , n576 );
nand ( n30586 , n30584 , n30585 );
buf ( n30587 , n30586 );
buf ( n30588 , n30587 );
xor ( n30589 , n30576 , n30588 );
buf ( n30590 , n30589 );
buf ( n30591 , n30590 );
buf ( n30592 , n18392 );
not ( n30593 , n30592 );
buf ( n30594 , n580 );
not ( n30595 , n30594 );
not ( n30596 , n17981 );
not ( n30597 , n30596 );
not ( n30598 , n30597 );
buf ( n30599 , n30598 );
not ( n30600 , n30599 );
or ( n30601 , n30595 , n30600 );
buf ( n30602 , n30597 );
buf ( n30603 , n18402 );
nand ( n30604 , n30602 , n30603 );
buf ( n30605 , n30604 );
buf ( n30606 , n30605 );
nand ( n30607 , n30601 , n30606 );
buf ( n30608 , n30607 );
buf ( n30609 , n30608 );
not ( n30610 , n30609 );
or ( n30611 , n30593 , n30610 );
buf ( n30612 , n580 );
not ( n30613 , n30612 );
buf ( n30614 , n18170 );
not ( n30615 , n30614 );
or ( n30616 , n30613 , n30615 );
buf ( n30617 , n18167 );
buf ( n30618 , n18402 );
nand ( n30619 , n30617 , n30618 );
buf ( n30620 , n30619 );
buf ( n30621 , n30620 );
nand ( n30622 , n30616 , n30621 );
buf ( n30623 , n30622 );
buf ( n30624 , n30623 );
buf ( n30625 , n18418 );
nand ( n30626 , n30624 , n30625 );
buf ( n30627 , n30626 );
buf ( n30628 , n30627 );
nand ( n30629 , n30611 , n30628 );
buf ( n30630 , n30629 );
buf ( n30631 , n30630 );
buf ( n30632 , n18340 );
not ( n30633 , n30632 );
buf ( n30634 , n30525 );
not ( n30635 , n30634 );
or ( n30636 , n30633 , n30635 );
and ( n30637 , n30582 , n576 );
not ( n30638 , n30582 );
and ( n30639 , n30638 , n7809 );
or ( n30640 , n30637 , n30639 );
buf ( n30641 , n30640 );
buf ( n30642 , n30529 );
nand ( n30643 , n30641 , n30642 );
buf ( n30644 , n30643 );
buf ( n30645 , n30644 );
nand ( n30646 , n30636 , n30645 );
buf ( n30647 , n30646 );
buf ( n30648 , n30647 );
buf ( n30649 , n19167 );
buf ( n30650 , n576 );
and ( n30651 , n30649 , n30650 );
buf ( n30652 , n30651 );
buf ( n30653 , n30652 );
xor ( n30654 , n30648 , n30653 );
or ( n30655 , n18316 , n18657 );
buf ( n30656 , n582 );
not ( n30657 , n30656 );
buf ( n30658 , n18170 );
not ( n30659 , n30658 );
or ( n30660 , n30657 , n30659 );
buf ( n30661 , n18167 );
buf ( n30662 , n18303 );
nand ( n30663 , n30661 , n30662 );
buf ( n30664 , n30663 );
buf ( n30665 , n30664 );
nand ( n30666 , n30660 , n30665 );
buf ( n30667 , n30666 );
nand ( n30668 , n30655 , n30667 );
buf ( n30669 , n30668 );
and ( n30670 , n30654 , n30669 );
and ( n30671 , n30648 , n30653 );
or ( n30672 , n30670 , n30671 );
buf ( n30673 , n30672 );
buf ( n30674 , n30673 );
xor ( n30675 , n30631 , n30674 );
buf ( n30676 , n18219 );
not ( n30677 , n30676 );
buf ( n30678 , n30555 );
not ( n30679 , n30678 );
or ( n30680 , n30677 , n30679 );
buf ( n30681 , n578 );
not ( n30682 , n30681 );
buf ( n30683 , n28661 );
not ( n30684 , n30683 );
or ( n30685 , n30682 , n30684 );
buf ( n30686 , n30497 );
buf ( n30687 , n18233 );
nand ( n30688 , n30686 , n30687 );
buf ( n30689 , n30688 );
buf ( n30690 , n30689 );
nand ( n30691 , n30685 , n30690 );
buf ( n30692 , n30691 );
buf ( n30693 , n30692 );
buf ( n30694 , n18264 );
nand ( n30695 , n30693 , n30694 );
buf ( n30696 , n30695 );
buf ( n30697 , n30696 );
nand ( n30698 , n30680 , n30697 );
buf ( n30699 , n30698 );
buf ( n30700 , n30699 );
buf ( n30701 , n18418 );
not ( n30702 , n30701 );
buf ( n30703 , n30608 );
not ( n30704 , n30703 );
or ( n30705 , n30702 , n30704 );
buf ( n30706 , n580 );
not ( n30707 , n30706 );
buf ( n30708 , n30019 );
not ( n30709 , n30708 );
or ( n30710 , n30707 , n30709 );
buf ( n30711 , n30562 );
buf ( n30712 , n18402 );
nand ( n30713 , n30711 , n30712 );
buf ( n30714 , n30713 );
buf ( n30715 , n30714 );
nand ( n30716 , n30710 , n30715 );
buf ( n30717 , n30716 );
buf ( n30718 , n30717 );
buf ( n30719 , n18392 );
nand ( n30720 , n30718 , n30719 );
buf ( n30721 , n30720 );
buf ( n30722 , n30721 );
nand ( n30723 , n30705 , n30722 );
buf ( n30724 , n30723 );
buf ( n30725 , n30724 );
xor ( n30726 , n30700 , n30725 );
not ( n30727 , n24218 );
nand ( n30728 , n30727 , n576 );
buf ( n30729 , n30728 );
not ( n30730 , n30729 );
buf ( n30731 , n30730 );
buf ( n30732 , n30731 );
and ( n30733 , n30726 , n30732 );
and ( n30734 , n30700 , n30725 );
or ( n30735 , n30733 , n30734 );
buf ( n30736 , n30735 );
buf ( n30737 , n30736 );
xor ( n30738 , n30675 , n30737 );
buf ( n30739 , n30738 );
buf ( n30740 , n30739 );
xor ( n30741 , n30591 , n30740 );
xor ( n30742 , n30648 , n30653 );
xor ( n30743 , n30742 , n30669 );
buf ( n30744 , n30743 );
buf ( n30745 , n30744 );
buf ( n30746 , n30529 );
not ( n30747 , n30746 );
buf ( n30748 , n576 );
not ( n30749 , n30748 );
buf ( n30750 , n24324 );
not ( n30751 , n30750 );
or ( n30752 , n30749 , n30751 );
buf ( n30753 , n19167 );
buf ( n30754 , n7809 );
nand ( n30755 , n30753 , n30754 );
buf ( n30756 , n30755 );
buf ( n30757 , n30756 );
nand ( n30758 , n30752 , n30757 );
buf ( n30759 , n30758 );
buf ( n30760 , n30759 );
not ( n30761 , n30760 );
or ( n30762 , n30747 , n30761 );
buf ( n30763 , n30640 );
buf ( n30764 , n18340 );
nand ( n30765 , n30763 , n30764 );
buf ( n30766 , n30765 );
buf ( n30767 , n30766 );
nand ( n30768 , n30762 , n30767 );
buf ( n30769 , n30768 );
buf ( n30770 , n30769 );
buf ( n30771 , n18219 );
not ( n30772 , n30771 );
buf ( n30773 , n30692 );
not ( n30774 , n30773 );
or ( n30775 , n30772 , n30774 );
buf ( n30776 , n578 );
not ( n30777 , n30776 );
buf ( n30778 , n24346 );
not ( n30779 , n30778 );
or ( n30780 , n30777 , n30779 );
buf ( n30781 , n19209 );
buf ( n30782 , n18233 );
nand ( n30783 , n30781 , n30782 );
buf ( n30784 , n30783 );
buf ( n30785 , n30784 );
nand ( n30786 , n30780 , n30785 );
buf ( n30787 , n30786 );
buf ( n30788 , n30787 );
buf ( n30789 , n18264 );
nand ( n30790 , n30788 , n30789 );
buf ( n30791 , n30790 );
buf ( n30792 , n30791 );
nand ( n30793 , n30775 , n30792 );
buf ( n30794 , n30793 );
buf ( n30795 , n30794 );
xor ( n30796 , n30770 , n30795 );
buf ( n30797 , n18316 );
not ( n30798 , n30797 );
buf ( n30799 , n582 );
not ( n30800 , n30799 );
buf ( n30801 , n30016 );
not ( n30802 , n30801 );
or ( n30803 , n30800 , n30802 );
buf ( n30804 , n18303 );
buf ( n30805 , n30015 );
nand ( n30806 , n30804 , n30805 );
buf ( n30807 , n30806 );
buf ( n30808 , n30807 );
nand ( n30809 , n30803 , n30808 );
buf ( n30810 , n30809 );
buf ( n30811 , n30810 );
not ( n30812 , n30811 );
or ( n30813 , n30798 , n30812 );
buf ( n30814 , n30667 );
buf ( n30815 , n18657 );
nand ( n30816 , n30814 , n30815 );
buf ( n30817 , n30816 );
buf ( n30818 , n30817 );
nand ( n30819 , n30813 , n30818 );
buf ( n30820 , n30819 );
buf ( n30821 , n30820 );
and ( n30822 , n30796 , n30821 );
and ( n30823 , n30770 , n30795 );
or ( n30824 , n30822 , n30823 );
buf ( n30825 , n30824 );
buf ( n30826 , n30825 );
xor ( n30827 , n30745 , n30826 );
buf ( n30828 , n18418 );
not ( n30829 , n30828 );
buf ( n30830 , n30717 );
not ( n30831 , n30830 );
or ( n30832 , n30829 , n30831 );
buf ( n30833 , n580 );
not ( n30834 , n30833 );
buf ( n30835 , n24462 );
not ( n30836 , n30835 );
or ( n30837 , n30834 , n30836 );
buf ( n30838 , n19398 );
buf ( n30839 , n18402 );
nand ( n30840 , n30838 , n30839 );
buf ( n30841 , n30840 );
buf ( n30842 , n30841 );
nand ( n30843 , n30837 , n30842 );
buf ( n30844 , n30843 );
buf ( n30845 , n30844 );
buf ( n30846 , n18392 );
nand ( n30847 , n30845 , n30846 );
buf ( n30848 , n30847 );
buf ( n30849 , n30848 );
nand ( n30850 , n30832 , n30849 );
buf ( n30851 , n30850 );
buf ( n30852 , n30851 );
buf ( n30853 , n30728 );
xor ( n30854 , n30852 , n30853 );
buf ( n30855 , n20389 );
buf ( n30856 , n576 );
and ( n30857 , n30855 , n30856 );
buf ( n30858 , n30857 );
buf ( n30859 , n30858 );
buf ( n30860 , n18861 );
buf ( n30861 , n576 );
nand ( n30862 , n30860 , n30861 );
buf ( n30863 , n30862 );
buf ( n30864 , n30863 );
not ( n30865 , n30864 );
buf ( n30866 , n30865 );
buf ( n30867 , n30866 );
xor ( n30868 , n30859 , n30867 );
buf ( n30869 , n18219 );
not ( n30870 , n30869 );
buf ( n30871 , n30787 );
not ( n30872 , n30871 );
or ( n30873 , n30870 , n30872 );
buf ( n30874 , n578 );
not ( n30875 , n30874 );
buf ( n30876 , n30582 );
not ( n30877 , n30876 );
or ( n30878 , n30875 , n30877 );
buf ( n30879 , n30579 );
buf ( n30880 , n18233 );
nand ( n30881 , n30879 , n30880 );
buf ( n30882 , n30881 );
buf ( n30883 , n30882 );
nand ( n30884 , n30878 , n30883 );
buf ( n30885 , n30884 );
buf ( n30886 , n30885 );
buf ( n30887 , n18264 );
nand ( n30888 , n30886 , n30887 );
buf ( n30889 , n30888 );
buf ( n30890 , n30889 );
nand ( n30891 , n30873 , n30890 );
buf ( n30892 , n30891 );
buf ( n30893 , n30892 );
and ( n30894 , n30868 , n30893 );
and ( n30895 , n30859 , n30867 );
or ( n30896 , n30894 , n30895 );
buf ( n30897 , n30896 );
buf ( n30898 , n30897 );
and ( n30899 , n30854 , n30898 );
and ( n30900 , n30852 , n30853 );
or ( n30901 , n30899 , n30900 );
buf ( n30902 , n30901 );
buf ( n30903 , n30902 );
and ( n30904 , n30827 , n30903 );
and ( n30905 , n30745 , n30826 );
or ( n30906 , n30904 , n30905 );
buf ( n30907 , n30906 );
buf ( n30908 , n30907 );
xor ( n30909 , n30741 , n30908 );
buf ( n30910 , n30909 );
not ( n30911 , n30910 );
xor ( n30912 , n30700 , n30725 );
xor ( n30913 , n30912 , n30732 );
buf ( n30914 , n30913 );
buf ( n30915 , n30914 );
xor ( n30916 , n30745 , n30826 );
xor ( n30917 , n30916 , n30903 );
buf ( n30918 , n30917 );
buf ( n30919 , n30918 );
xor ( n30920 , n30915 , n30919 );
buf ( n30921 , n30529 );
not ( n30922 , n30921 );
buf ( n30923 , n576 );
not ( n30924 , n30923 );
buf ( n30925 , n19254 );
not ( n30926 , n30925 );
or ( n30927 , n30924 , n30926 );
nand ( n30928 , n20137 , n7809 );
buf ( n30929 , n30928 );
nand ( n30930 , n30927 , n30929 );
buf ( n30931 , n30930 );
buf ( n30932 , n30931 );
not ( n30933 , n30932 );
or ( n30934 , n30922 , n30933 );
buf ( n30935 , n30759 );
buf ( n30936 , n18340 );
nand ( n30937 , n30935 , n30936 );
buf ( n30938 , n30937 );
buf ( n30939 , n30938 );
nand ( n30940 , n30934 , n30939 );
buf ( n30941 , n30940 );
buf ( n30942 , n30941 );
buf ( n30943 , n18392 );
not ( n30944 , n30943 );
buf ( n30945 , n580 );
not ( n30946 , n30945 );
buf ( n30947 , n30500 );
not ( n30948 , n30947 );
or ( n30949 , n30946 , n30948 );
buf ( n30950 , n28661 );
not ( n30951 , n30950 );
buf ( n30952 , n18402 );
nand ( n30953 , n30951 , n30952 );
buf ( n30954 , n30953 );
buf ( n30955 , n30954 );
nand ( n30956 , n30949 , n30955 );
buf ( n30957 , n30956 );
buf ( n30958 , n30957 );
not ( n30959 , n30958 );
or ( n30960 , n30944 , n30959 );
buf ( n30961 , n30844 );
buf ( n30962 , n18418 );
nand ( n30963 , n30961 , n30962 );
buf ( n30964 , n30963 );
buf ( n30965 , n30964 );
nand ( n30966 , n30960 , n30965 );
buf ( n30967 , n30966 );
buf ( n30968 , n30967 );
xor ( n30969 , n30942 , n30968 );
not ( n30970 , n584 );
not ( n30971 , n18170 );
or ( n30972 , n30970 , n30971 );
buf ( n30973 , n18167 );
buf ( n30974 , n18277 );
nand ( n30975 , n30973 , n30974 );
buf ( n30976 , n30975 );
nand ( n30977 , n30972 , n30976 );
not ( n30978 , n18479 );
nand ( n30979 , n30978 , n18912 );
nand ( n30980 , n30977 , n30979 );
buf ( n30981 , n30980 );
and ( n30982 , n30969 , n30981 );
and ( n30983 , n30942 , n30968 );
or ( n30984 , n30982 , n30983 );
buf ( n30985 , n30984 );
buf ( n30986 , n30985 );
xor ( n30987 , n30770 , n30795 );
xor ( n30988 , n30987 , n30821 );
buf ( n30989 , n30988 );
buf ( n30990 , n30989 );
xor ( n30991 , n30986 , n30990 );
buf ( n30992 , n18316 );
not ( n30993 , n30992 );
buf ( n30994 , n582 );
not ( n30995 , n30994 );
buf ( n30996 , n30565 );
not ( n30997 , n30996 );
or ( n30998 , n30995 , n30997 );
buf ( n30999 , n30019 );
not ( n31000 , n30999 );
buf ( n31001 , n18303 );
nand ( n31002 , n31000 , n31001 );
buf ( n31003 , n31002 );
buf ( n31004 , n31003 );
nand ( n31005 , n30998 , n31004 );
buf ( n31006 , n31005 );
buf ( n31007 , n31006 );
not ( n31008 , n31007 );
or ( n31009 , n30993 , n31008 );
buf ( n31010 , n30810 );
buf ( n31011 , n18657 );
nand ( n31012 , n31010 , n31011 );
buf ( n31013 , n31012 );
buf ( n31014 , n31013 );
nand ( n31015 , n31009 , n31014 );
buf ( n31016 , n31015 );
buf ( n31017 , n31016 );
buf ( n31018 , n30863 );
buf ( n31019 , n18264 );
not ( n31020 , n31019 );
buf ( n31021 , n18233 );
not ( n31022 , n31021 );
buf ( n31023 , n19783 );
not ( n31024 , n31023 );
or ( n31025 , n31022 , n31024 );
buf ( n31026 , n24324 );
buf ( n31027 , n578 );
nand ( n31028 , n31026 , n31027 );
buf ( n31029 , n31028 );
buf ( n31030 , n31029 );
nand ( n31031 , n31025 , n31030 );
buf ( n31032 , n31031 );
buf ( n31033 , n31032 );
not ( n31034 , n31033 );
or ( n31035 , n31020 , n31034 );
buf ( n31036 , n30885 );
buf ( n31037 , n18219 );
nand ( n31038 , n31036 , n31037 );
buf ( n31039 , n31038 );
buf ( n31040 , n31039 );
nand ( n31041 , n31035 , n31040 );
buf ( n31042 , n31041 );
buf ( n31043 , n31042 );
xor ( n31044 , n31018 , n31043 );
buf ( n31045 , n18340 );
not ( n31046 , n31045 );
buf ( n31047 , n30931 );
not ( n31048 , n31047 );
or ( n31049 , n31046 , n31048 );
buf ( n31050 , n576 );
not ( n31051 , n31050 );
buf ( n31052 , n24135 );
not ( n31053 , n31052 );
or ( n31054 , n31051 , n31053 );
buf ( n31055 , n18725 );
buf ( n31056 , n7809 );
nand ( n31057 , n31055 , n31056 );
buf ( n31058 , n31057 );
buf ( n31059 , n31058 );
nand ( n31060 , n31054 , n31059 );
buf ( n31061 , n31060 );
buf ( n31062 , n31061 );
buf ( n31063 , n31062 );
buf ( n31064 , n30529 );
nand ( n31065 , n31063 , n31064 );
buf ( n31066 , n31065 );
buf ( n31067 , n31066 );
nand ( n31068 , n31049 , n31067 );
buf ( n31069 , n31068 );
buf ( n31070 , n31069 );
and ( n31071 , n31044 , n31070 );
and ( n31072 , n31018 , n31043 );
or ( n31073 , n31071 , n31072 );
buf ( n31074 , n31073 );
buf ( n31075 , n31074 );
xor ( n31076 , n31017 , n31075 );
xor ( n31077 , n30859 , n30867 );
xor ( n31078 , n31077 , n30893 );
buf ( n31079 , n31078 );
buf ( n31080 , n31079 );
and ( n31081 , n31076 , n31080 );
and ( n31082 , n31017 , n31075 );
or ( n31083 , n31081 , n31082 );
buf ( n31084 , n31083 );
buf ( n31085 , n31084 );
and ( n31086 , n30991 , n31085 );
and ( n31087 , n30986 , n30990 );
or ( n31088 , n31086 , n31087 );
buf ( n31089 , n31088 );
buf ( n31090 , n31089 );
and ( n31091 , n30920 , n31090 );
and ( n31092 , n30915 , n30919 );
or ( n31093 , n31091 , n31092 );
buf ( n31094 , n31093 );
not ( n31095 , n31094 );
and ( n31096 , n30911 , n31095 );
xor ( n31097 , n30852 , n30853 );
xor ( n31098 , n31097 , n30898 );
buf ( n31099 , n31098 );
buf ( n31100 , n31099 );
xor ( n31101 , n30986 , n30990 );
xor ( n31102 , n31101 , n31085 );
buf ( n31103 , n31102 );
buf ( n31104 , n31103 );
xor ( n31105 , n31100 , n31104 );
and ( n31106 , n576 , n20160 );
buf ( n31107 , n31106 );
not ( n31108 , n18340 );
not ( n31109 , n31061 );
or ( n31110 , n31108 , n31109 );
buf ( n31111 , n576 );
not ( n31112 , n31111 );
buf ( n31113 , n18442 );
not ( n31114 , n31113 );
or ( n31115 , n31112 , n31114 );
buf ( n31116 , n18861 );
buf ( n31117 , n7809 );
nand ( n31118 , n31116 , n31117 );
buf ( n31119 , n31118 );
buf ( n31120 , n31119 );
nand ( n31121 , n31115 , n31120 );
buf ( n31122 , n31121 );
nand ( n31123 , n31122 , n18365 );
nand ( n31124 , n31110 , n31123 );
buf ( n31125 , n31124 );
xor ( n31126 , n31107 , n31125 );
buf ( n31127 , n18909 );
buf ( n31128 , n31127 );
buf ( n31129 , n576 );
nand ( n31130 , n31128 , n31129 );
buf ( n31131 , n31130 );
buf ( n31132 , n31131 );
not ( n31133 , n31132 );
buf ( n31134 , n31133 );
buf ( n31135 , n31134 );
and ( n31136 , n31126 , n31135 );
and ( n31137 , n31107 , n31125 );
or ( n31138 , n31136 , n31137 );
buf ( n31139 , n31138 );
buf ( n31140 , n31139 );
buf ( n31141 , n18418 );
not ( n31142 , n31141 );
buf ( n31143 , n30957 );
not ( n31144 , n31143 );
or ( n31145 , n31142 , n31144 );
not ( n31146 , n580 );
not ( n31147 , n24346 );
or ( n31148 , n31146 , n31147 );
buf ( n31149 , n19209 );
buf ( n31150 , n18402 );
nand ( n31151 , n31149 , n31150 );
buf ( n31152 , n31151 );
nand ( n31153 , n31148 , n31152 );
buf ( n31154 , n31153 );
buf ( n31155 , n18392 );
nand ( n31156 , n31154 , n31155 );
buf ( n31157 , n31156 );
buf ( n31158 , n31157 );
nand ( n31159 , n31145 , n31158 );
buf ( n31160 , n31159 );
buf ( n31161 , n31160 );
xor ( n31162 , n31140 , n31161 );
not ( n31163 , n18431 );
not ( n31164 , n30977 );
or ( n31165 , n31163 , n31164 );
not ( n31166 , n584 );
not ( n31167 , n24498 );
or ( n31168 , n31166 , n31167 );
not ( n31169 , n30596 );
nand ( n31170 , n31169 , n18277 );
nand ( n31171 , n31168 , n31170 );
buf ( n31172 , n31171 );
buf ( n31173 , n18479 );
nand ( n31174 , n31172 , n31173 );
buf ( n31175 , n31174 );
nand ( n31176 , n31165 , n31175 );
buf ( n31177 , n31176 );
and ( n31178 , n31162 , n31177 );
and ( n31179 , n31140 , n31161 );
or ( n31180 , n31178 , n31179 );
buf ( n31181 , n31180 );
buf ( n31182 , n31181 );
xor ( n31183 , n30942 , n30968 );
xor ( n31184 , n31183 , n30981 );
buf ( n31185 , n31184 );
buf ( n31186 , n31185 );
xor ( n31187 , n31182 , n31186 );
xor ( n31188 , n31017 , n31075 );
xor ( n31189 , n31188 , n31080 );
buf ( n31190 , n31189 );
buf ( n31191 , n31190 );
and ( n31192 , n31187 , n31191 );
and ( n31193 , n31182 , n31186 );
or ( n31194 , n31192 , n31193 );
buf ( n31195 , n31194 );
buf ( n31196 , n31195 );
and ( n31197 , n31105 , n31196 );
and ( n31198 , n31100 , n31104 );
or ( n31199 , n31197 , n31198 );
buf ( n31200 , n31199 );
xor ( n31201 , n30915 , n30919 );
xor ( n31202 , n31201 , n31090 );
buf ( n31203 , n31202 );
nor ( n31204 , n31200 , n31203 );
nor ( n31205 , n31096 , n31204 );
buf ( n31206 , n31205 );
xor ( n31207 , n30591 , n30740 );
and ( n31208 , n31207 , n30908 );
and ( n31209 , n30591 , n30740 );
or ( n31210 , n31208 , n31209 );
buf ( n31211 , n31210 );
buf ( n31212 , n31211 );
not ( n31213 , n31212 );
buf ( n31214 , n31213 );
buf ( n31215 , n31214 );
xor ( n31216 , n30536 , n30575 );
and ( n31217 , n31216 , n30588 );
and ( n31218 , n30536 , n30575 );
or ( n31219 , n31217 , n31218 );
buf ( n31220 , n31219 );
buf ( n31221 , n31220 );
buf ( n31222 , n18264 );
not ( n31223 , n31222 );
buf ( n31224 , n30572 );
not ( n31225 , n31224 );
or ( n31226 , n31223 , n31225 );
buf ( n31227 , n578 );
not ( n31228 , n31227 );
buf ( n31229 , n30598 );
not ( n31230 , n31229 );
or ( n31231 , n31228 , n31230 );
buf ( n31232 , n30597 );
buf ( n31233 , n31232 );
buf ( n31234 , n18233 );
nand ( n31235 , n31233 , n31234 );
buf ( n31236 , n31235 );
buf ( n31237 , n31236 );
nand ( n31238 , n31231 , n31237 );
buf ( n31239 , n31238 );
buf ( n31240 , n31239 );
buf ( n31241 , n18219 );
nand ( n31242 , n31240 , n31241 );
buf ( n31243 , n31242 );
buf ( n31244 , n31243 );
nand ( n31245 , n31226 , n31244 );
buf ( n31246 , n31245 );
buf ( n31247 , n31246 );
buf ( n31248 , n30587 );
not ( n31249 , n31248 );
buf ( n31250 , n31249 );
buf ( n31251 , n31250 );
xor ( n31252 , n31247 , n31251 );
not ( n31253 , n28238 );
buf ( n31254 , n31253 );
buf ( n31255 , n576 );
and ( n31256 , n31254 , n31255 );
buf ( n31257 , n31256 );
buf ( n31258 , n31257 );
buf ( n31259 , n18525 );
not ( n31260 , n31259 );
buf ( n31261 , n18392 );
not ( n31262 , n31261 );
buf ( n31263 , n31262 );
buf ( n31264 , n31263 );
not ( n31265 , n31264 );
or ( n31266 , n31260 , n31265 );
buf ( n31267 , n30623 );
nand ( n31268 , n31266 , n31267 );
buf ( n31269 , n31268 );
buf ( n31270 , n31269 );
xor ( n31271 , n31258 , n31270 );
buf ( n31272 , n18340 );
not ( n31273 , n31272 );
buf ( n31274 , n576 );
buf ( n31275 , n19398 );
xor ( n31276 , n31274 , n31275 );
buf ( n31277 , n31276 );
buf ( n31278 , n31277 );
not ( n31279 , n31278 );
or ( n31280 , n31273 , n31279 );
buf ( n31281 , n30510 );
buf ( n31282 , n30529 );
nand ( n31283 , n31281 , n31282 );
buf ( n31284 , n31283 );
buf ( n31285 , n31284 );
nand ( n31286 , n31280 , n31285 );
buf ( n31287 , n31286 );
buf ( n31288 , n31287 );
xor ( n31289 , n31271 , n31288 );
buf ( n31290 , n31289 );
buf ( n31291 , n31290 );
xor ( n31292 , n31252 , n31291 );
buf ( n31293 , n31292 );
buf ( n31294 , n31293 );
xor ( n31295 , n31221 , n31294 );
xor ( n31296 , n30631 , n30674 );
and ( n31297 , n31296 , n30737 );
and ( n31298 , n30631 , n30674 );
or ( n31299 , n31297 , n31298 );
buf ( n31300 , n31299 );
buf ( n31301 , n31300 );
xor ( n31302 , n31295 , n31301 );
buf ( n31303 , n31302 );
buf ( n31304 , n31303 );
not ( n31305 , n31304 );
buf ( n31306 , n31305 );
buf ( n31307 , n31306 );
nand ( n31308 , n31215 , n31307 );
buf ( n31309 , n31308 );
buf ( n31310 , n31309 );
nand ( n31311 , n31206 , n31310 );
buf ( n31312 , n31311 );
buf ( n31313 , n31312 );
not ( n31314 , n31313 );
buf ( n31315 , n31314 );
not ( n31316 , n31315 );
buf ( n31317 , n18657 );
not ( n31318 , n31317 );
buf ( n31319 , n31006 );
not ( n31320 , n31319 );
or ( n31321 , n31318 , n31320 );
buf ( n31322 , n582 );
not ( n31323 , n31322 );
buf ( n31324 , n30542 );
not ( n31325 , n31324 );
or ( n31326 , n31323 , n31325 );
buf ( n31327 , n30548 );
buf ( n31328 , n18303 );
nand ( n31329 , n31327 , n31328 );
buf ( n31330 , n31329 );
buf ( n31331 , n31330 );
nand ( n31332 , n31326 , n31331 );
buf ( n31333 , n31332 );
buf ( n31334 , n31333 );
buf ( n31335 , n18316 );
nand ( n31336 , n31334 , n31335 );
buf ( n31337 , n31336 );
buf ( n31338 , n31337 );
nand ( n31339 , n31321 , n31338 );
buf ( n31340 , n31339 );
buf ( n31341 , n31340 );
buf ( n31342 , n18418 );
not ( n31343 , n31342 );
buf ( n31344 , n31153 );
not ( n31345 , n31344 );
or ( n31346 , n31343 , n31345 );
buf ( n31347 , n30579 );
buf ( n31348 , n18402 );
nand ( n31349 , n31347 , n31348 );
buf ( n31350 , n31349 );
not ( n31351 , n31350 );
nand ( n31352 , n30582 , n580 );
not ( n31353 , n31352 );
or ( n31354 , n31351 , n31353 );
nand ( n31355 , n31354 , n18392 );
buf ( n31356 , n31355 );
nand ( n31357 , n31346 , n31356 );
buf ( n31358 , n31357 );
buf ( n31359 , n31358 );
buf ( n31360 , n18264 );
not ( n31361 , n31360 );
buf ( n31362 , n578 );
not ( n31363 , n31362 );
buf ( n31364 , n24218 );
not ( n31365 , n31364 );
or ( n31366 , n31363 , n31365 );
buf ( n31367 , n19254 );
not ( n31368 , n31367 );
buf ( n31369 , n18233 );
nand ( n31370 , n31368 , n31369 );
buf ( n31371 , n31370 );
buf ( n31372 , n31371 );
nand ( n31373 , n31366 , n31372 );
buf ( n31374 , n31373 );
buf ( n31375 , n31374 );
not ( n31376 , n31375 );
or ( n31377 , n31361 , n31376 );
buf ( n31378 , n31032 );
buf ( n31379 , n18219 );
nand ( n31380 , n31378 , n31379 );
buf ( n31381 , n31380 );
buf ( n31382 , n31381 );
nand ( n31383 , n31377 , n31382 );
buf ( n31384 , n31383 );
buf ( n31385 , n31384 );
xor ( n31386 , n31359 , n31385 );
buf ( n31387 , n18316 );
not ( n31388 , n31387 );
buf ( n31389 , n582 );
not ( n31390 , n31389 );
buf ( n31391 , n28661 );
not ( n31392 , n31391 );
or ( n31393 , n31390 , n31392 );
buf ( n31394 , n24450 );
not ( n31395 , n31394 );
buf ( n31396 , n18303 );
nand ( n31397 , n31395 , n31396 );
buf ( n31398 , n31397 );
buf ( n31399 , n31398 );
nand ( n31400 , n31393 , n31399 );
buf ( n31401 , n31400 );
buf ( n31402 , n31401 );
not ( n31403 , n31402 );
or ( n31404 , n31388 , n31403 );
buf ( n31405 , n31333 );
buf ( n31406 , n18657 );
nand ( n31407 , n31405 , n31406 );
buf ( n31408 , n31407 );
buf ( n31409 , n31408 );
nand ( n31410 , n31404 , n31409 );
buf ( n31411 , n31410 );
buf ( n31412 , n31411 );
and ( n31413 , n31386 , n31412 );
and ( n31414 , n31359 , n31385 );
or ( n31415 , n31413 , n31414 );
buf ( n31416 , n31415 );
buf ( n31417 , n31416 );
xor ( n31418 , n31341 , n31417 );
xor ( n31419 , n31018 , n31043 );
xor ( n31420 , n31419 , n31070 );
buf ( n31421 , n31420 );
buf ( n31422 , n31421 );
xor ( n31423 , n31418 , n31422 );
buf ( n31424 , n31423 );
buf ( n31425 , n31424 );
buf ( n31426 , n586 );
not ( n31427 , n31426 );
buf ( n31428 , n18163 );
not ( n31429 , n31428 );
or ( n31430 , n31427 , n31429 );
buf ( n31431 , n18164 );
buf ( n31432 , n18840 );
nand ( n31433 , n31431 , n31432 );
buf ( n31434 , n31433 );
buf ( n31435 , n31434 );
nand ( n31436 , n31430 , n31435 );
buf ( n31437 , n31436 );
nand ( n31438 , n18856 , n23249 );
nand ( n31439 , n31437 , n31438 );
buf ( n31440 , n31439 );
buf ( n31441 , n18479 );
not ( n31442 , n31441 );
not ( n31443 , n584 );
not ( n31444 , n24512 );
or ( n31445 , n31443 , n31444 );
buf ( n31446 , n30007 );
buf ( n31447 , n18277 );
nand ( n31448 , n31446 , n31447 );
buf ( n31449 , n31448 );
nand ( n31450 , n31445 , n31449 );
buf ( n31451 , n31450 );
not ( n31452 , n31451 );
or ( n31453 , n31442 , n31452 );
buf ( n31454 , n31171 );
buf ( n31455 , n18431 );
nand ( n31456 , n31454 , n31455 );
buf ( n31457 , n31456 );
buf ( n31458 , n31457 );
nand ( n31459 , n31453 , n31458 );
buf ( n31460 , n31459 );
buf ( n31461 , n31460 );
xor ( n31462 , n31440 , n31461 );
xor ( n31463 , n31107 , n31125 );
xor ( n31464 , n31463 , n31135 );
buf ( n31465 , n31464 );
buf ( n31466 , n31465 );
and ( n31467 , n31462 , n31466 );
and ( n31468 , n31440 , n31461 );
or ( n31469 , n31467 , n31468 );
buf ( n31470 , n31469 );
buf ( n31471 , n31470 );
xor ( n31472 , n31140 , n31161 );
xor ( n31473 , n31472 , n31177 );
buf ( n31474 , n31473 );
buf ( n31475 , n31474 );
xor ( n31476 , n31471 , n31475 );
buf ( n31477 , n18340 );
not ( n31478 , n31477 );
buf ( n31479 , n31122 );
not ( n31480 , n31479 );
or ( n31481 , n31478 , n31480 );
xor ( n31482 , n576 , n20160 );
nand ( n31483 , n31482 , n30529 );
buf ( n31484 , n31483 );
nand ( n31485 , n31481 , n31484 );
buf ( n31486 , n31485 );
buf ( n31487 , n31486 );
buf ( n31488 , n31131 );
xor ( n31489 , n31487 , n31488 );
and ( n31490 , n576 , n13592 );
buf ( n31491 , n31490 );
buf ( n31492 , n18340 );
not ( n31493 , n31492 );
buf ( n31494 , n31493 );
buf ( n31495 , n31494 );
buf ( n31496 , n7809 );
nor ( n31497 , n31495 , n31496 );
buf ( n31498 , n31497 );
nand ( n31499 , n20163 , n31498 );
buf ( n31500 , n31494 );
buf ( n31501 , n576 );
nor ( n31502 , n31500 , n31501 );
buf ( n31503 , n31502 );
nand ( n31504 , n20160 , n31503 );
xor ( n31505 , n576 , n18203 );
nand ( n31506 , n31505 , n18365 );
nand ( n31507 , n31499 , n31504 , n31506 );
buf ( n31508 , n31507 );
xor ( n31509 , n31491 , n31508 );
buf ( n31510 , n10822 );
buf ( n31511 , n576 );
nand ( n31512 , n31510 , n31511 );
buf ( n31513 , n31512 );
buf ( n31514 , n31513 );
not ( n31515 , n31514 );
buf ( n31516 , n31515 );
buf ( n31517 , n31516 );
and ( n31518 , n31509 , n31517 );
and ( n31519 , n31491 , n31508 );
or ( n31520 , n31518 , n31519 );
buf ( n31521 , n31520 );
buf ( n31522 , n31521 );
and ( n31523 , n31489 , n31522 );
and ( n31524 , n31487 , n31488 );
or ( n31525 , n31523 , n31524 );
buf ( n31526 , n31525 );
buf ( n31527 , n31526 );
xor ( n31528 , n31359 , n31385 );
xor ( n31529 , n31528 , n31412 );
buf ( n31530 , n31529 );
buf ( n31531 , n31530 );
xor ( n31532 , n31527 , n31531 );
buf ( n31533 , n18392 );
not ( n31534 , n31533 );
buf ( n31535 , n18402 );
not ( n31536 , n31535 );
buf ( n31537 , n19783 );
not ( n31538 , n31537 );
or ( n31539 , n31536 , n31538 );
buf ( n31540 , n24324 );
buf ( n31541 , n580 );
nand ( n31542 , n31540 , n31541 );
buf ( n31543 , n31542 );
buf ( n31544 , n31543 );
nand ( n31545 , n31539 , n31544 );
buf ( n31546 , n31545 );
buf ( n31547 , n31546 );
not ( n31548 , n31547 );
or ( n31549 , n31534 , n31548 );
buf ( n31550 , n580 );
not ( n31551 , n31550 );
buf ( n31552 , n30582 );
not ( n31553 , n31552 );
or ( n31554 , n31551 , n31553 );
buf ( n31555 , n31350 );
nand ( n31556 , n31554 , n31555 );
buf ( n31557 , n31556 );
buf ( n31558 , n31557 );
buf ( n31559 , n18418 );
nand ( n31560 , n31558 , n31559 );
buf ( n31561 , n31560 );
buf ( n31562 , n31561 );
nand ( n31563 , n31549 , n31562 );
buf ( n31564 , n31563 );
buf ( n31565 , n31564 );
buf ( n31566 , n18219 );
not ( n31567 , n31566 );
buf ( n31568 , n31374 );
not ( n31569 , n31568 );
or ( n31570 , n31567 , n31569 );
buf ( n31571 , n578 );
not ( n31572 , n31571 );
buf ( n31573 , n18726 );
not ( n31574 , n31573 );
or ( n31575 , n31572 , n31574 );
buf ( n31576 , n18725 );
buf ( n31577 , n18233 );
nand ( n31578 , n31576 , n31577 );
buf ( n31579 , n31578 );
buf ( n31580 , n31579 );
nand ( n31581 , n31575 , n31580 );
buf ( n31582 , n31581 );
buf ( n31583 , n31582 );
buf ( n31584 , n18264 );
nand ( n31585 , n31583 , n31584 );
buf ( n31586 , n31585 );
buf ( n31587 , n31586 );
nand ( n31588 , n31570 , n31587 );
buf ( n31589 , n31588 );
buf ( n31590 , n31589 );
xor ( n31591 , n31565 , n31590 );
buf ( n31592 , n18316 );
not ( n31593 , n31592 );
buf ( n31594 , n582 );
not ( n31595 , n31594 );
buf ( n31596 , n24346 );
not ( n31597 , n31596 );
or ( n31598 , n31595 , n31597 );
buf ( n31599 , n19209 );
buf ( n31600 , n18303 );
nand ( n31601 , n31599 , n31600 );
buf ( n31602 , n31601 );
buf ( n31603 , n31602 );
nand ( n31604 , n31598 , n31603 );
buf ( n31605 , n31604 );
buf ( n31606 , n31605 );
not ( n31607 , n31606 );
or ( n31608 , n31593 , n31607 );
buf ( n31609 , n31401 );
buf ( n31610 , n18657 );
nand ( n31611 , n31609 , n31610 );
buf ( n31612 , n31611 );
buf ( n31613 , n31612 );
nand ( n31614 , n31608 , n31613 );
buf ( n31615 , n31614 );
buf ( n31616 , n31615 );
and ( n31617 , n31591 , n31616 );
and ( n31618 , n31565 , n31590 );
or ( n31619 , n31617 , n31618 );
buf ( n31620 , n31619 );
buf ( n31621 , n31620 );
and ( n31622 , n31532 , n31621 );
and ( n31623 , n31527 , n31531 );
or ( n31624 , n31622 , n31623 );
buf ( n31625 , n31624 );
buf ( n31626 , n31625 );
xor ( n31627 , n31476 , n31626 );
buf ( n31628 , n31627 );
buf ( n31629 , n31628 );
xor ( n31630 , n31425 , n31629 );
xor ( n31631 , n31440 , n31461 );
xor ( n31632 , n31631 , n31466 );
buf ( n31633 , n31632 );
buf ( n31634 , n31633 );
buf ( n31635 , n18881 );
not ( n31636 , n31635 );
buf ( n31637 , n586 );
not ( n31638 , n31637 );
buf ( n31639 , n30596 );
not ( n31640 , n31639 );
or ( n31641 , n31638 , n31640 );
buf ( n31642 , n24497 );
buf ( n31643 , n18840 );
nand ( n31644 , n31642 , n31643 );
buf ( n31645 , n31644 );
buf ( n31646 , n31645 );
nand ( n31647 , n31641 , n31646 );
buf ( n31648 , n31647 );
buf ( n31649 , n31648 );
not ( n31650 , n31649 );
or ( n31651 , n31636 , n31650 );
buf ( n31652 , n31437 );
buf ( n31653 , n18857 );
nand ( n31654 , n31652 , n31653 );
buf ( n31655 , n31654 );
buf ( n31656 , n31655 );
nand ( n31657 , n31651 , n31656 );
buf ( n31658 , n31657 );
buf ( n31659 , n31658 );
buf ( n31660 , n18431 );
not ( n31661 , n31660 );
buf ( n31662 , n31450 );
not ( n31663 , n31662 );
or ( n31664 , n31661 , n31663 );
buf ( n31665 , n584 );
not ( n31666 , n31665 );
buf ( n31667 , n30542 );
not ( n31668 , n31667 );
or ( n31669 , n31666 , n31668 );
buf ( n31670 , n30548 );
buf ( n31671 , n18277 );
nand ( n31672 , n31670 , n31671 );
buf ( n31673 , n31672 );
buf ( n31674 , n31673 );
nand ( n31675 , n31669 , n31674 );
buf ( n31676 , n31675 );
buf ( n31677 , n31676 );
buf ( n31678 , n18479 );
nand ( n31679 , n31677 , n31678 );
buf ( n31680 , n31679 );
buf ( n31681 , n31680 );
nand ( n31682 , n31664 , n31681 );
buf ( n31683 , n31682 );
buf ( n31684 , n31683 );
xor ( n31685 , n31659 , n31684 );
buf ( n31686 , n18219 );
not ( n31687 , n31686 );
buf ( n31688 , n31582 );
not ( n31689 , n31688 );
or ( n31690 , n31687 , n31689 );
buf ( n31691 , n578 );
not ( n31692 , n31691 );
buf ( n31693 , n18442 );
not ( n31694 , n31693 );
or ( n31695 , n31692 , n31694 );
buf ( n31696 , n20629 );
buf ( n31697 , n18233 );
nand ( n31698 , n31696 , n31697 );
buf ( n31699 , n31698 );
buf ( n31700 , n31699 );
nand ( n31701 , n31695 , n31700 );
buf ( n31702 , n31701 );
buf ( n31703 , n31702 );
buf ( n31704 , n18264 );
nand ( n31705 , n31703 , n31704 );
buf ( n31706 , n31705 );
buf ( n31707 , n31706 );
nand ( n31708 , n31690 , n31707 );
buf ( n31709 , n31708 );
buf ( n31710 , n31709 );
buf ( n31711 , n18392 );
not ( n31712 , n31711 );
and ( n31713 , n18082 , n18402 );
not ( n31714 , n18082 );
and ( n31715 , n31714 , n580 );
or ( n31716 , n31713 , n31715 );
buf ( n31717 , n31716 );
not ( n31718 , n31717 );
or ( n31719 , n31712 , n31718 );
buf ( n31720 , n31546 );
buf ( n31721 , n18418 );
nand ( n31722 , n31720 , n31721 );
buf ( n31723 , n31722 );
buf ( n31724 , n31723 );
nand ( n31725 , n31719 , n31724 );
buf ( n31726 , n31725 );
buf ( n31727 , n31726 );
xor ( n31728 , n31710 , n31727 );
buf ( n31729 , n18657 );
not ( n31730 , n31729 );
buf ( n31731 , n31605 );
not ( n31732 , n31731 );
or ( n31733 , n31730 , n31732 );
buf ( n31734 , n582 );
not ( n31735 , n31734 );
not ( n31736 , n19181 );
buf ( n31737 , n31736 );
not ( n31738 , n31737 );
or ( n31739 , n31735 , n31738 );
buf ( n31740 , n18184 );
buf ( n31741 , n18303 );
nand ( n31742 , n31740 , n31741 );
buf ( n31743 , n31742 );
buf ( n31744 , n31743 );
nand ( n31745 , n31739 , n31744 );
buf ( n31746 , n31745 );
buf ( n31747 , n31746 );
buf ( n31748 , n18316 );
nand ( n31749 , n31747 , n31748 );
buf ( n31750 , n31749 );
buf ( n31751 , n31750 );
nand ( n31752 , n31733 , n31751 );
buf ( n31753 , n31752 );
buf ( n31754 , n31753 );
and ( n31755 , n31728 , n31754 );
and ( n31756 , n31710 , n31727 );
or ( n31757 , n31755 , n31756 );
buf ( n31758 , n31757 );
buf ( n31759 , n31758 );
and ( n31760 , n31685 , n31759 );
and ( n31761 , n31659 , n31684 );
or ( n31762 , n31760 , n31761 );
buf ( n31763 , n31762 );
buf ( n31764 , n31763 );
xor ( n31765 , n31634 , n31764 );
xor ( n31766 , n31487 , n31488 );
xor ( n31767 , n31766 , n31522 );
buf ( n31768 , n31767 );
buf ( n31769 , n31768 );
not ( n31770 , n18340 );
not ( n31771 , n31505 );
or ( n31772 , n31770 , n31771 );
xor ( n31773 , n576 , n13592 );
nand ( n31774 , n31773 , n18365 );
nand ( n31775 , n31772 , n31774 );
buf ( n31776 , n31775 );
not ( n31777 , n18365 );
buf ( n31778 , n576 );
not ( n31779 , n31778 );
buf ( n31780 , n18397 );
not ( n31781 , n31780 );
or ( n31782 , n31779 , n31781 );
buf ( n31783 , n10819 );
buf ( n31784 , n7809 );
nand ( n31785 , n31783 , n31784 );
buf ( n31786 , n31785 );
buf ( n31787 , n31786 );
nand ( n31788 , n31782 , n31787 );
buf ( n31789 , n31788 );
not ( n31790 , n31789 );
or ( n31791 , n31777 , n31790 );
nand ( n31792 , n31773 , n18340 );
nand ( n31793 , n31791 , n31792 );
buf ( n31794 , n31793 );
xor ( n31795 , n31776 , n31794 );
buf ( n31796 , n31513 );
and ( n31797 , n31795 , n31796 );
and ( n31798 , n31776 , n31794 );
or ( n31799 , n31797 , n31798 );
buf ( n31800 , n31799 );
buf ( n31801 , n31800 );
xor ( n31802 , n31491 , n31508 );
xor ( n31803 , n31802 , n31517 );
buf ( n31804 , n31803 );
buf ( n31805 , n31804 );
xor ( n31806 , n31801 , n31805 );
buf ( n31807 , n18431 );
not ( n31808 , n31807 );
buf ( n31809 , n31676 );
not ( n31810 , n31809 );
or ( n31811 , n31808 , n31810 );
and ( n31812 , n19403 , n18277 );
not ( n31813 , n19403 );
and ( n31814 , n31813 , n584 );
or ( n31815 , n31812 , n31814 );
buf ( n31816 , n31815 );
buf ( n31817 , n18479 );
nand ( n31818 , n31816 , n31817 );
buf ( n31819 , n31818 );
buf ( n31820 , n31819 );
nand ( n31821 , n31811 , n31820 );
buf ( n31822 , n31821 );
buf ( n31823 , n31822 );
and ( n31824 , n31806 , n31823 );
and ( n31825 , n31801 , n31805 );
or ( n31826 , n31824 , n31825 );
buf ( n31827 , n31826 );
buf ( n31828 , n31827 );
xor ( n31829 , n31769 , n31828 );
xor ( n31830 , n31565 , n31590 );
xor ( n31831 , n31830 , n31616 );
buf ( n31832 , n31831 );
buf ( n31833 , n31832 );
and ( n31834 , n31829 , n31833 );
and ( n31835 , n31769 , n31828 );
or ( n31836 , n31834 , n31835 );
buf ( n31837 , n31836 );
buf ( n31838 , n31837 );
and ( n31839 , n31765 , n31838 );
and ( n31840 , n31634 , n31764 );
or ( n31841 , n31839 , n31840 );
buf ( n31842 , n31841 );
buf ( n31843 , n31842 );
xor ( n31844 , n31630 , n31843 );
buf ( n31845 , n31844 );
not ( n31846 , n31845 );
xor ( n31847 , n31527 , n31531 );
xor ( n31848 , n31847 , n31621 );
buf ( n31849 , n31848 );
buf ( n31850 , n31849 );
xor ( n31851 , n31634 , n31764 );
xor ( n31852 , n31851 , n31838 );
buf ( n31853 , n31852 );
buf ( n31854 , n31853 );
xor ( n31855 , n31850 , n31854 );
xor ( n31856 , n31659 , n31684 );
xor ( n31857 , n31856 , n31759 );
buf ( n31858 , n31857 );
buf ( n31859 , n31858 );
buf ( n31860 , n21813 );
not ( n31861 , n31860 );
buf ( n31862 , n19151 );
not ( n31863 , n31862 );
or ( n31864 , n31861 , n31863 );
buf ( n31865 , n588 );
not ( n31866 , n31865 );
buf ( n31867 , n18163 );
not ( n31868 , n31867 );
or ( n31869 , n31866 , n31868 );
buf ( n31870 , n588 );
not ( n31871 , n31870 );
buf ( n31872 , n18164 );
nand ( n31873 , n31871 , n31872 );
buf ( n31874 , n31873 );
buf ( n31875 , n31874 );
nand ( n31876 , n31869 , n31875 );
buf ( n31877 , n31876 );
buf ( n31878 , n31877 );
nand ( n31879 , n31864 , n31878 );
buf ( n31880 , n31879 );
buf ( n31881 , n31880 );
buf ( n31882 , n18881 );
not ( n31883 , n31882 );
buf ( n31884 , n586 );
not ( n31885 , n31884 );
buf ( n31886 , n30019 );
not ( n31887 , n31886 );
or ( n31888 , n31885 , n31887 );
buf ( n31889 , n30007 );
buf ( n31890 , n18840 );
nand ( n31891 , n31889 , n31890 );
buf ( n31892 , n31891 );
buf ( n31893 , n31892 );
nand ( n31894 , n31888 , n31893 );
buf ( n31895 , n31894 );
buf ( n31896 , n31895 );
not ( n31897 , n31896 );
or ( n31898 , n31883 , n31897 );
buf ( n31899 , n31648 );
buf ( n31900 , n18857 );
nand ( n31901 , n31899 , n31900 );
buf ( n31902 , n31901 );
buf ( n31903 , n31902 );
nand ( n31904 , n31898 , n31903 );
buf ( n31905 , n31904 );
buf ( n31906 , n31905 );
xor ( n31907 , n31881 , n31906 );
buf ( n31908 , n18219 );
not ( n31909 , n31908 );
buf ( n31910 , n31702 );
not ( n31911 , n31910 );
or ( n31912 , n31909 , n31911 );
and ( n31913 , n15680 , n18233 );
not ( n31914 , n15680 );
and ( n31915 , n31914 , n578 );
or ( n31916 , n31913 , n31915 );
buf ( n31917 , n31916 );
buf ( n31918 , n18264 );
nand ( n31919 , n31917 , n31918 );
buf ( n31920 , n31919 );
buf ( n31921 , n31920 );
nand ( n31922 , n31912 , n31921 );
buf ( n31923 , n31922 );
buf ( n31924 , n31923 );
buf ( n31925 , n18418 );
not ( n31926 , n31925 );
buf ( n31927 , n31716 );
not ( n31928 , n31927 );
or ( n31929 , n31926 , n31928 );
buf ( n31930 , n580 );
not ( n31931 , n31930 );
buf ( n31932 , n19761 );
not ( n31933 , n31932 );
or ( n31934 , n31931 , n31933 );
buf ( n31935 , n18725 );
buf ( n31936 , n18402 );
nand ( n31937 , n31935 , n31936 );
buf ( n31938 , n31937 );
buf ( n31939 , n31938 );
nand ( n31940 , n31934 , n31939 );
buf ( n31941 , n31940 );
buf ( n31942 , n31941 );
buf ( n31943 , n18392 );
nand ( n31944 , n31942 , n31943 );
buf ( n31945 , n31944 );
buf ( n31946 , n31945 );
nand ( n31947 , n31929 , n31946 );
buf ( n31948 , n31947 );
buf ( n31949 , n31948 );
xor ( n31950 , n31924 , n31949 );
buf ( n31951 , n10854 );
buf ( n31952 , n576 );
and ( n31953 , n31951 , n31952 );
buf ( n31954 , n31953 );
buf ( n31955 , n31954 );
not ( n31956 , n31793 );
buf ( n31957 , n31956 );
xor ( n31958 , n31955 , n31957 );
buf ( n31959 , n18219 );
not ( n31960 , n31959 );
buf ( n31961 , n31916 );
not ( n31962 , n31961 );
or ( n31963 , n31960 , n31962 );
buf ( n31964 , n578 );
not ( n31965 , n31964 );
buf ( n31966 , n18296 );
not ( n31967 , n31966 );
or ( n31968 , n31965 , n31967 );
buf ( n31969 , n18203 );
buf ( n31970 , n18233 );
nand ( n31971 , n31969 , n31970 );
buf ( n31972 , n31971 );
buf ( n31973 , n31972 );
nand ( n31974 , n31968 , n31973 );
buf ( n31975 , n31974 );
buf ( n31976 , n31975 );
buf ( n31977 , n18264 );
nand ( n31978 , n31976 , n31977 );
buf ( n31979 , n31978 );
buf ( n31980 , n31979 );
nand ( n31981 , n31963 , n31980 );
buf ( n31982 , n31981 );
buf ( n31983 , n31982 );
and ( n31984 , n31958 , n31983 );
and ( n31985 , n31955 , n31957 );
or ( n31986 , n31984 , n31985 );
buf ( n31987 , n31986 );
buf ( n31988 , n31987 );
and ( n31989 , n31950 , n31988 );
and ( n31990 , n31924 , n31949 );
or ( n31991 , n31989 , n31990 );
buf ( n31992 , n31991 );
buf ( n31993 , n31992 );
and ( n31994 , n31907 , n31993 );
and ( n31995 , n31881 , n31906 );
or ( n31996 , n31994 , n31995 );
buf ( n31997 , n31996 );
buf ( n31998 , n31997 );
xor ( n31999 , n31859 , n31998 );
not ( n32000 , n18316 );
buf ( n32001 , n18303 );
not ( n32002 , n32001 );
buf ( n32003 , n18137 );
not ( n32004 , n32003 );
or ( n32005 , n32002 , n32004 );
buf ( n32006 , n24324 );
buf ( n32007 , n582 );
nand ( n32008 , n32006 , n32007 );
buf ( n32009 , n32008 );
buf ( n32010 , n32009 );
nand ( n32011 , n32005 , n32010 );
buf ( n32012 , n32011 );
not ( n32013 , n32012 );
or ( n32014 , n32000 , n32013 );
not ( n32015 , n31743 );
nand ( n32016 , n31736 , n582 );
not ( n32017 , n32016 );
or ( n32018 , n32015 , n32017 );
nand ( n32019 , n32018 , n18657 );
nand ( n32020 , n32014 , n32019 );
buf ( n32021 , n32020 );
xor ( n32022 , n31776 , n31794 );
xor ( n32023 , n32022 , n31796 );
buf ( n32024 , n32023 );
buf ( n32025 , n32024 );
xor ( n32026 , n32021 , n32025 );
buf ( n32027 , n18431 );
not ( n32028 , n32027 );
buf ( n32029 , n31815 );
not ( n32030 , n32029 );
or ( n32031 , n32028 , n32030 );
buf ( n32032 , n19209 );
not ( n32033 , n32032 );
buf ( n32034 , n584 );
nand ( n32035 , n32033 , n32034 );
buf ( n32036 , n32035 );
buf ( n32037 , n32036 );
not ( n32038 , n32037 );
buf ( n32039 , n24346 );
not ( n32040 , n32039 );
buf ( n32041 , n18277 );
nand ( n32042 , n32040 , n32041 );
buf ( n32043 , n32042 );
buf ( n32044 , n32043 );
not ( n32045 , n32044 );
or ( n32046 , n32038 , n32045 );
buf ( n32047 , n18479 );
nand ( n32048 , n32046 , n32047 );
buf ( n32049 , n32048 );
buf ( n32050 , n32049 );
nand ( n32051 , n32031 , n32050 );
buf ( n32052 , n32051 );
buf ( n32053 , n32052 );
and ( n32054 , n32026 , n32053 );
and ( n32055 , n32021 , n32025 );
or ( n32056 , n32054 , n32055 );
buf ( n32057 , n32056 );
buf ( n32058 , n32057 );
xor ( n32059 , n31710 , n31727 );
xor ( n32060 , n32059 , n31754 );
buf ( n32061 , n32060 );
buf ( n32062 , n32061 );
xor ( n32063 , n32058 , n32062 );
xor ( n32064 , n31801 , n31805 );
xor ( n32065 , n32064 , n31823 );
buf ( n32066 , n32065 );
buf ( n32067 , n32066 );
and ( n32068 , n32063 , n32067 );
and ( n32069 , n32058 , n32062 );
or ( n32070 , n32068 , n32069 );
buf ( n32071 , n32070 );
buf ( n32072 , n32071 );
and ( n32073 , n31999 , n32072 );
and ( n32074 , n31859 , n31998 );
or ( n32075 , n32073 , n32074 );
buf ( n32076 , n32075 );
buf ( n32077 , n32076 );
and ( n32078 , n31855 , n32077 );
and ( n32079 , n31850 , n31854 );
or ( n32080 , n32078 , n32079 );
buf ( n32081 , n32080 );
not ( n32082 , n32081 );
and ( n32083 , n31846 , n32082 );
xor ( n32084 , n31850 , n31854 );
xor ( n32085 , n32084 , n32077 );
buf ( n32086 , n32085 );
xor ( n32087 , n31769 , n31828 );
xor ( n32088 , n32087 , n31833 );
buf ( n32089 , n32088 );
buf ( n32090 , n32089 );
xor ( n32091 , n31859 , n31998 );
xor ( n32092 , n32091 , n32072 );
buf ( n32093 , n32092 );
buf ( n32094 , n32093 );
xor ( n32095 , n32090 , n32094 );
xor ( n32096 , n31881 , n31906 );
xor ( n32097 , n32096 , n31993 );
buf ( n32098 , n32097 );
buf ( n32099 , n32098 );
buf ( n32100 , n19152 );
not ( n32101 , n32100 );
and ( n32102 , n588 , n30596 );
not ( n32103 , n588 );
and ( n32104 , n32103 , n24497 );
or ( n32105 , n32102 , n32104 );
buf ( n32106 , n32105 );
not ( n32107 , n32106 );
or ( n32108 , n32101 , n32107 );
buf ( n32109 , n31877 );
buf ( n32110 , n19143 );
nand ( n32111 , n32109 , n32110 );
buf ( n32112 , n32111 );
buf ( n32113 , n32112 );
nand ( n32114 , n32108 , n32113 );
buf ( n32115 , n32114 );
buf ( n32116 , n32115 );
buf ( n32117 , n18857 );
not ( n32118 , n32117 );
buf ( n32119 , n31895 );
not ( n32120 , n32119 );
or ( n32121 , n32118 , n32120 );
buf ( n32122 , n19398 );
not ( n32123 , n32122 );
buf ( n32124 , n18840 );
not ( n32125 , n32124 );
and ( n32126 , n32123 , n32125 );
buf ( n32127 , n24462 );
not ( n32128 , n32127 );
buf ( n32129 , n32128 );
buf ( n32130 , n32129 );
buf ( n32131 , n18840 );
and ( n32132 , n32130 , n32131 );
nor ( n32133 , n32126 , n32132 );
buf ( n32134 , n32133 );
buf ( n32135 , n32134 );
not ( n32136 , n32135 );
buf ( n32137 , n18881 );
nand ( n32138 , n32136 , n32137 );
buf ( n32139 , n32138 );
buf ( n32140 , n32139 );
nand ( n32141 , n32121 , n32140 );
buf ( n32142 , n32141 );
buf ( n32143 , n32142 );
xor ( n32144 , n32116 , n32143 );
buf ( n32145 , n18418 );
not ( n32146 , n32145 );
buf ( n32147 , n31941 );
not ( n32148 , n32147 );
or ( n32149 , n32146 , n32148 );
buf ( n32150 , n580 );
not ( n32151 , n32150 );
buf ( n32152 , n18442 );
not ( n32153 , n32152 );
or ( n32154 , n32151 , n32153 );
buf ( n32155 , n18861 );
buf ( n32156 , n18402 );
nand ( n32157 , n32155 , n32156 );
buf ( n32158 , n32157 );
buf ( n32159 , n32158 );
nand ( n32160 , n32154 , n32159 );
buf ( n32161 , n32160 );
buf ( n32162 , n32161 );
buf ( n32163 , n18392 );
nand ( n32164 , n32162 , n32163 );
buf ( n32165 , n32164 );
buf ( n32166 , n32165 );
nand ( n32167 , n32149 , n32166 );
buf ( n32168 , n32167 );
buf ( n32169 , n32168 );
buf ( n32170 , n18340 );
not ( n32171 , n32170 );
buf ( n32172 , n31789 );
not ( n32173 , n32172 );
or ( n32174 , n32171 , n32173 );
nand ( n32175 , n24295 , n18365 );
buf ( n32176 , n32175 );
nand ( n32177 , n32174 , n32176 );
buf ( n32178 , n32177 );
buf ( n32179 , n32178 );
and ( n32180 , n24188 , n24189 );
buf ( n32181 , n32180 );
buf ( n32182 , n32181 );
xor ( n32183 , n32179 , n32182 );
buf ( n32184 , n18219 );
not ( n32185 , n32184 );
buf ( n32186 , n31975 );
not ( n32187 , n32186 );
or ( n32188 , n32185 , n32187 );
not ( n32189 , n24278 );
not ( n32190 , n24273 );
or ( n32191 , n32189 , n32190 );
nand ( n32192 , n32191 , n18264 );
buf ( n32193 , n32192 );
nand ( n32194 , n32188 , n32193 );
buf ( n32195 , n32194 );
buf ( n32196 , n32195 );
and ( n32197 , n32183 , n32196 );
and ( n32198 , n32179 , n32182 );
or ( n32199 , n32197 , n32198 );
buf ( n32200 , n32199 );
buf ( n32201 , n32200 );
xor ( n32202 , n32169 , n32201 );
buf ( n32203 , n18316 );
not ( n32204 , n32203 );
nand ( n32205 , n582 , n24218 );
buf ( n32206 , n18303 );
buf ( n32207 , n18082 );
nand ( n32208 , n32206 , n32207 );
buf ( n32209 , n32208 );
nand ( n32210 , n32205 , n32209 );
buf ( n32211 , n32210 );
not ( n32212 , n32211 );
or ( n32213 , n32204 , n32212 );
buf ( n32214 , n32012 );
buf ( n32215 , n18657 );
nand ( n32216 , n32214 , n32215 );
buf ( n32217 , n32216 );
buf ( n32218 , n32217 );
nand ( n32219 , n32213 , n32218 );
buf ( n32220 , n32219 );
buf ( n32221 , n32220 );
and ( n32222 , n32202 , n32221 );
and ( n32223 , n32169 , n32201 );
or ( n32224 , n32222 , n32223 );
buf ( n32225 , n32224 );
buf ( n32226 , n32225 );
and ( n32227 , n32144 , n32226 );
and ( n32228 , n32116 , n32143 );
or ( n32229 , n32227 , n32228 );
buf ( n32230 , n32229 );
buf ( n32231 , n32230 );
xor ( n32232 , n32099 , n32231 );
buf ( n32233 , n19387 );
not ( n32234 , n32233 );
buf ( n32235 , n18916 );
nand ( n32236 , n32234 , n32235 );
buf ( n32237 , n32236 );
buf ( n32238 , n32237 );
buf ( n32239 , n19181 );
not ( n32240 , n32239 );
buf ( n32241 , n23060 );
nand ( n32242 , n32240 , n32241 );
buf ( n32243 , n32242 );
buf ( n32244 , n32243 );
buf ( n32245 , n19181 );
buf ( n32246 , n24312 );
nand ( n32247 , n32245 , n32246 );
buf ( n32248 , n32247 );
buf ( n32249 , n32248 );
buf ( n32250 , n19387 );
buf ( n32251 , n18936 );
nand ( n32252 , n32250 , n32251 );
buf ( n32253 , n32252 );
buf ( n32254 , n32253 );
nand ( n32255 , n32238 , n32244 , n32249 , n32254 );
buf ( n32256 , n32255 );
buf ( n32257 , n32256 );
xor ( n32258 , n31955 , n31957 );
xor ( n32259 , n32258 , n31983 );
buf ( n32260 , n32259 );
buf ( n32261 , n32260 );
xor ( n32262 , n32257 , n32261 );
buf ( n32263 , n18881 );
not ( n32264 , n32263 );
buf ( n32265 , n19403 );
buf ( n32266 , n586 );
and ( n32267 , n32265 , n32266 );
not ( n32268 , n32265 );
buf ( n32269 , n18840 );
and ( n32270 , n32268 , n32269 );
nor ( n32271 , n32267 , n32270 );
buf ( n32272 , n32271 );
buf ( n32273 , n32272 );
not ( n32274 , n32273 );
or ( n32275 , n32264 , n32274 );
buf ( n32276 , n32134 );
buf ( n32277 , n18856 );
or ( n32278 , n32276 , n32277 );
nand ( n32279 , n32275 , n32278 );
buf ( n32280 , n32279 );
buf ( n32281 , n32280 );
and ( n32282 , n32262 , n32281 );
and ( n32283 , n32257 , n32261 );
or ( n32284 , n32282 , n32283 );
buf ( n32285 , n32284 );
buf ( n32286 , n32285 );
xor ( n32287 , n31924 , n31949 );
xor ( n32288 , n32287 , n31988 );
buf ( n32289 , n32288 );
buf ( n32290 , n32289 );
xor ( n32291 , n32286 , n32290 );
xor ( n32292 , n32021 , n32025 );
xor ( n32293 , n32292 , n32053 );
buf ( n32294 , n32293 );
buf ( n32295 , n32294 );
and ( n32296 , n32291 , n32295 );
and ( n32297 , n32286 , n32290 );
or ( n32298 , n32296 , n32297 );
buf ( n32299 , n32298 );
buf ( n32300 , n32299 );
and ( n32301 , n32232 , n32300 );
and ( n32302 , n32099 , n32231 );
or ( n32303 , n32301 , n32302 );
buf ( n32304 , n32303 );
buf ( n32305 , n32304 );
and ( n32306 , n32095 , n32305 );
and ( n32307 , n32090 , n32094 );
or ( n32308 , n32306 , n32307 );
buf ( n32309 , n32308 );
nor ( n32310 , n32086 , n32309 );
nor ( n32311 , n32083 , n32310 );
xor ( n32312 , n31341 , n31417 );
and ( n32313 , n32312 , n31422 );
and ( n32314 , n31341 , n31417 );
or ( n32315 , n32313 , n32314 );
buf ( n32316 , n32315 );
buf ( n32317 , n32316 );
xor ( n32318 , n31182 , n31186 );
xor ( n32319 , n32318 , n31191 );
buf ( n32320 , n32319 );
buf ( n32321 , n32320 );
xor ( n32322 , n32317 , n32321 );
xor ( n32323 , n31471 , n31475 );
and ( n32324 , n32323 , n31626 );
and ( n32325 , n31471 , n31475 );
or ( n32326 , n32324 , n32325 );
buf ( n32327 , n32326 );
buf ( n32328 , n32327 );
xor ( n32329 , n32322 , n32328 );
buf ( n32330 , n32329 );
not ( n32331 , n32330 );
xor ( n32332 , n31425 , n31629 );
and ( n32333 , n32332 , n31843 );
and ( n32334 , n31425 , n31629 );
or ( n32335 , n32333 , n32334 );
buf ( n32336 , n32335 );
not ( n32337 , n32336 );
and ( n32338 , n32331 , n32337 );
xor ( n32339 , n31100 , n31104 );
xor ( n32340 , n32339 , n31196 );
buf ( n32341 , n32340 );
not ( n32342 , n32341 );
xor ( n32343 , n32317 , n32321 );
and ( n32344 , n32343 , n32328 );
and ( n32345 , n32317 , n32321 );
or ( n32346 , n32344 , n32345 );
buf ( n32347 , n32346 );
not ( n32348 , n32347 );
and ( n32349 , n32342 , n32348 );
nor ( n32350 , n32338 , n32349 );
nand ( n32351 , n32311 , n32350 );
buf ( n32352 , n32351 );
not ( n32353 , n32352 );
buf ( n32354 , n32353 );
not ( n32355 , n32354 );
xor ( n32356 , n32286 , n32290 );
xor ( n32357 , n32356 , n32295 );
buf ( n32358 , n32357 );
buf ( n32359 , n32358 );
buf ( n32360 , n18857 );
not ( n32361 , n32360 );
buf ( n32362 , n32272 );
not ( n32363 , n32362 );
or ( n32364 , n32361 , n32363 );
buf ( n32365 , n24356 );
buf ( n32366 , n18881 );
nand ( n32367 , n32365 , n32366 );
buf ( n32368 , n32367 );
buf ( n32369 , n32368 );
nand ( n32370 , n32364 , n32369 );
buf ( n32371 , n32370 );
buf ( n32372 , n32371 );
buf ( n32373 , n19143 );
not ( n32374 , n32373 );
xor ( n32375 , n588 , n30007 );
buf ( n32376 , n32375 );
not ( n32377 , n32376 );
or ( n32378 , n32374 , n32377 );
buf ( n32379 , n24473 );
buf ( n32380 , n19152 );
nand ( n32381 , n32379 , n32380 );
buf ( n32382 , n32381 );
buf ( n32383 , n32382 );
nand ( n32384 , n32378 , n32383 );
buf ( n32385 , n32384 );
buf ( n32386 , n32385 );
xor ( n32387 , n32372 , n32386 );
buf ( n32388 , n19244 );
not ( n32389 , n32388 );
buf ( n32390 , n24506 );
not ( n32391 , n32390 );
or ( n32392 , n32389 , n32391 );
xor ( n32393 , n590 , n18164 );
buf ( n32394 , n32393 );
buf ( n32395 , n591 );
nand ( n32396 , n32394 , n32395 );
buf ( n32397 , n32396 );
buf ( n32398 , n32397 );
nand ( n32399 , n32392 , n32398 );
buf ( n32400 , n32399 );
buf ( n32401 , n32400 );
and ( n32402 , n32387 , n32401 );
and ( n32403 , n32372 , n32386 );
or ( n32404 , n32402 , n32403 );
buf ( n32405 , n32404 );
buf ( n32406 , n32405 );
buf ( n32407 , n23568 );
not ( n32408 , n32407 );
buf ( n32409 , n20622 );
not ( n32410 , n32409 );
or ( n32411 , n32408 , n32410 );
buf ( n32412 , n32393 );
nand ( n32413 , n32411 , n32412 );
buf ( n32414 , n32413 );
buf ( n32415 , n32414 );
buf ( n32416 , n18418 );
not ( n32417 , n32416 );
buf ( n32418 , n32161 );
not ( n32419 , n32418 );
or ( n32420 , n32417 , n32419 );
buf ( n32421 , n24106 );
buf ( n32422 , n18392 );
nand ( n32423 , n32421 , n32422 );
buf ( n32424 , n32423 );
buf ( n32425 , n32424 );
nand ( n32426 , n32420 , n32425 );
buf ( n32427 , n32426 );
buf ( n32428 , n32427 );
xor ( n32429 , n24267 , n24285 );
and ( n32430 , n32429 , n24303 );
and ( n32431 , n24267 , n24285 );
or ( n32432 , n32430 , n32431 );
buf ( n32433 , n32432 );
buf ( n32434 , n32433 );
xor ( n32435 , n32428 , n32434 );
xor ( n32436 , n32179 , n32182 );
xor ( n32437 , n32436 , n32196 );
buf ( n32438 , n32437 );
buf ( n32439 , n32438 );
and ( n32440 , n32435 , n32439 );
and ( n32441 , n32428 , n32434 );
or ( n32442 , n32440 , n32441 );
buf ( n32443 , n32442 );
buf ( n32444 , n32443 );
xor ( n32445 , n32415 , n32444 );
buf ( n32446 , n19143 );
not ( n32447 , n32446 );
buf ( n32448 , n32105 );
not ( n32449 , n32448 );
or ( n32450 , n32447 , n32449 );
buf ( n32451 , n32375 );
buf ( n32452 , n19152 );
nand ( n32453 , n32451 , n32452 );
buf ( n32454 , n32453 );
buf ( n32455 , n32454 );
nand ( n32456 , n32450 , n32455 );
buf ( n32457 , n32456 );
buf ( n32458 , n32457 );
xor ( n32459 , n32445 , n32458 );
buf ( n32460 , n32459 );
buf ( n32461 , n32460 );
xor ( n32462 , n32406 , n32461 );
xor ( n32463 , n32428 , n32434 );
xor ( n32464 , n32463 , n32439 );
buf ( n32465 , n32464 );
buf ( n32466 , n32465 );
xor ( n32467 , n24306 , n24338 );
and ( n32468 , n32467 , n24359 );
and ( n32469 , n24306 , n24338 );
or ( n32470 , n32468 , n32469 );
buf ( n32471 , n32470 );
buf ( n32472 , n32471 );
xor ( n32473 , n32466 , n32472 );
buf ( n32474 , n18479 );
not ( n32475 , n32474 );
buf ( n32476 , n18277 );
buf ( n32477 , n24324 );
and ( n32478 , n32476 , n32477 );
not ( n32479 , n32476 );
buf ( n32480 , n19783 );
and ( n32481 , n32479 , n32480 );
nor ( n32482 , n32478 , n32481 );
buf ( n32483 , n32482 );
buf ( n32484 , n32483 );
not ( n32485 , n32484 );
or ( n32486 , n32475 , n32485 );
buf ( n32487 , n584 );
not ( n32488 , n32487 );
buf ( n32489 , n31736 );
not ( n32490 , n32489 );
or ( n32491 , n32488 , n32490 );
buf ( n32492 , n18277 );
buf ( n32493 , n18184 );
nand ( n32494 , n32492 , n32493 );
buf ( n32495 , n32494 );
buf ( n32496 , n32495 );
nand ( n32497 , n32491 , n32496 );
buf ( n32498 , n32497 );
buf ( n32499 , n32498 );
buf ( n32500 , n18431 );
nand ( n32501 , n32499 , n32500 );
buf ( n32502 , n32501 );
buf ( n32503 , n32502 );
nand ( n32504 , n32486 , n32503 );
buf ( n32505 , n32504 );
buf ( n32506 , n32505 );
not ( n32507 , n18657 );
not ( n32508 , n32210 );
or ( n32509 , n32507 , n32508 );
and ( n32510 , n26807 , n18303 );
not ( n32511 , n26807 );
and ( n32512 , n32511 , n582 );
or ( n32513 , n32510 , n32512 );
nand ( n32514 , n32513 , n18316 );
nand ( n32515 , n32509 , n32514 );
buf ( n32516 , n32515 );
xor ( n32517 , n32506 , n32516 );
xor ( n32518 , n24122 , n24163 );
and ( n32519 , n32518 , n24207 );
and ( n32520 , n24122 , n24163 );
or ( n32521 , n32519 , n32520 );
buf ( n32522 , n32521 );
buf ( n32523 , n32522 );
xor ( n32524 , n32517 , n32523 );
buf ( n32525 , n32524 );
buf ( n32526 , n32525 );
and ( n32527 , n32473 , n32526 );
and ( n32528 , n32466 , n32472 );
or ( n32529 , n32527 , n32528 );
buf ( n32530 , n32529 );
buf ( n32531 , n32530 );
and ( n32532 , n32462 , n32531 );
and ( n32533 , n32406 , n32461 );
or ( n32534 , n32532 , n32533 );
buf ( n32535 , n32534 );
buf ( n32536 , n32535 );
xor ( n32537 , n32359 , n32536 );
xor ( n32538 , n32415 , n32444 );
and ( n32539 , n32538 , n32458 );
and ( n32540 , n32415 , n32444 );
or ( n32541 , n32539 , n32540 );
buf ( n32542 , n32541 );
buf ( n32543 , n32542 );
xor ( n32544 , n32116 , n32143 );
xor ( n32545 , n32544 , n32226 );
buf ( n32546 , n32545 );
buf ( n32547 , n32546 );
xor ( n32548 , n32543 , n32547 );
xor ( n32549 , n32169 , n32201 );
xor ( n32550 , n32549 , n32221 );
buf ( n32551 , n32550 );
buf ( n32552 , n32551 );
xor ( n32553 , n32506 , n32516 );
and ( n32554 , n32553 , n32523 );
and ( n32555 , n32506 , n32516 );
or ( n32556 , n32554 , n32555 );
buf ( n32557 , n32556 );
buf ( n32558 , n32557 );
xor ( n32559 , n32552 , n32558 );
xor ( n32560 , n32257 , n32261 );
xor ( n32561 , n32560 , n32281 );
buf ( n32562 , n32561 );
buf ( n32563 , n32562 );
and ( n32564 , n32559 , n32563 );
and ( n32565 , n32552 , n32558 );
or ( n32566 , n32564 , n32565 );
buf ( n32567 , n32566 );
buf ( n32568 , n32567 );
xor ( n32569 , n32548 , n32568 );
buf ( n32570 , n32569 );
buf ( n32571 , n32570 );
xor ( n32572 , n32537 , n32571 );
buf ( n32573 , n32572 );
buf ( n32574 , n32573 );
xor ( n32575 , n32552 , n32558 );
xor ( n32576 , n32575 , n32563 );
buf ( n32577 , n32576 );
buf ( n32578 , n32577 );
xor ( n32579 , n32406 , n32461 );
xor ( n32580 , n32579 , n32531 );
buf ( n32581 , n32580 );
buf ( n32582 , n32581 );
xor ( n32583 , n32578 , n32582 );
xor ( n32584 , n24481 , n24487 );
and ( n32585 , n32584 , n24522 );
and ( n32586 , n24481 , n24487 );
or ( n32587 , n32585 , n32586 );
buf ( n32588 , n32587 );
buf ( n32589 , n32588 );
xor ( n32590 , n32372 , n32386 );
xor ( n32591 , n32590 , n32401 );
buf ( n32592 , n32591 );
buf ( n32593 , n32592 );
xor ( n32594 , n32589 , n32593 );
xor ( n32595 , n24210 , n24263 );
and ( n32596 , n32595 , n24362 );
and ( n32597 , n24210 , n24263 );
or ( n32598 , n32596 , n32597 );
buf ( n32599 , n32598 );
buf ( n32600 , n32599 );
and ( n32601 , n32594 , n32600 );
and ( n32602 , n32589 , n32593 );
or ( n32603 , n32601 , n32602 );
buf ( n32604 , n32603 );
buf ( n32605 , n32604 );
and ( n32606 , n32583 , n32605 );
and ( n32607 , n32578 , n32582 );
or ( n32608 , n32606 , n32607 );
buf ( n32609 , n32608 );
buf ( n32610 , n32609 );
nor ( n32611 , n32574 , n32610 );
buf ( n32612 , n32611 );
xor ( n32613 , n32578 , n32582 );
xor ( n32614 , n32613 , n32605 );
buf ( n32615 , n32614 );
buf ( n32616 , n32615 );
xor ( n32617 , n32466 , n32472 );
xor ( n32618 , n32617 , n32526 );
buf ( n32619 , n32618 );
buf ( n32620 , n32619 );
xor ( n32621 , n32589 , n32593 );
xor ( n32622 , n32621 , n32600 );
buf ( n32623 , n32622 );
buf ( n32624 , n32623 );
xor ( n32625 , n32620 , n32624 );
xor ( n32626 , n24441 , n24525 );
and ( n32627 , n32626 , n24555 );
and ( n32628 , n24441 , n24525 );
or ( n32629 , n32627 , n32628 );
buf ( n32630 , n32629 );
buf ( n32631 , n32630 );
and ( n32632 , n32625 , n32631 );
and ( n32633 , n32620 , n32624 );
or ( n32634 , n32632 , n32633 );
buf ( n32635 , n32634 );
buf ( n32636 , n32635 );
nand ( n32637 , n32616 , n32636 );
buf ( n32638 , n32637 );
or ( n32639 , n32612 , n32638 );
buf ( n32640 , n32609 );
buf ( n32641 , n32573 );
nand ( n32642 , n32640 , n32641 );
buf ( n32643 , n32642 );
nand ( n32644 , n32639 , n32643 );
xor ( n32645 , n32058 , n32062 );
xor ( n32646 , n32645 , n32067 );
buf ( n32647 , n32646 );
buf ( n32648 , n32647 );
xor ( n32649 , n32099 , n32231 );
xor ( n32650 , n32649 , n32300 );
buf ( n32651 , n32650 );
buf ( n32652 , n32651 );
xor ( n32653 , n32648 , n32652 );
xor ( n32654 , n32543 , n32547 );
and ( n32655 , n32654 , n32568 );
and ( n32656 , n32543 , n32547 );
or ( n32657 , n32655 , n32656 );
buf ( n32658 , n32657 );
buf ( n32659 , n32658 );
xor ( n32660 , n32653 , n32659 );
buf ( n32661 , n32660 );
not ( n32662 , n32661 );
xor ( n32663 , n32359 , n32536 );
and ( n32664 , n32663 , n32571 );
and ( n32665 , n32359 , n32536 );
or ( n32666 , n32664 , n32665 );
buf ( n32667 , n32666 );
buf ( n32668 , n32667 );
not ( n32669 , n32668 );
buf ( n32670 , n32669 );
nand ( n32671 , n32662 , n32670 );
xor ( n32672 , n32090 , n32094 );
xor ( n32673 , n32672 , n32305 );
buf ( n32674 , n32673 );
not ( n32675 , n32674 );
xor ( n32676 , n32648 , n32652 );
and ( n32677 , n32676 , n32659 );
and ( n32678 , n32648 , n32652 );
or ( n32679 , n32677 , n32678 );
buf ( n32680 , n32679 );
not ( n32681 , n32680 );
nand ( n32682 , n32675 , n32681 );
nand ( n32683 , n32644 , n32671 , n32682 );
nor ( n32684 , n32674 , n32680 );
not ( n32685 , n32684 );
nand ( n32686 , n32661 , n32667 );
not ( n32687 , n32686 );
and ( n32688 , n32685 , n32687 );
buf ( n32689 , n32681 );
not ( n32690 , n32689 );
buf ( n32691 , n32690 );
not ( n32692 , n32675 );
and ( n32693 , n32691 , n32692 );
nor ( n32694 , n32688 , n32693 );
nand ( n32695 , n32683 , n32694 );
not ( n32696 , n32695 );
or ( n32697 , n32355 , n32696 );
buf ( n32698 , n32661 );
not ( n32699 , n32698 );
buf ( n32700 , n32699 );
nand ( n32701 , n32670 , n32700 );
not ( n32702 , n32615 );
not ( n32703 , n32635 );
and ( n32704 , n32702 , n32703 );
nor ( n32705 , n32573 , n32609 );
nor ( n32706 , n32704 , n32705 );
nand ( n32707 , n32681 , n32675 );
nand ( n32708 , n32701 , n32706 , n32707 );
nor ( n32709 , n32351 , n32708 );
not ( n32710 , n24560 );
not ( n32711 , n24580 );
and ( n32712 , n32710 , n32711 );
xor ( n32713 , n32620 , n32624 );
xor ( n32714 , n32713 , n32631 );
buf ( n32715 , n32714 );
buf ( n32716 , n32715 );
xor ( n32717 , n24365 , n24434 );
and ( n32718 , n32717 , n24558 );
and ( n32719 , n24365 , n24434 );
or ( n32720 , n32718 , n32719 );
buf ( n32721 , n32720 );
buf ( n32722 , n32721 );
nor ( n32723 , n32716 , n32722 );
buf ( n32724 , n32723 );
nor ( n32725 , n32712 , n32724 );
not ( n32726 , n32725 );
not ( n32727 , n24634 );
or ( n32728 , n32726 , n32727 );
buf ( n32729 , n32724 );
not ( n32730 , n32729 );
buf ( n32731 , n24587 );
not ( n32732 , n32731 );
and ( n32733 , n32730 , n32732 );
buf ( n32734 , n32715 );
buf ( n32735 , n32721 );
and ( n32736 , n32734 , n32735 );
buf ( n32737 , n32736 );
buf ( n32738 , n32737 );
nor ( n32739 , n32733 , n32738 );
buf ( n32740 , n32739 );
nand ( n32741 , n32728 , n32740 );
nand ( n32742 , n32709 , n32741 );
nand ( n32743 , n32697 , n32742 );
buf ( n32744 , n32743 );
not ( n32745 , n32744 );
buf ( n32746 , n32745 );
buf ( n32747 , n32746 );
not ( n32748 , n32350 );
buf ( n32749 , n31845 );
buf ( n32750 , n32749 );
buf ( n32751 , n32750 );
buf ( n32752 , n32751 );
buf ( n32753 , n32081 );
buf ( n32754 , n32753 );
buf ( n32755 , n32754 );
buf ( n32756 , n32755 );
nor ( n32757 , n32752 , n32756 );
buf ( n32758 , n32757 );
buf ( n32759 , n32086 );
buf ( n32760 , n32759 );
buf ( n32761 , n32760 );
nand ( n32762 , n32761 , n32309 );
or ( n32763 , n32758 , n32762 );
buf ( n32764 , n32751 );
buf ( n32765 , n32755 );
nand ( n32766 , n32764 , n32765 );
buf ( n32767 , n32766 );
nand ( n32768 , n32763 , n32767 );
not ( n32769 , n32768 );
or ( n32770 , n32748 , n32769 );
buf ( n32771 , n32341 );
buf ( n32772 , n32771 );
buf ( n32773 , n32772 );
buf ( n32774 , n32773 );
not ( n32775 , n32774 );
buf ( n32776 , n32775 );
not ( n32777 , n32776 );
buf ( n32778 , n32347 );
buf ( n32779 , n32778 );
buf ( n32780 , n32779 );
buf ( n32781 , n32780 );
not ( n32782 , n32781 );
buf ( n32783 , n32782 );
not ( n32784 , n32783 );
and ( n32785 , n32777 , n32784 );
buf ( n32786 , n32330 );
buf ( n32787 , n32786 );
buf ( n32788 , n32787 );
buf ( n32789 , n32788 );
buf ( n32790 , n32336 );
buf ( n32791 , n32790 );
nand ( n32792 , n32789 , n32791 );
buf ( n32793 , n32792 );
buf ( n32794 , n32793 );
not ( n32795 , n32794 );
buf ( n32796 , n32795 );
buf ( n32797 , n32776 );
buf ( n32798 , n32783 );
nand ( n32799 , n32797 , n32798 );
buf ( n32800 , n32799 );
and ( n32801 , n32796 , n32800 );
nor ( n32802 , n32785 , n32801 );
nand ( n32803 , n32770 , n32802 );
buf ( n32804 , n32803 );
not ( n32805 , n32804 );
buf ( n32806 , n32805 );
buf ( n32807 , n32806 );
nand ( n32808 , n32747 , n32807 );
buf ( n32809 , n32808 );
not ( n32810 , n32809 );
or ( n32811 , n31316 , n32810 );
buf ( n32812 , n31214 );
buf ( n32813 , n31306 );
nand ( n32814 , n32812 , n32813 );
buf ( n32815 , n32814 );
buf ( n32816 , n32815 );
not ( n32817 , n32816 );
buf ( n32818 , n31094 );
buf ( n32819 , n30910 );
nor ( n32820 , n32818 , n32819 );
buf ( n32821 , n32820 );
buf ( n32822 , n31200 );
buf ( n32823 , n31203 );
nand ( n32824 , n32822 , n32823 );
buf ( n32825 , n32824 );
or ( n32826 , n32821 , n32825 );
buf ( n32827 , n31094 );
buf ( n32828 , n30910 );
nand ( n32829 , n32827 , n32828 );
buf ( n32830 , n32829 );
nand ( n32831 , n32826 , n32830 );
buf ( n32832 , n32831 );
not ( n32833 , n32832 );
or ( n32834 , n32817 , n32833 );
buf ( n32835 , n31306 );
not ( n32836 , n32835 );
buf ( n32837 , n31211 );
nand ( n32838 , n32836 , n32837 );
buf ( n32839 , n32838 );
buf ( n32840 , n32839 );
nand ( n32841 , n32834 , n32840 );
buf ( n32842 , n32841 );
buf ( n32843 , n32842 );
not ( n32844 , n32843 );
buf ( n32845 , n32844 );
nand ( n32846 , n32811 , n32845 );
xor ( n32847 , n31221 , n31294 );
and ( n32848 , n32847 , n31301 );
and ( n32849 , n31221 , n31294 );
or ( n32850 , n32848 , n32849 );
buf ( n32851 , n32850 );
buf ( n32852 , n32851 );
xor ( n32853 , n31258 , n31270 );
and ( n32854 , n32853 , n31288 );
and ( n32855 , n31258 , n31270 );
or ( n32856 , n32854 , n32855 );
buf ( n32857 , n32856 );
buf ( n32858 , n32857 );
buf ( n32859 , n18340 );
not ( n32860 , n32859 );
buf ( n32861 , n576 );
not ( n32862 , n32861 );
buf ( n32863 , n30565 );
not ( n32864 , n32863 );
or ( n32865 , n32862 , n32864 );
buf ( n32866 , n30562 );
buf ( n32867 , n7809 );
nand ( n32868 , n32866 , n32867 );
buf ( n32869 , n32868 );
buf ( n32870 , n32869 );
nand ( n32871 , n32865 , n32870 );
buf ( n32872 , n32871 );
buf ( n32873 , n32872 );
not ( n32874 , n32873 );
or ( n32875 , n32860 , n32874 );
buf ( n32876 , n31277 );
buf ( n32877 , n30529 );
nand ( n32878 , n32876 , n32877 );
buf ( n32879 , n32878 );
buf ( n32880 , n32879 );
nand ( n32881 , n32875 , n32880 );
buf ( n32882 , n32881 );
buf ( n32883 , n32882 );
buf ( n32884 , n18264 );
not ( n32885 , n32884 );
buf ( n32886 , n31239 );
not ( n32887 , n32886 );
or ( n32888 , n32885 , n32887 );
buf ( n32889 , n578 );
not ( n32890 , n32889 );
buf ( n32891 , n18170 );
not ( n32892 , n32891 );
or ( n32893 , n32890 , n32892 );
buf ( n32894 , n18167 );
buf ( n32895 , n18233 );
nand ( n32896 , n32894 , n32895 );
buf ( n32897 , n32896 );
buf ( n32898 , n32897 );
nand ( n32899 , n32893 , n32898 );
buf ( n32900 , n32899 );
buf ( n32901 , n32900 );
buf ( n32902 , n18219 );
nand ( n32903 , n32901 , n32902 );
buf ( n32904 , n32903 );
buf ( n32905 , n32904 );
nand ( n32906 , n32888 , n32905 );
buf ( n32907 , n32906 );
buf ( n32908 , n32907 );
xor ( n32909 , n32883 , n32908 );
buf ( n32910 , n30497 );
buf ( n32911 , n576 );
nand ( n32912 , n32910 , n32911 );
buf ( n32913 , n32912 );
buf ( n32914 , n32913 );
xor ( n32915 , n32909 , n32914 );
buf ( n32916 , n32915 );
buf ( n32917 , n32916 );
xor ( n32918 , n32858 , n32917 );
xor ( n32919 , n31247 , n31251 );
and ( n32920 , n32919 , n31291 );
and ( n32921 , n31247 , n31251 );
or ( n32922 , n32920 , n32921 );
buf ( n32923 , n32922 );
buf ( n32924 , n32923 );
xor ( n32925 , n32918 , n32924 );
buf ( n32926 , n32925 );
buf ( n32927 , n32926 );
nor ( n32928 , n32852 , n32927 );
buf ( n32929 , n32928 );
buf ( n32930 , n32929 );
not ( n32931 , n32930 );
buf ( n32932 , n32931 );
not ( n32933 , n32932 );
buf ( n32934 , n32851 );
buf ( n32935 , n32926 );
and ( n32936 , n32934 , n32935 );
buf ( n32937 , n32936 );
nor ( n32938 , n32933 , n32937 );
and ( n32939 , n32846 , n32938 );
not ( n32940 , n32846 );
not ( n32941 , n32938 );
and ( n32942 , n32940 , n32941 );
nor ( n32943 , n32939 , n32942 );
not ( n32944 , n32943 );
not ( n32945 , n31205 );
nand ( n32946 , n32746 , n32806 );
not ( n32947 , n32946 );
or ( n32948 , n32945 , n32947 );
not ( n32949 , n32831 );
nand ( n32950 , n32948 , n32949 );
buf ( n32951 , n32839 );
nand ( n32952 , n32951 , n31309 );
not ( n32953 , n32952 );
and ( n32954 , n32950 , n32953 );
not ( n32955 , n32950 );
and ( n32956 , n32955 , n32952 );
nor ( n32957 , n32954 , n32956 );
not ( n32958 , n32957 );
or ( n32959 , n32944 , n32958 );
not ( n32960 , n32957 );
not ( n32961 , n32943 );
nand ( n32962 , n32960 , n32961 );
nand ( n32963 , n32959 , n32962 );
buf ( n32964 , n32963 );
buf ( n32965 , n32964 );
buf ( n32966 , n32965 );
buf ( n32967 , n32966 );
not ( n32968 , n32967 );
buf ( n32969 , n32968 );
buf ( n32970 , n32969 );
buf ( n32971 , n32970 );
buf ( n32972 , n32971 );
buf ( n32973 , n32972 );
not ( n32974 , n32973 );
buf ( n32975 , n32913 );
not ( n32976 , n32975 );
buf ( n32977 , n32976 );
buf ( n32978 , n32977 );
buf ( n32979 , n18219 );
not ( n32980 , n32979 );
buf ( n32981 , n32980 );
buf ( n32982 , n32981 );
not ( n32983 , n32982 );
buf ( n32984 , n18263 );
not ( n32985 , n32984 );
or ( n32986 , n32983 , n32985 );
buf ( n32987 , n32900 );
nand ( n32988 , n32986 , n32987 );
buf ( n32989 , n32988 );
buf ( n32990 , n32989 );
and ( n32991 , n31274 , n31275 );
buf ( n32992 , n32991 );
buf ( n32993 , n32992 );
xor ( n32994 , n32990 , n32993 );
buf ( n32995 , n18340 );
not ( n32996 , n32995 );
buf ( n32997 , n576 );
buf ( n32998 , n30597 );
xor ( n32999 , n32997 , n32998 );
buf ( n33000 , n32999 );
buf ( n33001 , n33000 );
not ( n33002 , n33001 );
or ( n33003 , n32996 , n33002 );
buf ( n33004 , n32872 );
buf ( n33005 , n30529 );
nand ( n33006 , n33004 , n33005 );
buf ( n33007 , n33006 );
buf ( n33008 , n33007 );
nand ( n33009 , n33003 , n33008 );
buf ( n33010 , n33009 );
buf ( n33011 , n33010 );
xor ( n33012 , n32994 , n33011 );
buf ( n33013 , n33012 );
buf ( n33014 , n33013 );
xor ( n33015 , n32978 , n33014 );
xor ( n33016 , n32883 , n32908 );
and ( n33017 , n33016 , n32914 );
and ( n33018 , n32883 , n32908 );
or ( n33019 , n33017 , n33018 );
buf ( n33020 , n33019 );
buf ( n33021 , n33020 );
xor ( n33022 , n33015 , n33021 );
buf ( n33023 , n33022 );
xor ( n33024 , n32858 , n32917 );
and ( n33025 , n33024 , n32924 );
and ( n33026 , n32858 , n32917 );
or ( n33027 , n33025 , n33026 );
buf ( n33028 , n33027 );
or ( n33029 , n33023 , n33028 );
buf ( n33030 , n33028 );
buf ( n33031 , n33023 );
nand ( n33032 , n33030 , n33031 );
buf ( n33033 , n33032 );
nand ( n33034 , n33029 , n33033 );
buf ( n33035 , n33034 );
not ( n33036 , n33035 );
buf ( n33037 , n33036 );
not ( n33038 , n33037 );
buf ( n33039 , n32743 );
buf ( n33040 , n32803 );
or ( n33041 , n33039 , n33040 );
buf ( n33042 , n31312 );
buf ( n33043 , n32929 );
nor ( n33044 , n33042 , n33043 );
buf ( n33045 , n33044 );
buf ( n33046 , n33045 );
buf ( n33047 , n33046 );
buf ( n33048 , n33047 );
buf ( n33049 , n33048 );
nand ( n33050 , n33041 , n33049 );
buf ( n33051 , n33050 );
buf ( n33052 , n33051 );
buf ( n33053 , n32842 );
buf ( n33054 , n32937 );
or ( n33055 , n33053 , n33054 );
buf ( n33056 , n32932 );
nand ( n33057 , n33055 , n33056 );
buf ( n33058 , n33057 );
buf ( n33059 , n33058 );
buf ( n33060 , n33059 );
buf ( n33061 , n33060 );
buf ( n33062 , n33061 );
nand ( n33063 , n33052 , n33062 );
buf ( n33064 , n33063 );
buf ( n33065 , n33064 );
not ( n33066 , n33065 );
buf ( n33067 , n33066 );
not ( n33068 , n33067 );
or ( n33069 , n33038 , n33068 );
buf ( n33070 , n33064 );
buf ( n33071 , n33034 );
nand ( n33072 , n33070 , n33071 );
buf ( n33073 , n33072 );
nand ( n33074 , n33069 , n33073 );
not ( n33075 , n33074 );
not ( n33076 , n33075 );
buf ( n33077 , n33076 );
buf ( n33078 , n33077 );
not ( n33079 , n33078 );
buf ( n33080 , n33079 );
buf ( n33081 , n33080 );
not ( n33082 , n33081 );
buf ( n33083 , n33082 );
buf ( n33084 , n33083 );
not ( n33085 , n33084 );
buf ( n33086 , n5430 );
not ( n33087 , n33086 );
buf ( n33088 , n600 );
not ( n33089 , n33088 );
buf ( n33090 , n18175 );
not ( n33091 , n33090 );
buf ( n33092 , n33091 );
buf ( n33093 , n33092 );
not ( n33094 , n33093 );
or ( n33095 , n33089 , n33094 );
buf ( n33096 , n18175 );
buf ( n33097 , n5383 );
nand ( n33098 , n33096 , n33097 );
buf ( n33099 , n33098 );
buf ( n33100 , n33099 );
nand ( n33101 , n33095 , n33100 );
buf ( n33102 , n33101 );
buf ( n33103 , n33102 );
not ( n33104 , n33103 );
or ( n33105 , n33087 , n33104 );
buf ( n33106 , n600 );
not ( n33107 , n33106 );
buf ( n33108 , n18177 );
buf ( n33109 , n33108 );
buf ( n33110 , n33109 );
buf ( n33111 , n33110 );
not ( n33112 , n33111 );
buf ( n33113 , n33112 );
buf ( n33114 , n33113 );
not ( n33115 , n33114 );
or ( n33116 , n33107 , n33115 );
buf ( n33117 , n33110 );
buf ( n33118 , n5383 );
nand ( n33119 , n33117 , n33118 );
buf ( n33120 , n33119 );
buf ( n33121 , n33120 );
nand ( n33122 , n33116 , n33121 );
buf ( n33123 , n33122 );
buf ( n33124 , n33123 );
buf ( n33125 , n10945 );
nand ( n33126 , n33124 , n33125 );
buf ( n33127 , n33126 );
buf ( n33128 , n33127 );
nand ( n33129 , n33105 , n33128 );
buf ( n33130 , n33129 );
buf ( n33131 , n33130 );
buf ( n33132 , n26278 );
not ( n33133 , n33132 );
buf ( n33134 , n596 );
not ( n33135 , n33134 );
buf ( n33136 , n28907 );
not ( n33137 , n33136 );
or ( n33138 , n33135 , n33137 );
buf ( n33139 , n28247 );
buf ( n33140 , n2371 );
nand ( n33141 , n33139 , n33140 );
buf ( n33142 , n33141 );
buf ( n33143 , n33142 );
nand ( n33144 , n33138 , n33143 );
buf ( n33145 , n33144 );
buf ( n33146 , n33145 );
not ( n33147 , n33146 );
or ( n33148 , n33133 , n33147 );
buf ( n33149 , n596 );
not ( n33150 , n33149 );
buf ( n33151 , n28664 );
not ( n33152 , n33151 );
buf ( n33153 , n33152 );
buf ( n33154 , n33153 );
not ( n33155 , n33154 );
or ( n33156 , n33150 , n33155 );
buf ( n33157 , n28664 );
buf ( n33158 , n2371 );
nand ( n33159 , n33157 , n33158 );
buf ( n33160 , n33159 );
buf ( n33161 , n33160 );
nand ( n33162 , n33156 , n33161 );
buf ( n33163 , n33162 );
buf ( n33164 , n33163 );
buf ( n33165 , n825 );
nand ( n33166 , n33164 , n33165 );
buf ( n33167 , n33166 );
buf ( n33168 , n33167 );
nand ( n33169 , n33148 , n33168 );
buf ( n33170 , n33169 );
buf ( n33171 , n33170 );
buf ( n33172 , n28180 );
buf ( n33173 , n592 );
nand ( n33174 , n33172 , n33173 );
buf ( n33175 , n33174 );
buf ( n33176 , n33175 );
not ( n33177 , n33176 );
buf ( n33178 , n33177 );
buf ( n33179 , n33178 );
xor ( n33180 , n33171 , n33179 );
buf ( n33181 , n602 );
not ( n33182 , n33181 );
buf ( n33183 , n18177 );
not ( n33184 , n33183 );
buf ( n33185 , n33184 );
buf ( n33186 , n33185 );
not ( n33187 , n33186 );
or ( n33188 , n33182 , n33187 );
buf ( n33189 , n18177 );
buf ( n33190 , n2912 );
nand ( n33191 , n33189 , n33190 );
buf ( n33192 , n33191 );
buf ( n33193 , n33192 );
nand ( n33194 , n33188 , n33193 );
buf ( n33195 , n33194 );
buf ( n33196 , n33195 );
buf ( n33197 , n7619 );
not ( n33198 , n33197 );
buf ( n33199 , n5652 );
nand ( n33200 , n33198 , n33199 );
buf ( n33201 , n33200 );
buf ( n33202 , n33201 );
nand ( n33203 , n33196 , n33202 );
buf ( n33204 , n33203 );
buf ( n33205 , n33204 );
and ( n33206 , n33180 , n33205 );
and ( n33207 , n33171 , n33179 );
or ( n33208 , n33206 , n33207 );
buf ( n33209 , n33208 );
buf ( n33210 , n33209 );
xor ( n33211 , n33131 , n33210 );
not ( n33212 , n2452 );
buf ( n33213 , n592 );
not ( n33214 , n33213 );
buf ( n33215 , n26088 );
not ( n33216 , n33215 );
or ( n33217 , n33214 , n33216 );
buf ( n33218 , n26088 );
not ( n33219 , n33218 );
buf ( n33220 , n33219 );
buf ( n33221 , n33220 );
buf ( n33222 , n2416 );
nand ( n33223 , n33221 , n33222 );
buf ( n33224 , n33223 );
buf ( n33225 , n33224 );
nand ( n33226 , n33217 , n33225 );
buf ( n33227 , n33226 );
not ( n33228 , n33227 );
or ( n33229 , n33212 , n33228 );
buf ( n33230 , n592 );
not ( n33231 , n33230 );
buf ( n33232 , n28611 );
not ( n33233 , n33232 );
or ( n33234 , n33231 , n33233 );
buf ( n33235 , n28611 );
not ( n33236 , n33235 );
buf ( n33237 , n33236 );
buf ( n33238 , n33237 );
buf ( n33239 , n2416 );
nand ( n33240 , n33238 , n33239 );
buf ( n33241 , n33240 );
buf ( n33242 , n33241 );
nand ( n33243 , n33234 , n33242 );
buf ( n33244 , n33243 );
nand ( n33245 , n33244 , n28544 );
nand ( n33246 , n33229 , n33245 );
buf ( n33247 , n33246 );
buf ( n33248 , n2592 );
not ( n33249 , n33248 );
buf ( n33250 , n594 );
not ( n33251 , n33250 );
buf ( n33252 , n18191 );
not ( n33253 , n33252 );
buf ( n33254 , n33253 );
buf ( n33255 , n33254 );
not ( n33256 , n33255 );
or ( n33257 , n33251 , n33256 );
buf ( n33258 , n18191 );
buf ( n33259 , n2481 );
nand ( n33260 , n33258 , n33259 );
buf ( n33261 , n33260 );
buf ( n33262 , n33261 );
nand ( n33263 , n33257 , n33262 );
buf ( n33264 , n33263 );
buf ( n33265 , n33264 );
not ( n33266 , n33265 );
or ( n33267 , n33249 , n33266 );
not ( n33268 , n594 );
not ( n33269 , n28907 );
or ( n33270 , n33268 , n33269 );
buf ( n33271 , n28247 );
buf ( n33272 , n2481 );
nand ( n33273 , n33271 , n33272 );
buf ( n33274 , n33273 );
nand ( n33275 , n33270 , n33274 );
nand ( n33276 , n33275 , n2541 );
buf ( n33277 , n33276 );
nand ( n33278 , n33267 , n33277 );
buf ( n33279 , n33278 );
buf ( n33280 , n33279 );
xor ( n33281 , n33247 , n33280 );
buf ( n33282 , n28626 );
buf ( n33283 , n592 );
nand ( n33284 , n33282 , n33283 );
buf ( n33285 , n33284 );
buf ( n33286 , n33285 );
xor ( n33287 , n33281 , n33286 );
buf ( n33288 , n33287 );
buf ( n33289 , n33288 );
xor ( n33290 , n33211 , n33289 );
buf ( n33291 , n33290 );
buf ( n33292 , n33291 );
buf ( n33293 , n5550 );
not ( n33294 , n33293 );
buf ( n33295 , n598 );
not ( n33296 , n33295 );
buf ( n33297 , n30026 );
not ( n33298 , n33297 );
buf ( n33299 , n33298 );
buf ( n33300 , n33299 );
not ( n33301 , n33300 );
or ( n33302 , n33296 , n33301 );
buf ( n33303 , n30032 );
not ( n33304 , n33303 );
buf ( n33305 , n33304 );
buf ( n33306 , n33305 );
buf ( n33307 , n818 );
nand ( n33308 , n33306 , n33307 );
buf ( n33309 , n33308 );
buf ( n33310 , n33309 );
nand ( n33311 , n33302 , n33310 );
buf ( n33312 , n33311 );
buf ( n33313 , n33312 );
not ( n33314 , n33313 );
or ( n33315 , n33294 , n33314 );
buf ( n33316 , n598 );
not ( n33317 , n33316 );
not ( n33318 , n29202 );
buf ( n33319 , n33318 );
not ( n33320 , n33319 );
or ( n33321 , n33317 , n33320 );
buf ( n33322 , n29202 );
buf ( n33323 , n818 );
nand ( n33324 , n33322 , n33323 );
buf ( n33325 , n33324 );
buf ( n33326 , n33325 );
nand ( n33327 , n33321 , n33326 );
buf ( n33328 , n33327 );
buf ( n33329 , n33328 );
buf ( n33330 , n5631 );
nand ( n33331 , n33329 , n33330 );
buf ( n33332 , n33331 );
buf ( n33333 , n33332 );
nand ( n33334 , n33315 , n33333 );
buf ( n33335 , n33334 );
buf ( n33336 , n33335 );
not ( n33337 , n825 );
nand ( n33338 , n28947 , n2371 );
nand ( n33339 , n596 , n28941 );
nand ( n33340 , n33338 , n33339 );
not ( n33341 , n33340 );
or ( n33342 , n33337 , n33341 );
buf ( n33343 , n33163 );
buf ( n33344 , n26278 );
nand ( n33345 , n33343 , n33344 );
buf ( n33346 , n33345 );
nand ( n33347 , n33342 , n33346 );
buf ( n33348 , n33347 );
xor ( n33349 , n33336 , n33348 );
buf ( n33350 , n26789 );
buf ( n33351 , n592 );
and ( n33352 , n33350 , n33351 );
buf ( n33353 , n33352 );
buf ( n33354 , n33353 );
buf ( n33355 , n2452 );
not ( n33356 , n33355 );
buf ( n33357 , n33244 );
not ( n33358 , n33357 );
or ( n33359 , n33356 , n33358 );
buf ( n33360 , n592 );
not ( n33361 , n33360 );
buf ( n33362 , n26813 );
not ( n33363 , n33362 );
or ( n33364 , n33361 , n33363 );
buf ( n33365 , n26810 );
buf ( n33366 , n2416 );
nand ( n33367 , n33365 , n33366 );
buf ( n33368 , n33367 );
buf ( n33369 , n33368 );
nand ( n33370 , n33364 , n33369 );
buf ( n33371 , n33370 );
buf ( n33372 , n33371 );
buf ( n33373 , n28544 );
nand ( n33374 , n33372 , n33373 );
buf ( n33375 , n33374 );
buf ( n33376 , n33375 );
nand ( n33377 , n33359 , n33376 );
buf ( n33378 , n33377 );
buf ( n33379 , n33378 );
xor ( n33380 , n33354 , n33379 );
buf ( n33381 , n2541 );
not ( n33382 , n33381 );
buf ( n33383 , n33264 );
not ( n33384 , n33383 );
or ( n33385 , n33382 , n33384 );
buf ( n33386 , n594 );
not ( n33387 , n33386 );
buf ( n33388 , n26094 );
not ( n33389 , n33388 );
buf ( n33390 , n33389 );
buf ( n33391 , n33390 );
not ( n33392 , n33391 );
or ( n33393 , n33387 , n33392 );
buf ( n33394 , n26094 );
buf ( n33395 , n2481 );
nand ( n33396 , n33394 , n33395 );
buf ( n33397 , n33396 );
buf ( n33398 , n33397 );
nand ( n33399 , n33393 , n33398 );
buf ( n33400 , n33399 );
buf ( n33401 , n33400 );
buf ( n33402 , n2592 );
nand ( n33403 , n33401 , n33402 );
buf ( n33404 , n33403 );
buf ( n33405 , n33404 );
nand ( n33406 , n33385 , n33405 );
buf ( n33407 , n33406 );
buf ( n33408 , n33407 );
and ( n33409 , n33380 , n33408 );
and ( n33410 , n33354 , n33379 );
or ( n33411 , n33409 , n33410 );
buf ( n33412 , n33411 );
buf ( n33413 , n33412 );
xor ( n33414 , n33349 , n33413 );
buf ( n33415 , n33414 );
buf ( n33416 , n33415 );
buf ( n33417 , n5550 );
not ( n33418 , n33417 );
buf ( n33419 , n33328 );
not ( n33420 , n33419 );
or ( n33421 , n33418 , n33420 );
buf ( n33422 , n598 );
not ( n33423 , n33422 );
buf ( n33424 , n28941 );
not ( n33425 , n33424 );
or ( n33426 , n33423 , n33425 );
buf ( n33427 , n28947 );
buf ( n33428 , n818 );
nand ( n33429 , n33427 , n33428 );
buf ( n33430 , n33429 );
buf ( n33431 , n33430 );
nand ( n33432 , n33426 , n33431 );
buf ( n33433 , n33432 );
buf ( n33434 , n33433 );
buf ( n33435 , n5631 );
nand ( n33436 , n33434 , n33435 );
buf ( n33437 , n33436 );
buf ( n33438 , n33437 );
nand ( n33439 , n33421 , n33438 );
buf ( n33440 , n33439 );
buf ( n33441 , n33440 );
buf ( n33442 , n10945 );
not ( n33443 , n33442 );
buf ( n33444 , n33102 );
not ( n33445 , n33444 );
or ( n33446 , n33443 , n33445 );
buf ( n33447 , n33299 );
not ( n33448 , n33447 );
buf ( n33449 , n33448 );
buf ( n33450 , n33449 );
buf ( n33451 , n11561 );
and ( n33452 , n33450 , n33451 );
buf ( n33453 , n33305 );
not ( n33454 , n33453 );
buf ( n33455 , n33454 );
buf ( n33456 , n33455 );
buf ( n33457 , n11571 );
and ( n33458 , n33456 , n33457 );
nor ( n33459 , n33452 , n33458 );
buf ( n33460 , n33459 );
buf ( n33461 , n33460 );
nand ( n33462 , n33446 , n33461 );
buf ( n33463 , n33462 );
buf ( n33464 , n33463 );
xor ( n33465 , n33441 , n33464 );
not ( n33466 , n2452 );
not ( n33467 , n33371 );
or ( n33468 , n33466 , n33467 );
buf ( n33469 , n592 );
not ( n33470 , n33469 );
buf ( n33471 , n26786 );
not ( n33472 , n33471 );
or ( n33473 , n33470 , n33472 );
buf ( n33474 , n26782 );
buf ( n33475 , n2416 );
nand ( n33476 , n33474 , n33475 );
buf ( n33477 , n33476 );
buf ( n33478 , n33477 );
nand ( n33479 , n33473 , n33478 );
buf ( n33480 , n33479 );
buf ( n33481 , n33480 );
buf ( n33482 , n28544 );
nand ( n33483 , n33481 , n33482 );
buf ( n33484 , n33483 );
nand ( n33485 , n33468 , n33484 );
buf ( n33486 , n33485 );
buf ( n33487 , n2592 );
not ( n33488 , n33487 );
buf ( n33489 , n594 );
not ( n33490 , n33489 );
buf ( n33491 , n28611 );
not ( n33492 , n33491 );
or ( n33493 , n33490 , n33492 );
buf ( n33494 , n26053 );
buf ( n33495 , n2481 );
nand ( n33496 , n33494 , n33495 );
buf ( n33497 , n33496 );
buf ( n33498 , n33497 );
nand ( n33499 , n33493 , n33498 );
buf ( n33500 , n33499 );
buf ( n33501 , n33500 );
not ( n33502 , n33501 );
or ( n33503 , n33488 , n33502 );
buf ( n33504 , n33400 );
buf ( n33505 , n2541 );
nand ( n33506 , n33504 , n33505 );
buf ( n33507 , n33506 );
buf ( n33508 , n33507 );
nand ( n33509 , n33503 , n33508 );
buf ( n33510 , n33509 );
buf ( n33511 , n33510 );
xor ( n33512 , n33486 , n33511 );
buf ( n33513 , n26278 );
not ( n33514 , n33513 );
buf ( n33515 , n596 );
not ( n33516 , n33515 );
buf ( n33517 , n33254 );
not ( n33518 , n33517 );
or ( n33519 , n33516 , n33518 );
buf ( n33520 , n18191 );
buf ( n33521 , n2371 );
nand ( n33522 , n33520 , n33521 );
buf ( n33523 , n33522 );
buf ( n33524 , n33523 );
nand ( n33525 , n33519 , n33524 );
buf ( n33526 , n33525 );
buf ( n33527 , n33526 );
not ( n33528 , n33527 );
or ( n33529 , n33514 , n33528 );
buf ( n33530 , n33145 );
buf ( n33531 , n825 );
nand ( n33532 , n33530 , n33531 );
buf ( n33533 , n33532 );
buf ( n33534 , n33533 );
nand ( n33535 , n33529 , n33534 );
buf ( n33536 , n33535 );
buf ( n33537 , n33536 );
and ( n33538 , n33512 , n33537 );
and ( n33539 , n33486 , n33511 );
or ( n33540 , n33538 , n33539 );
buf ( n33541 , n33540 );
buf ( n33542 , n33541 );
and ( n33543 , n33465 , n33542 );
and ( n33544 , n33441 , n33464 );
or ( n33545 , n33543 , n33544 );
buf ( n33546 , n33545 );
buf ( n33547 , n33546 );
xor ( n33548 , n33416 , n33547 );
xor ( n33549 , n33354 , n33379 );
xor ( n33550 , n33549 , n33408 );
buf ( n33551 , n33550 );
buf ( n33552 , n33551 );
xor ( n33553 , n33171 , n33179 );
xor ( n33554 , n33553 , n33205 );
buf ( n33555 , n33554 );
buf ( n33556 , n33555 );
xor ( n33557 , n33552 , n33556 );
buf ( n33558 , n33175 );
buf ( n33559 , n600 );
not ( n33560 , n33559 );
buf ( n33561 , n29203 );
not ( n33562 , n33561 );
or ( n33563 , n33560 , n33562 );
buf ( n33564 , n600 );
not ( n33565 , n33564 );
buf ( n33566 , n29202 );
nand ( n33567 , n33565 , n33566 );
buf ( n33568 , n33567 );
buf ( n33569 , n33568 );
nand ( n33570 , n33563 , n33569 );
buf ( n33571 , n33570 );
buf ( n33572 , n33571 );
buf ( n33573 , n5430 );
nand ( n33574 , n33572 , n33573 );
buf ( n33575 , n33574 );
buf ( n33576 , n33575 );
buf ( n33577 , n33299 );
buf ( n33578 , n26763 );
nand ( n33579 , n33577 , n33578 );
buf ( n33580 , n33579 );
buf ( n33581 , n33580 );
buf ( n33582 , n33449 );
buf ( n33583 , n26757 );
nand ( n33584 , n33582 , n33583 );
buf ( n33585 , n33584 );
buf ( n33586 , n33585 );
nand ( n33587 , n33576 , n33581 , n33586 );
buf ( n33588 , n33587 );
buf ( n33589 , n33588 );
xor ( n33590 , n33558 , n33589 );
buf ( n33591 , n5550 );
not ( n33592 , n33591 );
buf ( n33593 , n33433 );
not ( n33594 , n33593 );
or ( n33595 , n33592 , n33594 );
buf ( n33596 , n598 );
not ( n33597 , n33596 );
buf ( n33598 , n33153 );
not ( n33599 , n33598 );
or ( n33600 , n33597 , n33599 );
buf ( n33601 , n28664 );
buf ( n33602 , n818 );
nand ( n33603 , n33601 , n33602 );
buf ( n33604 , n33603 );
buf ( n33605 , n33604 );
nand ( n33606 , n33600 , n33605 );
buf ( n33607 , n33606 );
buf ( n33608 , n33607 );
buf ( n33609 , n5631 );
nand ( n33610 , n33608 , n33609 );
buf ( n33611 , n33610 );
buf ( n33612 , n33611 );
nand ( n33613 , n33595 , n33612 );
buf ( n33614 , n33613 );
buf ( n33615 , n33614 );
and ( n33616 , n33590 , n33615 );
and ( n33617 , n33558 , n33589 );
or ( n33618 , n33616 , n33617 );
buf ( n33619 , n33618 );
buf ( n33620 , n33619 );
and ( n33621 , n33557 , n33620 );
and ( n33622 , n33552 , n33556 );
or ( n33623 , n33621 , n33622 );
buf ( n33624 , n33623 );
buf ( n33625 , n33624 );
xor ( n33626 , n33548 , n33625 );
buf ( n33627 , n33626 );
buf ( n33628 , n33627 );
xor ( n33629 , n33292 , n33628 );
xor ( n33630 , n33441 , n33464 );
xor ( n33631 , n33630 , n33542 );
buf ( n33632 , n33631 );
buf ( n33633 , n33632 );
not ( n33634 , n33195 );
not ( n33635 , n5655 );
or ( n33636 , n33634 , n33635 );
and ( n33637 , n33092 , n11930 );
not ( n33638 , n33092 );
and ( n33639 , n33638 , n11923 );
nor ( n33640 , n33637 , n33639 );
nand ( n33641 , n33636 , n33640 );
buf ( n33642 , n33641 );
buf ( n33643 , n2452 );
not ( n33644 , n33643 );
buf ( n33645 , n33480 );
not ( n33646 , n33645 );
or ( n33647 , n33644 , n33646 );
not ( n33648 , n592 );
not ( n33649 , n26973 );
or ( n33650 , n33648 , n33649 );
buf ( n33651 , n26737 );
buf ( n33652 , n2416 );
nand ( n33653 , n33651 , n33652 );
buf ( n33654 , n33653 );
nand ( n33655 , n33650 , n33654 );
buf ( n33656 , n33655 );
buf ( n33657 , n28544 );
nand ( n33658 , n33656 , n33657 );
buf ( n33659 , n33658 );
buf ( n33660 , n33659 );
nand ( n33661 , n33647 , n33660 );
buf ( n33662 , n33661 );
buf ( n33663 , n33662 );
buf ( n33664 , n592 );
buf ( n33665 , n27312 );
and ( n33666 , n33664 , n33665 );
buf ( n33667 , n33666 );
buf ( n33668 , n33667 );
xor ( n33669 , n33663 , n33668 );
buf ( n33670 , n2541 );
not ( n33671 , n33670 );
buf ( n33672 , n33500 );
not ( n33673 , n33672 );
or ( n33674 , n33671 , n33673 );
buf ( n33675 , n594 );
not ( n33676 , n33675 );
buf ( n33677 , n26813 );
not ( n33678 , n33677 );
or ( n33679 , n33676 , n33678 );
buf ( n33680 , n26810 );
buf ( n33681 , n2481 );
nand ( n33682 , n33680 , n33681 );
buf ( n33683 , n33682 );
buf ( n33684 , n33683 );
nand ( n33685 , n33679 , n33684 );
buf ( n33686 , n33685 );
buf ( n33687 , n33686 );
buf ( n33688 , n2592 );
nand ( n33689 , n33687 , n33688 );
buf ( n33690 , n33689 );
buf ( n33691 , n33690 );
nand ( n33692 , n33674 , n33691 );
buf ( n33693 , n33692 );
buf ( n33694 , n33693 );
and ( n33695 , n33669 , n33694 );
and ( n33696 , n33663 , n33668 );
or ( n33697 , n33695 , n33696 );
buf ( n33698 , n33697 );
buf ( n33699 , n33698 );
xor ( n33700 , n33642 , n33699 );
buf ( n33701 , n825 );
not ( n33702 , n33701 );
buf ( n33703 , n33526 );
not ( n33704 , n33703 );
or ( n33705 , n33702 , n33704 );
buf ( n33706 , n596 );
not ( n33707 , n33706 );
buf ( n33708 , n26088 );
not ( n33709 , n33708 );
or ( n33710 , n33707 , n33709 );
buf ( n33711 , n33220 );
buf ( n33712 , n2371 );
nand ( n33713 , n33711 , n33712 );
buf ( n33714 , n33713 );
buf ( n33715 , n33714 );
nand ( n33716 , n33710 , n33715 );
buf ( n33717 , n33716 );
buf ( n33718 , n33717 );
buf ( n33719 , n26278 );
nand ( n33720 , n33718 , n33719 );
buf ( n33721 , n33720 );
buf ( n33722 , n33721 );
nand ( n33723 , n33705 , n33722 );
buf ( n33724 , n33723 );
buf ( n33725 , n33724 );
not ( n33726 , n2592 );
not ( n33727 , n594 );
not ( n33728 , n26786 );
or ( n33729 , n33727 , n33728 );
buf ( n33730 , n26782 );
buf ( n33731 , n2481 );
nand ( n33732 , n33730 , n33731 );
buf ( n33733 , n33732 );
nand ( n33734 , n33729 , n33733 );
not ( n33735 , n33734 );
or ( n33736 , n33726 , n33735 );
buf ( n33737 , n33686 );
buf ( n33738 , n2541 );
nand ( n33739 , n33737 , n33738 );
buf ( n33740 , n33739 );
nand ( n33741 , n33736 , n33740 );
buf ( n33742 , n33741 );
xor ( n33743 , n33725 , n33742 );
not ( n33744 , n5550 );
not ( n33745 , n33607 );
or ( n33746 , n33744 , n33745 );
buf ( n33747 , n28247 );
buf ( n33748 , n818 );
nand ( n33749 , n33747 , n33748 );
buf ( n33750 , n33749 );
nand ( n33751 , n28907 , n598 );
nand ( n33752 , n33750 , n33751 );
nand ( n33753 , n33752 , n5631 );
nand ( n33754 , n33746 , n33753 );
buf ( n33755 , n33754 );
and ( n33756 , n33743 , n33755 );
and ( n33757 , n33725 , n33742 );
or ( n33758 , n33756 , n33757 );
buf ( n33759 , n33758 );
buf ( n33760 , n33759 );
and ( n33761 , n33700 , n33760 );
and ( n33762 , n33642 , n33699 );
or ( n33763 , n33761 , n33762 );
buf ( n33764 , n33763 );
buf ( n33765 , n33764 );
xor ( n33766 , n33633 , n33765 );
xor ( n33767 , n33486 , n33511 );
xor ( n33768 , n33767 , n33537 );
buf ( n33769 , n33768 );
buf ( n33770 , n33769 );
xor ( n33771 , n33558 , n33589 );
xor ( n33772 , n33771 , n33615 );
buf ( n33773 , n33772 );
buf ( n33774 , n33773 );
xor ( n33775 , n33770 , n33774 );
buf ( n33776 , n5430 );
not ( n33777 , n33776 );
and ( n33778 , n600 , n28941 );
not ( n33779 , n600 );
and ( n33780 , n33779 , n30073 );
or ( n33781 , n33778 , n33780 );
buf ( n33782 , n33781 );
not ( n33783 , n33782 );
or ( n33784 , n33777 , n33783 );
and ( n33785 , n29202 , n26757 );
not ( n33786 , n29202 );
and ( n33787 , n33786 , n26763 );
nor ( n33788 , n33785 , n33787 );
buf ( n33789 , n33788 );
nand ( n33790 , n33784 , n33789 );
buf ( n33791 , n33790 );
buf ( n33792 , n33791 );
xor ( n33793 , n604 , n18177 );
buf ( n33794 , n33793 );
buf ( n33795 , n8581 );
not ( n33796 , n33795 );
buf ( n33797 , n12443 );
nand ( n33798 , n33796 , n33797 );
buf ( n33799 , n33798 );
buf ( n33800 , n33799 );
nand ( n33801 , n33794 , n33800 );
buf ( n33802 , n33801 );
buf ( n33803 , n33802 );
xor ( n33804 , n33792 , n33803 );
xor ( n33805 , n33663 , n33668 );
xor ( n33806 , n33805 , n33694 );
buf ( n33807 , n33806 );
buf ( n33808 , n33807 );
and ( n33809 , n33804 , n33808 );
and ( n33810 , n33792 , n33803 );
or ( n33811 , n33809 , n33810 );
buf ( n33812 , n33811 );
buf ( n33813 , n33812 );
and ( n33814 , n33775 , n33813 );
and ( n33815 , n33770 , n33774 );
or ( n33816 , n33814 , n33815 );
buf ( n33817 , n33816 );
buf ( n33818 , n33817 );
and ( n33819 , n33766 , n33818 );
and ( n33820 , n33633 , n33765 );
or ( n33821 , n33819 , n33820 );
buf ( n33822 , n33821 );
buf ( n33823 , n33822 );
xor ( n33824 , n33629 , n33823 );
buf ( n33825 , n33824 );
not ( n33826 , n33825 );
xor ( n33827 , n33552 , n33556 );
xor ( n33828 , n33827 , n33620 );
buf ( n33829 , n33828 );
buf ( n33830 , n33829 );
xor ( n33831 , n33633 , n33765 );
xor ( n33832 , n33831 , n33818 );
buf ( n33833 , n33832 );
buf ( n33834 , n33833 );
xor ( n33835 , n33830 , n33834 );
xor ( n33836 , n33642 , n33699 );
xor ( n33837 , n33836 , n33760 );
buf ( n33838 , n33837 );
buf ( n33839 , n33838 );
buf ( n33840 , n602 );
not ( n33841 , n33840 );
buf ( n33842 , n33299 );
not ( n33843 , n33842 );
or ( n33844 , n33841 , n33843 );
buf ( n33845 , n30026 );
buf ( n33846 , n2912 );
nand ( n33847 , n33845 , n33846 );
buf ( n33848 , n33847 );
buf ( n33849 , n33848 );
nand ( n33850 , n33844 , n33849 );
buf ( n33851 , n33850 );
buf ( n33852 , n33851 );
buf ( n33853 , n7619 );
nand ( n33854 , n33852 , n33853 );
buf ( n33855 , n33854 );
buf ( n33856 , n33855 );
buf ( n33857 , n18175 );
not ( n33858 , n33857 );
buf ( n33859 , n33858 );
buf ( n33860 , n33859 );
buf ( n33861 , n26682 );
nand ( n33862 , n33860 , n33861 );
buf ( n33863 , n33862 );
buf ( n33864 , n33863 );
buf ( n33865 , n18175 );
not ( n33866 , n33865 );
buf ( n33867 , n33866 );
buf ( n33868 , n33867 );
not ( n33869 , n33868 );
buf ( n33870 , n33869 );
buf ( n33871 , n33870 );
buf ( n33872 , n26693 );
nand ( n33873 , n33871 , n33872 );
buf ( n33874 , n33873 );
buf ( n33875 , n33874 );
nand ( n33876 , n33856 , n33864 , n33875 );
buf ( n33877 , n33876 );
buf ( n33878 , n33877 );
buf ( n33879 , n28544 );
not ( n33880 , n33879 );
xor ( n33881 , n33664 , n33665 );
buf ( n33882 , n33881 );
buf ( n33883 , n33882 );
not ( n33884 , n33883 );
or ( n33885 , n33880 , n33884 );
buf ( n33886 , n33655 );
buf ( n33887 , n2452 );
nand ( n33888 , n33886 , n33887 );
buf ( n33889 , n33888 );
buf ( n33890 , n33889 );
nand ( n33891 , n33885 , n33890 );
buf ( n33892 , n33891 );
buf ( n33893 , n33892 );
buf ( n33894 , n592 );
buf ( n33895 , n28162 );
and ( n33896 , n33894 , n33895 );
buf ( n33897 , n33896 );
buf ( n33898 , n33897 );
xor ( n33899 , n33893 , n33898 );
buf ( n33900 , n26278 );
not ( n33901 , n33900 );
and ( n33902 , n26056 , n596 );
not ( n33903 , n26056 );
and ( n33904 , n33903 , n2371 );
or ( n33905 , n33902 , n33904 );
buf ( n33906 , n33905 );
not ( n33907 , n33906 );
or ( n33908 , n33901 , n33907 );
buf ( n33909 , n33717 );
buf ( n33910 , n825 );
nand ( n33911 , n33909 , n33910 );
buf ( n33912 , n33911 );
buf ( n33913 , n33912 );
nand ( n33914 , n33908 , n33913 );
buf ( n33915 , n33914 );
buf ( n33916 , n33915 );
and ( n33917 , n33899 , n33916 );
and ( n33918 , n33893 , n33898 );
or ( n33919 , n33917 , n33918 );
buf ( n33920 , n33919 );
buf ( n33921 , n33920 );
xor ( n33922 , n33878 , n33921 );
not ( n33923 , n10831 );
nand ( n33924 , n33923 , n592 );
buf ( n33925 , n33924 );
not ( n33926 , n33925 );
buf ( n33927 , n33926 );
buf ( n33928 , n33927 );
buf ( n33929 , n33741 );
not ( n33930 , n33929 );
buf ( n33931 , n33930 );
buf ( n33932 , n33931 );
xor ( n33933 , n33928 , n33932 );
buf ( n33934 , n5550 );
not ( n33935 , n33934 );
buf ( n33936 , n33752 );
not ( n33937 , n33936 );
or ( n33938 , n33935 , n33937 );
buf ( n33939 , n598 );
not ( n33940 , n33939 );
buf ( n33941 , n33254 );
not ( n33942 , n33941 );
or ( n33943 , n33940 , n33942 );
buf ( n33944 , n18191 );
buf ( n33945 , n818 );
nand ( n33946 , n33944 , n33945 );
buf ( n33947 , n33946 );
buf ( n33948 , n33947 );
nand ( n33949 , n33943 , n33948 );
buf ( n33950 , n33949 );
buf ( n33951 , n33950 );
buf ( n33952 , n5631 );
nand ( n33953 , n33951 , n33952 );
buf ( n33954 , n33953 );
buf ( n33955 , n33954 );
nand ( n33956 , n33938 , n33955 );
buf ( n33957 , n33956 );
buf ( n33958 , n33957 );
and ( n33959 , n33933 , n33958 );
and ( n33960 , n33928 , n33932 );
or ( n33961 , n33959 , n33960 );
buf ( n33962 , n33961 );
buf ( n33963 , n33962 );
and ( n33964 , n33922 , n33963 );
and ( n33965 , n33878 , n33921 );
or ( n33966 , n33964 , n33965 );
buf ( n33967 , n33966 );
buf ( n33968 , n33967 );
xor ( n33969 , n33839 , n33968 );
xor ( n33970 , n33725 , n33742 );
xor ( n33971 , n33970 , n33755 );
buf ( n33972 , n33971 );
buf ( n33973 , n33972 );
xor ( n33974 , n33792 , n33803 );
xor ( n33975 , n33974 , n33808 );
buf ( n33976 , n33975 );
buf ( n33977 , n33976 );
xor ( n33978 , n33973 , n33977 );
buf ( n33979 , n5655 );
not ( n33980 , n33979 );
buf ( n33981 , n33851 );
not ( n33982 , n33981 );
or ( n33983 , n33980 , n33982 );
buf ( n33984 , n602 );
not ( n33985 , n33984 );
buf ( n33986 , n33318 );
not ( n33987 , n33986 );
or ( n33988 , n33985 , n33987 );
buf ( n33989 , n29202 );
buf ( n33990 , n2912 );
nand ( n33991 , n33989 , n33990 );
buf ( n33992 , n33991 );
buf ( n33993 , n33992 );
nand ( n33994 , n33988 , n33993 );
buf ( n33995 , n33994 );
buf ( n33996 , n33995 );
buf ( n33997 , n7619 );
nand ( n33998 , n33996 , n33997 );
buf ( n33999 , n33998 );
buf ( n34000 , n33999 );
nand ( n34001 , n33983 , n34000 );
buf ( n34002 , n34001 );
buf ( n34003 , n34002 );
buf ( n34004 , n2915 );
not ( n34005 , n34004 );
buf ( n34006 , n33781 );
not ( n34007 , n34006 );
or ( n34008 , n34005 , n34007 );
buf ( n34009 , n600 );
not ( n34010 , n34009 );
buf ( n34011 , n28667 );
not ( n34012 , n34011 );
or ( n34013 , n34010 , n34012 );
buf ( n34014 , n28664 );
buf ( n34015 , n5383 );
nand ( n34016 , n34014 , n34015 );
buf ( n34017 , n34016 );
buf ( n34018 , n34017 );
nand ( n34019 , n34013 , n34018 );
buf ( n34020 , n34019 );
buf ( n34021 , n34020 );
buf ( n34022 , n5430 );
nand ( n34023 , n34021 , n34022 );
buf ( n34024 , n34023 );
buf ( n34025 , n34024 );
nand ( n34026 , n34008 , n34025 );
buf ( n34027 , n34026 );
buf ( n34028 , n34027 );
xor ( n34029 , n34003 , n34028 );
xor ( n34030 , n33893 , n33898 );
xor ( n34031 , n34030 , n33916 );
buf ( n34032 , n34031 );
buf ( n34033 , n34032 );
and ( n34034 , n34029 , n34033 );
and ( n34035 , n34003 , n34028 );
or ( n34036 , n34034 , n34035 );
buf ( n34037 , n34036 );
buf ( n34038 , n34037 );
and ( n34039 , n33978 , n34038 );
and ( n34040 , n33973 , n33977 );
or ( n34041 , n34039 , n34040 );
buf ( n34042 , n34041 );
buf ( n34043 , n34042 );
and ( n34044 , n33969 , n34043 );
and ( n34045 , n33839 , n33968 );
or ( n34046 , n34044 , n34045 );
buf ( n34047 , n34046 );
buf ( n34048 , n34047 );
and ( n34049 , n33835 , n34048 );
and ( n34050 , n33830 , n33834 );
or ( n34051 , n34049 , n34050 );
buf ( n34052 , n34051 );
not ( n34053 , n34052 );
and ( n34054 , n33826 , n34053 );
xor ( n34055 , n33770 , n33774 );
xor ( n34056 , n34055 , n33813 );
buf ( n34057 , n34056 );
buf ( n34058 , n34057 );
xor ( n34059 , n33839 , n33968 );
xor ( n34060 , n34059 , n34043 );
buf ( n34061 , n34060 );
buf ( n34062 , n34061 );
xor ( n34063 , n34058 , n34062 );
xor ( n34064 , n33878 , n33921 );
xor ( n34065 , n34064 , n33963 );
buf ( n34066 , n34065 );
buf ( n34067 , n34066 );
buf ( n34068 , n8581 );
not ( n34069 , n34068 );
buf ( n34070 , n604 );
buf ( n34071 , n18175 );
and ( n34072 , n34070 , n34071 );
not ( n34073 , n34070 );
buf ( n34074 , n33867 );
and ( n34075 , n34073 , n34074 );
nor ( n34076 , n34072 , n34075 );
buf ( n34077 , n34076 );
buf ( n34078 , n34077 );
not ( n34079 , n34078 );
or ( n34080 , n34069 , n34079 );
buf ( n34081 , n33793 );
buf ( n34082 , n7790 );
nand ( n34083 , n34081 , n34082 );
buf ( n34084 , n34083 );
buf ( n34085 , n34084 );
nand ( n34086 , n34080 , n34085 );
buf ( n34087 , n34086 );
buf ( n34088 , n34087 );
buf ( n34089 , n2592 );
not ( n34090 , n34089 );
buf ( n34091 , n594 );
not ( n34092 , n34091 );
buf ( n34093 , n27548 );
not ( n34094 , n34093 );
or ( n34095 , n34092 , n34094 );
buf ( n34096 , n26737 );
buf ( n34097 , n2481 );
nand ( n34098 , n34096 , n34097 );
buf ( n34099 , n34098 );
buf ( n34100 , n34099 );
nand ( n34101 , n34095 , n34100 );
buf ( n34102 , n34101 );
buf ( n34103 , n34102 );
not ( n34104 , n34103 );
or ( n34105 , n34090 , n34104 );
nand ( n34106 , n33734 , n2541 );
buf ( n34107 , n34106 );
nand ( n34108 , n34105 , n34107 );
buf ( n34109 , n34108 );
buf ( n34110 , n34109 );
buf ( n34111 , n2452 );
not ( n34112 , n34111 );
buf ( n34113 , n33882 );
not ( n34114 , n34113 );
or ( n34115 , n34112 , n34114 );
xor ( n34116 , n33894 , n33895 );
buf ( n34117 , n34116 );
buf ( n34118 , n34117 );
buf ( n34119 , n28544 );
nand ( n34120 , n34118 , n34119 );
buf ( n34121 , n34120 );
buf ( n34122 , n34121 );
nand ( n34123 , n34115 , n34122 );
buf ( n34124 , n34123 );
buf ( n34125 , n34124 );
xor ( n34126 , n34110 , n34125 );
buf ( n34127 , n825 );
not ( n34128 , n34127 );
buf ( n34129 , n33905 );
not ( n34130 , n34129 );
or ( n34131 , n34128 , n34130 );
buf ( n34132 , n596 );
not ( n34133 , n34132 );
buf ( n34134 , n26851 );
not ( n34135 , n34134 );
or ( n34136 , n34133 , n34135 );
buf ( n34137 , n26810 );
buf ( n34138 , n2371 );
nand ( n34139 , n34137 , n34138 );
buf ( n34140 , n34139 );
buf ( n34141 , n34140 );
nand ( n34142 , n34136 , n34141 );
buf ( n34143 , n34142 );
buf ( n34144 , n34143 );
buf ( n34145 , n26278 );
nand ( n34146 , n34144 , n34145 );
buf ( n34147 , n34146 );
buf ( n34148 , n34147 );
nand ( n34149 , n34131 , n34148 );
buf ( n34150 , n34149 );
buf ( n34151 , n34150 );
and ( n34152 , n34126 , n34151 );
and ( n34153 , n34110 , n34125 );
or ( n34154 , n34152 , n34153 );
buf ( n34155 , n34154 );
buf ( n34156 , n34155 );
xor ( n34157 , n34088 , n34156 );
buf ( n34158 , n33924 );
buf ( n34159 , n5550 );
not ( n34160 , n34159 );
buf ( n34161 , n33950 );
not ( n34162 , n34161 );
or ( n34163 , n34160 , n34162 );
buf ( n34164 , n598 );
not ( n34165 , n34164 );
buf ( n34166 , n33390 );
not ( n34167 , n34166 );
or ( n34168 , n34165 , n34167 );
buf ( n34169 , n33220 );
buf ( n34170 , n818 );
nand ( n34171 , n34169 , n34170 );
buf ( n34172 , n34171 );
buf ( n34173 , n34172 );
nand ( n34174 , n34168 , n34173 );
buf ( n34175 , n34174 );
buf ( n34176 , n34175 );
buf ( n34177 , n5631 );
nand ( n34178 , n34176 , n34177 );
buf ( n34179 , n34178 );
buf ( n34180 , n34179 );
nand ( n34181 , n34163 , n34180 );
buf ( n34182 , n34181 );
buf ( n34183 , n34182 );
xor ( n34184 , n34158 , n34183 );
buf ( n34185 , n5430 );
not ( n34186 , n34185 );
and ( n34187 , n600 , n28244 );
not ( n34188 , n600 );
and ( n34189 , n34188 , n28247 );
or ( n34190 , n34187 , n34189 );
buf ( n34191 , n34190 );
not ( n34192 , n34191 );
or ( n34193 , n34186 , n34192 );
buf ( n34194 , n34020 );
buf ( n34195 , n10945 );
nand ( n34196 , n34194 , n34195 );
buf ( n34197 , n34196 );
buf ( n34198 , n34197 );
nand ( n34199 , n34193 , n34198 );
buf ( n34200 , n34199 );
buf ( n34201 , n34200 );
and ( n34202 , n34184 , n34201 );
and ( n34203 , n34158 , n34183 );
or ( n34204 , n34202 , n34203 );
buf ( n34205 , n34204 );
buf ( n34206 , n34205 );
and ( n34207 , n34157 , n34206 );
and ( n34208 , n34088 , n34156 );
or ( n34209 , n34207 , n34208 );
buf ( n34210 , n34209 );
buf ( n34211 , n34210 );
xor ( n34212 , n34067 , n34211 );
xor ( n34213 , n33928 , n33932 );
xor ( n34214 , n34213 , n33958 );
buf ( n34215 , n34214 );
buf ( n34216 , n34215 );
buf ( n34217 , n7619 );
not ( n34218 , n34217 );
xor ( n34219 , n28941 , n2912 );
buf ( n34220 , n34219 );
not ( n34221 , n34220 );
or ( n34222 , n34218 , n34221 );
buf ( n34223 , n602 );
not ( n34224 , n34223 );
buf ( n34225 , n29203 );
not ( n34226 , n34225 );
or ( n34227 , n34224 , n34226 );
buf ( n34228 , n33992 );
nand ( n34229 , n34227 , n34228 );
buf ( n34230 , n34229 );
buf ( n34231 , n34230 );
buf ( n34232 , n5655 );
nand ( n34233 , n34231 , n34232 );
buf ( n34234 , n34233 );
buf ( n34235 , n34234 );
nand ( n34236 , n34222 , n34235 );
buf ( n34237 , n34236 );
buf ( n34238 , n34237 );
buf ( n34239 , n10858 );
buf ( n34240 , n592 );
and ( n34241 , n34239 , n34240 );
buf ( n34242 , n34241 );
buf ( n34243 , n34242 );
buf ( n34244 , n26278 );
not ( n34245 , n34244 );
buf ( n34246 , n596 );
not ( n34247 , n34246 );
buf ( n34248 , n26786 );
not ( n34249 , n34248 );
or ( n34250 , n34247 , n34249 );
buf ( n34251 , n26782 );
buf ( n34252 , n2371 );
nand ( n34253 , n34251 , n34252 );
buf ( n34254 , n34253 );
buf ( n34255 , n34254 );
nand ( n34256 , n34250 , n34255 );
buf ( n34257 , n34256 );
buf ( n34258 , n34257 );
not ( n34259 , n34258 );
or ( n34260 , n34245 , n34259 );
buf ( n34261 , n34143 );
buf ( n34262 , n825 );
nand ( n34263 , n34261 , n34262 );
buf ( n34264 , n34263 );
buf ( n34265 , n34264 );
nand ( n34266 , n34260 , n34265 );
buf ( n34267 , n34266 );
buf ( n34268 , n34267 );
xor ( n34269 , n34243 , n34268 );
buf ( n34270 , n2452 );
not ( n34271 , n34270 );
buf ( n34272 , n34117 );
not ( n34273 , n34272 );
or ( n34274 , n34271 , n34273 );
buf ( n34275 , n592 );
not ( n34276 , n34275 );
buf ( n34277 , n10831 );
not ( n34278 , n34277 );
or ( n34279 , n34276 , n34278 );
buf ( n34280 , n10830 );
buf ( n34281 , n2416 );
nand ( n34282 , n34280 , n34281 );
buf ( n34283 , n34282 );
buf ( n34284 , n34283 );
nand ( n34285 , n34279 , n34284 );
buf ( n34286 , n34285 );
buf ( n34287 , n34286 );
buf ( n34288 , n28544 );
nand ( n34289 , n34287 , n34288 );
buf ( n34290 , n34289 );
buf ( n34291 , n34290 );
nand ( n34292 , n34274 , n34291 );
buf ( n34293 , n34292 );
buf ( n34294 , n34293 );
and ( n34295 , n34269 , n34294 );
and ( n34296 , n34243 , n34268 );
or ( n34297 , n34295 , n34296 );
buf ( n34298 , n34297 );
buf ( n34299 , n34298 );
xor ( n34300 , n34238 , n34299 );
buf ( n34301 , n606 );
not ( n34302 , n34301 );
buf ( n34303 , n33185 );
not ( n34304 , n34303 );
or ( n34305 , n34302 , n34304 );
buf ( n34306 , n18177 );
buf ( n34307 , n10836 );
nand ( n34308 , n34306 , n34307 );
buf ( n34309 , n34308 );
buf ( n34310 , n34309 );
nand ( n34311 , n34305 , n34310 );
buf ( n34312 , n34311 );
buf ( n34313 , n34312 );
buf ( n34314 , n10882 );
not ( n34315 , n34314 );
buf ( n34316 , n12475 );
nand ( n34317 , n34315 , n34316 );
buf ( n34318 , n34317 );
buf ( n34319 , n34318 );
nand ( n34320 , n34313 , n34319 );
buf ( n34321 , n34320 );
buf ( n34322 , n34321 );
and ( n34323 , n34300 , n34322 );
and ( n34324 , n34238 , n34299 );
or ( n34325 , n34323 , n34324 );
buf ( n34326 , n34325 );
buf ( n34327 , n34326 );
xor ( n34328 , n34216 , n34327 );
xor ( n34329 , n34003 , n34028 );
xor ( n34330 , n34329 , n34033 );
buf ( n34331 , n34330 );
buf ( n34332 , n34331 );
and ( n34333 , n34328 , n34332 );
and ( n34334 , n34216 , n34327 );
or ( n34335 , n34333 , n34334 );
buf ( n34336 , n34335 );
buf ( n34337 , n34336 );
and ( n34338 , n34212 , n34337 );
and ( n34339 , n34067 , n34211 );
or ( n34340 , n34338 , n34339 );
buf ( n34341 , n34340 );
buf ( n34342 , n34341 );
and ( n34343 , n34063 , n34342 );
and ( n34344 , n34058 , n34062 );
or ( n34345 , n34343 , n34344 );
buf ( n34346 , n34345 );
buf ( n34347 , n34346 );
xor ( n34348 , n33830 , n33834 );
xor ( n34349 , n34348 , n34048 );
buf ( n34350 , n34349 );
buf ( n34351 , n34350 );
nor ( n34352 , n34347 , n34351 );
buf ( n34353 , n34352 );
nor ( n34354 , n34054 , n34353 );
xor ( n34355 , n33131 , n33210 );
and ( n34356 , n34355 , n33289 );
and ( n34357 , n33131 , n33210 );
or ( n34358 , n34356 , n34357 );
buf ( n34359 , n34358 );
buf ( n34360 , n34359 );
xor ( n34361 , n33336 , n33348 );
and ( n34362 , n34361 , n33413 );
and ( n34363 , n33336 , n33348 );
or ( n34364 , n34362 , n34363 );
buf ( n34365 , n34364 );
buf ( n34366 , n34365 );
buf ( n34367 , n2541 );
not ( n34368 , n34367 );
buf ( n34369 , n594 );
not ( n34370 , n34369 );
buf ( n34371 , n33153 );
not ( n34372 , n34371 );
or ( n34373 , n34370 , n34372 );
buf ( n34374 , n28664 );
buf ( n34375 , n2481 );
nand ( n34376 , n34374 , n34375 );
buf ( n34377 , n34376 );
buf ( n34378 , n34377 );
nand ( n34379 , n34373 , n34378 );
buf ( n34380 , n34379 );
buf ( n34381 , n34380 );
not ( n34382 , n34381 );
or ( n34383 , n34368 , n34382 );
nand ( n34384 , n33275 , n2592 );
buf ( n34385 , n34384 );
nand ( n34386 , n34383 , n34385 );
buf ( n34387 , n34386 );
buf ( n34388 , n34387 );
buf ( n34389 , n11547 );
not ( n34390 , n34389 );
buf ( n34391 , n5430 );
not ( n34392 , n34391 );
buf ( n34393 , n34392 );
buf ( n34394 , n34393 );
not ( n34395 , n34394 );
or ( n34396 , n34390 , n34395 );
buf ( n34397 , n33123 );
nand ( n34398 , n34396 , n34397 );
buf ( n34399 , n34398 );
buf ( n34400 , n34399 );
xor ( n34401 , n34388 , n34400 );
buf ( n34402 , n26278 );
not ( n34403 , n34402 );
buf ( n34404 , n33340 );
not ( n34405 , n34404 );
or ( n34406 , n34403 , n34405 );
buf ( n34407 , n596 );
not ( n34408 , n34407 );
buf ( n34409 , n33318 );
not ( n34410 , n34409 );
or ( n34411 , n34408 , n34410 );
not ( n34412 , n33318 );
buf ( n34413 , n34412 );
buf ( n34414 , n2371 );
nand ( n34415 , n34413 , n34414 );
buf ( n34416 , n34415 );
buf ( n34417 , n34416 );
nand ( n34418 , n34411 , n34417 );
buf ( n34419 , n34418 );
buf ( n34420 , n34419 );
buf ( n34421 , n825 );
nand ( n34422 , n34420 , n34421 );
buf ( n34423 , n34422 );
buf ( n34424 , n34423 );
nand ( n34425 , n34406 , n34424 );
buf ( n34426 , n34425 );
buf ( n34427 , n34426 );
xor ( n34428 , n34401 , n34427 );
buf ( n34429 , n34428 );
buf ( n34430 , n34429 );
xor ( n34431 , n34366 , n34430 );
buf ( n34432 , n5550 );
not ( n34433 , n34432 );
buf ( n34434 , n598 );
not ( n34435 , n34434 );
buf ( n34436 , n33092 );
not ( n34437 , n34436 );
or ( n34438 , n34435 , n34437 );
buf ( n34439 , n33870 );
buf ( n34440 , n818 );
nand ( n34441 , n34439 , n34440 );
buf ( n34442 , n34441 );
buf ( n34443 , n34442 );
nand ( n34444 , n34438 , n34443 );
buf ( n34445 , n34444 );
buf ( n34446 , n34445 );
not ( n34447 , n34446 );
or ( n34448 , n34433 , n34447 );
buf ( n34449 , n33312 );
buf ( n34450 , n5631 );
nand ( n34451 , n34449 , n34450 );
buf ( n34452 , n34451 );
buf ( n34453 , n34452 );
nand ( n34454 , n34448 , n34453 );
buf ( n34455 , n34454 );
buf ( n34456 , n34455 );
xor ( n34457 , n33247 , n33280 );
and ( n34458 , n34457 , n33286 );
and ( n34459 , n33247 , n33280 );
or ( n34460 , n34458 , n34459 );
buf ( n34461 , n34460 );
buf ( n34462 , n34461 );
xor ( n34463 , n34456 , n34462 );
buf ( n34464 , n2452 );
not ( n34465 , n34464 );
buf ( n34466 , n592 );
buf ( n34467 , n33254 );
not ( n34468 , n34467 );
buf ( n34469 , n34468 );
buf ( n34470 , n34469 );
xor ( n34471 , n34466 , n34470 );
buf ( n34472 , n34471 );
buf ( n34473 , n34472 );
not ( n34474 , n34473 );
or ( n34475 , n34465 , n34474 );
buf ( n34476 , n33227 );
buf ( n34477 , n28544 );
nand ( n34478 , n34476 , n34477 );
buf ( n34479 , n34478 );
buf ( n34480 , n34479 );
nand ( n34481 , n34475 , n34480 );
buf ( n34482 , n34481 );
buf ( n34483 , n34482 );
buf ( n34484 , n33237 );
buf ( n34485 , n592 );
and ( n34486 , n34484 , n34485 );
buf ( n34487 , n34486 );
buf ( n34488 , n34487 );
xor ( n34489 , n34483 , n34488 );
buf ( n34490 , n33285 );
not ( n34491 , n34490 );
buf ( n34492 , n34491 );
buf ( n34493 , n34492 );
xor ( n34494 , n34489 , n34493 );
buf ( n34495 , n34494 );
buf ( n34496 , n34495 );
xor ( n34497 , n34463 , n34496 );
buf ( n34498 , n34497 );
buf ( n34499 , n34498 );
xor ( n34500 , n34431 , n34499 );
buf ( n34501 , n34500 );
buf ( n34502 , n34501 );
xor ( n34503 , n34360 , n34502 );
xor ( n34504 , n33416 , n33547 );
and ( n34505 , n34504 , n33625 );
and ( n34506 , n33416 , n33547 );
or ( n34507 , n34505 , n34506 );
buf ( n34508 , n34507 );
buf ( n34509 , n34508 );
xor ( n34510 , n34503 , n34509 );
buf ( n34511 , n34510 );
not ( n34512 , n34511 );
xor ( n34513 , n33292 , n33628 );
and ( n34514 , n34513 , n33823 );
and ( n34515 , n33292 , n33628 );
or ( n34516 , n34514 , n34515 );
buf ( n34517 , n34516 );
not ( n34518 , n34517 );
nand ( n34519 , n34512 , n34518 );
nand ( n34520 , n34354 , n34519 );
buf ( n34521 , n825 );
not ( n34522 , n34521 );
buf ( n34523 , n596 );
not ( n34524 , n34523 );
buf ( n34525 , n33455 );
not ( n34526 , n34525 );
or ( n34527 , n34524 , n34526 );
buf ( n34528 , n33455 );
not ( n34529 , n34528 );
buf ( n34530 , n34529 );
buf ( n34531 , n34530 );
buf ( n34532 , n2371 );
nand ( n34533 , n34531 , n34532 );
buf ( n34534 , n34533 );
buf ( n34535 , n34534 );
nand ( n34536 , n34527 , n34535 );
buf ( n34537 , n34536 );
buf ( n34538 , n34537 );
not ( n34539 , n34538 );
or ( n34540 , n34522 , n34539 );
buf ( n34541 , n34419 );
buf ( n34542 , n26278 );
nand ( n34543 , n34541 , n34542 );
buf ( n34544 , n34543 );
buf ( n34545 , n34544 );
nand ( n34546 , n34540 , n34545 );
buf ( n34547 , n34546 );
buf ( n34548 , n34547 );
buf ( n34549 , n5631 );
not ( n34550 , n34549 );
buf ( n34551 , n34445 );
not ( n34552 , n34551 );
or ( n34553 , n34550 , n34552 );
buf ( n34554 , n598 );
not ( n34555 , n34554 );
buf ( n34556 , n33113 );
not ( n34557 , n34556 );
or ( n34558 , n34555 , n34557 );
buf ( n34559 , n33110 );
buf ( n34560 , n818 );
nand ( n34561 , n34559 , n34560 );
buf ( n34562 , n34561 );
buf ( n34563 , n34562 );
nand ( n34564 , n34558 , n34563 );
buf ( n34565 , n34564 );
buf ( n34566 , n34565 );
buf ( n34567 , n5550 );
nand ( n34568 , n34566 , n34567 );
buf ( n34569 , n34568 );
buf ( n34570 , n34569 );
nand ( n34571 , n34553 , n34570 );
buf ( n34572 , n34571 );
buf ( n34573 , n34572 );
xor ( n34574 , n34548 , n34573 );
xor ( n34575 , n34483 , n34488 );
and ( n34576 , n34575 , n34493 );
and ( n34577 , n34483 , n34488 );
or ( n34578 , n34576 , n34577 );
buf ( n34579 , n34578 );
buf ( n34580 , n34579 );
xor ( n34581 , n34574 , n34580 );
buf ( n34582 , n34581 );
buf ( n34583 , n34582 );
xor ( n34584 , n34388 , n34400 );
and ( n34585 , n34584 , n34427 );
and ( n34586 , n34388 , n34400 );
or ( n34587 , n34585 , n34586 );
buf ( n34588 , n34587 );
buf ( n34589 , n34588 );
buf ( n34590 , n2452 );
not ( n34591 , n34590 );
buf ( n34592 , n592 );
not ( n34593 , n34592 );
buf ( n34594 , n28907 );
not ( n34595 , n34594 );
or ( n34596 , n34593 , n34595 );
buf ( n34597 , n28247 );
buf ( n34598 , n2416 );
nand ( n34599 , n34597 , n34598 );
buf ( n34600 , n34599 );
buf ( n34601 , n34600 );
nand ( n34602 , n34596 , n34601 );
buf ( n34603 , n34602 );
buf ( n34604 , n34603 );
not ( n34605 , n34604 );
or ( n34606 , n34591 , n34605 );
buf ( n34607 , n34472 );
buf ( n34608 , n28544 );
nand ( n34609 , n34607 , n34608 );
buf ( n34610 , n34609 );
buf ( n34611 , n34610 );
nand ( n34612 , n34606 , n34611 );
buf ( n34613 , n34612 );
buf ( n34614 , n34613 );
not ( n34615 , n2541 );
buf ( n34616 , n28947 );
buf ( n34617 , n34616 );
buf ( n34618 , n34617 );
and ( n34619 , n34618 , n594 );
not ( n34620 , n34618 );
and ( n34621 , n34620 , n2481 );
nor ( n34622 , n34619 , n34621 );
not ( n34623 , n34622 );
or ( n34624 , n34615 , n34623 );
nand ( n34625 , n34380 , n2592 );
nand ( n34626 , n34624 , n34625 );
buf ( n34627 , n34626 );
xor ( n34628 , n34614 , n34627 );
buf ( n34629 , n33220 );
buf ( n34630 , n592 );
and ( n34631 , n34629 , n34630 );
buf ( n34632 , n34631 );
buf ( n34633 , n34632 );
not ( n34634 , n34633 );
buf ( n34635 , n34634 );
buf ( n34636 , n34635 );
xor ( n34637 , n34628 , n34636 );
buf ( n34638 , n34637 );
buf ( n34639 , n34638 );
xor ( n34640 , n34589 , n34639 );
xor ( n34641 , n34456 , n34462 );
and ( n34642 , n34641 , n34496 );
and ( n34643 , n34456 , n34462 );
or ( n34644 , n34642 , n34643 );
buf ( n34645 , n34644 );
buf ( n34646 , n34645 );
xor ( n34647 , n34640 , n34646 );
buf ( n34648 , n34647 );
buf ( n34649 , n34648 );
xor ( n34650 , n34583 , n34649 );
xor ( n34651 , n34366 , n34430 );
and ( n34652 , n34651 , n34499 );
and ( n34653 , n34366 , n34430 );
or ( n34654 , n34652 , n34653 );
buf ( n34655 , n34654 );
buf ( n34656 , n34655 );
xor ( n34657 , n34650 , n34656 );
buf ( n34658 , n34657 );
xor ( n34659 , n34360 , n34502 );
and ( n34660 , n34659 , n34509 );
and ( n34661 , n34360 , n34502 );
or ( n34662 , n34660 , n34661 );
buf ( n34663 , n34662 );
nor ( n34664 , n34658 , n34663 );
buf ( n34665 , n34664 );
nor ( n34666 , n34520 , n34665 );
not ( n34667 , n34666 );
buf ( n34668 , n592 );
buf ( n34669 , n28664 );
and ( n34670 , n34668 , n34669 );
buf ( n34671 , n34670 );
buf ( n34672 , n34671 );
buf ( n34673 , n11218 );
not ( n34674 , n34673 );
buf ( n34675 , n26278 );
not ( n34676 , n34675 );
buf ( n34677 , n34676 );
buf ( n34678 , n34677 );
not ( n34679 , n34678 );
or ( n34680 , n34674 , n34679 );
buf ( n34681 , n596 );
not ( n34682 , n34681 );
buf ( n34683 , n33113 );
not ( n34684 , n34683 );
or ( n34685 , n34682 , n34684 );
buf ( n34686 , n33110 );
buf ( n34687 , n2371 );
nand ( n34688 , n34686 , n34687 );
buf ( n34689 , n34688 );
buf ( n34690 , n34689 );
nand ( n34691 , n34685 , n34690 );
buf ( n34692 , n34691 );
buf ( n34693 , n34692 );
nand ( n34694 , n34680 , n34693 );
buf ( n34695 , n34694 );
buf ( n34696 , n34695 );
xor ( n34697 , n34672 , n34696 );
buf ( n34698 , n2452 );
not ( n34699 , n34698 );
buf ( n34700 , n592 );
buf ( n34701 , n34412 );
xor ( n34702 , n34700 , n34701 );
buf ( n34703 , n34702 );
buf ( n34704 , n34703 );
not ( n34705 , n34704 );
or ( n34706 , n34699 , n34705 );
buf ( n34707 , n592 );
not ( n34708 , n34707 );
buf ( n34709 , n28941 );
not ( n34710 , n34709 );
or ( n34711 , n34708 , n34710 );
buf ( n34712 , n34618 );
buf ( n34713 , n2416 );
nand ( n34714 , n34712 , n34713 );
buf ( n34715 , n34714 );
buf ( n34716 , n34715 );
nand ( n34717 , n34711 , n34716 );
buf ( n34718 , n34717 );
buf ( n34719 , n34718 );
buf ( n34720 , n28544 );
nand ( n34721 , n34719 , n34720 );
buf ( n34722 , n34721 );
buf ( n34723 , n34722 );
nand ( n34724 , n34706 , n34723 );
buf ( n34725 , n34724 );
buf ( n34726 , n34725 );
and ( n34727 , n34697 , n34726 );
and ( n34728 , n34672 , n34696 );
or ( n34729 , n34727 , n34728 );
buf ( n34730 , n34729 );
buf ( n34731 , n34730 );
buf ( n34732 , n2452 );
not ( n34733 , n34732 );
and ( n34734 , n34530 , n2416 );
not ( n34735 , n34530 );
and ( n34736 , n34735 , n592 );
or ( n34737 , n34734 , n34736 );
buf ( n34738 , n34737 );
not ( n34739 , n34738 );
or ( n34740 , n34733 , n34739 );
buf ( n34741 , n34703 );
buf ( n34742 , n28544 );
nand ( n34743 , n34741 , n34742 );
buf ( n34744 , n34743 );
buf ( n34745 , n34744 );
nand ( n34746 , n34740 , n34745 );
buf ( n34747 , n34746 );
buf ( n34748 , n34747 );
buf ( n34749 , n2592 );
not ( n34750 , n34749 );
buf ( n34751 , n594 );
not ( n34752 , n34751 );
buf ( n34753 , n33859 );
not ( n34754 , n34753 );
or ( n34755 , n34752 , n34754 );
buf ( n34756 , n33859 );
not ( n34757 , n34756 );
buf ( n34758 , n34757 );
buf ( n34759 , n34758 );
buf ( n34760 , n2481 );
nand ( n34761 , n34759 , n34760 );
buf ( n34762 , n34761 );
buf ( n34763 , n34762 );
nand ( n34764 , n34755 , n34763 );
buf ( n34765 , n34764 );
buf ( n34766 , n34765 );
not ( n34767 , n34766 );
or ( n34768 , n34750 , n34767 );
buf ( n34769 , n594 );
not ( n34770 , n34769 );
buf ( n34771 , n33113 );
not ( n34772 , n34771 );
or ( n34773 , n34770 , n34772 );
buf ( n34774 , n33110 );
buf ( n34775 , n2481 );
nand ( n34776 , n34774 , n34775 );
buf ( n34777 , n34776 );
buf ( n34778 , n34777 );
nand ( n34779 , n34773 , n34778 );
buf ( n34780 , n34779 );
buf ( n34781 , n34780 );
buf ( n34782 , n2541 );
nand ( n34783 , n34781 , n34782 );
buf ( n34784 , n34783 );
buf ( n34785 , n34784 );
nand ( n34786 , n34768 , n34785 );
buf ( n34787 , n34786 );
buf ( n34788 , n34787 );
xor ( n34789 , n34748 , n34788 );
buf ( n34790 , n34618 );
buf ( n34791 , n592 );
nand ( n34792 , n34790 , n34791 );
buf ( n34793 , n34792 );
buf ( n34794 , n34793 );
xor ( n34795 , n34789 , n34794 );
buf ( n34796 , n34795 );
buf ( n34797 , n34796 );
xor ( n34798 , n34731 , n34797 );
buf ( n34799 , n2541 );
not ( n34800 , n34799 );
buf ( n34801 , n34765 );
not ( n34802 , n34801 );
or ( n34803 , n34800 , n34802 );
not ( n34804 , n594 );
not ( n34805 , n33299 );
or ( n34806 , n34804 , n34805 );
buf ( n34807 , n33305 );
buf ( n34808 , n2481 );
nand ( n34809 , n34807 , n34808 );
buf ( n34810 , n34809 );
nand ( n34811 , n34806 , n34810 );
nand ( n34812 , n34811 , n2592 );
buf ( n34813 , n34812 );
nand ( n34814 , n34803 , n34813 );
buf ( n34815 , n34814 );
buf ( n34816 , n34815 );
buf ( n34817 , n28247 );
buf ( n34818 , n592 );
nand ( n34819 , n34817 , n34818 );
buf ( n34820 , n34819 );
buf ( n34821 , n34820 );
not ( n34822 , n34821 );
buf ( n34823 , n34822 );
buf ( n34824 , n34823 );
xor ( n34825 , n34816 , n34824 );
xor ( n34826 , n34672 , n34696 );
xor ( n34827 , n34826 , n34726 );
buf ( n34828 , n34827 );
buf ( n34829 , n34828 );
and ( n34830 , n34825 , n34829 );
and ( n34831 , n34816 , n34824 );
or ( n34832 , n34830 , n34831 );
buf ( n34833 , n34832 );
buf ( n34834 , n34833 );
xor ( n34835 , n34798 , n34834 );
buf ( n34836 , n34835 );
not ( n34837 , n34836 );
buf ( n34838 , n2452 );
not ( n34839 , n34838 );
buf ( n34840 , n34718 );
not ( n34841 , n34840 );
or ( n34842 , n34839 , n34841 );
xor ( n34843 , n34668 , n34669 );
buf ( n34844 , n34843 );
buf ( n34845 , n34844 );
buf ( n34846 , n28544 );
nand ( n34847 , n34845 , n34846 );
buf ( n34848 , n34847 );
buf ( n34849 , n34848 );
nand ( n34850 , n34842 , n34849 );
buf ( n34851 , n34850 );
buf ( n34852 , n34851 );
buf ( n34853 , n594 );
not ( n34854 , n34853 );
buf ( n34855 , n33318 );
not ( n34856 , n34855 );
or ( n34857 , n34854 , n34856 );
buf ( n34858 , n29202 );
buf ( n34859 , n2481 );
nand ( n34860 , n34858 , n34859 );
buf ( n34861 , n34860 );
buf ( n34862 , n34861 );
nand ( n34863 , n34857 , n34862 );
buf ( n34864 , n34863 );
and ( n34865 , n34864 , n2592 );
not ( n34866 , n34865 );
nand ( n34867 , n2541 , n594 , n33299 );
not ( n34868 , n34810 );
nand ( n34869 , n34868 , n2541 );
nand ( n34870 , n34866 , n34867 , n34869 );
buf ( n34871 , n34870 );
xor ( n34872 , n34852 , n34871 );
buf ( n34873 , n26278 );
not ( n34874 , n34873 );
buf ( n34875 , n596 );
not ( n34876 , n34875 );
buf ( n34877 , n33859 );
not ( n34878 , n34877 );
or ( n34879 , n34876 , n34878 );
buf ( n34880 , n33870 );
buf ( n34881 , n2371 );
nand ( n34882 , n34880 , n34881 );
buf ( n34883 , n34882 );
buf ( n34884 , n34883 );
nand ( n34885 , n34879 , n34884 );
buf ( n34886 , n34885 );
buf ( n34887 , n34886 );
not ( n34888 , n34887 );
or ( n34889 , n34874 , n34888 );
buf ( n34890 , n34692 );
buf ( n34891 , n825 );
nand ( n34892 , n34890 , n34891 );
buf ( n34893 , n34892 );
buf ( n34894 , n34893 );
nand ( n34895 , n34889 , n34894 );
buf ( n34896 , n34895 );
buf ( n34897 , n34896 );
and ( n34898 , n34872 , n34897 );
and ( n34899 , n34852 , n34871 );
or ( n34900 , n34898 , n34899 );
buf ( n34901 , n34900 );
buf ( n34902 , n34901 );
xor ( n34903 , n34816 , n34824 );
xor ( n34904 , n34903 , n34829 );
buf ( n34905 , n34904 );
buf ( n34906 , n34905 );
xor ( n34907 , n34902 , n34906 );
buf ( n34908 , n34820 );
and ( n34909 , n34466 , n34470 );
buf ( n34910 , n34909 );
buf ( n34911 , n34910 );
buf ( n34912 , n28544 );
not ( n34913 , n34912 );
buf ( n34914 , n34603 );
not ( n34915 , n34914 );
or ( n34916 , n34913 , n34915 );
buf ( n34917 , n34844 );
buf ( n34918 , n2452 );
nand ( n34919 , n34917 , n34918 );
buf ( n34920 , n34919 );
buf ( n34921 , n34920 );
nand ( n34922 , n34916 , n34921 );
buf ( n34923 , n34922 );
buf ( n34924 , n34923 );
xor ( n34925 , n34911 , n34924 );
buf ( n34926 , n34565 );
buf ( n34927 , n5631 );
not ( n34928 , n34927 );
buf ( n34929 , n5618 );
nand ( n34930 , n34928 , n34929 );
buf ( n34931 , n34930 );
buf ( n34932 , n34931 );
nand ( n34933 , n34926 , n34932 );
buf ( n34934 , n34933 );
buf ( n34935 , n34934 );
and ( n34936 , n34925 , n34935 );
and ( n34937 , n34911 , n34924 );
or ( n34938 , n34936 , n34937 );
buf ( n34939 , n34938 );
buf ( n34940 , n34939 );
xor ( n34941 , n34908 , n34940 );
xor ( n34942 , n34852 , n34871 );
xor ( n34943 , n34942 , n34897 );
buf ( n34944 , n34943 );
buf ( n34945 , n34944 );
and ( n34946 , n34941 , n34945 );
and ( n34947 , n34908 , n34940 );
or ( n34948 , n34946 , n34947 );
buf ( n34949 , n34948 );
buf ( n34950 , n34949 );
and ( n34951 , n34907 , n34950 );
and ( n34952 , n34902 , n34906 );
or ( n34953 , n34951 , n34952 );
buf ( n34954 , n34953 );
not ( n34955 , n34954 );
and ( n34956 , n34837 , n34955 );
xor ( n34957 , n34583 , n34649 );
and ( n34958 , n34957 , n34656 );
and ( n34959 , n34583 , n34649 );
or ( n34960 , n34958 , n34959 );
buf ( n34961 , n34960 );
xor ( n34962 , n34548 , n34573 );
and ( n34963 , n34962 , n34580 );
and ( n34964 , n34548 , n34573 );
or ( n34965 , n34963 , n34964 );
buf ( n34966 , n34965 );
buf ( n34967 , n34966 );
xor ( n34968 , n34911 , n34924 );
xor ( n34969 , n34968 , n34935 );
buf ( n34970 , n34969 );
buf ( n34971 , n34970 );
xor ( n34972 , n34614 , n34627 );
and ( n34973 , n34972 , n34636 );
and ( n34974 , n34614 , n34627 );
or ( n34975 , n34973 , n34974 );
buf ( n34976 , n34975 );
buf ( n34977 , n34976 );
xor ( n34978 , n34971 , n34977 );
buf ( n34979 , n34632 );
not ( n34980 , n2592 );
not ( n34981 , n34622 );
or ( n34982 , n34980 , n34981 );
buf ( n34983 , n34864 );
buf ( n34984 , n2541 );
nand ( n34985 , n34983 , n34984 );
buf ( n34986 , n34985 );
nand ( n34987 , n34982 , n34986 );
buf ( n34988 , n34987 );
xor ( n34989 , n34979 , n34988 );
buf ( n34990 , n825 );
not ( n34991 , n34990 );
buf ( n34992 , n34886 );
not ( n34993 , n34992 );
or ( n34994 , n34991 , n34993 );
buf ( n34995 , n34537 );
buf ( n34996 , n26278 );
nand ( n34997 , n34995 , n34996 );
buf ( n34998 , n34997 );
buf ( n34999 , n34998 );
nand ( n35000 , n34994 , n34999 );
buf ( n35001 , n35000 );
buf ( n35002 , n35001 );
xor ( n35003 , n34989 , n35002 );
buf ( n35004 , n35003 );
buf ( n35005 , n35004 );
xor ( n35006 , n34978 , n35005 );
buf ( n35007 , n35006 );
buf ( n35008 , n35007 );
xor ( n35009 , n34967 , n35008 );
xor ( n35010 , n34589 , n34639 );
and ( n35011 , n35010 , n34646 );
and ( n35012 , n34589 , n34639 );
or ( n35013 , n35011 , n35012 );
buf ( n35014 , n35013 );
buf ( n35015 , n35014 );
xor ( n35016 , n35009 , n35015 );
buf ( n35017 , n35016 );
nor ( n35018 , n34961 , n35017 );
buf ( n35019 , n35018 );
xor ( n35020 , n34967 , n35008 );
and ( n35021 , n35020 , n35015 );
and ( n35022 , n34967 , n35008 );
or ( n35023 , n35021 , n35022 );
buf ( n35024 , n35023 );
buf ( n35025 , n35024 );
xor ( n35026 , n34979 , n34988 );
and ( n35027 , n35026 , n35002 );
and ( n35028 , n34979 , n34988 );
or ( n35029 , n35027 , n35028 );
buf ( n35030 , n35029 );
buf ( n35031 , n35030 );
xor ( n35032 , n34908 , n34940 );
xor ( n35033 , n35032 , n34945 );
buf ( n35034 , n35033 );
buf ( n35035 , n35034 );
xor ( n35036 , n35031 , n35035 );
xor ( n35037 , n34971 , n34977 );
and ( n35038 , n35037 , n35005 );
and ( n35039 , n34971 , n34977 );
or ( n35040 , n35038 , n35039 );
buf ( n35041 , n35040 );
buf ( n35042 , n35041 );
xor ( n35043 , n35036 , n35042 );
buf ( n35044 , n35043 );
buf ( n35045 , n35044 );
nor ( n35046 , n35025 , n35045 );
buf ( n35047 , n35046 );
buf ( n35048 , n35047 );
nor ( n35049 , n35019 , n35048 );
buf ( n35050 , n35049 );
buf ( n35051 , n35050 );
xor ( n35052 , n35031 , n35035 );
and ( n35053 , n35052 , n35042 );
and ( n35054 , n35031 , n35035 );
or ( n35055 , n35053 , n35054 );
buf ( n35056 , n35055 );
xor ( n35057 , n34902 , n34906 );
xor ( n35058 , n35057 , n34950 );
buf ( n35059 , n35058 );
or ( n35060 , n35056 , n35059 );
buf ( n35061 , n35060 );
nand ( n35062 , n35051 , n35061 );
buf ( n35063 , n35062 );
nor ( n35064 , n34956 , n35063 );
buf ( n35065 , n35064 );
not ( n35066 , n35065 );
buf ( n35067 , n35066 );
nor ( n35068 , n34667 , n35067 );
xor ( n35069 , n34058 , n34062 );
xor ( n35070 , n35069 , n34342 );
buf ( n35071 , n35070 );
buf ( n35072 , n35071 );
xor ( n35073 , n33973 , n33977 );
xor ( n35074 , n35073 , n34038 );
buf ( n35075 , n35074 );
buf ( n35076 , n35075 );
xor ( n35077 , n34067 , n34211 );
xor ( n35078 , n35077 , n34337 );
buf ( n35079 , n35078 );
buf ( n35080 , n35079 );
xor ( n35081 , n35076 , n35080 );
xor ( n35082 , n34088 , n34156 );
xor ( n35083 , n35082 , n34206 );
buf ( n35084 , n35083 );
buf ( n35085 , n35084 );
xor ( n35086 , n34110 , n34125 );
xor ( n35087 , n35086 , n34151 );
buf ( n35088 , n35087 );
buf ( n35089 , n35088 );
buf ( n35090 , n7790 );
not ( n35091 , n35090 );
buf ( n35092 , n34077 );
not ( n35093 , n35092 );
or ( n35094 , n35091 , n35093 );
buf ( n35095 , n604 );
not ( n35096 , n35095 );
buf ( n35097 , n30032 );
not ( n35098 , n35097 );
or ( n35099 , n35096 , n35098 );
buf ( n35100 , n30026 );
buf ( n35101 , n12329 );
nand ( n35102 , n35100 , n35101 );
buf ( n35103 , n35102 );
buf ( n35104 , n35103 );
nand ( n35105 , n35099 , n35104 );
buf ( n35106 , n35105 );
buf ( n35107 , n35106 );
buf ( n35108 , n8581 );
nand ( n35109 , n35107 , n35108 );
buf ( n35110 , n35109 );
buf ( n35111 , n35110 );
nand ( n35112 , n35094 , n35111 );
buf ( n35113 , n35112 );
buf ( n35114 , n35113 );
xor ( n35115 , n35089 , n35114 );
buf ( n35116 , n2592 );
not ( n35117 , n35116 );
buf ( n35118 , n594 );
not ( n35119 , n35118 );
buf ( n35120 , n26921 );
not ( n35121 , n35120 );
or ( n35122 , n35119 , n35121 );
buf ( n35123 , n26676 );
buf ( n35124 , n2481 );
nand ( n35125 , n35123 , n35124 );
buf ( n35126 , n35125 );
buf ( n35127 , n35126 );
nand ( n35128 , n35122 , n35127 );
buf ( n35129 , n35128 );
buf ( n35130 , n35129 );
not ( n35131 , n35130 );
or ( n35132 , n35117 , n35131 );
buf ( n35133 , n34102 );
buf ( n35134 , n2541 );
nand ( n35135 , n35133 , n35134 );
buf ( n35136 , n35135 );
buf ( n35137 , n35136 );
nand ( n35138 , n35132 , n35137 );
buf ( n35139 , n35138 );
buf ( n35140 , n35139 );
buf ( n35141 , n5631 );
not ( n35142 , n35141 );
and ( n35143 , n26053 , n818 );
not ( n35144 , n26053 );
and ( n35145 , n35144 , n598 );
or ( n35146 , n35143 , n35145 );
buf ( n35147 , n35146 );
not ( n35148 , n35147 );
or ( n35149 , n35142 , n35148 );
buf ( n35150 , n34175 );
buf ( n35151 , n5550 );
nand ( n35152 , n35150 , n35151 );
buf ( n35153 , n35152 );
buf ( n35154 , n35153 );
nand ( n35155 , n35149 , n35154 );
buf ( n35156 , n35155 );
buf ( n35157 , n35156 );
xor ( n35158 , n35140 , n35157 );
buf ( n35159 , n5430 );
not ( n35160 , n35159 );
buf ( n35161 , n600 );
not ( n35162 , n35161 );
buf ( n35163 , n27000 );
not ( n35164 , n35163 );
or ( n35165 , n35162 , n35164 );
buf ( n35166 , n18191 );
buf ( n35167 , n7650 );
nand ( n35168 , n35166 , n35167 );
buf ( n35169 , n35168 );
buf ( n35170 , n35169 );
nand ( n35171 , n35165 , n35170 );
buf ( n35172 , n35171 );
buf ( n35173 , n35172 );
not ( n35174 , n35173 );
or ( n35175 , n35160 , n35174 );
buf ( n35176 , n34190 );
buf ( n35177 , n2915 );
nand ( n35178 , n35176 , n35177 );
buf ( n35179 , n35178 );
buf ( n35180 , n35179 );
nand ( n35181 , n35175 , n35180 );
buf ( n35182 , n35181 );
buf ( n35183 , n35182 );
and ( n35184 , n35158 , n35183 );
and ( n35185 , n35140 , n35157 );
or ( n35186 , n35184 , n35185 );
buf ( n35187 , n35186 );
buf ( n35188 , n35187 );
and ( n35189 , n35115 , n35188 );
and ( n35190 , n35089 , n35114 );
or ( n35191 , n35189 , n35190 );
buf ( n35192 , n35191 );
buf ( n35193 , n35192 );
xor ( n35194 , n35085 , n35193 );
xor ( n35195 , n34158 , n34183 );
xor ( n35196 , n35195 , n34201 );
buf ( n35197 , n35196 );
buf ( n35198 , n35197 );
buf ( n35199 , n28868 );
buf ( n35200 , n592 );
and ( n35201 , n35199 , n35200 );
buf ( n35202 , n35201 );
buf ( n35203 , n35202 );
buf ( n35204 , n28544 );
not ( n35205 , n35204 );
buf ( n35206 , n30105 );
not ( n35207 , n35206 );
or ( n35208 , n35205 , n35207 );
and ( n35209 , n10829 , n2416 );
not ( n35210 , n10829 );
and ( n35211 , n35210 , n592 );
or ( n35212 , n35209 , n35211 );
nand ( n35213 , n35212 , n2452 );
buf ( n35214 , n35213 );
nand ( n35215 , n35208 , n35214 );
buf ( n35216 , n35215 );
buf ( n35217 , n35216 );
xor ( n35218 , n35203 , n35217 );
not ( n35219 , n26278 );
not ( n35220 , n30127 );
or ( n35221 , n35219 , n35220 );
nand ( n35222 , n34257 , n825 );
nand ( n35223 , n35221 , n35222 );
buf ( n35224 , n35223 );
and ( n35225 , n35218 , n35224 );
and ( n35226 , n35203 , n35217 );
or ( n35227 , n35225 , n35226 );
buf ( n35228 , n35227 );
buf ( n35229 , n35228 );
buf ( n35230 , n7790 );
not ( n35231 , n35230 );
buf ( n35232 , n35106 );
not ( n35233 , n35232 );
or ( n35234 , n35231 , n35233 );
and ( n35235 , n604 , n29203 );
not ( n35236 , n604 );
and ( n35237 , n35236 , n29202 );
or ( n35238 , n35235 , n35237 );
buf ( n35239 , n35238 );
buf ( n35240 , n8581 );
nand ( n35241 , n35239 , n35240 );
buf ( n35242 , n35241 );
buf ( n35243 , n35242 );
nand ( n35244 , n35234 , n35243 );
buf ( n35245 , n35244 );
buf ( n35246 , n35245 );
xor ( n35247 , n35229 , n35246 );
buf ( n35248 , n5655 );
not ( n35249 , n35248 );
buf ( n35250 , n34219 );
not ( n35251 , n35250 );
or ( n35252 , n35249 , n35251 );
buf ( n35253 , n28664 );
not ( n35254 , n35253 );
buf ( n35255 , n26971 );
not ( n35256 , n35255 );
and ( n35257 , n35254 , n35256 );
buf ( n35258 , n28664 );
buf ( n35259 , n11923 );
and ( n35260 , n35258 , n35259 );
nor ( n35261 , n35257 , n35260 );
buf ( n35262 , n35261 );
buf ( n35263 , n35262 );
nand ( n35264 , n35252 , n35263 );
buf ( n35265 , n35264 );
buf ( n35266 , n35265 );
and ( n35267 , n35247 , n35266 );
and ( n35268 , n35229 , n35246 );
or ( n35269 , n35267 , n35268 );
buf ( n35270 , n35269 );
buf ( n35271 , n35270 );
xor ( n35272 , n35198 , n35271 );
xor ( n35273 , n34238 , n34299 );
xor ( n35274 , n35273 , n34322 );
buf ( n35275 , n35274 );
buf ( n35276 , n35275 );
and ( n35277 , n35272 , n35276 );
and ( n35278 , n35198 , n35271 );
or ( n35279 , n35277 , n35278 );
buf ( n35280 , n35279 );
buf ( n35281 , n35280 );
and ( n35282 , n35194 , n35281 );
and ( n35283 , n35085 , n35193 );
or ( n35284 , n35282 , n35283 );
buf ( n35285 , n35284 );
buf ( n35286 , n35285 );
and ( n35287 , n35081 , n35286 );
and ( n35288 , n35076 , n35080 );
or ( n35289 , n35287 , n35288 );
buf ( n35290 , n35289 );
buf ( n35291 , n35290 );
nor ( n35292 , n35072 , n35291 );
buf ( n35293 , n35292 );
buf ( n35294 , n35293 );
xor ( n35295 , n35076 , n35080 );
xor ( n35296 , n35295 , n35286 );
buf ( n35297 , n35296 );
buf ( n35298 , n35297 );
xor ( n35299 , n34216 , n34327 );
xor ( n35300 , n35299 , n34332 );
buf ( n35301 , n35300 );
buf ( n35302 , n35301 );
xor ( n35303 , n35085 , n35193 );
xor ( n35304 , n35303 , n35281 );
buf ( n35305 , n35304 );
buf ( n35306 , n35305 );
xor ( n35307 , n35302 , n35306 );
xor ( n35308 , n34243 , n34268 );
xor ( n35309 , n35308 , n34294 );
buf ( n35310 , n35309 );
buf ( n35311 , n35310 );
buf ( n35312 , n10882 );
not ( n35313 , n35312 );
buf ( n35314 , n10836 );
buf ( n35315 , n33092 );
and ( n35316 , n35314 , n35315 );
not ( n35317 , n35314 );
buf ( n35318 , n18175 );
and ( n35319 , n35317 , n35318 );
nor ( n35320 , n35316 , n35319 );
buf ( n35321 , n35320 );
buf ( n35322 , n35321 );
not ( n35323 , n35322 );
or ( n35324 , n35313 , n35323 );
buf ( n35325 , n34312 );
buf ( n35326 , n607 );
nand ( n35327 , n35325 , n35326 );
buf ( n35328 , n35327 );
buf ( n35329 , n35328 );
nand ( n35330 , n35324 , n35329 );
buf ( n35331 , n35330 );
buf ( n35332 , n35331 );
xor ( n35333 , n35311 , n35332 );
buf ( n35334 , n2541 );
not ( n35335 , n35334 );
buf ( n35336 , n35129 );
not ( n35337 , n35336 );
or ( n35338 , n35335 , n35337 );
buf ( n35339 , n29921 );
buf ( n35340 , n2592 );
nand ( n35341 , n35339 , n35340 );
buf ( n35342 , n35341 );
buf ( n35343 , n35342 );
nand ( n35344 , n35338 , n35343 );
buf ( n35345 , n35344 );
buf ( n35346 , n35345 );
buf ( n35347 , n5550 );
not ( n35348 , n35347 );
buf ( n35349 , n35146 );
not ( n35350 , n35349 );
or ( n35351 , n35348 , n35350 );
nand ( n35352 , n29902 , n5631 );
buf ( n35353 , n35352 );
nand ( n35354 , n35351 , n35353 );
buf ( n35355 , n35354 );
buf ( n35356 , n35355 );
xor ( n35357 , n35346 , n35356 );
buf ( n35358 , n2915 );
not ( n35359 , n35358 );
buf ( n35360 , n35172 );
not ( n35361 , n35360 );
or ( n35362 , n35359 , n35361 );
buf ( n35363 , n29952 );
buf ( n35364 , n5430 );
nand ( n35365 , n35363 , n35364 );
buf ( n35366 , n35365 );
buf ( n35367 , n35366 );
nand ( n35368 , n35362 , n35367 );
buf ( n35369 , n35368 );
buf ( n35370 , n35369 );
and ( n35371 , n35357 , n35370 );
and ( n35372 , n35346 , n35356 );
or ( n35373 , n35371 , n35372 );
buf ( n35374 , n35373 );
buf ( n35375 , n35374 );
and ( n35376 , n35333 , n35375 );
and ( n35377 , n35311 , n35332 );
or ( n35378 , n35376 , n35377 );
buf ( n35379 , n35378 );
buf ( n35380 , n35379 );
xor ( n35381 , n35089 , n35114 );
xor ( n35382 , n35381 , n35188 );
buf ( n35383 , n35382 );
buf ( n35384 , n35383 );
xor ( n35385 , n35380 , n35384 );
xor ( n35386 , n35140 , n35157 );
xor ( n35387 , n35386 , n35183 );
buf ( n35388 , n35387 );
buf ( n35389 , n35388 );
buf ( n35390 , n7619 );
not ( n35391 , n35390 );
buf ( n35392 , n28247 );
buf ( n35393 , n602 );
and ( n35394 , n35392 , n35393 );
not ( n35395 , n35392 );
buf ( n35396 , n2912 );
and ( n35397 , n35395 , n35396 );
nor ( n35398 , n35394 , n35397 );
buf ( n35399 , n35398 );
buf ( n35400 , n35399 );
not ( n35401 , n35400 );
or ( n35402 , n35391 , n35401 );
buf ( n35403 , n28664 );
buf ( n35404 , n26693 );
and ( n35405 , n35403 , n35404 );
buf ( n35406 , n28667 );
buf ( n35407 , n26682 );
and ( n35408 , n35406 , n35407 );
nor ( n35409 , n35405 , n35408 );
buf ( n35410 , n35409 );
buf ( n35411 , n35410 );
nand ( n35412 , n35402 , n35411 );
buf ( n35413 , n35412 );
buf ( n35414 , n35413 );
xor ( n35415 , n35203 , n35217 );
xor ( n35416 , n35415 , n35224 );
buf ( n35417 , n35416 );
buf ( n35418 , n35417 );
xor ( n35419 , n35414 , n35418 );
buf ( n35420 , n8581 );
not ( n35421 , n35420 );
buf ( n35422 , n30075 );
not ( n35423 , n35422 );
or ( n35424 , n35421 , n35423 );
buf ( n35425 , n35238 );
buf ( n35426 , n7790 );
nand ( n35427 , n35425 , n35426 );
buf ( n35428 , n35427 );
buf ( n35429 , n35428 );
nand ( n35430 , n35424 , n35429 );
buf ( n35431 , n35430 );
buf ( n35432 , n35431 );
and ( n35433 , n35419 , n35432 );
and ( n35434 , n35414 , n35418 );
or ( n35435 , n35433 , n35434 );
buf ( n35436 , n35435 );
buf ( n35437 , n35436 );
xor ( n35438 , n35389 , n35437 );
xor ( n35439 , n35229 , n35246 );
xor ( n35440 , n35439 , n35266 );
buf ( n35441 , n35440 );
buf ( n35442 , n35441 );
and ( n35443 , n35438 , n35442 );
and ( n35444 , n35389 , n35437 );
or ( n35445 , n35443 , n35444 );
buf ( n35446 , n35445 );
buf ( n35447 , n35446 );
and ( n35448 , n35385 , n35447 );
and ( n35449 , n35380 , n35384 );
or ( n35450 , n35448 , n35449 );
buf ( n35451 , n35450 );
buf ( n35452 , n35451 );
and ( n35453 , n35307 , n35452 );
and ( n35454 , n35302 , n35306 );
or ( n35455 , n35453 , n35454 );
buf ( n35456 , n35455 );
buf ( n35457 , n35456 );
nor ( n35458 , n35298 , n35457 );
buf ( n35459 , n35458 );
buf ( n35460 , n35459 );
nor ( n35461 , n35294 , n35460 );
buf ( n35462 , n35461 );
not ( n35463 , n35462 );
xor ( n35464 , n35302 , n35306 );
xor ( n35465 , n35464 , n35452 );
buf ( n35466 , n35465 );
buf ( n35467 , n35466 );
xor ( n35468 , n35198 , n35271 );
xor ( n35469 , n35468 , n35276 );
buf ( n35470 , n35469 );
buf ( n35471 , n35470 );
xor ( n35472 , n35380 , n35384 );
xor ( n35473 , n35472 , n35447 );
buf ( n35474 , n35473 );
buf ( n35475 , n35474 );
xor ( n35476 , n35471 , n35475 );
xor ( n35477 , n30091 , n30116 );
and ( n35478 , n35477 , n30135 );
and ( n35479 , n30091 , n30116 );
or ( n35480 , n35478 , n35479 );
buf ( n35481 , n35480 );
buf ( n35482 , n35481 );
xor ( n35483 , n29907 , n29934 );
and ( n35484 , n35483 , n29960 );
and ( n35485 , n29907 , n29934 );
or ( n35486 , n35484 , n35485 );
buf ( n35487 , n35486 );
buf ( n35488 , n35487 );
xor ( n35489 , n35482 , n35488 );
buf ( n35490 , n607 );
not ( n35491 , n35490 );
buf ( n35492 , n35321 );
not ( n35493 , n35492 );
or ( n35494 , n35491 , n35493 );
buf ( n35495 , n33305 );
not ( n35496 , n35495 );
buf ( n35497 , n10882 );
nand ( n35498 , n35496 , n35497 );
buf ( n35499 , n35498 );
buf ( n35500 , n35499 );
nand ( n35501 , n35494 , n35500 );
buf ( n35502 , n35501 );
buf ( n35503 , n35502 );
and ( n35504 , n35489 , n35503 );
and ( n35505 , n35482 , n35488 );
or ( n35506 , n35504 , n35505 );
buf ( n35507 , n35506 );
buf ( n35508 , n35507 );
xor ( n35509 , n35311 , n35332 );
xor ( n35510 , n35509 , n35375 );
buf ( n35511 , n35510 );
buf ( n35512 , n35511 );
xor ( n35513 , n35508 , n35512 );
xor ( n35514 , n35346 , n35356 );
xor ( n35515 , n35514 , n35370 );
buf ( n35516 , n35515 );
buf ( n35517 , n35516 );
xor ( n35518 , n29995 , n30001 );
and ( n35519 , n35518 , n30047 );
and ( n35520 , n29995 , n30001 );
or ( n35521 , n35519 , n35520 );
buf ( n35522 , n35521 );
buf ( n35523 , n35522 );
xor ( n35524 , n35517 , n35523 );
xor ( n35525 , n35414 , n35418 );
xor ( n35526 , n35525 , n35432 );
buf ( n35527 , n35526 );
buf ( n35528 , n35527 );
and ( n35529 , n35524 , n35528 );
and ( n35530 , n35517 , n35523 );
or ( n35531 , n35529 , n35530 );
buf ( n35532 , n35531 );
buf ( n35533 , n35532 );
and ( n35534 , n35513 , n35533 );
and ( n35535 , n35508 , n35512 );
or ( n35536 , n35534 , n35535 );
buf ( n35537 , n35536 );
buf ( n35538 , n35537 );
and ( n35539 , n35476 , n35538 );
and ( n35540 , n35471 , n35475 );
or ( n35541 , n35539 , n35540 );
buf ( n35542 , n35541 );
buf ( n35543 , n35542 );
nand ( n35544 , n35467 , n35543 );
buf ( n35545 , n35544 );
buf ( n35546 , n35545 );
xor ( n35547 , n35471 , n35475 );
xor ( n35548 , n35547 , n35538 );
buf ( n35549 , n35548 );
buf ( n35550 , n35549 );
xor ( n35551 , n35389 , n35437 );
xor ( n35552 , n35551 , n35442 );
buf ( n35553 , n35552 );
buf ( n35554 , n35553 );
xor ( n35555 , n30086 , n30138 );
and ( n35556 , n35555 , n30145 );
and ( n35557 , n30086 , n30138 );
or ( n35558 , n35556 , n35557 );
buf ( n35559 , n35558 );
buf ( n35560 , n35559 );
xor ( n35561 , n35482 , n35488 );
xor ( n35562 , n35561 , n35503 );
buf ( n35563 , n35562 );
buf ( n35564 , n35563 );
xor ( n35565 , n35560 , n35564 );
xor ( n35566 , n29963 , n29969 );
and ( n35567 , n35566 , n30050 );
and ( n35568 , n29963 , n29969 );
or ( n35569 , n35567 , n35568 );
buf ( n35570 , n35569 );
buf ( n35571 , n35570 );
and ( n35572 , n35565 , n35571 );
and ( n35573 , n35560 , n35564 );
or ( n35574 , n35572 , n35573 );
buf ( n35575 , n35574 );
buf ( n35576 , n35575 );
xor ( n35577 , n35554 , n35576 );
xor ( n35578 , n35508 , n35512 );
xor ( n35579 , n35578 , n35533 );
buf ( n35580 , n35579 );
buf ( n35581 , n35580 );
and ( n35582 , n35577 , n35581 );
and ( n35583 , n35554 , n35576 );
or ( n35584 , n35582 , n35583 );
buf ( n35585 , n35584 );
buf ( n35586 , n35585 );
nand ( n35587 , n35550 , n35586 );
buf ( n35588 , n35587 );
buf ( n35589 , n35588 );
and ( n35590 , n35546 , n35589 );
buf ( n35591 , n35466 );
buf ( n35592 , n35542 );
nor ( n35593 , n35591 , n35592 );
buf ( n35594 , n35593 );
buf ( n35595 , n35594 );
nor ( n35596 , n35590 , n35595 );
buf ( n35597 , n35596 );
not ( n35598 , n35597 );
or ( n35599 , n35463 , n35598 );
buf ( n35600 , n35071 );
buf ( n35601 , n35290 );
nor ( n35602 , n35600 , n35601 );
buf ( n35603 , n35602 );
buf ( n35604 , n35603 );
not ( n35605 , n35604 );
nand ( n35606 , n35456 , n35297 );
buf ( n35607 , n35606 );
not ( n35608 , n35607 );
and ( n35609 , n35605 , n35608 );
buf ( n35610 , n35071 );
buf ( n35611 , n35290 );
and ( n35612 , n35610 , n35611 );
buf ( n35613 , n35612 );
buf ( n35614 , n35613 );
nor ( n35615 , n35609 , n35614 );
buf ( n35616 , n35615 );
nand ( n35617 , n35599 , n35616 );
not ( n35618 , n35617 );
nor ( n35619 , n35542 , n35466 );
buf ( n35620 , n35549 );
buf ( n35621 , n35585 );
nor ( n35622 , n35620 , n35621 );
buf ( n35623 , n35622 );
nor ( n35624 , n35619 , n35623 );
and ( n35625 , n35462 , n35624 );
xor ( n35626 , n35517 , n35523 );
xor ( n35627 , n35626 , n35528 );
buf ( n35628 , n35627 );
buf ( n35629 , n35628 );
xor ( n35630 , n35560 , n35564 );
xor ( n35631 , n35630 , n35571 );
buf ( n35632 , n35631 );
buf ( n35633 , n35632 );
xor ( n35634 , n35629 , n35633 );
xor ( n35635 , n30066 , n30148 );
and ( n35636 , n35635 , n30155 );
and ( n35637 , n30066 , n30148 );
or ( n35638 , n35636 , n35637 );
buf ( n35639 , n35638 );
buf ( n35640 , n35639 );
xor ( n35641 , n35634 , n35640 );
buf ( n35642 , n35641 );
buf ( n35643 , n35642 );
not ( n35644 , n35643 );
buf ( n35645 , n35644 );
buf ( n35646 , n35645 );
xor ( n35647 , n30053 , n30059 );
and ( n35648 , n35647 , n30158 );
and ( n35649 , n30053 , n30059 );
or ( n35650 , n35648 , n35649 );
buf ( n35651 , n35650 );
buf ( n35652 , n35651 );
not ( n35653 , n35652 );
buf ( n35654 , n35653 );
buf ( n35655 , n35654 );
nand ( n35656 , n35646 , n35655 );
buf ( n35657 , n35656 );
xor ( n35658 , n35554 , n35576 );
xor ( n35659 , n35658 , n35581 );
buf ( n35660 , n35659 );
buf ( n35661 , n35660 );
not ( n35662 , n35661 );
xor ( n35663 , n35629 , n35633 );
and ( n35664 , n35663 , n35640 );
and ( n35665 , n35629 , n35633 );
or ( n35666 , n35664 , n35665 );
buf ( n35667 , n35666 );
buf ( n35668 , n35667 );
not ( n35669 , n35668 );
buf ( n35670 , n35669 );
buf ( n35671 , n35670 );
nand ( n35672 , n35662 , n35671 );
buf ( n35673 , n35672 );
nand ( n35674 , n35657 , n35673 );
not ( n35675 , n35674 );
not ( n35676 , n28980 );
not ( n35677 , n28985 );
or ( n35678 , n35676 , n35677 );
buf ( n35679 , n29242 );
buf ( n35680 , n29248 );
nand ( n35681 , n35679 , n35680 );
buf ( n35682 , n35681 );
nand ( n35683 , n35678 , n35682 );
not ( n35684 , n35683 );
buf ( n35685 , n30160 );
buf ( n35686 , n30167 );
nor ( n35687 , n35685 , n35686 );
buf ( n35688 , n35687 );
buf ( n35689 , n35688 );
buf ( n35690 , n29251 );
nor ( n35691 , n35689 , n35690 );
buf ( n35692 , n35691 );
not ( n35693 , n35692 );
or ( n35694 , n35684 , n35693 );
buf ( n35695 , n35642 );
buf ( n35696 , n35651 );
nand ( n35697 , n35695 , n35696 );
buf ( n35698 , n35697 );
buf ( n35699 , n35698 );
buf ( n35700 , n30160 );
buf ( n35701 , n30167 );
nand ( n35702 , n35700 , n35701 );
buf ( n35703 , n35702 );
buf ( n35704 , n35703 );
and ( n35705 , n35699 , n35704 );
buf ( n35706 , n35705 );
nand ( n35707 , n35694 , n35706 );
nand ( n35708 , n35675 , n35707 );
not ( n35709 , n35674 );
and ( n35710 , n29878 , n30173 );
nand ( n35711 , n35709 , n29013 , n35710 );
buf ( n35712 , n35667 );
buf ( n35713 , n35660 );
buf ( n35714 , n35713 );
buf ( n35715 , n35714 );
nand ( n35716 , n35712 , n35715 );
nand ( n35717 , n35708 , n35711 , n35716 );
nand ( n35718 , n35625 , n35717 );
nand ( n35719 , n35618 , n35718 );
nand ( n35720 , n35068 , n35719 );
not ( n35721 , n35720 );
buf ( n35722 , n33825 );
buf ( n35723 , n34052 );
nand ( n35724 , n35722 , n35723 );
buf ( n35725 , n35724 );
not ( n35726 , n35725 );
buf ( n35727 , n34346 );
buf ( n35728 , n34350 );
nand ( n35729 , n35727 , n35728 );
buf ( n35730 , n35729 );
not ( n35731 , n35730 );
or ( n35732 , n35726 , n35731 );
not ( n35733 , n33825 );
buf ( n35734 , n34052 );
not ( n35735 , n35734 );
buf ( n35736 , n35735 );
nand ( n35737 , n35733 , n35736 );
nand ( n35738 , n35732 , n35737 );
not ( n35739 , n35738 );
nand ( n35740 , n34658 , n34663 );
nand ( n35741 , n34511 , n34517 );
and ( n35742 , n35740 , n35741 );
not ( n35743 , n35742 );
or ( n35744 , n35739 , n35743 );
not ( n35745 , n34511 );
nand ( n35746 , n35745 , n34518 );
not ( n35747 , n34658 );
not ( n35748 , n34663 );
nand ( n35749 , n35747 , n35748 );
nand ( n35750 , n35746 , n35749 );
nand ( n35751 , n35740 , n35750 );
nand ( n35752 , n35744 , n35751 );
not ( n35753 , n35752 );
buf ( n35754 , n35067 );
not ( n35755 , n35754 );
buf ( n35756 , n35755 );
and ( n35757 , n35753 , n35756 );
or ( n35758 , n34836 , n34954 );
nand ( n35759 , n34961 , n35017 );
nor ( n35760 , n35044 , n35024 );
or ( n35761 , n35759 , n35760 );
nand ( n35762 , n35044 , n35024 );
nand ( n35763 , n35761 , n35762 );
nand ( n35764 , n35758 , n35763 , n35060 );
nand ( n35765 , n35059 , n35056 );
not ( n35766 , n35765 );
nand ( n35767 , n35758 , n35766 );
nand ( n35768 , n34836 , n34954 );
nand ( n35769 , n35764 , n35767 , n35768 );
nor ( n35770 , n35757 , n35769 );
buf ( n35771 , n35770 );
not ( n35772 , n35771 );
buf ( n35773 , n28544 );
not ( n35774 , n35773 );
buf ( n35775 , n592 );
buf ( n35776 , n34758 );
xor ( n35777 , n35775 , n35776 );
buf ( n35778 , n35777 );
buf ( n35779 , n35778 );
not ( n35780 , n35779 );
or ( n35781 , n35774 , n35780 );
buf ( n35782 , n592 );
not ( n35783 , n35782 );
buf ( n35784 , n33113 );
not ( n35785 , n35784 );
or ( n35786 , n35783 , n35785 );
buf ( n35787 , n33110 );
buf ( n35788 , n2416 );
nand ( n35789 , n35787 , n35788 );
buf ( n35790 , n35789 );
buf ( n35791 , n35790 );
nand ( n35792 , n35786 , n35791 );
buf ( n35793 , n35792 );
buf ( n35794 , n35793 );
buf ( n35795 , n2452 );
nand ( n35796 , n35794 , n35795 );
buf ( n35797 , n35796 );
buf ( n35798 , n35797 );
nand ( n35799 , n35781 , n35798 );
buf ( n35800 , n35799 );
buf ( n35801 , n35800 );
buf ( n35802 , n34530 );
buf ( n35803 , n592 );
nand ( n35804 , n35802 , n35803 );
buf ( n35805 , n35804 );
buf ( n35806 , n35805 );
xor ( n35807 , n35801 , n35806 );
buf ( n35808 , n2540 );
not ( n35809 , n35808 );
buf ( n35810 , n2591 );
not ( n35811 , n35810 );
or ( n35812 , n35809 , n35811 );
buf ( n35813 , n34780 );
nand ( n35814 , n35812 , n35813 );
buf ( n35815 , n35814 );
buf ( n35816 , n35815 );
and ( n35817 , n34700 , n34701 );
buf ( n35818 , n35817 );
buf ( n35819 , n35818 );
xor ( n35820 , n35816 , n35819 );
buf ( n35821 , n2452 );
not ( n35822 , n35821 );
buf ( n35823 , n35778 );
not ( n35824 , n35823 );
or ( n35825 , n35822 , n35824 );
buf ( n35826 , n34737 );
buf ( n35827 , n28544 );
nand ( n35828 , n35826 , n35827 );
buf ( n35829 , n35828 );
buf ( n35830 , n35829 );
nand ( n35831 , n35825 , n35830 );
buf ( n35832 , n35831 );
buf ( n35833 , n35832 );
and ( n35834 , n35820 , n35833 );
and ( n35835 , n35816 , n35819 );
or ( n35836 , n35834 , n35835 );
buf ( n35837 , n35836 );
buf ( n35838 , n35837 );
and ( n35839 , n35807 , n35838 );
and ( n35840 , n35801 , n35806 );
or ( n35841 , n35839 , n35840 );
buf ( n35842 , n35841 );
buf ( n35843 , n2519 );
not ( n35844 , n35843 );
buf ( n35845 , n28544 );
not ( n35846 , n35845 );
buf ( n35847 , n35846 );
buf ( n35848 , n35847 );
not ( n35849 , n35848 );
or ( n35850 , n35844 , n35849 );
buf ( n35851 , n35793 );
nand ( n35852 , n35850 , n35851 );
buf ( n35853 , n35852 );
buf ( n35854 , n35853 );
and ( n35855 , n35775 , n35776 );
buf ( n35856 , n35855 );
buf ( n35857 , n35856 );
xor ( n35858 , n35854 , n35857 );
buf ( n35859 , n35805 );
not ( n35860 , n35859 );
buf ( n35861 , n35860 );
buf ( n35862 , n35861 );
xor ( n35863 , n35858 , n35862 );
buf ( n35864 , n35863 );
or ( n35865 , n35842 , n35864 );
not ( n35866 , n35865 );
buf ( n35867 , n35866 );
xor ( n35868 , n35854 , n35857 );
and ( n35869 , n35868 , n35862 );
and ( n35870 , n35854 , n35857 );
or ( n35871 , n35869 , n35870 );
buf ( n35872 , n35871 );
buf ( n35873 , n33110 );
buf ( n35874 , n592 );
nand ( n35875 , n35873 , n35874 );
buf ( n35876 , n35875 );
buf ( n35877 , C0 );
buf ( n35878 , n35877 );
nor ( n35879 , n35867 , n35878 );
buf ( n35880 , n35879 );
buf ( n35881 , n35880 );
not ( n35882 , n35881 );
buf ( n35883 , n34793 );
not ( n35884 , n35883 );
buf ( n35885 , n35884 );
buf ( n35886 , n35885 );
xor ( n35887 , n35816 , n35819 );
xor ( n35888 , n35887 , n35833 );
buf ( n35889 , n35888 );
buf ( n35890 , n35889 );
xor ( n35891 , n35886 , n35890 );
xor ( n35892 , n34748 , n34788 );
and ( n35893 , n35892 , n34794 );
and ( n35894 , n34748 , n34788 );
or ( n35895 , n35893 , n35894 );
buf ( n35896 , n35895 );
buf ( n35897 , n35896 );
xor ( n35898 , n35891 , n35897 );
buf ( n35899 , n35898 );
xor ( n35900 , n34731 , n34797 );
and ( n35901 , n35900 , n34834 );
and ( n35902 , n34731 , n34797 );
or ( n35903 , n35901 , n35902 );
buf ( n35904 , n35903 );
nand ( n35905 , n35899 , n35904 );
buf ( n35906 , n35905 );
xor ( n35907 , n35886 , n35890 );
and ( n35908 , n35907 , n35897 );
and ( n35909 , n35886 , n35890 );
or ( n35910 , n35908 , n35909 );
buf ( n35911 , n35910 );
buf ( n35912 , n35911 );
xor ( n35913 , n35801 , n35806 );
xor ( n35914 , n35913 , n35838 );
buf ( n35915 , n35914 );
buf ( n35916 , n35915 );
nor ( n35917 , n35912 , n35916 );
buf ( n35918 , n35917 );
buf ( n35919 , n35918 );
or ( n35920 , n35906 , n35919 );
buf ( n35921 , n35911 );
buf ( n35922 , n35915 );
nand ( n35923 , n35921 , n35922 );
buf ( n35924 , n35923 );
buf ( n35925 , n35924 );
nand ( n35926 , n35920 , n35925 );
buf ( n35927 , n35926 );
buf ( n35928 , n35927 );
not ( n35929 , n35928 );
or ( n35930 , n35882 , n35929 );
nand ( n35931 , n35842 , n35864 );
buf ( n35932 , n35931 );
buf ( n35933 , n35877 );
nor ( n35934 , n35932 , n35933 );
buf ( n35935 , n35934 );
buf ( n35936 , n35935 );
buf ( n35937 , n35872 );
buf ( n35938 , n35876 );
and ( n35939 , n35937 , n35938 );
buf ( n35940 , n35939 );
buf ( n35941 , n35940 );
nor ( n35942 , n35936 , n35941 );
buf ( n35943 , n35942 );
buf ( n35944 , n35943 );
nand ( n35945 , n35930 , n35944 );
buf ( n35946 , n35945 );
buf ( n35947 , n35946 );
nor ( n35948 , n35772 , n35947 );
buf ( n35949 , n35948 );
not ( n35950 , n35949 );
or ( n35951 , n35721 , n35950 );
buf ( n35952 , n35880 );
not ( n35953 , n35952 );
nor ( n35954 , n35904 , n35899 );
buf ( n35955 , n35954 );
buf ( n35956 , n35918 );
nor ( n35957 , n35955 , n35956 );
buf ( n35958 , n35957 );
buf ( n35959 , n35958 );
not ( n35960 , n35959 );
or ( n35961 , n35953 , n35960 );
buf ( n35962 , n35946 );
not ( n35963 , n35962 );
buf ( n35964 , n35963 );
buf ( n35965 , n35964 );
nand ( n35966 , n35961 , n35965 );
buf ( n35967 , n35966 );
nand ( n35968 , n35951 , n35967 );
not ( n35969 , n35968 );
not ( n35970 , n35969 );
not ( n35971 , n35970 );
not ( n35972 , n35971 );
not ( n35973 , n35972 );
buf ( n35974 , n35973 );
not ( n35975 , n35974 );
or ( n35976 , n33085 , n35975 );
buf ( n35977 , n35973 );
not ( n35978 , n35977 );
buf ( n35979 , n35978 );
buf ( n35980 , n35979 );
buf ( n35981 , n33080 );
nand ( n35982 , n35980 , n35981 );
buf ( n35983 , n35982 );
buf ( n35984 , n35983 );
nand ( n35985 , n35976 , n35984 );
buf ( n35986 , n35985 );
buf ( n35987 , n35986 );
not ( n35988 , n35987 );
or ( n35989 , n32974 , n35988 );
buf ( n35990 , n33083 );
not ( n35991 , n35990 );
not ( n35992 , n35958 );
not ( n35993 , n35769 );
or ( n35994 , n35992 , n35993 );
buf ( n35995 , n35927 );
not ( n35996 , n35995 );
buf ( n35997 , n35996 );
nand ( n35998 , n35994 , n35997 );
and ( n35999 , n35998 , n35865 );
not ( n36000 , n35931 );
nor ( n36001 , n35999 , n36000 );
nand ( n36002 , n34666 , n35625 , n35717 );
not ( n36003 , n36002 );
buf ( n36004 , n35064 );
buf ( n36005 , n35958 );
nand ( n36006 , n36004 , n36005 );
buf ( n36007 , n36006 );
nor ( n36008 , n35866 , n36007 );
nand ( n36009 , n36003 , n36008 );
not ( n36010 , n34354 );
not ( n36011 , n34664 );
nand ( n36012 , n36011 , n34519 );
nor ( n36013 , n36010 , n36012 );
not ( n36014 , n36013 );
not ( n36015 , n35617 );
or ( n36016 , n36014 , n36015 );
not ( n36017 , n35742 );
not ( n36018 , n35738 );
or ( n36019 , n36017 , n36018 );
nand ( n36020 , n35740 , n35750 );
nand ( n36021 , n36019 , n36020 );
nand ( n36022 , n36016 , n36021 );
nand ( n36023 , n36022 , n36008 );
nand ( n36024 , n36001 , n36009 , n36023 );
buf ( n36025 , n35877 );
buf ( n36026 , n35940 );
nor ( n36027 , n36025 , n36026 );
buf ( n36028 , n36027 );
xor ( n36029 , n36024 , n36028 );
buf ( n36030 , n36029 );
not ( n36031 , n36030 );
buf ( n36032 , n36031 );
buf ( n36033 , n36032 );
buf ( n36034 , n36033 );
buf ( n36035 , n36034 );
buf ( n36036 , n36035 );
not ( n36037 , n36036 );
buf ( n36038 , n36037 );
buf ( n36039 , n36038 );
not ( n36040 , n36039 );
buf ( n36041 , n36040 );
buf ( n36042 , n36041 );
buf ( n36043 , n36042 );
buf ( n36044 , n36043 );
buf ( n36045 , n36044 );
not ( n36046 , n36045 );
or ( n36047 , n35991 , n36046 );
buf ( n36048 , n33080 );
buf ( n36049 , n36032 );
not ( n36050 , n36049 );
buf ( n36051 , n36050 );
buf ( n36052 , n36051 );
not ( n36053 , n36052 );
buf ( n36054 , n36053 );
buf ( n36055 , n36054 );
not ( n36056 , n36055 );
buf ( n36057 , n36056 );
buf ( n36058 , n36057 );
nand ( n36059 , n36048 , n36058 );
buf ( n36060 , n36059 );
buf ( n36061 , n36060 );
nand ( n36062 , n36047 , n36061 );
buf ( n36063 , n36062 );
buf ( n36064 , n36063 );
buf ( n36065 , n32963 );
buf ( n36066 , n33037 );
not ( n36067 , n36066 );
buf ( n36068 , n33067 );
not ( n36069 , n36068 );
or ( n36070 , n36067 , n36069 );
buf ( n36071 , n33073 );
nand ( n36072 , n36070 , n36071 );
buf ( n36073 , n36072 );
buf ( n36074 , n36073 );
not ( n36075 , n36074 );
buf ( n36076 , n36075 );
buf ( n36077 , n36076 );
not ( n36078 , n36077 );
buf ( n36079 , n32943 );
not ( n36080 , n36079 );
or ( n36081 , n36078 , n36080 );
and ( n36082 , n32846 , n32938 );
not ( n36083 , n32846 );
and ( n36084 , n36083 , n32941 );
or ( n36085 , n36082 , n36084 );
buf ( n36086 , n36085 );
buf ( n36087 , n36073 );
nand ( n36088 , n36086 , n36087 );
buf ( n36089 , n36088 );
buf ( n36090 , n36089 );
nand ( n36091 , n36081 , n36090 );
buf ( n36092 , n36091 );
buf ( n36093 , n36092 );
nand ( n36094 , n36065 , n36093 );
buf ( n36095 , n36094 );
buf ( n36096 , n36095 );
buf ( n36097 , n36096 );
buf ( n36098 , n36097 );
buf ( n36099 , n36098 );
not ( n36100 , n36099 );
buf ( n36101 , n36100 );
buf ( n36102 , n36101 );
buf ( n36103 , n36102 );
buf ( n36104 , n36103 );
buf ( n36105 , n36104 );
buf ( n36106 , n36105 );
buf ( n36107 , n36106 );
buf ( n36108 , n36107 );
not ( n36109 , n36108 );
buf ( n36110 , n36109 );
buf ( n36111 , n36110 );
not ( n36112 , n36111 );
buf ( n36113 , n36112 );
buf ( n36114 , n36113 );
nand ( n36115 , n36064 , n36114 );
buf ( n36116 , n36115 );
buf ( n36117 , n36116 );
nand ( n36118 , n35989 , n36117 );
buf ( n36119 , n36118 );
buf ( n36120 , n36119 );
not ( n36121 , n36120 );
buf ( n36122 , n32354 );
not ( n36123 , n36122 );
buf ( n36124 , n33045 );
xor ( n36125 , n32978 , n33014 );
and ( n36126 , n36125 , n33021 );
and ( n36127 , n32978 , n33014 );
or ( n36128 , n36126 , n36127 );
buf ( n36129 , n36128 );
buf ( n36130 , n36129 );
buf ( n36131 , n30529 );
not ( n36132 , n36131 );
buf ( n36133 , n33000 );
not ( n36134 , n36133 );
or ( n36135 , n36132 , n36134 );
buf ( n36136 , n576 );
not ( n36137 , n36136 );
buf ( n36138 , n18170 );
not ( n36139 , n36138 );
or ( n36140 , n36137 , n36139 );
buf ( n36141 , n18167 );
buf ( n36142 , n7809 );
nand ( n36143 , n36141 , n36142 );
buf ( n36144 , n36143 );
buf ( n36145 , n36144 );
nand ( n36146 , n36140 , n36145 );
buf ( n36147 , n36146 );
buf ( n36148 , n36147 );
buf ( n36149 , n18340 );
nand ( n36150 , n36148 , n36149 );
buf ( n36151 , n36150 );
buf ( n36152 , n36151 );
nand ( n36153 , n36135 , n36152 );
buf ( n36154 , n36153 );
buf ( n36155 , n36154 );
buf ( n36156 , n30562 );
buf ( n36157 , n576 );
nand ( n36158 , n36156 , n36157 );
buf ( n36159 , n36158 );
buf ( n36160 , n36159 );
xor ( n36161 , n36155 , n36160 );
xor ( n36162 , n32990 , n32993 );
and ( n36163 , n36162 , n33011 );
and ( n36164 , n32990 , n32993 );
or ( n36165 , n36163 , n36164 );
buf ( n36166 , n36165 );
buf ( n36167 , n36166 );
xor ( n36168 , n36161 , n36167 );
buf ( n36169 , n36168 );
buf ( n36170 , n36169 );
or ( n36171 , n36130 , n36170 );
buf ( n36172 , n36171 );
nand ( n36173 , n36172 , n33029 );
buf ( n36174 , n36173 );
xor ( n36175 , n36155 , n36160 );
and ( n36176 , n36175 , n36167 );
and ( n36177 , n36155 , n36160 );
or ( n36178 , n36176 , n36177 );
buf ( n36179 , n36178 );
buf ( n36180 , n36179 );
buf ( n36181 , n31494 );
not ( n36182 , n36181 );
buf ( n36183 , n30529 );
not ( n36184 , n36183 );
buf ( n36185 , n36184 );
buf ( n36186 , n36185 );
not ( n36187 , n36186 );
or ( n36188 , n36182 , n36187 );
buf ( n36189 , n36147 );
nand ( n36190 , n36188 , n36189 );
buf ( n36191 , n36190 );
buf ( n36192 , n36191 );
and ( n36193 , n32997 , n32998 );
buf ( n36194 , n36193 );
buf ( n36195 , n36194 );
xor ( n36196 , n36192 , n36195 );
buf ( n36197 , n36159 );
not ( n36198 , n36197 );
buf ( n36199 , n36198 );
buf ( n36200 , n36199 );
xor ( n36201 , n36196 , n36200 );
buf ( n36202 , n36201 );
buf ( n36203 , n36202 );
nor ( n36204 , n36180 , n36203 );
buf ( n36205 , n36204 );
buf ( n36206 , n36205 );
nor ( n36207 , n36174 , n36206 );
buf ( n36208 , n36207 );
buf ( n36209 , n36208 );
nand ( n36210 , n36124 , n36209 );
buf ( n36211 , n36210 );
buf ( n36212 , n36211 );
nor ( n36213 , n36123 , n36212 );
buf ( n36214 , n36213 );
not ( n36215 , n36214 );
not ( n36216 , n32708 );
not ( n36217 , n36216 );
buf ( n36218 , n32725 );
not ( n36219 , n36218 );
buf ( n36220 , n24634 );
not ( n36221 , n36220 );
or ( n36222 , n36219 , n36221 );
buf ( n36223 , n32740 );
nand ( n36224 , n36222 , n36223 );
buf ( n36225 , n36224 );
not ( n36226 , n36225 );
or ( n36227 , n36217 , n36226 );
not ( n36228 , n32683 );
not ( n36229 , n32694 );
nor ( n36230 , n36228 , n36229 );
nand ( n36231 , n36227 , n36230 );
not ( n36232 , n36231 );
or ( n36233 , n36215 , n36232 );
not ( n36234 , n36211 );
nand ( n36235 , n36234 , n32803 );
nand ( n36236 , n36233 , n36235 );
not ( n36237 , n36236 );
not ( n36238 , n36237 );
buf ( n36239 , n36205 );
not ( n36240 , n36239 );
buf ( n36241 , n36240 );
buf ( n36242 , n36241 );
not ( n36243 , n36242 );
buf ( n36244 , n33058 );
buf ( n36245 , n36173 );
or ( n36246 , n36244 , n36245 );
buf ( n36247 , n36172 );
not ( n36248 , n36247 );
buf ( n36249 , n36248 );
buf ( n36250 , n36249 );
buf ( n36251 , n33033 );
or ( n36252 , n36250 , n36251 );
buf ( n36253 , n36129 );
buf ( n36254 , n36169 );
nand ( n36255 , n36253 , n36254 );
buf ( n36256 , n36255 );
buf ( n36257 , n36256 );
nand ( n36258 , n36252 , n36257 );
buf ( n36259 , n36258 );
buf ( n36260 , n36259 );
not ( n36261 , n36260 );
buf ( n36262 , n36261 );
buf ( n36263 , n36262 );
nand ( n36264 , n36246 , n36263 );
buf ( n36265 , n36264 );
buf ( n36266 , n36265 );
not ( n36267 , n36266 );
or ( n36268 , n36243 , n36267 );
buf ( n36269 , n36179 );
buf ( n36270 , n36202 );
nand ( n36271 , n36269 , n36270 );
buf ( n36272 , n36271 );
buf ( n36273 , n36272 );
nand ( n36274 , n36268 , n36273 );
buf ( n36275 , n36274 );
xor ( n36276 , n36192 , n36195 );
and ( n36277 , n36276 , n36200 );
and ( n36278 , n36192 , n36195 );
or ( n36279 , n36277 , n36278 );
buf ( n36280 , n36279 );
buf ( n36281 , n36280 );
buf ( n36282 , n18170 );
not ( n36283 , n36282 );
buf ( n36284 , n576 );
nand ( n36285 , n36283 , n36284 );
buf ( n36286 , n36285 );
buf ( n36287 , n36286 );
and ( n36288 , n36281 , n36287 );
buf ( n36289 , n36288 );
not ( n36290 , n36289 );
buf ( n36291 , n36280 );
buf ( n36292 , n36286 );
or ( n36293 , n36291 , n36292 );
buf ( n36294 , n36293 );
nand ( n36295 , n36290 , n36294 );
nor ( n36296 , n36275 , n36295 );
not ( n36297 , n36296 );
or ( n36298 , n36238 , n36297 );
or ( n36299 , n36236 , n36275 );
nand ( n36300 , n36299 , n36295 );
nand ( n36301 , n36298 , n36300 );
not ( n36302 , n36301 );
buf ( n36303 , n33048 );
not ( n36304 , n36303 );
buf ( n36305 , n36173 );
nor ( n36306 , n36304 , n36305 );
buf ( n36307 , n36306 );
buf ( n36308 , n36307 );
not ( n36309 , n36308 );
buf ( n36310 , n32809 );
not ( n36311 , n36310 );
or ( n36312 , n36309 , n36311 );
buf ( n36313 , n36265 );
not ( n36314 , n36313 );
buf ( n36315 , n36314 );
buf ( n36316 , n36315 );
nand ( n36317 , n36312 , n36316 );
buf ( n36318 , n36317 );
buf ( n36319 , n36241 );
buf ( n36320 , n36272 );
nand ( n36321 , n36319 , n36320 );
buf ( n36322 , n36321 );
buf ( n36323 , n36322 );
not ( n36324 , n36323 );
buf ( n36325 , n36324 );
and ( n36326 , n36318 , n36325 );
not ( n36327 , n36318 );
and ( n36328 , n36327 , n36322 );
nor ( n36329 , n36326 , n36328 );
buf ( n36330 , n36329 );
not ( n36331 , n36330 );
buf ( n36332 , n36331 );
not ( n36333 , n36332 );
or ( n36334 , n36302 , n36333 );
not ( n36335 , n36301 );
nand ( n36336 , n36329 , n36335 );
nand ( n36337 , n36334 , n36336 );
and ( n36338 , n36208 , n36294 );
not ( n36339 , n36338 );
not ( n36340 , n33064 );
or ( n36341 , n36339 , n36340 );
buf ( n36342 , n36241 );
not ( n36343 , n36342 );
buf ( n36344 , n36259 );
not ( n36345 , n36344 );
or ( n36346 , n36343 , n36345 );
buf ( n36347 , n36272 );
nand ( n36348 , n36346 , n36347 );
buf ( n36349 , n36348 );
buf ( n36350 , n36349 );
buf ( n36351 , n36294 );
and ( n36352 , n36350 , n36351 );
buf ( n36353 , n36289 );
nor ( n36354 , n36352 , n36353 );
buf ( n36355 , n36354 );
nand ( n36356 , n36341 , n36355 );
not ( n36357 , n36356 );
buf ( n36358 , n36357 );
buf ( n36359 , n36358 );
buf ( n36360 , n36359 );
buf ( n36361 , n36360 );
buf ( n36362 , n36361 );
buf ( n36363 , n36362 );
buf ( n36364 , n36363 );
not ( n36365 , n36364 );
not ( n36366 , n36022 );
nand ( n36367 , n36366 , n36002 );
buf ( n36368 , n36367 );
not ( n36369 , n36368 );
buf ( n36370 , n36369 );
buf ( n36371 , n36370 );
not ( n36372 , n36371 );
buf ( n36373 , n36372 );
not ( n36374 , n36373 );
buf ( n36375 , n35763 );
and ( n36376 , n36375 , n35060 );
nor ( n36377 , n36376 , n35766 );
not ( n36378 , n36377 );
nand ( n36379 , n35758 , n35768 );
nor ( n36380 , n36378 , n36379 );
nand ( n36381 , n36374 , n36380 );
buf ( n36382 , n35063 );
not ( n36383 , n36382 );
buf ( n36384 , n36383 );
not ( n36385 , n36384 );
not ( n36386 , n36379 );
nor ( n36387 , n36385 , n36386 );
nand ( n36388 , n36373 , n36387 );
not ( n36389 , n36386 );
not ( n36390 , n36377 );
and ( n36391 , n36389 , n36390 );
nor ( n36392 , n36379 , n36384 );
and ( n36393 , n36377 , n36392 );
nor ( n36394 , n36391 , n36393 );
nand ( n36395 , n36381 , n36388 , n36394 );
buf ( n36396 , n36395 );
buf ( n36397 , n36396 );
buf ( n36398 , n36397 );
buf ( n36399 , n36398 );
buf ( n36400 , n36399 );
not ( n36401 , n36400 );
buf ( n36402 , n36401 );
buf ( n36403 , n36402 );
not ( n36404 , n36403 );
or ( n36405 , n36365 , n36404 );
buf ( n36406 , n36399 );
buf ( n36407 , n36363 );
not ( n36408 , n36407 );
buf ( n36409 , n36408 );
buf ( n36410 , n36409 );
nand ( n36411 , n36406 , n36410 );
buf ( n36412 , n36411 );
buf ( n36413 , n36412 );
nand ( n36414 , n36405 , n36413 );
buf ( n36415 , n36414 );
buf ( n36416 , n36363 );
not ( n36417 , n36416 );
and ( n36418 , n35904 , n35899 );
nor ( n36419 , n36418 , n35954 );
not ( n36420 , n35068 );
not ( n36421 , n35719 );
or ( n36422 , n36420 , n36421 );
nand ( n36423 , n36422 , n35770 );
xor ( n36424 , n36419 , n36423 );
buf ( n36425 , n36424 );
buf ( n36426 , n36425 );
buf ( n36427 , n36426 );
buf ( n36428 , n36427 );
not ( n36429 , n36428 );
buf ( n36430 , n36429 );
buf ( n36431 , n36430 );
not ( n36432 , n36431 );
or ( n36433 , n36417 , n36432 );
buf ( n36434 , n36427 );
buf ( n36435 , n36409 );
nand ( n36436 , n36434 , n36435 );
buf ( n36437 , n36436 );
buf ( n36438 , n36437 );
nand ( n36439 , n36433 , n36438 );
buf ( n36440 , n36439 );
buf ( n36441 , n36440 );
buf ( n36442 , n36337 );
buf ( n36443 , n36442 );
buf ( n36444 , n36443 );
buf ( n36445 , n36444 );
not ( n36446 , n36445 );
buf ( n36447 , n36446 );
buf ( n36448 , n36447 );
buf ( n36449 , n36448 );
buf ( n36450 , n36449 );
buf ( n36451 , n36450 );
not ( n36452 , n36451 );
buf ( n36453 , n36452 );
buf ( n36454 , n36453 );
buf ( n36455 , n36454 );
buf ( n36456 , n36455 );
buf ( n36457 , n36456 );
nand ( n36458 , n36441 , n36457 );
buf ( n36459 , n36458 );
buf ( n36460 , n36459 );
nand ( n36461 , C1 , n36460 );
buf ( n36462 , n36461 );
buf ( n36463 , n36462 );
not ( n36464 , n36463 );
buf ( n36465 , n36464 );
buf ( n36466 , n36465 );
not ( n36467 , n36466 );
or ( n36468 , n36121 , n36467 );
buf ( n36469 , n36329 );
not ( n36470 , n33029 );
not ( n36471 , n33064 );
or ( n36472 , n36470 , n36471 );
nand ( n36473 , n36472 , n33033 );
buf ( n36474 , n36172 );
buf ( n36475 , n36256 );
nand ( n36476 , n36474 , n36475 );
buf ( n36477 , n36476 );
buf ( n36478 , n36477 );
not ( n36479 , n36478 );
buf ( n36480 , n36479 );
and ( n36481 , n36473 , n36480 );
not ( n36482 , n36473 );
and ( n36483 , n36482 , n36477 );
nor ( n36484 , n36481 , n36483 );
buf ( n36485 , n36484 );
not ( n36486 , n36485 );
buf ( n36487 , n36486 );
buf ( n36488 , n36487 );
not ( n36489 , n36488 );
buf ( n36490 , n36489 );
and ( n36491 , n36469 , n36490 );
buf ( n36492 , n36329 );
buf ( n36493 , n36492 );
not ( n36494 , n36493 );
buf ( n36495 , n36494 );
and ( n36496 , n36495 , n36487 );
nor ( n36497 , n36491 , n36496 );
buf ( n36498 , n33074 );
not ( n36499 , n36498 );
buf ( n36500 , n36499 );
buf ( n36501 , n36500 );
buf ( n36502 , n36473 );
buf ( n36503 , n36480 );
and ( n36504 , n36502 , n36503 );
not ( n36505 , n36502 );
buf ( n36506 , n36477 );
and ( n36507 , n36505 , n36506 );
nor ( n36508 , n36504 , n36507 );
buf ( n36509 , n36508 );
buf ( n36510 , n36509 );
and ( n36511 , n36501 , n36510 );
not ( n36512 , n36501 );
buf ( n36513 , n36487 );
and ( n36514 , n36512 , n36513 );
nor ( n36515 , n36511 , n36514 );
buf ( n36516 , n36515 );
nand ( n36517 , n36497 , n36516 );
buf ( n36518 , n36517 );
buf ( n36519 , n36518 );
buf ( n36520 , n36519 );
buf ( n36521 , n36520 );
not ( n36522 , n36521 );
buf ( n36523 , n36522 );
buf ( n36524 , n36523 );
buf ( n36525 , n36524 );
not ( n36526 , n36525 );
buf ( n36527 , n36492 );
buf ( n36528 , n36527 );
not ( n36529 , n36528 );
buf ( n36530 , n36529 );
buf ( n36531 , n36530 );
not ( n36532 , n36531 );
buf ( n36533 , n36532 );
buf ( n36534 , n36533 );
not ( n36535 , n36534 );
not ( n36536 , n35954 );
nand ( n36537 , n36423 , n36536 );
buf ( n36538 , n35918 );
not ( n36539 , n36538 );
buf ( n36540 , n35924 );
nand ( n36541 , n36539 , n36540 );
buf ( n36542 , n36541 );
not ( n36543 , n36542 );
or ( n36544 , n36537 , n36543 );
not ( n36545 , n35905 );
nand ( n36546 , n36545 , n36542 );
and ( n36547 , n36546 , n36536 );
not ( n36548 , n36547 );
not ( n36549 , n36423 );
or ( n36550 , n36548 , n36549 );
not ( n36551 , n35905 );
nor ( n36552 , n36551 , n36542 );
not ( n36553 , n36552 );
nand ( n36554 , n36553 , n36546 );
nand ( n36555 , n36550 , n36554 );
nand ( n36556 , n36544 , n36555 );
buf ( n36557 , n36556 );
buf ( n36558 , n36557 );
buf ( n36559 , n36558 );
buf ( n36560 , n36559 );
buf ( n36561 , n36560 );
buf ( n36562 , n36561 );
buf ( n36563 , n36562 );
not ( n36564 , n36563 );
buf ( n36565 , n36564 );
buf ( n36566 , n36565 );
buf ( n36567 , n36566 );
buf ( n36568 , n36567 );
buf ( n36569 , n36568 );
not ( n36570 , n36569 );
or ( n36571 , n36535 , n36570 );
buf ( n36572 , n36568 );
not ( n36573 , n36572 );
buf ( n36574 , n36573 );
buf ( n36575 , n36574 );
buf ( n36576 , n36533 );
not ( n36577 , n36576 );
buf ( n36578 , n36577 );
buf ( n36579 , n36578 );
nand ( n36580 , n36575 , n36579 );
buf ( n36581 , n36580 );
buf ( n36582 , n36581 );
nand ( n36583 , n36571 , n36582 );
buf ( n36584 , n36583 );
buf ( n36585 , n36584 );
not ( n36586 , n36585 );
or ( n36587 , n36526 , n36586 );
buf ( n36588 , n36533 );
not ( n36589 , n36588 );
not ( n36590 , n36002 );
nand ( n36591 , n36013 , n35617 );
not ( n36592 , n36591 );
or ( n36593 , n36590 , n36592 );
buf ( n36594 , n36007 );
not ( n36595 , n36594 );
buf ( n36596 , n36595 );
nand ( n36597 , n36593 , n36596 );
buf ( n36598 , n35753 );
buf ( n36599 , n36596 );
and ( n36600 , n36598 , n36599 );
buf ( n36601 , n35998 );
nor ( n36602 , n36600 , n36601 );
buf ( n36603 , n36602 );
nand ( n36604 , n36597 , n36603 );
nand ( n36605 , n35865 , n35931 );
not ( n36606 , n36605 );
and ( n36607 , n36604 , n36606 );
not ( n36608 , n36604 );
and ( n36609 , n36608 , n36605 );
nor ( n36610 , n36607 , n36609 );
buf ( n36611 , n36610 );
buf ( n36612 , n36611 );
not ( n36613 , n36612 );
buf ( n36614 , n36613 );
buf ( n36615 , n36614 );
not ( n36616 , n36615 );
buf ( n36617 , n36616 );
buf ( n36618 , n36617 );
not ( n36619 , n36618 );
buf ( n36620 , n36619 );
buf ( n36621 , n36620 );
buf ( n36622 , n36621 );
buf ( n36623 , n36622 );
buf ( n36624 , n36623 );
not ( n36625 , n36624 );
or ( n36626 , n36589 , n36625 );
buf ( n36627 , n36623 );
not ( n36628 , n36627 );
buf ( n36629 , n36628 );
buf ( n36630 , n36629 );
buf ( n36631 , n36578 );
nand ( n36632 , n36630 , n36631 );
buf ( n36633 , n36632 );
buf ( n36634 , n36633 );
nand ( n36635 , n36626 , n36634 );
buf ( n36636 , n36635 );
buf ( n36637 , n36636 );
buf ( n36638 , n36516 );
buf ( n36639 , n36638 );
buf ( n36640 , n36639 );
buf ( n36641 , n36640 );
not ( n36642 , n36641 );
buf ( n36643 , n36642 );
buf ( n36644 , n36643 );
nand ( n36645 , n36637 , n36644 );
buf ( n36646 , n36645 );
buf ( n36647 , n36646 );
nand ( n36648 , n36587 , n36647 );
buf ( n36649 , n36648 );
buf ( n36650 , n36649 );
nand ( n36651 , n36468 , n36650 );
buf ( n36652 , n36651 );
buf ( n36653 , n36652 );
buf ( n36654 , n36462 );
buf ( n36655 , n36119 );
not ( n36656 , n36655 );
buf ( n36657 , n36656 );
buf ( n36658 , n36657 );
nand ( n36659 , n36654 , n36658 );
buf ( n36660 , n36659 );
buf ( n36661 , n36660 );
and ( n36662 , n36653 , n36661 );
buf ( n36663 , n36662 );
buf ( n36664 , n36663 );
not ( n36665 , n36664 );
buf ( n36666 , n36665 );
buf ( n36667 , n36666 );
buf ( n36668 , n36119 );
nand ( n36669 , n36667 , n36668 );
buf ( n36670 , n36669 );
not ( n36671 , n36670 );
buf ( n36672 , n36533 );
not ( n36673 , n36672 );
buf ( n36674 , n36044 );
not ( n36675 , n36674 );
or ( n36676 , n36673 , n36675 );
buf ( n36677 , n36057 );
buf ( n36678 , n36578 );
nand ( n36679 , n36677 , n36678 );
buf ( n36680 , n36679 );
buf ( n36681 , n36680 );
nand ( n36682 , n36676 , n36681 );
buf ( n36683 , n36682 );
buf ( n36684 , n36683 );
not ( n36685 , n36684 );
buf ( n36686 , n36523 );
not ( n36687 , n36686 );
buf ( n36688 , n36687 );
buf ( n36689 , n36688 );
nor ( n36690 , n36685 , n36689 );
buf ( n36691 , n36690 );
buf ( n36692 , n36691 );
buf ( n36693 , n35979 );
not ( n36694 , n36693 );
buf ( n36695 , n36578 );
not ( n36696 , n36695 );
and ( n36697 , n36694 , n36696 );
buf ( n36698 , n35979 );
buf ( n36699 , n36578 );
and ( n36700 , n36698 , n36699 );
nor ( n36701 , n36697 , n36700 );
buf ( n36702 , n36701 );
buf ( n36703 , n36702 );
buf ( n36704 , n36643 );
not ( n36705 , n36704 );
buf ( n36706 , n36705 );
buf ( n36707 , n36706 );
nor ( n36708 , n36703 , n36707 );
buf ( n36709 , n36708 );
buf ( n36710 , n36709 );
nor ( n36711 , n36692 , n36710 );
buf ( n36712 , n36711 );
buf ( n36713 , n36712 );
buf ( n36714 , n36409 );
buf ( n36715 , n36568 );
xnor ( n36716 , n36714 , n36715 );
buf ( n36717 , n36716 );
buf ( n36718 , n36409 );
buf ( n36719 , n36623 );
and ( n36720 , n36718 , n36719 );
not ( n36721 , n36718 );
buf ( n36722 , n36629 );
and ( n36723 , n36721 , n36722 );
nor ( n36724 , n36720 , n36723 );
buf ( n36725 , n36724 );
buf ( n36726 , n36725 );
buf ( n36727 , n36456 );
nand ( n36728 , n36726 , n36727 );
buf ( n36729 , n36728 );
buf ( n36730 , n36729 );
nand ( n36731 , C1 , n36730 );
buf ( n36732 , n36731 );
buf ( n36733 , n36732 );
xor ( n36734 , n36713 , n36733 );
buf ( n36735 , n36643 );
not ( n36736 , n36735 );
buf ( n36737 , n36683 );
not ( n36738 , n36737 );
or ( n36739 , n36736 , n36738 );
buf ( n36740 , n36636 );
buf ( n36741 , n36523 );
nand ( n36742 , n36740 , n36741 );
buf ( n36743 , n36742 );
buf ( n36744 , n36743 );
nand ( n36745 , n36739 , n36744 );
buf ( n36746 , n36745 );
buf ( n36747 , n36746 );
not ( n36748 , n36747 );
buf ( n36749 , n32972 );
not ( n36750 , n36749 );
buf ( n36751 , n36750 );
buf ( n36752 , n36751 );
not ( n36753 , n36752 );
buf ( n36754 , n36110 );
not ( n36755 , n36754 );
or ( n36756 , n36753 , n36755 );
buf ( n36757 , n35986 );
nand ( n36758 , n36756 , n36757 );
buf ( n36759 , n36758 );
buf ( n36760 , n36759 );
not ( n36761 , n36760 );
buf ( n36762 , n36761 );
buf ( n36763 , n36762 );
nand ( n36764 , n36748 , n36763 );
buf ( n36765 , n36764 );
buf ( n36766 , n36765 );
not ( n36767 , n36766 );
buf ( n36768 , n36717 );
not ( n36769 , n36768 );
buf ( n36770 , n36456 );
not ( n36771 , n36770 );
buf ( n36772 , n36771 );
buf ( n36773 , n36772 );
not ( n36774 , n36773 );
and ( n36775 , n36769 , n36774 );
nor ( n36776 , n36775 , C0 );
buf ( n36777 , n36776 );
buf ( n36778 , n36777 );
not ( n36779 , n36778 );
buf ( n36780 , n36779 );
buf ( n36781 , n36780 );
not ( n36782 , n36781 );
or ( n36783 , n36767 , n36782 );
buf ( n36784 , n36759 );
buf ( n36785 , n36746 );
nand ( n36786 , n36784 , n36785 );
buf ( n36787 , n36786 );
buf ( n36788 , n36787 );
nand ( n36789 , n36783 , n36788 );
buf ( n36790 , n36789 );
buf ( n36791 , n36790 );
xor ( n36792 , n36734 , n36791 );
buf ( n36793 , n36792 );
not ( n36794 , n36793 );
buf ( n36795 , n36657 );
not ( n36796 , n36795 );
buf ( n36797 , n36663 );
not ( n36798 , n36797 );
or ( n36799 , n36796 , n36798 );
buf ( n36800 , n36777 );
not ( n36801 , n36800 );
buf ( n36802 , n36762 );
not ( n36803 , n36802 );
buf ( n36804 , n36746 );
not ( n36805 , n36804 );
or ( n36806 , n36803 , n36805 );
buf ( n36807 , n36746 );
buf ( n36808 , n36762 );
or ( n36809 , n36807 , n36808 );
nand ( n36810 , n36806 , n36809 );
buf ( n36811 , n36810 );
buf ( n36812 , n36811 );
not ( n36813 , n36812 );
and ( n36814 , n36801 , n36813 );
buf ( n36815 , n36777 );
buf ( n36816 , n36811 );
and ( n36817 , n36815 , n36816 );
nor ( n36818 , n36814 , n36817 );
buf ( n36819 , n36818 );
buf ( n36820 , n36819 );
not ( n36821 , n36820 );
buf ( n36822 , n36821 );
buf ( n36823 , n36822 );
nand ( n36824 , n36799 , n36823 );
buf ( n36825 , n36824 );
nand ( n36826 , n36794 , n36825 );
nor ( n36827 , n36671 , n36826 );
buf ( n36828 , n36827 );
not ( n36829 , n36828 );
nand ( n36830 , n36825 , n36670 );
buf ( n36831 , n36830 );
buf ( n36832 , n36793 );
nand ( n36833 , n36831 , n36832 );
buf ( n36834 , n36833 );
buf ( n36835 , n36834 );
nand ( n36836 , n36829 , n36835 );
buf ( n36837 , n36836 );
buf ( n36838 , n36837 );
buf ( n36839 , n36837 );
not ( n36840 , n36839 );
buf ( n36841 , n36840 );
buf ( n36842 , n36841 );
buf ( n36843 , n32972 );
not ( n36844 , n36843 );
buf ( n36845 , n36063 );
not ( n36846 , n36845 );
or ( n36847 , n36844 , n36846 );
buf ( n36848 , n36629 );
not ( n36849 , n36848 );
buf ( n36850 , n33080 );
not ( n36851 , n36850 );
and ( n36852 , n36849 , n36851 );
buf ( n36853 , n36629 );
buf ( n36854 , n33080 );
and ( n36855 , n36853 , n36854 );
nor ( n36856 , n36852 , n36855 );
buf ( n36857 , n36856 );
buf ( n36858 , n36857 );
not ( n36859 , n36858 );
buf ( n36860 , n36113 );
nand ( n36861 , n36859 , n36860 );
buf ( n36862 , n36861 );
buf ( n36863 , n36862 );
nand ( n36864 , n36847 , n36863 );
buf ( n36865 , n36864 );
buf ( n36866 , n36865 );
not ( n36867 , n36866 );
or ( n36868 , n31200 , n31203 );
buf ( n36869 , n32825 );
buf ( n36870 , n36869 );
buf ( n36871 , n36870 );
nand ( n36872 , n36868 , n36871 );
and ( n36873 , n32946 , n36872 );
not ( n36874 , n32946 );
not ( n36875 , n36872 );
and ( n36876 , n36874 , n36875 );
nor ( n36877 , n36873 , n36876 );
buf ( n36878 , n36877 );
not ( n36879 , n36878 );
not ( n36880 , n36879 );
nor ( n36881 , n31094 , n30910 );
buf ( n36882 , n36881 );
not ( n36883 , n36882 );
buf ( n36884 , n32830 );
nand ( n36885 , n36883 , n36884 );
buf ( n36886 , n36885 );
not ( n36887 , n36886 );
not ( n36888 , n36887 );
buf ( n36889 , n36868 );
not ( n36890 , n36889 );
buf ( n36891 , n32946 );
not ( n36892 , n36891 );
or ( n36893 , n36890 , n36892 );
buf ( n36894 , n36871 );
nand ( n36895 , n36893 , n36894 );
buf ( n36896 , n36895 );
not ( n36897 , n36896 );
not ( n36898 , n36897 );
or ( n36899 , n36888 , n36898 );
nand ( n36900 , n36896 , n36886 );
nand ( n36901 , n36899 , n36900 );
not ( n36902 , n36901 );
or ( n36903 , n36880 , n36902 );
not ( n36904 , n36901 );
nand ( n36905 , n36904 , n36878 );
nand ( n36906 , n36903 , n36905 );
buf ( n36907 , n36906 );
buf ( n36908 , n36907 );
buf ( n36909 , n36908 );
buf ( n36910 , n36909 );
not ( n36911 , n36910 );
buf ( n36912 , n36911 );
buf ( n36913 , n36912 );
buf ( n36914 , n36913 );
buf ( n36915 , n36914 );
buf ( n36916 , n36915 );
not ( n36917 , n36916 );
buf ( n36918 , n32957 );
buf ( n36919 , n36918 );
buf ( n36920 , n36919 );
buf ( n36921 , n36920 );
not ( n36922 , n36921 );
buf ( n36923 , n36922 );
buf ( n36924 , n36923 );
buf ( n36925 , n36924 );
buf ( n36926 , n36925 );
buf ( n36927 , n36926 );
not ( n36928 , n36927 );
buf ( n36929 , n36928 );
buf ( n36930 , n36929 );
not ( n36931 , n36930 );
buf ( n36932 , n36931 );
buf ( n36933 , n36932 );
not ( n36934 , n36933 );
buf ( n36935 , n36934 );
and ( n36936 , n36935 , n35973 );
not ( n36937 , n36935 );
and ( n36938 , n36937 , n35979 );
or ( n36939 , n36936 , n36938 );
buf ( n36940 , n36939 );
not ( n36941 , n36940 );
or ( n36942 , n36917 , n36941 );
buf ( n36943 , n36935 );
not ( n36944 , n36943 );
buf ( n36945 , n36044 );
not ( n36946 , n36945 );
or ( n36947 , n36944 , n36946 );
buf ( n36948 , n36057 );
buf ( n36949 , n36935 );
not ( n36950 , n36949 );
buf ( n36951 , n36950 );
buf ( n36952 , n36951 );
nand ( n36953 , n36948 , n36952 );
buf ( n36954 , n36953 );
buf ( n36955 , n36954 );
nand ( n36956 , n36947 , n36955 );
buf ( n36957 , n36956 );
buf ( n36958 , n36957 );
buf ( n36959 , n36906 );
buf ( n36960 , n36901 );
buf ( n36961 , n36920 );
and ( n36962 , n36960 , n36961 );
not ( n36963 , n36960 );
buf ( n36964 , n36920 );
not ( n36965 , n36964 );
buf ( n36966 , n36965 );
buf ( n36967 , n36966 );
and ( n36968 , n36963 , n36967 );
nor ( n36969 , n36962 , n36968 );
buf ( n36970 , n36969 );
buf ( n36971 , n36970 );
nand ( n36972 , n36959 , n36971 );
buf ( n36973 , n36972 );
buf ( n36974 , n36973 );
not ( n36975 , n36974 );
buf ( n36976 , n36975 );
buf ( n36977 , n36976 );
buf ( n36978 , n36977 );
buf ( n36979 , n36978 );
buf ( n36980 , n36979 );
not ( n36981 , n36980 );
buf ( n36982 , n36981 );
buf ( n36983 , n36982 );
buf ( n36984 , n36983 );
buf ( n36985 , n36984 );
buf ( n36986 , n36985 );
not ( n36987 , n36986 );
buf ( n36988 , n36987 );
buf ( n36989 , n36988 );
nand ( n36990 , n36958 , n36989 );
buf ( n36991 , n36990 );
buf ( n36992 , n36991 );
nand ( n36993 , n36942 , n36992 );
buf ( n36994 , n36993 );
buf ( n36995 , n36994 );
not ( n36996 , n36995 );
or ( n36997 , n36867 , n36996 );
buf ( n36998 , n36994 );
buf ( n36999 , n36865 );
or ( n37000 , n36998 , n36999 );
buf ( n37001 , n36939 );
buf ( n37002 , n36985 );
buf ( n37003 , n36915 );
not ( n37004 , n37003 );
buf ( n37005 , n37004 );
buf ( n37006 , n37005 );
nand ( n37007 , n37002 , n37006 );
buf ( n37008 , n37007 );
buf ( n37009 , n37008 );
and ( n37010 , n37001 , n37009 );
buf ( n37011 , n37010 );
buf ( n37012 , n37011 );
not ( n37013 , n37012 );
buf ( n37014 , n37013 );
buf ( n37015 , n37014 );
nand ( n37016 , n37000 , n37015 );
buf ( n37017 , n37016 );
buf ( n37018 , n37017 );
nand ( n37019 , n36997 , n37018 );
buf ( n37020 , n37019 );
buf ( n37021 , n37020 );
buf ( n37022 , n36649 );
not ( n37023 , n37022 );
buf ( n37024 , n36119 );
not ( n37025 , n37024 );
and ( n37026 , n37023 , n37025 );
buf ( n37027 , n36649 );
buf ( n37028 , n36119 );
and ( n37029 , n37027 , n37028 );
nor ( n37030 , n37026 , n37029 );
buf ( n37031 , n37030 );
and ( n37032 , n37031 , n36462 );
not ( n37033 , n37031 );
and ( n37034 , n37033 , n36465 );
or ( n37035 , n37032 , n37034 );
buf ( n37036 , n37035 );
xor ( n37037 , n37021 , n37036 );
buf ( n37038 , n36524 );
not ( n37039 , n37038 );
buf ( n37040 , n36533 );
not ( n37041 , n37040 );
buf ( n37042 , n36430 );
not ( n37043 , n37042 );
or ( n37044 , n37041 , n37043 );
buf ( n37045 , n36427 );
buf ( n37046 , n36578 );
nand ( n37047 , n37045 , n37046 );
buf ( n37048 , n37047 );
buf ( n37049 , n37048 );
nand ( n37050 , n37044 , n37049 );
buf ( n37051 , n37050 );
buf ( n37052 , n37051 );
not ( n37053 , n37052 );
or ( n37054 , n37039 , n37053 );
buf ( n37055 , n36584 );
buf ( n37056 , n36643 );
nand ( n37057 , n37055 , n37056 );
buf ( n37058 , n37057 );
buf ( n37059 , n37058 );
nand ( n37060 , n37054 , n37059 );
buf ( n37061 , n37060 );
buf ( n37062 , n37061 );
not ( n37063 , n37062 );
and ( n37064 , n36415 , n36456 );
buf ( n37065 , n36363 );
not ( n37066 , n37065 );
not ( n37067 , n36367 );
not ( n37068 , n35050 );
or ( n37069 , n37067 , n37068 );
not ( n37070 , n36375 );
nand ( n37071 , n37069 , n37070 );
nand ( n37072 , n35060 , n35765 );
not ( n37073 , n37072 );
and ( n37074 , n37071 , n37073 );
not ( n37075 , n37071 );
and ( n37076 , n37075 , n37072 );
nor ( n37077 , n37074 , n37076 );
buf ( n37078 , n37077 );
buf ( n37079 , n37078 );
not ( n37080 , n37079 );
buf ( n37081 , n37080 );
buf ( n37082 , n37081 );
buf ( n37083 , n37082 );
buf ( n37084 , n37083 );
buf ( n37085 , n37084 );
not ( n37086 , n37085 );
or ( n37087 , n37066 , n37086 );
buf ( n37088 , n37084 );
not ( n37089 , n37088 );
buf ( n37090 , n37089 );
buf ( n37091 , n37090 );
buf ( n37092 , n36409 );
nand ( n37093 , n37091 , n37092 );
buf ( n37094 , n37093 );
buf ( n37095 , n37094 );
nand ( n37096 , n37087 , n37095 );
buf ( n37097 , n37096 );
nor ( n37098 , n37064 , C0 );
buf ( n37099 , n37098 );
nand ( n37100 , n37063 , n37099 );
buf ( n37101 , n37100 );
buf ( n37102 , n37101 );
not ( n37103 , n37102 );
not ( n37104 , n36857 );
not ( n37105 , n36751 );
and ( n37106 , n37104 , n37105 );
buf ( n37107 , n33083 );
not ( n37108 , n37107 );
buf ( n37109 , n36568 );
not ( n37110 , n37109 );
or ( n37111 , n37108 , n37110 );
buf ( n37112 , n36574 );
buf ( n37113 , n33080 );
nand ( n37114 , n37112 , n37113 );
buf ( n37115 , n37114 );
buf ( n37116 , n37115 );
nand ( n37117 , n37111 , n37116 );
buf ( n37118 , n37117 );
and ( n37119 , n37118 , n36113 );
nor ( n37120 , n37106 , n37119 );
buf ( n37121 , n37120 );
not ( n37122 , n37121 );
buf ( n37123 , n37122 );
buf ( n37124 , n37123 );
not ( n37125 , n37124 );
buf ( n37126 , n36456 );
not ( n37127 , n37126 );
buf ( n37128 , n37097 );
not ( n37129 , n37128 );
or ( n37130 , n37127 , n37129 );
buf ( n37131 , n36363 );
not ( n37132 , n37131 );
not ( n37133 , n35018 );
not ( n37134 , n37133 );
not ( n37135 , n36367 );
or ( n37136 , n37134 , n37135 );
buf ( n37137 , n35759 );
nand ( n37138 , n37136 , n37137 );
not ( n37139 , n35047 );
nand ( n37140 , n37139 , n35762 );
not ( n37141 , n37140 );
and ( n37142 , n37138 , n37141 );
not ( n37143 , n37138 );
and ( n37144 , n37143 , n37140 );
nor ( n37145 , n37142 , n37144 );
buf ( n37146 , n37145 );
not ( n37147 , n37146 );
not ( n37148 , n37147 );
not ( n37149 , n37148 );
buf ( n37150 , n37149 );
not ( n37151 , n37150 );
or ( n37152 , n37132 , n37151 );
not ( n37153 , n37149 );
buf ( n37154 , n37153 );
buf ( n37155 , n36409 );
nand ( n37156 , n37154 , n37155 );
buf ( n37157 , n37156 );
buf ( n37158 , n37157 );
nand ( n37159 , n37152 , n37158 );
buf ( n37160 , n37159 );
buf ( n37161 , C1 );
buf ( n37162 , n37161 );
nand ( n37163 , n37130 , n37162 );
buf ( n37164 , n37163 );
buf ( n37165 , n37164 );
not ( n37166 , n37165 );
or ( n37167 , n37125 , n37166 );
buf ( n37168 , n37164 );
not ( n37169 , n37168 );
buf ( n37170 , n37169 );
buf ( n37171 , n37170 );
buf ( n37172 , n37120 );
nand ( n37173 , n37171 , n37172 );
buf ( n37174 , n37173 );
buf ( n37175 , n37174 );
buf ( n37176 , n36523 );
not ( n37177 , n37176 );
buf ( n37178 , n36533 );
not ( n37179 , n37178 );
buf ( n37180 , n36402 );
not ( n37181 , n37180 );
or ( n37182 , n37179 , n37181 );
buf ( n37183 , n36399 );
buf ( n37184 , n36578 );
nand ( n37185 , n37183 , n37184 );
buf ( n37186 , n37185 );
buf ( n37187 , n37186 );
nand ( n37188 , n37182 , n37187 );
buf ( n37189 , n37188 );
buf ( n37190 , n37189 );
not ( n37191 , n37190 );
or ( n37192 , n37177 , n37191 );
buf ( n37193 , n37051 );
buf ( n37194 , n36643 );
nand ( n37195 , n37193 , n37194 );
buf ( n37196 , n37195 );
buf ( n37197 , n37196 );
nand ( n37198 , n37192 , n37197 );
buf ( n37199 , n37198 );
buf ( n37200 , n37199 );
nand ( n37201 , n37175 , n37200 );
buf ( n37202 , n37201 );
buf ( n37203 , n37202 );
nand ( n37204 , n37167 , n37203 );
buf ( n37205 , n37204 );
buf ( n37206 , n37205 );
not ( n37207 , n37206 );
or ( n37208 , n37103 , n37207 );
buf ( n37209 , n37098 );
not ( n37210 , n37209 );
buf ( n37211 , n37061 );
nand ( n37212 , n37210 , n37211 );
buf ( n37213 , n37212 );
buf ( n37214 , n37213 );
nand ( n37215 , n37208 , n37214 );
buf ( n37216 , n37215 );
buf ( n37217 , n37216 );
and ( n37218 , n37037 , n37217 );
and ( n37219 , n37021 , n37036 );
or ( n37220 , n37218 , n37219 );
buf ( n37221 , n37220 );
not ( n37222 , n37221 );
buf ( n37223 , n36657 );
not ( n37224 , n37223 );
buf ( n37225 , n36822 );
not ( n37226 , n37225 );
or ( n37227 , n37224 , n37226 );
buf ( n37228 , n36819 );
buf ( n37229 , n36119 );
nand ( n37230 , n37228 , n37229 );
buf ( n37231 , n37230 );
buf ( n37232 , n37231 );
nand ( n37233 , n37227 , n37232 );
buf ( n37234 , n37233 );
buf ( n37235 , n37234 );
buf ( n37236 , n36663 );
and ( n37237 , n37235 , n37236 );
not ( n37238 , n37235 );
buf ( n37239 , n36666 );
and ( n37240 , n37238 , n37239 );
nor ( n37241 , n37237 , n37240 );
buf ( n37242 , n37241 );
nand ( n37243 , n37222 , n37242 );
not ( n37244 , n37243 );
buf ( n37245 , n36578 );
buf ( n37246 , n34353 );
not ( n37247 , n37246 );
buf ( n37248 , n37247 );
not ( n37249 , n37248 );
not ( n37250 , n35719 );
or ( n37251 , n37249 , n37250 );
buf ( n37252 , n34346 );
buf ( n37253 , n34350 );
nand ( n37254 , n37252 , n37253 );
buf ( n37255 , n37254 );
buf ( n37256 , n37255 );
nand ( n37257 , n37251 , n37256 );
xor ( n37258 , n35733 , n35736 );
not ( n37259 , n37258 );
and ( n37260 , n37257 , n37259 );
not ( n37261 , n37257 );
and ( n37262 , n37261 , n37258 );
nor ( n37263 , n37260 , n37262 );
not ( n37264 , n37263 );
buf ( n37265 , n37264 );
buf ( n37266 , n37265 );
not ( n37267 , n37266 );
buf ( n37268 , n37267 );
buf ( n37269 , n37268 );
not ( n37270 , n37269 );
buf ( n37271 , n37270 );
buf ( n37272 , n37271 );
and ( n37273 , n37245 , n37272 );
not ( n37274 , n37245 );
buf ( n37275 , n37268 );
and ( n37276 , n37274 , n37275 );
nor ( n37277 , n37273 , n37276 );
buf ( n37278 , n37277 );
or ( n37279 , n37278 , n36706 );
not ( n37280 , n36578 );
buf ( n37281 , n35719 );
not ( n37282 , n37281 );
buf ( n37283 , n37282 );
buf ( n37284 , n37248 );
buf ( n37285 , n37255 );
and ( n37286 , n37284 , n37285 );
buf ( n37287 , n37286 );
not ( n37288 , n37287 );
and ( n37289 , n37283 , n37288 );
not ( n37290 , n37283 );
and ( n37291 , n37290 , n37287 );
nor ( n37292 , n37289 , n37291 );
buf ( n37293 , n37292 );
buf ( n37294 , n37293 );
not ( n37295 , n37294 );
not ( n37296 , n37295 );
or ( n37297 , n37280 , n37296 );
not ( n37298 , n37295 );
nand ( n37299 , n36533 , n37298 );
nand ( n37300 , n37297 , n37299 );
not ( n37301 , n37300 );
nand ( n37302 , n37301 , n36523 );
nand ( n37303 , n37279 , n37302 );
not ( n37304 , n37303 );
not ( n37305 , n37304 );
buf ( n37306 , n32671 );
buf ( n37307 , n32700 );
not ( n37308 , n37307 );
buf ( n37309 , n32667 );
nand ( n37310 , n37308 , n37309 );
buf ( n37311 , n37310 );
buf ( n37312 , n37311 );
and ( n37313 , n37306 , n37312 );
buf ( n37314 , n37313 );
not ( n37315 , n37314 );
not ( n37316 , n37315 );
not ( n37317 , n32706 );
not ( n37318 , n32741 );
or ( n37319 , n37317 , n37318 );
not ( n37320 , n32644 );
nand ( n37321 , n37319 , n37320 );
not ( n37322 , n37321 );
not ( n37323 , n37322 );
or ( n37324 , n37316 , n37323 );
nand ( n37325 , n37321 , n37314 );
nand ( n37326 , n37324 , n37325 );
not ( n37327 , n37326 );
not ( n37328 , n37327 );
buf ( n37329 , n37328 );
not ( n37330 , n37329 );
not ( n37331 , n37330 );
not ( n37332 , n35971 );
or ( n37333 , n37331 , n37332 );
or ( n37334 , n35971 , n37330 );
nand ( n37335 , n37333 , n37334 );
not ( n37336 , n37326 );
buf ( n37337 , n37336 );
not ( n37338 , n37337 );
buf ( n37339 , n32615 );
buf ( n37340 , n37339 );
buf ( n37341 , n37340 );
buf ( n37342 , n37341 );
buf ( n37343 , n32635 );
buf ( n37344 , n37343 );
buf ( n37345 , n37344 );
buf ( n37346 , n37345 );
or ( n37347 , n37342 , n37346 );
buf ( n37348 , n37347 );
not ( n37349 , n37348 );
not ( n37350 , n32741 );
or ( n37351 , n37349 , n37350 );
buf ( n37352 , n37341 );
buf ( n37353 , n37345 );
nand ( n37354 , n37352 , n37353 );
buf ( n37355 , n37354 );
nand ( n37356 , n37351 , n37355 );
buf ( n37357 , n32612 );
not ( n37358 , n37357 );
buf ( n37359 , n32573 );
buf ( n37360 , n32609 );
nand ( n37361 , n37359 , n37360 );
buf ( n37362 , n37361 );
buf ( n37363 , n37362 );
nand ( n37364 , n37358 , n37363 );
buf ( n37365 , n37364 );
xnor ( n37366 , n37356 , n37365 );
buf ( n37367 , n37366 );
not ( n37368 , n37367 );
buf ( n37369 , n37368 );
buf ( n37370 , n37369 );
nand ( n37371 , n37338 , n37370 );
buf ( n37372 , n37371 );
and ( n37373 , n37348 , n37355 );
not ( n37374 , n37373 );
not ( n37375 , n32741 );
not ( n37376 , n37375 );
or ( n37377 , n37374 , n37376 );
not ( n37378 , n37375 );
xnor ( n37379 , n37341 , n37345 );
nand ( n37380 , n37378 , n37379 );
nand ( n37381 , n37377 , n37380 );
not ( n37382 , n37381 );
and ( n37383 , n37382 , n37366 );
not ( n37384 , n37382 );
not ( n37385 , n37366 );
and ( n37386 , n37384 , n37385 );
nor ( n37387 , n37383 , n37386 );
buf ( n37388 , n37336 );
xnor ( n37389 , n37356 , n37365 );
buf ( n37390 , n37389 );
nand ( n37391 , n37388 , n37390 );
buf ( n37392 , n37391 );
nand ( n37393 , n37372 , n37387 , n37392 );
not ( n37394 , n37393 );
buf ( n37395 , n37394 );
buf ( n37396 , n37395 );
buf ( n37397 , n37396 );
buf ( n37398 , n37397 );
buf ( n37399 , n37398 );
buf ( n37400 , n37399 );
buf ( n37401 , n37400 );
buf ( n37402 , n37401 );
buf ( n37403 , n37402 );
buf ( n37404 , n37403 );
not ( n37405 , n37404 );
buf ( n37406 , n37405 );
not ( n37407 , n37387 );
buf ( n37408 , n37407 );
buf ( n37409 , n37408 );
buf ( n37410 , n37409 );
buf ( n37411 , n37410 );
buf ( n37412 , n37411 );
buf ( n37413 , n37412 );
buf ( n37414 , n37413 );
not ( n37415 , n37414 );
buf ( n37416 , n37415 );
nand ( n37417 , n37406 , n37416 );
and ( n37418 , n37335 , n37417 );
buf ( n37419 , n37336 );
not ( n37420 , n37419 );
buf ( n37421 , n37420 );
not ( n37422 , n37421 );
buf ( n37423 , n32671 );
not ( n37424 , n37423 );
not ( n37425 , n37321 );
or ( n37426 , n37424 , n37425 );
nand ( n37427 , n37426 , n37311 );
nand ( n37428 , n32691 , n32692 );
nand ( n37429 , n37428 , n32707 );
not ( n37430 , n37429 );
and ( n37431 , n37427 , n37430 );
not ( n37432 , n37427 );
and ( n37433 , n37432 , n37429 );
nor ( n37434 , n37431 , n37433 );
not ( n37435 , n37434 );
or ( n37436 , n37422 , n37435 );
not ( n37437 , n37434 );
nand ( n37438 , n37437 , n37336 );
nand ( n37439 , n37436 , n37438 );
buf ( n37440 , n37439 );
buf ( n37441 , n37440 );
not ( n37442 , n37441 );
buf ( n37443 , n37442 );
buf ( n37444 , n37443 );
not ( n37445 , n37444 );
buf ( n37446 , n37445 );
buf ( n37447 , n37446 );
not ( n37448 , n37447 );
buf ( n37449 , n37448 );
buf ( n37450 , n37449 );
not ( n37451 , n37450 );
buf ( n37452 , n37451 );
not ( n37453 , n37452 );
or ( n37454 , n32086 , n32309 );
buf ( n37455 , n37454 );
buf ( n37456 , n32762 );
buf ( n37457 , n37456 );
nand ( n37458 , n37455 , n37457 );
buf ( n37459 , n37458 );
not ( n37460 , n37459 );
buf ( n37461 , n36231 );
buf ( n37462 , n37461 );
buf ( n37463 , n37462 );
not ( n37464 , n37463 );
or ( n37465 , n37460 , n37464 );
buf ( n37466 , n36231 );
buf ( n37467 , n37459 );
or ( n37468 , n37466 , n37467 );
buf ( n37469 , n37468 );
nand ( n37470 , n37465 , n37469 );
not ( n37471 , n37470 );
buf ( n37472 , n37471 );
not ( n37473 , n37472 );
buf ( n37474 , n37473 );
not ( n37475 , n37474 );
not ( n37476 , n37475 );
and ( n37477 , n37476 , n36041 );
not ( n37478 , n37476 );
buf ( n37479 , n36041 );
not ( n37480 , n37479 );
buf ( n37481 , n37480 );
and ( n37482 , n37478 , n37481 );
or ( n37483 , n37477 , n37482 );
not ( n37484 , n37483 );
or ( n37485 , n37453 , n37484 );
buf ( n37486 , n37476 );
not ( n37487 , n37486 );
buf ( n37488 , n36620 );
not ( n37489 , n37488 );
or ( n37490 , n37487 , n37489 );
buf ( n37491 , n36617 );
buf ( n37492 , n37475 );
nand ( n37493 , n37491 , n37492 );
buf ( n37494 , n37493 );
buf ( n37495 , n37494 );
nand ( n37496 , n37490 , n37495 );
buf ( n37497 , n37496 );
buf ( n37498 , n37497 );
not ( n37499 , n37437 );
not ( n37500 , n37499 );
buf ( n37501 , n37470 );
not ( n37502 , n37501 );
not ( n37503 , n37502 );
or ( n37504 , n37500 , n37503 );
nand ( n37505 , n37501 , n37437 );
nand ( n37506 , n37504 , n37505 );
buf ( n37507 , n37439 );
not ( n37508 , n37507 );
buf ( n37509 , n37508 );
nand ( n37510 , n37506 , n37509 );
buf ( n37511 , n37510 );
buf ( n37512 , n37511 );
buf ( n37513 , n37512 );
buf ( n37514 , n37513 );
buf ( n37515 , n37514 );
not ( n37516 , n37515 );
buf ( n37517 , n37516 );
buf ( n37518 , n37517 );
nand ( n37519 , n37498 , n37518 );
buf ( n37520 , n37519 );
nand ( n37521 , n37485 , n37520 );
xnor ( n37522 , n37418 , n37521 );
not ( n37523 , n37522 );
or ( n37524 , n37305 , n37523 );
not ( n37525 , n37521 );
nand ( n37526 , n37418 , n37525 );
not ( n37527 , n37526 );
not ( n37528 , n37418 );
and ( n37529 , n37521 , n37528 );
or ( n37530 , n37527 , n37529 );
nand ( n37531 , n37530 , n37303 );
nand ( n37532 , n37524 , n37531 );
not ( n37533 , n37532 );
buf ( n37534 , n37517 );
not ( n37535 , n37534 );
buf ( n37536 , n37476 );
not ( n37537 , n37536 );
buf ( n37538 , n36565 );
not ( n37539 , n37538 );
or ( n37540 , n37537 , n37539 );
buf ( n37541 , n36565 );
not ( n37542 , n37541 );
buf ( n37543 , n37542 );
buf ( n37544 , n37543 );
not ( n37545 , n37476 );
buf ( n37546 , n37545 );
nand ( n37547 , n37544 , n37546 );
buf ( n37548 , n37547 );
buf ( n37549 , n37548 );
nand ( n37550 , n37540 , n37549 );
buf ( n37551 , n37550 );
buf ( n37552 , n37551 );
not ( n37553 , n37552 );
or ( n37554 , n37535 , n37553 );
buf ( n37555 , n37497 );
buf ( n37556 , n37452 );
nand ( n37557 , n37555 , n37556 );
buf ( n37558 , n37557 );
buf ( n37559 , n37558 );
nand ( n37560 , n37554 , n37559 );
buf ( n37561 , n37560 );
buf ( n37562 , n37561 );
not ( n37563 , n36453 );
buf ( n37564 , n36360 );
not ( n37565 , n37564 );
buf ( n37566 , n35549 );
buf ( n37567 , n35585 );
nor ( n37568 , n37566 , n37567 );
buf ( n37569 , n37568 );
buf ( n37570 , n37569 );
not ( n37571 , n37570 );
buf ( n37572 , n35588 );
buf ( n37573 , n37572 );
buf ( n37574 , n37573 );
buf ( n37575 , n37574 );
nand ( n37576 , n37571 , n37575 );
buf ( n37577 , n37576 );
buf ( n37578 , n37577 );
not ( n37579 , n37578 );
buf ( n37580 , n37579 );
nand ( n37581 , n35715 , n35667 );
and ( n37582 , n35711 , n35708 , n37581 );
or ( n37583 , n37580 , n37582 );
nand ( n37584 , n37580 , n37582 );
nand ( n37585 , n37583 , n37584 );
buf ( n37586 , n37585 );
buf ( n37587 , n37586 );
not ( n37588 , n37587 );
buf ( n37589 , n37588 );
buf ( n37590 , n37589 );
not ( n37591 , n37590 );
or ( n37592 , n37565 , n37591 );
buf ( n37593 , n37586 );
not ( n37594 , n37593 );
buf ( n37595 , n37594 );
buf ( n37596 , n37595 );
not ( n37597 , n37596 );
buf ( n37598 , n37597 );
buf ( n37599 , n37598 );
buf ( n37600 , n36360 );
not ( n37601 , n37600 );
buf ( n37602 , n37601 );
buf ( n37603 , n37602 );
nand ( n37604 , n37599 , n37603 );
buf ( n37605 , n37604 );
buf ( n37606 , n37605 );
nand ( n37607 , n37592 , n37606 );
buf ( n37608 , n37607 );
not ( n37609 , n37608 );
or ( n37610 , n37563 , n37609 );
buf ( n37611 , n36360 );
not ( n37612 , n37611 );
buf ( n37613 , n35715 );
not ( n37614 , n37613 );
buf ( n37615 , n35670 );
nand ( n37616 , n37614 , n37615 );
buf ( n37617 , n37616 );
and ( n37618 , n37617 , n35716 );
buf ( n37619 , n35657 );
buf ( n37620 , n37619 );
buf ( n37621 , n37620 );
nand ( n37622 , n37621 , n35707 );
and ( n37623 , n37618 , n37622 );
not ( n37624 , n37623 );
not ( n37625 , n29278 );
buf ( n37626 , n37621 );
buf ( n37627 , n30176 );
nand ( n37628 , n37626 , n37627 );
buf ( n37629 , n37628 );
not ( n37630 , n37629 );
nand ( n37631 , n37625 , n37630 , n29881 );
buf ( n37632 , n37631 );
not ( n37633 , n37632 );
or ( n37634 , n37624 , n37633 );
not ( n37635 , n37622 );
not ( n37636 , n37631 );
or ( n37637 , n37635 , n37636 );
not ( n37638 , n37618 );
nand ( n37639 , n37637 , n37638 );
nand ( n37640 , n37634 , n37639 );
buf ( n37641 , n37640 );
not ( n37642 , n37641 );
buf ( n37643 , n37642 );
not ( n37644 , n37643 );
or ( n37645 , n37612 , n37644 );
buf ( n37646 , n37641 );
buf ( n37647 , n36357 );
not ( n37648 , n37647 );
buf ( n37649 , n37648 );
buf ( n37650 , n37649 );
nand ( n37651 , n37646 , n37650 );
buf ( n37652 , n37651 );
buf ( n37653 , n37652 );
nand ( n37654 , n37645 , n37653 );
buf ( n37655 , n37654 );
buf ( n37656 , C1 );
nand ( n37657 , n37610 , n37656 );
buf ( n37658 , n37657 );
buf ( n37659 , n36643 );
not ( n37660 , n37659 );
not ( n37661 , n36533 );
buf ( n37662 , n35624 );
or ( n37663 , n35297 , n35456 );
nand ( n37664 , n37662 , n37663 );
or ( n37665 , n37664 , n37582 );
buf ( n37666 , n35597 );
nand ( n37667 , n37666 , n37663 );
buf ( n37668 , n35606 );
nand ( n37669 , n37667 , n37668 );
not ( n37670 , n37669 );
nand ( n37671 , n37665 , n37670 );
buf ( n37672 , n35603 );
buf ( n37673 , n35613 );
nor ( n37674 , n37672 , n37673 );
not ( n37675 , n37674 );
nor ( n37676 , n37671 , n37675 );
buf ( n37677 , n37676 );
not ( n37678 , n37677 );
not ( n37679 , n37674 );
nand ( n37680 , n37679 , n37671 );
buf ( n37681 , n37680 );
nand ( n37682 , n37678 , n37681 );
buf ( n37683 , n37682 );
buf ( n37684 , n37683 );
buf ( n37685 , n37684 );
buf ( n37686 , n37685 );
buf ( n37687 , n37686 );
not ( n37688 , n37687 );
buf ( n37689 , n37688 );
buf ( n37690 , n37689 );
not ( n37691 , n37690 );
buf ( n37692 , n37691 );
buf ( n37693 , n37692 );
buf ( n37694 , n37693 );
buf ( n37695 , n37694 );
buf ( n37696 , n37695 );
not ( n37697 , n37696 );
buf ( n37698 , n37697 );
not ( n37699 , n37698 );
or ( n37700 , n37661 , n37699 );
buf ( n37701 , n37676 );
not ( n37702 , n37701 );
buf ( n37703 , n37680 );
nand ( n37704 , n37702 , n37703 );
buf ( n37705 , n37704 );
buf ( n37706 , n37705 );
not ( n37707 , n37706 );
buf ( n37708 , n37707 );
buf ( n37709 , n37708 );
not ( n37710 , n37709 );
buf ( n37711 , n37710 );
buf ( n37712 , n37711 );
not ( n37713 , n37712 );
buf ( n37714 , n37713 );
buf ( n37715 , n37714 );
buf ( n37716 , n37715 );
buf ( n37717 , n37716 );
buf ( n37718 , n37717 );
buf ( n37719 , n36533 );
or ( n37720 , n37718 , n37719 );
buf ( n37721 , n37720 );
nand ( n37722 , n37700 , n37721 );
buf ( n37723 , n37722 );
not ( n37724 , n37723 );
or ( n37725 , n37660 , n37724 );
buf ( n37726 , n36523 );
buf ( n37727 , n36533 );
not ( n37728 , n37727 );
and ( n37729 , n37668 , n37663 );
not ( n37730 , n37729 );
not ( n37731 , n37662 );
nand ( n37732 , n35711 , n35708 , n37581 );
not ( n37733 , n37732 );
or ( n37734 , n37731 , n37733 );
not ( n37735 , n37666 );
nand ( n37736 , n37734 , n37735 );
not ( n37737 , n37736 );
not ( n37738 , n37737 );
or ( n37739 , n37730 , n37738 );
not ( n37740 , n37729 );
nand ( n37741 , n37740 , n37736 );
nand ( n37742 , n37739 , n37741 );
buf ( n37743 , n37742 );
not ( n37744 , n37743 );
buf ( n37745 , n37744 );
buf ( n37746 , n37745 );
buf ( n37747 , n37746 );
not ( n37748 , n37747 );
or ( n37749 , n37728 , n37748 );
not ( n37750 , n37746 );
buf ( n37751 , n37750 );
buf ( n37752 , n36530 );
nand ( n37753 , n37751 , n37752 );
buf ( n37754 , n37753 );
buf ( n37755 , n37754 );
nand ( n37756 , n37749 , n37755 );
buf ( n37757 , n37756 );
buf ( n37758 , n37757 );
nand ( n37759 , n37726 , n37758 );
buf ( n37760 , n37759 );
buf ( n37761 , n37760 );
nand ( n37762 , n37725 , n37761 );
buf ( n37763 , n37762 );
buf ( n37764 , n37763 );
xor ( n37765 , n37658 , n37764 );
not ( n37766 , n36456 );
buf ( n37767 , n36360 );
not ( n37768 , n37767 );
not ( n37769 , n37569 );
not ( n37770 , n37769 );
not ( n37771 , n37732 );
or ( n37772 , n37770 , n37771 );
nand ( n37773 , n37772 , n37574 );
not ( n37774 , n35594 );
nand ( n37775 , n35542 , n35466 );
nand ( n37776 , n37774 , n37775 );
not ( n37777 , n37776 );
and ( n37778 , n37773 , n37777 );
not ( n37779 , n37773 );
and ( n37780 , n37779 , n37776 );
nor ( n37781 , n37778 , n37780 );
not ( n37782 , n37781 );
not ( n37783 , n37782 );
buf ( n37784 , n37783 );
not ( n37785 , n37784 );
buf ( n37786 , n37785 );
buf ( n37787 , n37786 );
not ( n37788 , n37787 );
or ( n37789 , n37768 , n37788 );
buf ( n37790 , n37786 );
not ( n37791 , n37790 );
buf ( n37792 , n37791 );
buf ( n37793 , n37792 );
buf ( n37794 , n37602 );
nand ( n37795 , n37793 , n37794 );
buf ( n37796 , n37795 );
buf ( n37797 , n37796 );
nand ( n37798 , n37789 , n37797 );
buf ( n37799 , n37798 );
not ( n37800 , n37799 );
or ( n37801 , n37766 , n37800 );
buf ( n37802 , C1 );
nand ( n37803 , n37801 , n37802 );
buf ( n37804 , n37803 );
and ( n37805 , n37765 , n37804 );
and ( n37806 , n37658 , n37764 );
or ( n37807 , n37805 , n37806 );
buf ( n37808 , n37807 );
buf ( n37809 , n37808 );
buf ( n37810 , n37809 );
xor ( n37811 , n37562 , n37810 );
not ( n37812 , n37454 );
not ( n37813 , n36231 );
or ( n37814 , n37812 , n37813 );
nand ( n37815 , n37814 , n37456 );
buf ( n37816 , n32751 );
buf ( n37817 , n32755 );
or ( n37818 , n37816 , n37817 );
buf ( n37819 , n37818 );
buf ( n37820 , n37819 );
buf ( n37821 , n32767 );
nand ( n37822 , n37820 , n37821 );
buf ( n37823 , n37822 );
and ( n37824 , n37815 , n37823 );
not ( n37825 , n37815 );
not ( n37826 , n37823 );
and ( n37827 , n37825 , n37826 );
nor ( n37828 , n37824 , n37827 );
not ( n37829 , n37828 );
not ( n37830 , n37829 );
nor ( n37831 , n32336 , n32330 );
buf ( n37832 , n37831 );
buf ( n37833 , n37832 );
buf ( n37834 , n37833 );
buf ( n37835 , n37834 );
not ( n37836 , n37835 );
buf ( n37837 , n32793 );
nand ( n37838 , n37836 , n37837 );
buf ( n37839 , n37838 );
not ( n37840 , n37839 );
not ( n37841 , n37840 );
not ( n37842 , n32311 );
not ( n37843 , n37842 );
not ( n37844 , n37843 );
not ( n37845 , n36231 );
or ( n37846 , n37844 , n37845 );
buf ( n37847 , n32768 );
not ( n37848 , n37847 );
buf ( n37849 , n37848 );
nand ( n37850 , n37846 , n37849 );
not ( n37851 , n37850 );
not ( n37852 , n37851 );
or ( n37853 , n37841 , n37852 );
buf ( n37854 , n37850 );
buf ( n37855 , n37839 );
nand ( n37856 , n37854 , n37855 );
buf ( n37857 , n37856 );
nand ( n37858 , n37853 , n37857 );
not ( n37859 , n37858 );
not ( n37860 , n37859 );
or ( n37861 , n37830 , n37860 );
nand ( n37862 , n37858 , n37828 );
nand ( n37863 , n37861 , n37862 );
not ( n37864 , n37828 );
not ( n37865 , n37470 );
or ( n37866 , n37864 , n37865 );
nand ( n37867 , n37471 , n37829 );
nand ( n37868 , n37866 , n37867 );
not ( n37869 , n37868 );
nand ( n37870 , n37863 , n37869 );
not ( n37871 , n37870 );
buf ( n37872 , n37871 );
buf ( n37873 , n37872 );
buf ( n37874 , n37873 );
buf ( n37875 , n37874 );
buf ( n37876 , n37875 );
not ( n37877 , n37876 );
or ( n37878 , n37850 , n37839 );
nand ( n37879 , n37878 , n37857 );
not ( n37880 , n37879 );
not ( n37881 , n37880 );
buf ( n37882 , n37881 );
buf ( n37883 , n37882 );
not ( n37884 , n37883 );
buf ( n37885 , n36399 );
not ( n37886 , n37885 );
buf ( n37887 , n37886 );
buf ( n37888 , n37887 );
not ( n37889 , n37888 );
or ( n37890 , n37884 , n37889 );
buf ( n37891 , n36399 );
not ( n37892 , n37880 );
not ( n37893 , n37892 );
buf ( n37894 , n37893 );
nand ( n37895 , n37891 , n37894 );
buf ( n37896 , n37895 );
buf ( n37897 , n37896 );
nand ( n37898 , n37890 , n37897 );
buf ( n37899 , n37898 );
buf ( n37900 , n37899 );
not ( n37901 , n37900 );
or ( n37902 , n37877 , n37901 );
buf ( n37903 , n37882 );
not ( n37904 , n37903 );
buf ( n37905 , n36430 );
not ( n37906 , n37905 );
or ( n37907 , n37904 , n37906 );
buf ( n37908 , n36427 );
buf ( n37909 , n37893 );
nand ( n37910 , n37908 , n37909 );
buf ( n37911 , n37910 );
buf ( n37912 , n37911 );
nand ( n37913 , n37907 , n37912 );
buf ( n37914 , n37913 );
buf ( n37915 , n37914 );
buf ( n37916 , n37869 );
buf ( n37917 , n37916 );
not ( n37918 , n37917 );
buf ( n37919 , n37918 );
buf ( n37920 , n37919 );
buf ( n37921 , n37920 );
buf ( n37922 , n37921 );
buf ( n37923 , n37922 );
nand ( n37924 , n37915 , n37923 );
buf ( n37925 , n37924 );
buf ( n37926 , n37925 );
nand ( n37927 , n37902 , n37926 );
buf ( n37928 , n37927 );
buf ( n37929 , n37928 );
and ( n37930 , n37811 , n37929 );
and ( n37931 , n37562 , n37810 );
or ( n37932 , n37930 , n37931 );
buf ( n37933 , n37932 );
xor ( n37934 , n37533 , n37933 );
buf ( n37935 , n36915 );
not ( n37936 , n37935 );
buf ( n37937 , n36935 );
not ( n37938 , n37937 );
buf ( n37939 , n37149 );
not ( n37940 , n37939 );
or ( n37941 , n37938 , n37940 );
buf ( n37942 , n37148 );
buf ( n37943 , n36951 );
nand ( n37944 , n37942 , n37943 );
buf ( n37945 , n37944 );
buf ( n37946 , n37945 );
nand ( n37947 , n37941 , n37946 );
buf ( n37948 , n37947 );
buf ( n37949 , n37948 );
not ( n37950 , n37949 );
or ( n37951 , n37936 , n37950 );
buf ( n37952 , n36935 );
not ( n37953 , n37952 );
buf ( n37954 , n37133 );
buf ( n37955 , n35759 );
nand ( n37956 , n37954 , n37955 );
buf ( n37957 , n37956 );
buf ( n37958 , n37957 );
not ( n37959 , n37958 );
buf ( n37960 , n37959 );
not ( n37961 , n37960 );
not ( n37962 , n36370 );
or ( n37963 , n37961 , n37962 );
buf ( n37964 , n36367 );
buf ( n37965 , n37957 );
nand ( n37966 , n37964 , n37965 );
buf ( n37967 , n37966 );
nand ( n37968 , n37963 , n37967 );
not ( n37969 , n37968 );
buf ( n37970 , n37969 );
buf ( n37971 , n37970 );
buf ( n37972 , n37971 );
not ( n37973 , n37972 );
or ( n37974 , n37953 , n37973 );
buf ( n37975 , n37971 );
not ( n37976 , n37975 );
buf ( n37977 , n37976 );
buf ( n37978 , n37977 );
buf ( n37979 , n36951 );
nand ( n37980 , n37978 , n37979 );
buf ( n37981 , n37980 );
buf ( n37982 , n37981 );
nand ( n37983 , n37974 , n37982 );
buf ( n37984 , n37983 );
buf ( n37985 , n37984 );
buf ( n37986 , n36988 );
nand ( n37987 , n37985 , n37986 );
buf ( n37988 , n37987 );
buf ( n37989 , n37988 );
nand ( n37990 , n37951 , n37989 );
buf ( n37991 , n37990 );
buf ( n37992 , n37991 );
buf ( n37993 , n37875 );
not ( n37994 , n37993 );
buf ( n37995 , n37914 );
not ( n37996 , n37995 );
or ( n37997 , n37994 , n37996 );
buf ( n37998 , n37882 );
not ( n37999 , n37998 );
buf ( n38000 , n36565 );
not ( n38001 , n38000 );
or ( n38002 , n37999 , n38001 );
buf ( n38003 , n37543 );
buf ( n38004 , n37893 );
nand ( n38005 , n38003 , n38004 );
buf ( n38006 , n38005 );
buf ( n38007 , n38006 );
nand ( n38008 , n38002 , n38007 );
buf ( n38009 , n38008 );
buf ( n38010 , n38009 );
buf ( n38011 , n37922 );
nand ( n38012 , n38010 , n38011 );
buf ( n38013 , n38012 );
buf ( n38014 , n38013 );
nand ( n38015 , n37997 , n38014 );
buf ( n38016 , n38015 );
buf ( n38017 , n38016 );
xor ( n38018 , n37992 , n38017 );
buf ( n38019 , n37858 );
nor ( n38020 , n37834 , n37842 );
nand ( n38021 , n38020 , n37463 );
not ( n38022 , n38021 );
or ( n38023 , n37849 , n37834 );
buf ( n38024 , n32793 );
nand ( n38025 , n38023 , n38024 );
buf ( n38026 , n32800 );
buf ( n38027 , n32773 );
buf ( n38028 , n32780 );
nand ( n38029 , n38027 , n38028 );
buf ( n38030 , n38029 );
buf ( n38031 , n38030 );
nand ( n38032 , n38026 , n38031 );
buf ( n38033 , n38032 );
nor ( n38034 , n38025 , n38033 );
not ( n38035 , n38034 );
or ( n38036 , n38022 , n38035 );
not ( n38037 , n38025 );
not ( n38038 , n38037 );
buf ( n38039 , n38033 );
not ( n38040 , n38039 );
buf ( n38041 , n38040 );
not ( n38042 , n38041 );
and ( n38043 , n38038 , n38042 );
not ( n38044 , n38020 );
nor ( n38045 , n38044 , n38041 );
and ( n38046 , n37463 , n38045 );
nor ( n38047 , n38043 , n38046 );
nand ( n38048 , n38036 , n38047 );
buf ( n38049 , n38048 );
xnor ( n38050 , n38019 , n38049 );
buf ( n38051 , n38050 );
buf ( n38052 , n38051 );
not ( n38053 , n38052 );
buf ( n38054 , n38053 );
buf ( n38055 , n38054 );
not ( n38056 , n38055 );
buf ( n38057 , n38056 );
buf ( n38058 , n38057 );
not ( n38059 , n38058 );
buf ( n38060 , n38059 );
buf ( n38061 , n38060 );
buf ( n38062 , n38061 );
buf ( n38063 , n38062 );
buf ( n38064 , n38063 );
not ( n38065 , n38064 );
buf ( n38066 , n36878 );
buf ( n38067 , n38066 );
buf ( n38068 , n38067 );
buf ( n38069 , n38068 );
buf ( n38070 , n38069 );
buf ( n38071 , n38070 );
buf ( n38072 , n38071 );
not ( n38073 , n38072 );
buf ( n38074 , n38073 );
buf ( n38075 , n38074 );
not ( n38076 , n38075 );
buf ( n38077 , n37887 );
not ( n38078 , n38077 );
or ( n38079 , n38076 , n38078 );
buf ( n38080 , n36399 );
buf ( n38081 , n38074 );
not ( n38082 , n38081 );
buf ( n38083 , n38082 );
buf ( n38084 , n38083 );
nand ( n38085 , n38080 , n38084 );
buf ( n38086 , n38085 );
buf ( n38087 , n38086 );
nand ( n38088 , n38079 , n38087 );
buf ( n38089 , n38088 );
buf ( n38090 , n38089 );
not ( n38091 , n38090 );
or ( n38092 , n38065 , n38091 );
buf ( n38093 , n38074 );
not ( n38094 , n38093 );
buf ( n38095 , n37084 );
not ( n38096 , n38095 );
or ( n38097 , n38094 , n38096 );
not ( n38098 , n37078 );
buf ( n38099 , n38098 );
not ( n38100 , n38099 );
buf ( n38101 , n38083 );
nand ( n38102 , n38100 , n38101 );
buf ( n38103 , n38102 );
buf ( n38104 , n38103 );
nand ( n38105 , n38097 , n38104 );
buf ( n38106 , n38105 );
buf ( n38107 , n38106 );
not ( n38108 , n36878 );
buf ( n38109 , n38108 );
buf ( n38110 , n38048 );
buf ( n38111 , n38110 );
buf ( n38112 , n38111 );
buf ( n38113 , n38112 );
nand ( n38114 , n38109 , n38113 );
buf ( n38115 , n38114 );
buf ( n38116 , n38115 );
buf ( n38117 , n38051 );
buf ( n38118 , n38112 );
not ( n38119 , n38118 );
buf ( n38120 , n38119 );
nand ( n38121 , n38120 , n36878 );
buf ( n38122 , n38121 );
nand ( n38123 , n38116 , n38117 , n38122 );
buf ( n38124 , n38123 );
buf ( n38125 , n38124 );
buf ( n38126 , n38125 );
buf ( n38127 , n38126 );
buf ( n38128 , n38127 );
not ( n38129 , n38128 );
buf ( n38130 , n38129 );
buf ( n38131 , n38130 );
buf ( n38132 , n38131 );
buf ( n38133 , n38132 );
buf ( n38134 , n38133 );
nand ( n38135 , n38107 , n38134 );
buf ( n38136 , n38135 );
buf ( n38137 , n38136 );
nand ( n38138 , n38092 , n38137 );
buf ( n38139 , n38138 );
buf ( n38140 , n38139 );
xnor ( n38141 , n38018 , n38140 );
buf ( n38142 , n38141 );
buf ( n38143 , n38142 );
not ( n38144 , n38143 );
buf ( n38145 , n38144 );
xor ( n38146 , n37934 , n38145 );
buf ( n38147 , n38146 );
buf ( n38148 , n37416 );
not ( n38149 , n38148 );
buf ( n38150 , n38149 );
buf ( n38151 , n38150 );
not ( n38152 , n38151 );
buf ( n38153 , n37330 );
not ( n38154 , n38153 );
buf ( n38155 , n36041 );
not ( n38156 , n38155 );
or ( n38157 , n38154 , n38156 );
buf ( n38158 , n36038 );
buf ( n38159 , n37329 );
nand ( n38160 , n38158 , n38159 );
buf ( n38161 , n38160 );
buf ( n38162 , n38161 );
nand ( n38163 , n38157 , n38162 );
buf ( n38164 , n38163 );
buf ( n38165 , n38164 );
not ( n38166 , n38165 );
or ( n38167 , n38152 , n38166 );
buf ( n38168 , n37406 );
not ( n38169 , n38168 );
buf ( n38170 , n37330 );
not ( n38171 , n38170 );
buf ( n38172 , n36620 );
not ( n38173 , n38172 );
or ( n38174 , n38171 , n38173 );
buf ( n38175 , n36617 );
buf ( n38176 , n37329 );
nand ( n38177 , n38175 , n38176 );
buf ( n38178 , n38177 );
buf ( n38179 , n38178 );
nand ( n38180 , n38174 , n38179 );
buf ( n38181 , n38180 );
buf ( n38182 , n38181 );
nand ( n38183 , n38169 , n38182 );
buf ( n38184 , n38183 );
buf ( n38185 , n38184 );
nand ( n38186 , n38167 , n38185 );
buf ( n38187 , n38186 );
buf ( n38188 , n38187 );
buf ( n38189 , n36915 );
not ( n38190 , n38189 );
buf ( n38191 , n36935 );
not ( n38192 , n38191 );
buf ( n38193 , n34354 );
buf ( n38194 , n38193 );
buf ( n38195 , n38194 );
not ( n38196 , n38195 );
not ( n38197 , n35617 );
or ( n38198 , n38196 , n38197 );
buf ( n38199 , n35738 );
buf ( n38200 , n38199 );
buf ( n38201 , n38200 );
nand ( n38202 , n38198 , n38201 );
buf ( n38203 , n35746 );
nand ( n38204 , n38202 , n38203 );
buf ( n38205 , n35718 );
buf ( n38206 , n34520 );
or ( n38207 , n38205 , n38206 );
buf ( n38208 , n38207 );
buf ( n38209 , n35740 );
nand ( n38210 , n38209 , n35749 );
and ( n38211 , n38210 , n35741 );
nand ( n38212 , n38204 , n38208 , n38211 );
or ( n38213 , n38204 , n38210 );
nor ( n38214 , n38208 , n38210 );
not ( n38215 , n38214 );
or ( n38216 , n38210 , n35741 );
nand ( n38217 , n38212 , n38213 , n38215 , n38216 );
buf ( n38218 , n38217 );
buf ( n38219 , n38218 );
buf ( n38220 , n38219 );
buf ( n38221 , n38220 );
buf ( n38222 , n38221 );
not ( n38223 , n38222 );
or ( n38224 , n38192 , n38223 );
buf ( n38225 , n38221 );
not ( n38226 , n38225 );
buf ( n38227 , n38226 );
buf ( n38228 , n38227 );
buf ( n38229 , n36951 );
nand ( n38230 , n38228 , n38229 );
buf ( n38231 , n38230 );
buf ( n38232 , n38231 );
nand ( n38233 , n38224 , n38232 );
buf ( n38234 , n38233 );
buf ( n38235 , n38234 );
not ( n38236 , n38235 );
or ( n38237 , n38190 , n38236 );
and ( n38238 , n38203 , n35741 );
not ( n38239 , n38195 );
not ( n38240 , n35719 );
or ( n38241 , n38239 , n38240 );
nand ( n38242 , n38241 , n38201 );
xor ( n38243 , n38238 , n38242 );
buf ( n38244 , n38243 );
buf ( n38245 , n38244 );
buf ( n38246 , n38245 );
buf ( n38247 , n38246 );
buf ( n38248 , n38247 );
not ( n38249 , n38248 );
buf ( n38250 , n38249 );
nand ( n38251 , n38250 , n36935 );
nand ( n38252 , n38247 , n36951 );
nand ( n38253 , n38251 , n38252 );
buf ( n38254 , n38253 );
buf ( n38255 , n36988 );
nand ( n38256 , n38254 , n38255 );
buf ( n38257 , n38256 );
buf ( n38258 , n38257 );
nand ( n38259 , n38237 , n38258 );
buf ( n38260 , n38259 );
buf ( n38261 , n38260 );
xor ( n38262 , n38188 , n38261 );
buf ( n38263 , n32972 );
not ( n38264 , n38263 );
buf ( n38265 , n33077 );
not ( n38266 , n38265 );
buf ( n38267 , n37268 );
not ( n38268 , n38267 );
or ( n38269 , n38266 , n38268 );
buf ( n38270 , n37271 );
buf ( n38271 , n33080 );
nand ( n38272 , n38270 , n38271 );
buf ( n38273 , n38272 );
buf ( n38274 , n38273 );
nand ( n38275 , n38269 , n38274 );
buf ( n38276 , n38275 );
buf ( n38277 , n38276 );
not ( n38278 , n38277 );
or ( n38279 , n38264 , n38278 );
buf ( n38280 , n33077 );
not ( n38281 , n38280 );
not ( n38282 , n37298 );
buf ( n38283 , n38282 );
not ( n38284 , n38283 );
or ( n38285 , n38281 , n38284 );
not ( n38286 , n37293 );
not ( n38287 , n38286 );
buf ( n38288 , n38287 );
buf ( n38289 , n33080 );
nand ( n38290 , n38288 , n38289 );
buf ( n38291 , n38290 );
buf ( n38292 , n38291 );
nand ( n38293 , n38285 , n38292 );
buf ( n38294 , n38293 );
buf ( n38295 , n38294 );
buf ( n38296 , n36107 );
nand ( n38297 , n38295 , n38296 );
buf ( n38298 , n38297 );
buf ( n38299 , n38298 );
nand ( n38300 , n38279 , n38299 );
buf ( n38301 , n38300 );
buf ( n38302 , n38301 );
and ( n38303 , n38262 , n38302 );
and ( n38304 , n38188 , n38261 );
or ( n38305 , n38303 , n38304 );
buf ( n38306 , n38305 );
buf ( n38307 , n38306 );
xnor ( n38308 , n36363 , n37746 );
buf ( n38309 , n38308 );
buf ( n38310 , n36456 );
nand ( n38311 , n38309 , n38310 );
buf ( n38312 , n38311 );
buf ( n38313 , n38312 );
nand ( n38314 , C1 , n38313 );
buf ( n38315 , n38314 );
buf ( n38316 , n38315 );
buf ( n38317 , n38150 );
not ( n38318 , n38317 );
buf ( n38319 , n37335 );
not ( n38320 , n38319 );
or ( n38321 , n38318 , n38320 );
buf ( n38322 , n38164 );
buf ( n38323 , n37403 );
nand ( n38324 , n38322 , n38323 );
buf ( n38325 , n38324 );
buf ( n38326 , n38325 );
nand ( n38327 , n38321 , n38326 );
buf ( n38328 , n38327 );
buf ( n38329 , n38328 );
xor ( n38330 , n38316 , n38329 );
buf ( n38331 , n36915 );
not ( n38332 , n38331 );
buf ( n38333 , n37984 );
not ( n38334 , n38333 );
or ( n38335 , n38332 , n38334 );
buf ( n38336 , n38234 );
buf ( n38337 , n36988 );
nand ( n38338 , n38336 , n38337 );
buf ( n38339 , n38338 );
buf ( n38340 , n38339 );
nand ( n38341 , n38335 , n38340 );
buf ( n38342 , n38341 );
buf ( n38343 , n38342 );
xor ( n38344 , n38330 , n38343 );
buf ( n38345 , n38344 );
buf ( n38346 , n38345 );
xor ( n38347 , n38307 , n38346 );
not ( n38348 , n24638 );
not ( n38349 , n38348 );
not ( n38350 , n38349 );
buf ( n38351 , n32724 );
buf ( n38352 , n32737 );
or ( n38353 , n38351 , n38352 );
buf ( n38354 , n38353 );
buf ( n38355 , n38354 );
not ( n38356 , n38355 );
buf ( n38357 , n38356 );
not ( n38358 , n38357 );
not ( n38359 , n38358 );
nand ( n38360 , n24637 , n24583 );
not ( n38361 , n38360 );
not ( n38362 , n38361 );
or ( n38363 , n38359 , n38362 );
not ( n38364 , n38357 );
not ( n38365 , n24587 );
and ( n38366 , n38364 , n38365 );
not ( n38367 , n24587 );
nor ( n38368 , n38367 , n38354 );
and ( n38369 , n38360 , n38368 );
nor ( n38370 , n38366 , n38369 );
nand ( n38371 , n38363 , n38370 );
buf ( n38372 , n38371 );
not ( n38373 , n38372 );
buf ( n38374 , n38373 );
not ( n38375 , n38374 );
not ( n38376 , n38375 );
or ( n38377 , n38350 , n38376 );
nand ( n38378 , n38374 , n38348 );
nand ( n38379 , n38377 , n38378 );
not ( n38380 , n38379 );
not ( n38381 , n38380 );
not ( n38382 , n38381 );
not ( n38383 , n38382 );
buf ( n38384 , n38383 );
not ( n38385 , n38384 );
buf ( n38386 , n37373 );
not ( n38387 , n38386 );
buf ( n38388 , n37375 );
not ( n38389 , n38388 );
or ( n38390 , n38387 , n38389 );
buf ( n38391 , n37380 );
nand ( n38392 , n38390 , n38391 );
buf ( n38393 , n38392 );
buf ( n38394 , n38393 );
buf ( n38395 , n38371 );
nand ( n38396 , n38394 , n38395 );
buf ( n38397 , n38396 );
not ( n38398 , n38397 );
nor ( n38399 , n37381 , n38371 );
nor ( n38400 , n38398 , n38399 );
or ( n38401 , n38374 , n38348 );
nand ( n38402 , n38401 , n38378 );
nand ( n38403 , n38400 , n38402 );
not ( n38404 , n38403 );
buf ( n38405 , n38404 );
not ( n38406 , n38405 );
buf ( n38407 , n38406 );
buf ( n38408 , n38407 );
not ( n38409 , n38408 );
or ( n38410 , n38385 , n38409 );
not ( n38411 , n37381 );
buf ( n38412 , n38411 );
not ( n38413 , n38412 );
buf ( n38414 , n38413 );
not ( n38415 , n38414 );
buf ( n38416 , n35973 );
not ( n38417 , n38416 );
or ( n38418 , n38415 , n38417 );
buf ( n38419 , n35972 );
not ( n38420 , n38413 );
buf ( n38421 , n38420 );
nand ( n38422 , n38419 , n38421 );
buf ( n38423 , n38422 );
buf ( n38424 , n38423 );
nand ( n38425 , n38418 , n38424 );
buf ( n38426 , n38425 );
buf ( n38427 , n38426 );
nand ( n38428 , n38410 , n38427 );
buf ( n38429 , n38428 );
buf ( n38430 , n38429 );
buf ( n38431 , n38063 );
not ( n38432 , n38431 );
and ( n38433 , n38074 , n37149 );
not ( n38434 , n38074 );
not ( n38435 , n37146 );
not ( n38436 , n38435 );
and ( n38437 , n38434 , n38436 );
or ( n38438 , n38433 , n38437 );
buf ( n38439 , n38438 );
not ( n38440 , n38439 );
or ( n38441 , n38432 , n38440 );
buf ( n38442 , n38074 );
not ( n38443 , n38442 );
buf ( n38444 , n37971 );
not ( n38445 , n38444 );
or ( n38446 , n38443 , n38445 );
not ( n38447 , n37970 );
buf ( n38448 , n38447 );
buf ( n38449 , n38071 );
nand ( n38450 , n38448 , n38449 );
buf ( n38451 , n38450 );
buf ( n38452 , n38451 );
nand ( n38453 , n38446 , n38452 );
buf ( n38454 , n38453 );
buf ( n38455 , n38454 );
buf ( n38456 , n38133 );
nand ( n38457 , n38455 , n38456 );
buf ( n38458 , n38457 );
buf ( n38459 , n38458 );
nand ( n38460 , n38441 , n38459 );
buf ( n38461 , n38460 );
buf ( n38462 , n38461 );
xor ( n38463 , n38430 , n38462 );
not ( n38464 , n37657 );
buf ( n38465 , n38464 );
buf ( n38466 , n36523 );
not ( n38467 , n38466 );
not ( n38468 , n36527 );
buf ( n38469 , n38468 );
not ( n38470 , n38469 );
buf ( n38471 , n38470 );
buf ( n38472 , n38471 );
not ( n38473 , n38472 );
buf ( n38474 , n37786 );
not ( n38475 , n38474 );
or ( n38476 , n38473 , n38475 );
not ( n38477 , n37782 );
buf ( n38478 , n38477 );
buf ( n38479 , n38478 );
buf ( n38480 , n38479 );
buf ( n38481 , n38480 );
buf ( n38482 , n36530 );
nand ( n38483 , n38481 , n38482 );
buf ( n38484 , n38483 );
buf ( n38485 , n38484 );
nand ( n38486 , n38476 , n38485 );
buf ( n38487 , n38486 );
buf ( n38488 , n38487 );
not ( n38489 , n38488 );
or ( n38490 , n38467 , n38489 );
buf ( n38491 , n37757 );
buf ( n38492 , n36643 );
nand ( n38493 , n38491 , n38492 );
buf ( n38494 , n38493 );
buf ( n38495 , n38494 );
nand ( n38496 , n38490 , n38495 );
buf ( n38497 , n38496 );
buf ( n38498 , n38497 );
xor ( n38499 , n38465 , n38498 );
buf ( n38500 , n32972 );
not ( n38501 , n38500 );
buf ( n38502 , n38294 );
not ( n38503 , n38502 );
or ( n38504 , n38501 , n38503 );
buf ( n38505 , n33077 );
buf ( n38506 , n37695 );
and ( n38507 , n38505 , n38506 );
not ( n38508 , n38505 );
buf ( n38509 , n37717 );
and ( n38510 , n38508 , n38509 );
nor ( n38511 , n38507 , n38510 );
buf ( n38512 , n38511 );
buf ( n38513 , n38512 );
buf ( n38514 , n36107 );
nand ( n38515 , n38513 , n38514 );
buf ( n38516 , n38515 );
buf ( n38517 , n38516 );
nand ( n38518 , n38504 , n38517 );
buf ( n38519 , n38518 );
buf ( n38520 , n38519 );
and ( n38521 , n38499 , n38520 );
and ( n38522 , n38465 , n38498 );
or ( n38523 , n38521 , n38522 );
buf ( n38524 , n38523 );
buf ( n38525 , n38524 );
and ( n38526 , n38463 , n38525 );
and ( n38527 , n38430 , n38462 );
or ( n38528 , n38526 , n38527 );
buf ( n38529 , n38528 );
buf ( n38530 , n38529 );
and ( n38531 , n38347 , n38530 );
and ( n38532 , n38307 , n38346 );
or ( n38533 , n38531 , n38532 );
buf ( n38534 , n38533 );
buf ( n38535 , n38534 );
not ( n38536 , n37300 );
not ( n38537 , n36706 );
and ( n38538 , n38536 , n38537 );
not ( n38539 , n36688 );
and ( n38540 , n37722 , n38539 );
nor ( n38541 , n38538 , n38540 );
buf ( n38542 , n38541 );
buf ( n38543 , n36107 );
not ( n38544 , n38543 );
buf ( n38545 , n38276 );
not ( n38546 , n38545 );
or ( n38547 , n38544 , n38546 );
buf ( n38548 , n33077 );
not ( n38549 , n38548 );
buf ( n38550 , n38250 );
not ( n38551 , n38550 );
or ( n38552 , n38549 , n38551 );
buf ( n38553 , n38247 );
buf ( n38554 , n33080 );
nand ( n38555 , n38553 , n38554 );
buf ( n38556 , n38555 );
buf ( n38557 , n38556 );
nand ( n38558 , n38552 , n38557 );
buf ( n38559 , n38558 );
buf ( n38560 , n38559 );
buf ( n38561 , n32972 );
nand ( n38562 , n38560 , n38561 );
buf ( n38563 , n38562 );
buf ( n38564 , n38563 );
nand ( n38565 , n38547 , n38564 );
buf ( n38566 , n38565 );
buf ( n38567 , n38566 );
xor ( n38568 , n38542 , n38567 );
buf ( n38569 , n38063 );
not ( n38570 , n38569 );
buf ( n38571 , n38106 );
not ( n38572 , n38571 );
or ( n38573 , n38570 , n38572 );
buf ( n38574 , n38438 );
buf ( n38575 , n38133 );
nand ( n38576 , n38574 , n38575 );
buf ( n38577 , n38576 );
buf ( n38578 , n38577 );
nand ( n38579 , n38573 , n38578 );
buf ( n38580 , n38579 );
buf ( n38581 , n38580 );
and ( n38582 , n38568 , n38581 );
and ( n38583 , n38542 , n38567 );
or ( n38584 , n38582 , n38583 );
buf ( n38585 , n38584 );
xor ( n38586 , n38316 , n38329 );
and ( n38587 , n38586 , n38343 );
and ( n38588 , n38316 , n38329 );
or ( n38589 , n38587 , n38588 );
buf ( n38590 , n38589 );
xor ( n38591 , n38585 , n38590 );
buf ( n38592 , n32972 );
not ( n38593 , n38592 );
buf ( n38594 , n33077 );
not ( n38595 , n38594 );
buf ( n38596 , n38221 );
not ( n38597 , n38596 );
or ( n38598 , n38595 , n38597 );
buf ( n38599 , n38227 );
buf ( n38600 , n33080 );
nand ( n38601 , n38599 , n38600 );
buf ( n38602 , n38601 );
buf ( n38603 , n38602 );
nand ( n38604 , n38598 , n38603 );
buf ( n38605 , n38604 );
buf ( n38606 , n38605 );
not ( n38607 , n38606 );
or ( n38608 , n38593 , n38607 );
buf ( n38609 , n38559 );
buf ( n38610 , n36107 );
nand ( n38611 , n38609 , n38610 );
buf ( n38612 , n38611 );
buf ( n38613 , n38612 );
nand ( n38614 , n38608 , n38613 );
buf ( n38615 , n38614 );
buf ( n38616 , n38615 );
buf ( n38617 , n38541 );
not ( n38618 , n38617 );
buf ( n38619 , n38618 );
buf ( n38620 , n38619 );
xor ( n38621 , n38616 , n38620 );
buf ( n38622 , n37698 );
buf ( n38623 , n38622 );
buf ( n38624 , n38623 );
not ( n38625 , n38624 );
xor ( n38626 , n36363 , n38625 );
not ( n38627 , n38626 );
not ( n38628 , n36456 );
or ( n38629 , n38627 , n38628 );
buf ( n38630 , C1 );
nand ( n38631 , n38629 , n38630 );
buf ( n38632 , n38631 );
xor ( n38633 , n38621 , n38632 );
buf ( n38634 , n38633 );
xor ( n38635 , n38591 , n38634 );
not ( n38636 , n38635 );
buf ( n38637 , n38636 );
and ( n38638 , n38535 , n38637 );
not ( n38639 , n38535 );
buf ( n38640 , n38635 );
and ( n38641 , n38639 , n38640 );
nor ( n38642 , n38638 , n38641 );
buf ( n38643 , n38642 );
buf ( n38644 , n38643 );
not ( n38645 , n38644 );
xor ( n38646 , n38542 , n38567 );
xor ( n38647 , n38646 , n38581 );
buf ( n38648 , n38647 );
buf ( n38649 , n38648 );
xor ( n38650 , n37562 , n37810 );
xor ( n38651 , n38650 , n37929 );
buf ( n38652 , n38651 );
buf ( n38653 , n38652 );
xor ( n38654 , n38649 , n38653 );
buf ( n38655 , n37922 );
not ( n38656 , n38655 );
buf ( n38657 , n37899 );
not ( n38658 , n38657 );
or ( n38659 , n38656 , n38658 );
not ( n38660 , n37882 );
not ( n38661 , n38660 );
not ( n38662 , n37090 );
or ( n38663 , n38661 , n38662 );
nand ( n38664 , n38098 , n37882 );
nand ( n38665 , n38663 , n38664 );
nand ( n38666 , n38665 , n37875 );
buf ( n38667 , n38666 );
nand ( n38668 , n38659 , n38667 );
buf ( n38669 , n38668 );
buf ( n38670 , n38669 );
buf ( n38671 , n37517 );
not ( n38672 , n38671 );
buf ( n38673 , n37476 );
not ( n38674 , n38673 );
buf ( n38675 , n36430 );
not ( n38676 , n38675 );
or ( n38677 , n38674 , n38676 );
buf ( n38678 , n36427 );
buf ( n38679 , n37545 );
nand ( n38680 , n38678 , n38679 );
buf ( n38681 , n38680 );
buf ( n38682 , n38681 );
nand ( n38683 , n38677 , n38682 );
buf ( n38684 , n38683 );
buf ( n38685 , n38684 );
not ( n38686 , n38685 );
or ( n38687 , n38672 , n38686 );
buf ( n38688 , n37551 );
buf ( n38689 , n37452 );
nand ( n38690 , n38688 , n38689 );
buf ( n38691 , n38690 );
buf ( n38692 , n38691 );
nand ( n38693 , n38687 , n38692 );
buf ( n38694 , n38693 );
buf ( n38695 , n38694 );
xor ( n38696 , n38670 , n38695 );
xor ( n38697 , n37658 , n37764 );
xor ( n38698 , n38697 , n37804 );
buf ( n38699 , n38698 );
buf ( n38700 , n38699 );
and ( n38701 , n38696 , n38700 );
and ( n38702 , n38670 , n38695 );
or ( n38703 , n38701 , n38702 );
buf ( n38704 , n38703 );
buf ( n38705 , n38704 );
and ( n38706 , n38654 , n38705 );
and ( n38707 , n38649 , n38653 );
or ( n38708 , n38706 , n38707 );
buf ( n38709 , n38708 );
buf ( n38710 , n38709 );
not ( n38711 , n38710 );
and ( n38712 , n38645 , n38711 );
buf ( n38713 , n38709 );
buf ( n38714 , n38643 );
and ( n38715 , n38713 , n38714 );
nor ( n38716 , n38712 , n38715 );
buf ( n38717 , n38716 );
buf ( n38718 , n38717 );
xor ( n38719 , n38147 , n38718 );
not ( n38720 , n38133 );
buf ( n38721 , n38071 );
buf ( n38722 , n38221 );
and ( n38723 , n38721 , n38722 );
not ( n38724 , n38721 );
buf ( n38725 , n38227 );
and ( n38726 , n38724 , n38725 );
nor ( n38727 , n38723 , n38726 );
buf ( n38728 , n38727 );
not ( n38729 , n38728 );
or ( n38730 , n38720 , n38729 );
buf ( n38731 , n38063 );
not ( n38732 , n38731 );
buf ( n38733 , n38732 );
not ( n38734 , n38733 );
nand ( n38735 , n38734 , n38454 );
nand ( n38736 , n38730 , n38735 );
buf ( n38737 , n38736 );
buf ( n38738 , n36988 );
not ( n38739 , n38738 );
and ( n38740 , n36935 , n37268 );
not ( n38741 , n36935 );
buf ( n38742 , n37263 );
not ( n38743 , n38742 );
and ( n38744 , n38741 , n38743 );
or ( n38745 , n38740 , n38744 );
buf ( n38746 , n38745 );
not ( n38747 , n38746 );
or ( n38748 , n38739 , n38747 );
buf ( n38749 , n38253 );
buf ( n38750 , n36915 );
nand ( n38751 , n38749 , n38750 );
buf ( n38752 , n38751 );
buf ( n38753 , n38752 );
nand ( n38754 , n38748 , n38753 );
buf ( n38755 , n38754 );
buf ( n38756 , n38755 );
xor ( n38757 , n38737 , n38756 );
not ( n38758 , n38383 );
buf ( n38759 , n38758 );
not ( n38760 , n38759 );
buf ( n38761 , n38426 );
not ( n38762 , n38761 );
or ( n38763 , n38760 , n38762 );
buf ( n38764 , n38413 );
buf ( n38765 , n37481 );
and ( n38766 , n38764 , n38765 );
not ( n38767 , n38764 );
buf ( n38768 , n36054 );
and ( n38769 , n38767 , n38768 );
nor ( n38770 , n38766 , n38769 );
buf ( n38771 , n38770 );
buf ( n38772 , n38771 );
buf ( n38773 , n38407 );
not ( n38774 , n38773 );
buf ( n38775 , n38774 );
buf ( n38776 , n38775 );
nand ( n38777 , n38772 , n38776 );
buf ( n38778 , n38777 );
buf ( n38779 , n38778 );
nand ( n38780 , n38763 , n38779 );
buf ( n38781 , n38780 );
buf ( n38782 , n38781 );
and ( n38783 , n38757 , n38782 );
and ( n38784 , n38737 , n38756 );
or ( n38785 , n38783 , n38784 );
buf ( n38786 , n38785 );
buf ( n38787 , n38786 );
xor ( n38788 , n38188 , n38261 );
xor ( n38789 , n38788 , n38302 );
buf ( n38790 , n38789 );
buf ( n38791 , n38790 );
xor ( n38792 , n38787 , n38791 );
not ( n38793 , n36453 );
not ( n38794 , n37655 );
or ( n38795 , n38793 , n38794 );
buf ( n38796 , n37649 );
not ( n38797 , n38796 );
buf ( n38798 , n38797 );
buf ( n38799 , n38798 );
not ( n38800 , n38799 );
not ( n38801 , n30180 );
nand ( n38802 , n29896 , n30176 );
not ( n38803 , n38802 );
or ( n38804 , n38801 , n38803 );
buf ( n38805 , n37621 );
buf ( n38806 , n35645 );
buf ( n38807 , n35654 );
or ( n38808 , n38806 , n38807 );
buf ( n38809 , n38808 );
buf ( n38810 , n38809 );
nand ( n38811 , n38805 , n38810 );
buf ( n38812 , n38811 );
nand ( n38813 , n38804 , n38812 );
not ( n38814 , n30176 );
not ( n38815 , n29896 );
or ( n38816 , n38814 , n38815 );
not ( n38817 , n30180 );
nor ( n38818 , n38817 , n38812 );
nand ( n38819 , n38816 , n38818 );
nand ( n38820 , n38813 , n38819 );
buf ( n38821 , n38820 );
buf ( n38822 , n38821 );
not ( n38823 , n38822 );
buf ( n38824 , n38823 );
buf ( n38825 , n38824 );
not ( n38826 , n38825 );
or ( n38827 , n38800 , n38826 );
buf ( n38828 , n38821 );
buf ( n38829 , n38828 );
buf ( n38830 , n38829 );
buf ( n38831 , n38830 );
buf ( n38832 , n36357 );
buf ( n38833 , n38832 );
buf ( n38834 , n38833 );
buf ( n38835 , n38834 );
not ( n38836 , n38835 );
buf ( n38837 , n38836 );
buf ( n38838 , n38837 );
nand ( n38839 , n38831 , n38838 );
buf ( n38840 , n38839 );
buf ( n38841 , n38840 );
nand ( n38842 , n38827 , n38841 );
buf ( n38843 , n38842 );
buf ( n38844 , C1 );
nand ( n38845 , n38795 , n38844 );
buf ( n38846 , n30187 );
buf ( n38847 , n38846 );
buf ( n38848 , n38847 );
buf ( n38849 , n38848 );
not ( n38850 , n38849 );
buf ( n38851 , n38850 );
buf ( n38852 , n38851 );
not ( n38853 , n38852 );
buf ( n38854 , n38853 );
buf ( n38855 , n38854 );
not ( n38856 , n38855 );
buf ( n38857 , n37649 );
not ( n38858 , n38857 );
and ( n38859 , n38856 , n38858 );
buf ( n38860 , n30187 );
not ( n38861 , n38860 );
buf ( n38862 , n38861 );
buf ( n38863 , n38862 );
not ( n38864 , n38863 );
buf ( n38865 , n38864 );
buf ( n38866 , n38865 );
buf ( n38867 , n37602 );
and ( n38868 , n38866 , n38867 );
nor ( n38869 , n38859 , n38868 );
buf ( n38870 , n38869 );
buf ( n38871 , n36453 );
buf ( n38872 , n38843 );
nand ( n38873 , n38871 , n38872 );
buf ( n38874 , n38873 );
nand ( n38875 , C1 , n38874 );
xor ( n38876 , n38845 , n38875 );
not ( n38877 , n38487 );
not ( n38878 , n36643 );
or ( n38879 , n38877 , n38878 );
buf ( n38880 , n36523 );
buf ( n38881 , n38471 );
not ( n38882 , n38881 );
buf ( n38883 , n37589 );
not ( n38884 , n38883 );
or ( n38885 , n38882 , n38884 );
buf ( n38886 , n37586 );
buf ( n38887 , n36530 );
nand ( n38888 , n38886 , n38887 );
buf ( n38889 , n38888 );
buf ( n38890 , n38889 );
nand ( n38891 , n38885 , n38890 );
buf ( n38892 , n38891 );
buf ( n38893 , n38892 );
nand ( n38894 , n38880 , n38893 );
buf ( n38895 , n38894 );
nand ( n38896 , n38879 , n38895 );
and ( n38897 , n38876 , n38896 );
and ( n38898 , n38845 , n38875 );
or ( n38899 , n38897 , n38898 );
not ( n38900 , n37922 );
not ( n38901 , n38665 );
or ( n38902 , n38900 , n38901 );
buf ( n38903 , n37882 );
not ( n38904 , n38903 );
buf ( n38905 , n37149 );
not ( n38906 , n38905 );
or ( n38907 , n38904 , n38906 );
buf ( n38908 , n38436 );
buf ( n38909 , n37893 );
nand ( n38910 , n38908 , n38909 );
buf ( n38911 , n38910 );
buf ( n38912 , n38911 );
nand ( n38913 , n38907 , n38912 );
buf ( n38914 , n38913 );
buf ( n38915 , n38914 );
buf ( n38916 , n37875 );
nand ( n38917 , n38915 , n38916 );
buf ( n38918 , n38917 );
nand ( n38919 , n38902 , n38918 );
xor ( n38920 , n38899 , n38919 );
not ( n38921 , n37403 );
buf ( n38922 , n37330 );
not ( n38923 , n38922 );
buf ( n38924 , n36565 );
not ( n38925 , n38924 );
or ( n38926 , n38923 , n38925 );
buf ( n38927 , n37543 );
buf ( n38928 , n37329 );
nand ( n38929 , n38927 , n38928 );
buf ( n38930 , n38929 );
buf ( n38931 , n38930 );
nand ( n38932 , n38926 , n38931 );
buf ( n38933 , n38932 );
not ( n38934 , n38933 );
or ( n38935 , n38921 , n38934 );
buf ( n38936 , n38181 );
buf ( n38937 , n38150 );
nand ( n38938 , n38936 , n38937 );
buf ( n38939 , n38938 );
nand ( n38940 , n38935 , n38939 );
and ( n38941 , n38920 , n38940 );
and ( n38942 , n38899 , n38919 );
or ( n38943 , n38941 , n38942 );
buf ( n38944 , n38943 );
and ( n38945 , n38792 , n38944 );
and ( n38946 , n38787 , n38791 );
or ( n38947 , n38945 , n38946 );
buf ( n38948 , n38947 );
buf ( n38949 , n38948 );
xor ( n38950 , n38307 , n38346 );
xor ( n38951 , n38950 , n38530 );
buf ( n38952 , n38951 );
buf ( n38953 , n38952 );
xor ( n38954 , n38949 , n38953 );
xor ( n38955 , n38430 , n38462 );
xor ( n38956 , n38955 , n38525 );
buf ( n38957 , n38956 );
buf ( n38958 , n38957 );
xor ( n38959 , n38465 , n38498 );
xor ( n38960 , n38959 , n38520 );
buf ( n38961 , n38960 );
buf ( n38962 , n38961 );
buf ( n38963 , n24091 );
or ( n38964 , n25139 , n38963 );
and ( n38965 , n25134 , n25129 );
not ( n38966 , n25134 );
not ( n38967 , n25129 );
and ( n38968 , n38966 , n38967 );
nor ( n38969 , n38965 , n38968 );
nand ( n38970 , n38969 , n38963 );
nand ( n38971 , n38964 , n38970 );
not ( n38972 , n38971 );
buf ( n38973 , n38972 );
buf ( n38974 , n38973 );
buf ( n38975 , n38974 );
not ( n38976 , n38975 );
buf ( n38977 , n24638 );
buf ( n38978 , n38977 );
buf ( n38979 , n38978 );
nand ( n38980 , n25140 , n38979 );
nand ( n38981 , n38969 , n38348 );
nand ( n38982 , n38980 , n38972 , n38981 );
buf ( n38983 , n38982 );
not ( n38984 , n38983 );
buf ( n38985 , n38984 );
buf ( n38986 , n38985 );
not ( n38987 , n38986 );
buf ( n38988 , n38987 );
buf ( n38989 , n38988 );
not ( n38990 , n38989 );
or ( n38991 , n38976 , n38990 );
buf ( n38992 , n38979 );
not ( n38993 , n38992 );
buf ( n38994 , n38993 );
buf ( n38995 , n38994 );
buf ( n38996 , n38995 );
buf ( n38997 , n38996 );
buf ( n38998 , n38997 );
not ( n38999 , n38998 );
buf ( n39000 , n38999 );
buf ( n39001 , n39000 );
not ( n39002 , n39001 );
buf ( n39003 , n35968 );
buf ( n39004 , n39003 );
buf ( n39005 , n39004 );
buf ( n39006 , n39005 );
not ( n39007 , n39006 );
buf ( n39008 , n39007 );
buf ( n39009 , n39008 );
not ( n39010 , n39009 );
or ( n39011 , n39002 , n39010 );
buf ( n39012 , n35970 );
buf ( n39013 , n38997 );
nand ( n39014 , n39012 , n39013 );
buf ( n39015 , n39014 );
buf ( n39016 , n39015 );
nand ( n39017 , n39011 , n39016 );
buf ( n39018 , n39017 );
buf ( n39019 , n39018 );
nand ( n39020 , n38991 , n39019 );
buf ( n39021 , n39020 );
not ( n39022 , n38512 );
not ( n39023 , n32972 );
or ( n39024 , n39022 , n39023 );
buf ( n39025 , n33077 );
not ( n39026 , n39025 );
buf ( n39027 , n37746 );
not ( n39028 , n39027 );
or ( n39029 , n39026 , n39028 );
buf ( n39030 , n37750 );
buf ( n39031 , n33080 );
nand ( n39032 , n39030 , n39031 );
buf ( n39033 , n39032 );
buf ( n39034 , n39033 );
nand ( n39035 , n39029 , n39034 );
buf ( n39036 , n39035 );
buf ( n39037 , n39036 );
buf ( n39038 , n36107 );
nand ( n39039 , n39037 , n39038 );
buf ( n39040 , n39039 );
nand ( n39041 , n39024 , n39040 );
xor ( n39042 , n39021 , n39041 );
buf ( n39043 , n38063 );
not ( n39044 , n39043 );
buf ( n39045 , n38728 );
not ( n39046 , n39045 );
or ( n39047 , n39044 , n39046 );
buf ( n39048 , n38074 );
buf ( n39049 , n38247 );
and ( n39050 , n39048 , n39049 );
not ( n39051 , n39048 );
buf ( n39052 , n38250 );
and ( n39053 , n39051 , n39052 );
nor ( n39054 , n39050 , n39053 );
buf ( n39055 , n39054 );
buf ( n39056 , n39055 );
buf ( n39057 , n38133 );
nand ( n39058 , n39056 , n39057 );
buf ( n39059 , n39058 );
buf ( n39060 , n39059 );
nand ( n39061 , n39047 , n39060 );
buf ( n39062 , n39061 );
and ( n39063 , n39042 , n39062 );
and ( n39064 , n39021 , n39041 );
or ( n39065 , n39063 , n39064 );
buf ( n39066 , n39065 );
xor ( n39067 , n38962 , n39066 );
not ( n39068 , n37476 );
not ( n39069 , n37887 );
or ( n39070 , n39068 , n39069 );
buf ( n39071 , n36399 );
buf ( n39072 , n37475 );
nand ( n39073 , n39071 , n39072 );
buf ( n39074 , n39073 );
nand ( n39075 , n39070 , n39074 );
not ( n39076 , n39075 );
not ( n39077 , n37517 );
or ( n39078 , n39076 , n39077 );
buf ( n39079 , n38684 );
buf ( n39080 , n37452 );
nand ( n39081 , n39079 , n39080 );
buf ( n39082 , n39081 );
nand ( n39083 , n39078 , n39082 );
buf ( n39084 , n39083 );
and ( n39085 , n39067 , n39084 );
and ( n39086 , n38962 , n39066 );
or ( n39087 , n39085 , n39086 );
buf ( n39088 , n39087 );
buf ( n39089 , n39088 );
xor ( n39090 , n38958 , n39089 );
xor ( n39091 , n38670 , n38695 );
xor ( n39092 , n39091 , n38700 );
buf ( n39093 , n39092 );
buf ( n39094 , n39093 );
and ( n39095 , n39090 , n39094 );
and ( n39096 , n38958 , n39089 );
or ( n39097 , n39095 , n39096 );
buf ( n39098 , n39097 );
buf ( n39099 , n39098 );
and ( n39100 , n38954 , n39099 );
and ( n39101 , n38949 , n38953 );
or ( n39102 , n39100 , n39101 );
buf ( n39103 , n39102 );
buf ( n39104 , n39103 );
not ( n39105 , n39104 );
buf ( n39106 , n39105 );
buf ( n39107 , n39106 );
xor ( n39108 , n38719 , n39107 );
buf ( n39109 , n39108 );
buf ( n39110 , n39109 );
xor ( n39111 , n38949 , n38953 );
xor ( n39112 , n39111 , n39099 );
buf ( n39113 , n39112 );
xor ( n39114 , n38649 , n38653 );
xor ( n39115 , n39114 , n38705 );
buf ( n39116 , n39115 );
nor ( n39117 , n39113 , n39116 );
not ( n39118 , n39117 );
xor ( n39119 , n38787 , n38791 );
xor ( n39120 , n39119 , n38944 );
buf ( n39121 , n39120 );
buf ( n39122 , n39121 );
buf ( n39123 , n36915 );
not ( n39124 , n39123 );
buf ( n39125 , n38745 );
not ( n39126 , n39125 );
or ( n39127 , n39124 , n39126 );
buf ( n39128 , n36935 );
not ( n39129 , n39128 );
buf ( n39130 , n37295 );
not ( n39131 , n39130 );
or ( n39132 , n39129 , n39131 );
buf ( n39133 , n37298 );
buf ( n39134 , n36966 );
not ( n39135 , n39134 );
buf ( n39136 , n39135 );
buf ( n39137 , n39136 );
not ( n39138 , n39137 );
buf ( n39139 , n39138 );
buf ( n39140 , n39139 );
nand ( n39141 , n39133 , n39140 );
buf ( n39142 , n39141 );
buf ( n39143 , n39142 );
nand ( n39144 , n39132 , n39143 );
buf ( n39145 , n39144 );
buf ( n39146 , n39145 );
buf ( n39147 , n36988 );
nand ( n39148 , n39146 , n39147 );
buf ( n39149 , n39148 );
buf ( n39150 , n39149 );
nand ( n39151 , n39127 , n39150 );
buf ( n39152 , n39151 );
buf ( n39153 , n39152 );
buf ( n39154 , n38758 );
not ( n39155 , n39154 );
buf ( n39156 , n38771 );
not ( n39157 , n39156 );
or ( n39158 , n39155 , n39157 );
buf ( n39159 , n38413 );
buf ( n39160 , n36617 );
and ( n39161 , n39159 , n39160 );
not ( n39162 , n39159 );
buf ( n39163 , n36614 );
and ( n39164 , n39162 , n39163 );
nor ( n39165 , n39161 , n39164 );
buf ( n39166 , n39165 );
buf ( n39167 , n39166 );
buf ( n39168 , n38775 );
nand ( n39169 , n39167 , n39168 );
buf ( n39170 , n39169 );
buf ( n39171 , n39170 );
nand ( n39172 , n39158 , n39171 );
buf ( n39173 , n39172 );
buf ( n39174 , n39173 );
xor ( n39175 , n39153 , n39174 );
xor ( n39176 , n38845 , n38875 );
xor ( n39177 , n39176 , n38896 );
buf ( n39178 , n39177 );
and ( n39179 , n39175 , n39178 );
and ( n39180 , n39153 , n39174 );
or ( n39181 , n39179 , n39180 );
buf ( n39182 , n39181 );
buf ( n39183 , n39182 );
xor ( n39184 , n38737 , n38756 );
xor ( n39185 , n39184 , n38782 );
buf ( n39186 , n39185 );
buf ( n39187 , n39186 );
xor ( n39188 , n39183 , n39187 );
xor ( n39189 , n38899 , n38919 );
xor ( n39190 , n39189 , n38940 );
buf ( n39191 , n39190 );
and ( n39192 , n39188 , n39191 );
and ( n39193 , n39183 , n39187 );
or ( n39194 , n39192 , n39193 );
buf ( n39195 , n39194 );
buf ( n39196 , n39195 );
xor ( n39197 , n39122 , n39196 );
buf ( n39198 , n38875 );
not ( n39199 , n39198 );
buf ( n39200 , n39199 );
buf ( n39201 , n39200 );
buf ( n39202 , n36533 );
nand ( n39203 , n37623 , n37632 );
nand ( n39204 , n37639 , n39203 );
buf ( n39205 , n39204 );
buf ( n39206 , n39205 );
and ( n39207 , n39202 , n39206 );
not ( n39208 , n39202 );
not ( n39209 , n39205 );
buf ( n39210 , n39209 );
and ( n39211 , n39208 , n39210 );
nor ( n39212 , n39207 , n39211 );
buf ( n39213 , n39212 );
buf ( n39214 , n39213 );
not ( n39215 , n39214 );
buf ( n39216 , n36523 );
not ( n39217 , n39216 );
or ( n39218 , n39215 , n39217 );
buf ( n39219 , n38892 );
buf ( n39220 , n36643 );
nand ( n39221 , n39219 , n39220 );
buf ( n39222 , n39221 );
buf ( n39223 , n39222 );
nand ( n39224 , n39218 , n39223 );
buf ( n39225 , n39224 );
buf ( n39226 , n39225 );
xor ( n39227 , n39201 , n39226 );
buf ( n39228 , n36915 );
not ( n39229 , n39228 );
buf ( n39230 , n39145 );
not ( n39231 , n39230 );
or ( n39232 , n39229 , n39231 );
buf ( n39233 , n39139 );
not ( n39234 , n39233 );
buf ( n39235 , n39234 );
buf ( n39236 , n39235 );
not ( n39237 , n39236 );
buf ( n39238 , n37708 );
buf ( n39239 , n39238 );
buf ( n39240 , n39239 );
buf ( n39241 , n39240 );
not ( n39242 , n39241 );
or ( n39243 , n39237 , n39242 );
buf ( n39244 , n39240 );
not ( n39245 , n39244 );
buf ( n39246 , n39245 );
buf ( n39247 , n39246 );
buf ( n39248 , n39139 );
nand ( n39249 , n39247 , n39248 );
buf ( n39250 , n39249 );
buf ( n39251 , n39250 );
nand ( n39252 , n39243 , n39251 );
buf ( n39253 , n39252 );
buf ( n39254 , n39253 );
buf ( n39255 , n36985 );
not ( n39256 , n39255 );
buf ( n39257 , n39256 );
buf ( n39258 , n39257 );
nand ( n39259 , n39254 , n39258 );
buf ( n39260 , n39259 );
buf ( n39261 , n39260 );
nand ( n39262 , n39232 , n39261 );
buf ( n39263 , n39262 );
buf ( n39264 , n39263 );
and ( n39265 , n39227 , n39264 );
and ( n39266 , n39201 , n39226 );
or ( n39267 , n39265 , n39266 );
buf ( n39268 , n39267 );
buf ( n39269 , n39268 );
buf ( n39270 , n37922 );
not ( n39271 , n39270 );
buf ( n39272 , n38914 );
not ( n39273 , n39272 );
or ( n39274 , n39271 , n39273 );
buf ( n39275 , n37882 );
not ( n39276 , n39275 );
not ( n39277 , n37969 );
buf ( n39278 , n39277 );
not ( n39279 , n39278 );
buf ( n39280 , n39279 );
buf ( n39281 , n39280 );
not ( n39282 , n39281 );
or ( n39283 , n39276 , n39282 );
buf ( n39284 , n38447 );
buf ( n39285 , n37893 );
nand ( n39286 , n39284 , n39285 );
buf ( n39287 , n39286 );
buf ( n39288 , n39287 );
nand ( n39289 , n39283 , n39288 );
buf ( n39290 , n39289 );
buf ( n39291 , n39290 );
buf ( n39292 , n37875 );
nand ( n39293 , n39291 , n39292 );
buf ( n39294 , n39293 );
buf ( n39295 , n39294 );
nand ( n39296 , n39274 , n39295 );
buf ( n39297 , n39296 );
buf ( n39298 , n39297 );
xor ( n39299 , n39269 , n39298 );
buf ( n39300 , n37403 );
not ( n39301 , n39300 );
buf ( n39302 , n37330 );
not ( n39303 , n39302 );
buf ( n39304 , n36430 );
not ( n39305 , n39304 );
or ( n39306 , n39303 , n39305 );
buf ( n39307 , n36427 );
buf ( n39308 , n37329 );
nand ( n39309 , n39307 , n39308 );
buf ( n39310 , n39309 );
buf ( n39311 , n39310 );
nand ( n39312 , n39306 , n39311 );
buf ( n39313 , n39312 );
buf ( n39314 , n39313 );
not ( n39315 , n39314 );
or ( n39316 , n39301 , n39315 );
buf ( n39317 , n38933 );
buf ( n39318 , n38150 );
nand ( n39319 , n39317 , n39318 );
buf ( n39320 , n39319 );
buf ( n39321 , n39320 );
nand ( n39322 , n39316 , n39321 );
buf ( n39323 , n39322 );
buf ( n39324 , n39323 );
and ( n39325 , n39299 , n39324 );
and ( n39326 , n39269 , n39298 );
or ( n39327 , n39325 , n39326 );
buf ( n39328 , n39327 );
buf ( n39329 , n39328 );
not ( n39330 , n37452 );
not ( n39331 , n39075 );
or ( n39332 , n39330 , n39331 );
buf ( n39333 , n37476 );
not ( n39334 , n39333 );
buf ( n39335 , n38098 );
not ( n39336 , n39335 );
or ( n39337 , n39334 , n39336 );
buf ( n39338 , n37081 );
not ( n39339 , n39338 );
buf ( n39340 , n39339 );
buf ( n39341 , n39340 );
buf ( n39342 , n37545 );
nand ( n39343 , n39341 , n39342 );
buf ( n39344 , n39343 );
buf ( n39345 , n39344 );
nand ( n39346 , n39337 , n39345 );
buf ( n39347 , n39346 );
buf ( n39348 , n39347 );
buf ( n39349 , n37517 );
nand ( n39350 , n39348 , n39349 );
buf ( n39351 , n39350 );
nand ( n39352 , n39332 , n39351 );
buf ( n39353 , n39352 );
buf ( n39354 , n36107 );
not ( n39355 , n39354 );
buf ( n39356 , n38480 );
not ( n39357 , n39356 );
buf ( n39358 , n39357 );
and ( n39359 , n33077 , n39358 );
not ( n39360 , n33077 );
and ( n39361 , n39360 , n38480 );
or ( n39362 , n39359 , n39361 );
buf ( n39363 , n39362 );
not ( n39364 , n39363 );
or ( n39365 , n39355 , n39364 );
buf ( n39366 , n39036 );
buf ( n39367 , n32972 );
nand ( n39368 , n39366 , n39367 );
buf ( n39369 , n39368 );
buf ( n39370 , n39369 );
nand ( n39371 , n39365 , n39370 );
buf ( n39372 , n39371 );
buf ( n39373 , n39372 );
not ( n39374 , n38974 );
buf ( n39375 , n39374 );
not ( n39376 , n39375 );
buf ( n39377 , n39018 );
not ( n39378 , n39377 );
or ( n39379 , n39376 , n39378 );
buf ( n39380 , n39000 );
not ( n39381 , n39380 );
buf ( n39382 , n36041 );
not ( n39383 , n39382 );
or ( n39384 , n39381 , n39383 );
buf ( n39385 , n36038 );
buf ( n39386 , n38997 );
nand ( n39387 , n39385 , n39386 );
buf ( n39388 , n39387 );
buf ( n39389 , n39388 );
nand ( n39390 , n39384 , n39389 );
buf ( n39391 , n39390 );
buf ( n39392 , n39391 );
buf ( n39393 , n38988 );
not ( n39394 , n39393 );
buf ( n39395 , n39394 );
buf ( n39396 , n39395 );
nand ( n39397 , n39392 , n39396 );
buf ( n39398 , n39397 );
buf ( n39399 , n39398 );
nand ( n39400 , n39379 , n39399 );
buf ( n39401 , n39400 );
buf ( n39402 , n39401 );
xor ( n39403 , n39373 , n39402 );
buf ( n39404 , n37875 );
not ( n39405 , n39404 );
buf ( n39406 , n38217 );
buf ( n39407 , n39406 );
and ( n39408 , n37892 , n39407 );
not ( n39409 , n37892 );
and ( n39410 , n39409 , n38227 );
or ( n39411 , n39408 , n39410 );
buf ( n39412 , n39411 );
not ( n39413 , n39412 );
or ( n39414 , n39405 , n39413 );
buf ( n39415 , n39290 );
buf ( n39416 , n37922 );
nand ( n39417 , n39415 , n39416 );
buf ( n39418 , n39417 );
buf ( n39419 , n39418 );
nand ( n39420 , n39414 , n39419 );
buf ( n39421 , n39420 );
buf ( n39422 , n39421 );
and ( n39423 , n39403 , n39422 );
and ( n39424 , n39373 , n39402 );
or ( n39425 , n39423 , n39424 );
buf ( n39426 , n39425 );
buf ( n39427 , n39426 );
xor ( n39428 , n39353 , n39427 );
xor ( n39429 , n39021 , n39041 );
xor ( n39430 , n39429 , n39062 );
buf ( n39431 , n39430 );
and ( n39432 , n39428 , n39431 );
and ( n39433 , n39353 , n39427 );
or ( n39434 , n39432 , n39433 );
buf ( n39435 , n39434 );
buf ( n39436 , n39435 );
xor ( n39437 , n39329 , n39436 );
xor ( n39438 , n38962 , n39066 );
xor ( n39439 , n39438 , n39084 );
buf ( n39440 , n39439 );
buf ( n39441 , n39440 );
and ( n39442 , n39437 , n39441 );
and ( n39443 , n39329 , n39436 );
or ( n39444 , n39442 , n39443 );
buf ( n39445 , n39444 );
buf ( n39446 , n39445 );
and ( n39447 , n39197 , n39446 );
and ( n39448 , n39122 , n39196 );
or ( n39449 , n39447 , n39448 );
buf ( n39450 , n39449 );
buf ( n39451 , n39450 );
not ( n39452 , n39451 );
buf ( n39453 , n39452 );
not ( n39454 , n39453 );
and ( n39455 , n39118 , n39454 );
buf ( n39456 , n39116 );
buf ( n39457 , n39113 );
and ( n39458 , n39456 , n39457 );
buf ( n39459 , n39458 );
nor ( n39460 , n39455 , n39459 );
buf ( n39461 , n39460 );
nand ( n39462 , n39110 , n39461 );
buf ( n39463 , n39462 );
buf ( n39464 , n39463 );
not ( n39465 , n39464 );
xor ( n39466 , n39269 , n39298 );
xor ( n39467 , n39466 , n39324 );
buf ( n39468 , n39467 );
buf ( n39469 , n39468 );
buf ( n39470 , n32972 );
not ( n39471 , n39470 );
buf ( n39472 , n39362 );
not ( n39473 , n39472 );
or ( n39474 , n39471 , n39473 );
not ( n39475 , n33075 );
buf ( n39476 , n39475 );
not ( n39477 , n39476 );
buf ( n39478 , n39477 );
buf ( n39479 , n39478 );
not ( n39480 , n39479 );
buf ( n39481 , n39480 );
buf ( n39482 , n39481 );
not ( n39483 , n39482 );
buf ( n39484 , n37595 );
not ( n39485 , n39484 );
or ( n39486 , n39483 , n39485 );
buf ( n39487 , n37586 );
buf ( n39488 , n39487 );
buf ( n39489 , n39488 );
buf ( n39490 , n39489 );
buf ( n39491 , n36076 );
buf ( n39492 , n39491 );
buf ( n39493 , n39492 );
buf ( n39494 , n39493 );
nand ( n39495 , n39490 , n39494 );
buf ( n39496 , n39495 );
buf ( n39497 , n39496 );
nand ( n39498 , n39486 , n39497 );
buf ( n39499 , n39498 );
buf ( n39500 , n39499 );
buf ( n39501 , n36104 );
nand ( n39502 , n39500 , n39501 );
buf ( n39503 , n39502 );
buf ( n39504 , n39503 );
nand ( n39505 , n39474 , n39504 );
buf ( n39506 , n39505 );
buf ( n39507 , n39506 );
buf ( n39508 , n36915 );
not ( n39509 , n39508 );
buf ( n39510 , n39253 );
not ( n39511 , n39510 );
or ( n39512 , n39509 , n39511 );
buf ( n39513 , n39257 );
buf ( n39514 , n36935 );
not ( n39515 , n39514 );
buf ( n39516 , n37745 );
buf ( n39517 , n39516 );
buf ( n39518 , n39517 );
buf ( n39519 , n39518 );
not ( n39520 , n39519 );
or ( n39521 , n39515 , n39520 );
not ( n39522 , n37745 );
buf ( n39523 , n39522 );
buf ( n39524 , n39139 );
nand ( n39525 , n39523 , n39524 );
buf ( n39526 , n39525 );
buf ( n39527 , n39526 );
nand ( n39528 , n39521 , n39527 );
buf ( n39529 , n39528 );
buf ( n39530 , n39529 );
nand ( n39531 , n39513 , n39530 );
buf ( n39532 , n39531 );
buf ( n39533 , n39532 );
nand ( n39534 , n39512 , n39533 );
buf ( n39535 , n39534 );
buf ( n39536 , n39535 );
xor ( n39537 , n39507 , n39536 );
buf ( n39538 , n37922 );
not ( n39539 , n39538 );
buf ( n39540 , n39411 );
not ( n39541 , n39540 );
or ( n39542 , n39539 , n39541 );
buf ( n39543 , n37892 );
not ( n39544 , n39543 );
buf ( n39545 , n38250 );
not ( n39546 , n39545 );
or ( n39547 , n39544 , n39546 );
nand ( n39548 , n38660 , n38247 );
buf ( n39549 , n39548 );
nand ( n39550 , n39547 , n39549 );
buf ( n39551 , n39550 );
buf ( n39552 , n39551 );
buf ( n39553 , n37875 );
nand ( n39554 , n39552 , n39553 );
buf ( n39555 , n39554 );
buf ( n39556 , n39555 );
nand ( n39557 , n39542 , n39556 );
buf ( n39558 , n39557 );
buf ( n39559 , n39558 );
and ( n39560 , n39537 , n39559 );
and ( n39561 , n39507 , n39536 );
or ( n39562 , n39560 , n39561 );
buf ( n39563 , n39562 );
buf ( n39564 , n39563 );
not ( n39565 , n39564 );
xor ( n39566 , n39373 , n39402 );
xor ( n39567 , n39566 , n39422 );
buf ( n39568 , n39567 );
buf ( n39569 , n39568 );
not ( n39570 , n39569 );
or ( n39571 , n39565 , n39570 );
buf ( n39572 , n39568 );
buf ( n39573 , n39563 );
or ( n39574 , n39572 , n39573 );
buf ( n39575 , n39374 );
not ( n39576 , n39575 );
buf ( n39577 , n39391 );
not ( n39578 , n39577 );
or ( n39579 , n39576 , n39578 );
buf ( n39580 , n39000 );
not ( n39581 , n39580 );
not ( n39582 , n36611 );
buf ( n39583 , n39582 );
not ( n39584 , n39583 );
or ( n39585 , n39581 , n39584 );
buf ( n39586 , n36617 );
buf ( n39587 , n38997 );
nand ( n39588 , n39586 , n39587 );
buf ( n39589 , n39588 );
buf ( n39590 , n39589 );
nand ( n39591 , n39585 , n39590 );
buf ( n39592 , n39591 );
buf ( n39593 , n39592 );
buf ( n39594 , n39395 );
nand ( n39595 , n39593 , n39594 );
buf ( n39596 , n39595 );
buf ( n39597 , n39596 );
nand ( n39598 , n39579 , n39597 );
buf ( n39599 , n39598 );
buf ( n39600 , n39599 );
not ( n39601 , n39600 );
buf ( n39602 , n38074 );
not ( n39603 , n39602 );
buf ( n39604 , n37268 );
not ( n39605 , n39604 );
or ( n39606 , n39603 , n39605 );
buf ( n39607 , n37271 );
buf ( n39608 , n38071 );
nand ( n39609 , n39607 , n39608 );
buf ( n39610 , n39609 );
buf ( n39611 , n39610 );
nand ( n39612 , n39606 , n39611 );
buf ( n39613 , n39612 );
buf ( n39614 , n39613 );
buf ( n39615 , n38063 );
and ( n39616 , n39614 , n39615 );
buf ( n39617 , n38074 );
not ( n39618 , n39617 );
buf ( n39619 , n37295 );
not ( n39620 , n39619 );
or ( n39621 , n39618 , n39620 );
buf ( n39622 , n38287 );
buf ( n39623 , n38071 );
nand ( n39624 , n39622 , n39623 );
buf ( n39625 , n39624 );
buf ( n39626 , n39625 );
nand ( n39627 , n39621 , n39626 );
buf ( n39628 , n39627 );
buf ( n39629 , n39628 );
not ( n39630 , n39629 );
buf ( n39631 , n38133 );
not ( n39632 , n39631 );
buf ( n39633 , n39632 );
buf ( n39634 , n39633 );
nor ( n39635 , n39630 , n39634 );
buf ( n39636 , n39635 );
buf ( n39637 , n39636 );
nor ( n39638 , n39616 , n39637 );
buf ( n39639 , n39638 );
buf ( n39640 , n39639 );
not ( n39641 , n39640 );
buf ( n39642 , n39641 );
buf ( n39643 , n39642 );
not ( n39644 , n39643 );
or ( n39645 , n39601 , n39644 );
buf ( n39646 , n39642 );
buf ( n39647 , n39599 );
or ( n39648 , n39646 , n39647 );
buf ( n39649 , n38798 );
not ( n39650 , n39649 );
buf ( n39651 , n29287 );
buf ( n39652 , n39651 );
buf ( n39653 , n39652 );
buf ( n39654 , n39653 );
not ( n39655 , n39654 );
buf ( n39656 , n39655 );
buf ( n39657 , n39656 );
not ( n39658 , n39657 );
and ( n39659 , n39650 , n39658 );
buf ( n39660 , n38798 );
buf ( n39661 , n39656 );
and ( n39662 , n39660 , n39661 );
nor ( n39663 , n39659 , n39662 );
buf ( n39664 , n39663 );
buf ( n39665 , n36444 );
not ( n39666 , n39665 );
buf ( n39667 , n39666 );
buf ( n39668 , n39667 );
buf ( n39669 , n38798 );
not ( n39670 , n39669 );
not ( n39671 , n29269 );
buf ( n39672 , n39671 );
buf ( n39673 , n39672 );
not ( n39674 , n39673 );
and ( n39675 , n39670 , n39674 );
buf ( n39676 , n37602 );
not ( n39677 , n39676 );
buf ( n39678 , n39677 );
buf ( n39679 , n39678 );
buf ( n39680 , n29269 );
not ( n39681 , n39680 );
buf ( n39682 , n39681 );
buf ( n39683 , n39682 );
buf ( n39684 , n39683 );
buf ( n39685 , n39684 );
buf ( n39686 , n39685 );
buf ( n39687 , n39686 );
buf ( n39688 , n39687 );
buf ( n39689 , n39688 );
and ( n39690 , n39679 , n39689 );
nor ( n39691 , n39675 , n39690 );
buf ( n39692 , n39691 );
buf ( n39693 , n39692 );
nor ( n39694 , n39668 , n39693 );
buf ( n39695 , n39694 );
buf ( n39696 , n39695 );
nor ( n39697 , C0 , n39696 );
buf ( n39698 , n39697 );
buf ( n39699 , n39698 );
not ( n39700 , n39481 );
not ( n39701 , n39205 );
not ( n39702 , n39701 );
or ( n39703 , n39700 , n39702 );
buf ( n39704 , n39205 );
buf ( n39705 , n39493 );
nand ( n39706 , n39704 , n39705 );
buf ( n39707 , n39706 );
nand ( n39708 , n39703 , n39707 );
not ( n39709 , n39708 );
not ( n39710 , n36104 );
or ( n39711 , n39709 , n39710 );
buf ( n39712 , n39499 );
buf ( n39713 , n32966 );
not ( n39714 , n39713 );
buf ( n39715 , n39714 );
buf ( n39716 , n39715 );
buf ( n39717 , n39716 );
buf ( n39718 , n39717 );
buf ( n39719 , n39718 );
nand ( n39720 , n39712 , n39719 );
buf ( n39721 , n39720 );
nand ( n39722 , n39711 , n39721 );
buf ( n39723 , n39722 );
xor ( n39724 , n39699 , n39723 );
buf ( n39725 , n36520 );
not ( n39726 , n36469 );
buf ( n39727 , n39726 );
not ( n39728 , n39727 );
buf ( n39729 , n39728 );
buf ( n39730 , n39729 );
buf ( n39731 , n38862 );
and ( n39732 , n39730 , n39731 );
not ( n39733 , n39730 );
buf ( n39734 , n38865 );
and ( n39735 , n39733 , n39734 );
nor ( n39736 , n39732 , n39735 );
buf ( n39737 , n39736 );
buf ( n39738 , n39737 );
or ( n39739 , n39725 , n39738 );
buf ( n39740 , n38830 );
not ( n39741 , n39740 );
buf ( n39742 , n39741 );
buf ( n39743 , n39742 );
buf ( n39744 , n39729 );
and ( n39745 , n39743 , n39744 );
buf ( n39746 , n38830 );
buf ( n39747 , n36530 );
and ( n39748 , n39746 , n39747 );
nor ( n39749 , n39745 , n39748 );
buf ( n39750 , n39749 );
buf ( n39751 , n39750 );
buf ( n39752 , n36640 );
or ( n39753 , n39751 , n39752 );
nand ( n39754 , n39739 , n39753 );
buf ( n39755 , n39754 );
buf ( n39756 , n39755 );
and ( n39757 , n39724 , n39756 );
and ( n39758 , n39699 , n39723 );
or ( n39759 , n39757 , n39758 );
buf ( n39760 , n39759 );
buf ( n39761 , n39760 );
nand ( n39762 , n39648 , n39761 );
buf ( n39763 , n39762 );
buf ( n39764 , n39763 );
nand ( n39765 , n39645 , n39764 );
buf ( n39766 , n39765 );
buf ( n39767 , n39766 );
nand ( n39768 , n39574 , n39767 );
buf ( n39769 , n39768 );
buf ( n39770 , n39769 );
nand ( n39771 , n39571 , n39770 );
buf ( n39772 , n39771 );
buf ( n39773 , n39772 );
xor ( n39774 , n39469 , n39773 );
xor ( n39775 , n39353 , n39427 );
xor ( n39776 , n39775 , n39431 );
buf ( n39777 , n39776 );
buf ( n39778 , n39777 );
xor ( n39779 , n39774 , n39778 );
buf ( n39780 , n39779 );
buf ( n39781 , n39780 );
not ( n39782 , n39781 );
xor ( n39783 , n39153 , n39174 );
xor ( n39784 , n39783 , n39178 );
buf ( n39785 , n39784 );
buf ( n39786 , n39785 );
buf ( n39787 , n36450 );
buf ( n39788 , n38870 );
or ( n39789 , n39787 , n39788 );
nand ( n39790 , C1 , n39789 );
buf ( n39791 , n39790 );
buf ( n39792 , n39791 );
buf ( n39793 , n39698 );
not ( n39794 , n39793 );
buf ( n39795 , n39794 );
buf ( n39796 , n39795 );
xor ( n39797 , n39792 , n39796 );
buf ( n39798 , n39750 );
not ( n39799 , n39798 );
buf ( n39800 , n39799 );
buf ( n39801 , n39800 );
not ( n39802 , n39801 );
not ( n39803 , n36517 );
buf ( n39804 , n39803 );
buf ( n39805 , n39804 );
buf ( n39806 , n39805 );
buf ( n39807 , n39806 );
not ( n39808 , n39807 );
or ( n39809 , n39802 , n39808 );
buf ( n39810 , n39213 );
buf ( n39811 , n36640 );
buf ( n39812 , n39811 );
buf ( n39813 , n39812 );
buf ( n39814 , n39813 );
not ( n39815 , n39814 );
buf ( n39816 , n39815 );
buf ( n39817 , n39816 );
nand ( n39818 , n39810 , n39817 );
buf ( n39819 , n39818 );
buf ( n39820 , n39819 );
nand ( n39821 , n39809 , n39820 );
buf ( n39822 , n39821 );
buf ( n39823 , n39822 );
and ( n39824 , n39797 , n39823 );
and ( n39825 , n39792 , n39796 );
or ( n39826 , n39824 , n39825 );
buf ( n39827 , n39826 );
buf ( n39828 , n39827 );
buf ( n39829 , n38133 );
not ( n39830 , n39829 );
buf ( n39831 , n39613 );
not ( n39832 , n39831 );
or ( n39833 , n39830 , n39832 );
buf ( n39834 , n39055 );
buf ( n39835 , n38063 );
nand ( n39836 , n39834 , n39835 );
buf ( n39837 , n39836 );
buf ( n39838 , n39837 );
nand ( n39839 , n39833 , n39838 );
buf ( n39840 , n39839 );
buf ( n39841 , n39840 );
xor ( n39842 , n39828 , n39841 );
xor ( n39843 , n39201 , n39226 );
xor ( n39844 , n39843 , n39264 );
buf ( n39845 , n39844 );
buf ( n39846 , n39845 );
and ( n39847 , n39842 , n39846 );
and ( n39848 , n39828 , n39841 );
or ( n39849 , n39847 , n39848 );
buf ( n39850 , n39849 );
buf ( n39851 , n39850 );
xor ( n39852 , n39786 , n39851 );
buf ( n39853 , n37452 );
not ( n39854 , n39853 );
buf ( n39855 , n39347 );
not ( n39856 , n39855 );
or ( n39857 , n39854 , n39856 );
buf ( n39858 , n37476 );
not ( n39859 , n39858 );
buf ( n39860 , n37146 );
not ( n39861 , n39860 );
buf ( n39862 , n39861 );
not ( n39863 , n39862 );
or ( n39864 , n39859 , n39863 );
buf ( n39865 , n38436 );
buf ( n39866 , n37475 );
nand ( n39867 , n39865 , n39866 );
buf ( n39868 , n39867 );
buf ( n39869 , n39868 );
nand ( n39870 , n39864 , n39869 );
buf ( n39871 , n39870 );
buf ( n39872 , n39871 );
buf ( n39873 , n37517 );
nand ( n39874 , n39872 , n39873 );
buf ( n39875 , n39874 );
buf ( n39876 , n39875 );
nand ( n39877 , n39857 , n39876 );
buf ( n39878 , n39877 );
buf ( n39879 , n39878 );
not ( n39880 , n39879 );
buf ( n39881 , n39880 );
buf ( n39882 , n39881 );
not ( n39883 , n39882 );
buf ( n39884 , n39313 );
buf ( n39885 , n38150 );
and ( n39886 , n39884 , n39885 );
buf ( n39887 , n37330 );
not ( n39888 , n39887 );
buf ( n39889 , n36396 );
not ( n39890 , n39889 );
buf ( n39891 , n39890 );
buf ( n39892 , n39891 );
not ( n39893 , n39892 );
or ( n39894 , n39888 , n39893 );
buf ( n39895 , n36396 );
not ( n39896 , n39895 );
buf ( n39897 , n39896 );
buf ( n39898 , n39897 );
not ( n39899 , n39898 );
buf ( n39900 , n37329 );
nand ( n39901 , n39899 , n39900 );
buf ( n39902 , n39901 );
buf ( n39903 , n39902 );
nand ( n39904 , n39894 , n39903 );
buf ( n39905 , n39904 );
buf ( n39906 , n39905 );
not ( n39907 , n39906 );
buf ( n39908 , n37406 );
nor ( n39909 , n39907 , n39908 );
buf ( n39910 , n39909 );
buf ( n39911 , n39910 );
nor ( n39912 , n39886 , n39911 );
buf ( n39913 , n39912 );
buf ( n39914 , n39913 );
not ( n39915 , n39914 );
or ( n39916 , n39883 , n39915 );
buf ( n39917 , n38413 );
not ( n39918 , n39917 );
buf ( n39919 , n36565 );
not ( n39920 , n39919 );
or ( n39921 , n39918 , n39920 );
buf ( n39922 , n36559 );
buf ( n39923 , n39922 );
buf ( n39924 , n39923 );
buf ( n39925 , n39924 );
not ( n39926 , n39925 );
buf ( n39927 , n39926 );
buf ( n39928 , n39927 );
buf ( n39929 , n39928 );
buf ( n39930 , n39929 );
buf ( n39931 , n39930 );
not ( n39932 , n39931 );
buf ( n39933 , n38420 );
nand ( n39934 , n39932 , n39933 );
buf ( n39935 , n39934 );
buf ( n39936 , n39935 );
nand ( n39937 , n39921 , n39936 );
buf ( n39938 , n39937 );
buf ( n39939 , n39938 );
buf ( n39940 , n38775 );
and ( n39941 , n39939 , n39940 );
buf ( n39942 , n39166 );
not ( n39943 , n39942 );
buf ( n39944 , n38383 );
nor ( n39945 , n39943 , n39944 );
buf ( n39946 , n39945 );
buf ( n39947 , n39946 );
nor ( n39948 , n39941 , n39947 );
buf ( n39949 , n39948 );
buf ( n39950 , n39949 );
not ( n39951 , n39950 );
buf ( n39952 , n39951 );
buf ( n39953 , n39952 );
nand ( n39954 , n39916 , n39953 );
buf ( n39955 , n39954 );
buf ( n39956 , n39955 );
buf ( n39957 , n39913 );
not ( n39958 , n39957 );
buf ( n39959 , n39958 );
buf ( n39960 , n39959 );
buf ( n39961 , n39878 );
nand ( n39962 , n39960 , n39961 );
buf ( n39963 , n39962 );
buf ( n39964 , n39963 );
nand ( n39965 , n39956 , n39964 );
buf ( n39966 , n39965 );
buf ( n39967 , n39966 );
xor ( n39968 , n39852 , n39967 );
buf ( n39969 , n39968 );
buf ( n39970 , n39969 );
not ( n39971 , n39970 );
not ( n39972 , n25098 );
buf ( n39973 , n25158 );
not ( n39974 , n39973 );
or ( n39975 , n39972 , n39974 );
or ( n39976 , n39973 , n25098 );
nand ( n39977 , n39975 , n39976 );
buf ( n39978 , n39977 );
buf ( n39979 , n39978 );
buf ( n39980 , n39979 );
buf ( n39981 , n39980 );
not ( n39982 , n39981 );
buf ( n39983 , n39982 );
buf ( n39984 , n39983 );
buf ( n39985 , n39984 );
buf ( n39986 , n39985 );
buf ( n39987 , n39986 );
not ( n39988 , n39987 );
buf ( n39989 , n39988 );
buf ( n39990 , n39989 );
not ( n39991 , n39990 );
and ( n39992 , n24091 , n25098 );
not ( n39993 , n24091 );
not ( n39994 , n25098 );
and ( n39995 , n39993 , n39994 );
nor ( n39996 , n39992 , n39995 );
nand ( n39997 , n39996 , n39977 );
buf ( n39998 , n39997 );
not ( n39999 , n39998 );
buf ( n40000 , n39999 );
buf ( n40001 , n40000 );
buf ( n40002 , n40001 );
buf ( n40003 , n40002 );
not ( n40004 , n40003 );
buf ( n40005 , n40004 );
buf ( n40006 , n40005 );
not ( n40007 , n40006 );
or ( n40008 , n39991 , n40007 );
not ( n40009 , n24092 );
not ( n40010 , n40009 );
buf ( n40011 , n40010 );
not ( n40012 , n40011 );
buf ( n40013 , n35971 );
not ( n40014 , n40013 );
or ( n40015 , n40012 , n40014 );
buf ( n40016 , n35970 );
buf ( n40017 , n40009 );
nand ( n40018 , n40016 , n40017 );
buf ( n40019 , n40018 );
buf ( n40020 , n40019 );
nand ( n40021 , n40015 , n40020 );
buf ( n40022 , n40021 );
buf ( n40023 , n40022 );
nand ( n40024 , n40008 , n40023 );
buf ( n40025 , n40024 );
buf ( n40026 , n40025 );
xor ( n40027 , n39792 , n39796 );
xor ( n40028 , n40027 , n39823 );
buf ( n40029 , n40028 );
buf ( n40030 , n40029 );
xor ( n40031 , n40026 , n40030 );
buf ( n40032 , n37452 );
not ( n40033 , n40032 );
buf ( n40034 , n39871 );
not ( n40035 , n40034 );
or ( n40036 , n40033 , n40035 );
buf ( n40037 , n37476 );
buf ( n40038 , n38447 );
and ( n40039 , n40037 , n40038 );
not ( n40040 , n40037 );
buf ( n40041 , n37971 );
and ( n40042 , n40040 , n40041 );
nor ( n40043 , n40039 , n40042 );
buf ( n40044 , n40043 );
buf ( n40045 , n40044 );
buf ( n40046 , n37517 );
nand ( n40047 , n40045 , n40046 );
buf ( n40048 , n40047 );
buf ( n40049 , n40048 );
nand ( n40050 , n40036 , n40049 );
buf ( n40051 , n40050 );
buf ( n40052 , n40051 );
and ( n40053 , n40031 , n40052 );
and ( n40054 , n40026 , n40030 );
or ( n40055 , n40053 , n40054 );
buf ( n40056 , n40055 );
buf ( n40057 , n40056 );
xor ( n40058 , n39828 , n39841 );
xor ( n40059 , n40058 , n39846 );
buf ( n40060 , n40059 );
buf ( n40061 , n40060 );
xor ( n40062 , n40057 , n40061 );
buf ( n40063 , n38775 );
not ( n40064 , n40063 );
buf ( n40065 , n36427 );
not ( n40066 , n40065 );
buf ( n40067 , n40066 );
and ( n40068 , n40067 , n38413 );
not ( n40069 , n40067 );
and ( n40070 , n40069 , n38420 );
or ( n40071 , n40068 , n40070 );
buf ( n40072 , n40071 );
not ( n40073 , n40072 );
or ( n40074 , n40064 , n40073 );
buf ( n40075 , n39938 );
buf ( n40076 , n38758 );
nand ( n40077 , n40075 , n40076 );
buf ( n40078 , n40077 );
buf ( n40079 , n40078 );
nand ( n40080 , n40074 , n40079 );
buf ( n40081 , n40080 );
buf ( n40082 , n40081 );
not ( n40083 , n40082 );
buf ( n40084 , n40083 );
buf ( n40085 , n40084 );
not ( n40086 , n40085 );
not ( n40087 , n37406 );
not ( n40088 , n37329 );
buf ( n40089 , n37078 );
not ( n40090 , n40089 );
or ( n40091 , n40088 , n40090 );
or ( n40092 , n40089 , n37329 );
nand ( n40093 , n40091 , n40092 );
not ( n40094 , n40093 );
not ( n40095 , n40094 );
and ( n40096 , n40087 , n40095 );
and ( n40097 , n39905 , n38150 );
nor ( n40098 , n40096 , n40097 );
buf ( n40099 , n40098 );
not ( n40100 , n40099 );
or ( n40101 , n40086 , n40100 );
xor ( n40102 , n39507 , n39536 );
xor ( n40103 , n40102 , n39559 );
buf ( n40104 , n40103 );
buf ( n40105 , n40104 );
nand ( n40106 , n40101 , n40105 );
buf ( n40107 , n40106 );
buf ( n40108 , n40107 );
not ( n40109 , n40098 );
buf ( n40110 , n40109 );
buf ( n40111 , n40081 );
nand ( n40112 , n40110 , n40111 );
buf ( n40113 , n40112 );
buf ( n40114 , n40113 );
nand ( n40115 , n40108 , n40114 );
buf ( n40116 , n40115 );
buf ( n40117 , n40116 );
and ( n40118 , n40062 , n40117 );
and ( n40119 , n40057 , n40061 );
or ( n40120 , n40118 , n40119 );
buf ( n40121 , n40120 );
buf ( n40122 , n40121 );
not ( n40123 , n40122 );
buf ( n40124 , n40123 );
buf ( n40125 , n40124 );
nand ( n40126 , n39971 , n40125 );
buf ( n40127 , n40126 );
buf ( n40128 , n40127 );
not ( n40129 , n40128 );
or ( n40130 , n39782 , n40129 );
buf ( n40131 , n39969 );
buf ( n40132 , n40121 );
nand ( n40133 , n40131 , n40132 );
buf ( n40134 , n40133 );
buf ( n40135 , n40134 );
nand ( n40136 , n40130 , n40135 );
buf ( n40137 , n40136 );
not ( n40138 , n40137 );
xor ( n40139 , n39183 , n39187 );
xor ( n40140 , n40139 , n39191 );
buf ( n40141 , n40140 );
buf ( n40142 , n40141 );
xor ( n40143 , n39786 , n39851 );
and ( n40144 , n40143 , n39967 );
and ( n40145 , n39786 , n39851 );
or ( n40146 , n40144 , n40145 );
buf ( n40147 , n40146 );
buf ( n40148 , n40147 );
xor ( n40149 , n40142 , n40148 );
xor ( n40150 , n39329 , n39436 );
xor ( n40151 , n40150 , n39441 );
buf ( n40152 , n40151 );
buf ( n40153 , n40152 );
xor ( n40154 , n40149 , n40153 );
buf ( n40155 , n40154 );
not ( n40156 , n40155 );
xor ( n40157 , n39469 , n39773 );
and ( n40158 , n40157 , n39778 );
and ( n40159 , n39469 , n39773 );
or ( n40160 , n40158 , n40159 );
buf ( n40161 , n40160 );
not ( n40162 , n40161 );
nand ( n40163 , n40156 , n40162 );
not ( n40164 , n40163 );
or ( n40165 , n40138 , n40164 );
buf ( n40166 , n40155 );
buf ( n40167 , n40161 );
nand ( n40168 , n40166 , n40167 );
buf ( n40169 , n40168 );
nand ( n40170 , n40165 , n40169 );
not ( n40171 , n40170 );
xor ( n40172 , n38958 , n39089 );
xor ( n40173 , n40172 , n39094 );
buf ( n40174 , n40173 );
xor ( n40175 , n40142 , n40148 );
and ( n40176 , n40175 , n40153 );
and ( n40177 , n40142 , n40148 );
or ( n40178 , n40176 , n40177 );
buf ( n40179 , n40178 );
xor ( n40180 , n40174 , n40179 );
xor ( n40181 , n39122 , n39196 );
xor ( n40182 , n40181 , n39446 );
buf ( n40183 , n40182 );
xor ( n40184 , n40180 , n40183 );
not ( n40185 , n40184 );
nand ( n40186 , n40171 , n40185 );
xor ( n40187 , n40174 , n40179 );
and ( n40188 , n40187 , n40183 );
and ( n40189 , n40174 , n40179 );
or ( n40190 , n40188 , n40189 );
xor ( n40191 , n39456 , n39457 );
buf ( n40192 , n40191 );
buf ( n40193 , n40192 );
buf ( n40194 , n39450 );
and ( n40195 , n40193 , n40194 );
not ( n40196 , n40193 );
buf ( n40197 , n39453 );
and ( n40198 , n40196 , n40197 );
nor ( n40199 , n40195 , n40198 );
buf ( n40200 , n40199 );
nor ( n40201 , n40190 , n40200 );
not ( n40202 , n40201 );
nand ( n40203 , n40186 , n40202 );
buf ( n40204 , n40203 );
nor ( n40205 , n39465 , n40204 );
buf ( n40206 , n40205 );
buf ( n40207 , n40206 );
buf ( n40208 , n38534 );
not ( n40209 , n40208 );
buf ( n40210 , n38636 );
nand ( n40211 , n40209 , n40210 );
buf ( n40212 , n40211 );
buf ( n40213 , n40212 );
not ( n40214 , n40213 );
buf ( n40215 , n38709 );
not ( n40216 , n40215 );
or ( n40217 , n40214 , n40216 );
buf ( n40218 , n38635 );
buf ( n40219 , n38534 );
nand ( n40220 , n40218 , n40219 );
buf ( n40221 , n40220 );
buf ( n40222 , n40221 );
nand ( n40223 , n40217 , n40222 );
buf ( n40224 , n40223 );
buf ( n40225 , n40224 );
not ( n40226 , n36456 );
and ( n40227 , n36363 , n37295 );
not ( n40228 , n36363 );
and ( n40229 , n40228 , n37298 );
or ( n40230 , n40227 , n40229 );
not ( n40231 , n40230 );
or ( n40232 , n40226 , n40231 );
buf ( n40233 , C1 );
nand ( n40234 , n40232 , n40233 );
not ( n40235 , n40234 );
buf ( n40236 , n36915 );
not ( n40237 , n40236 );
buf ( n40238 , n36935 );
not ( n40239 , n40238 );
buf ( n40240 , n37084 );
not ( n40241 , n40240 );
or ( n40242 , n40239 , n40241 );
buf ( n40243 , n37090 );
buf ( n40244 , n36951 );
nand ( n40245 , n40243 , n40244 );
buf ( n40246 , n40245 );
buf ( n40247 , n40246 );
nand ( n40248 , n40242 , n40247 );
buf ( n40249 , n40248 );
buf ( n40250 , n40249 );
not ( n40251 , n40250 );
or ( n40252 , n40237 , n40251 );
buf ( n40253 , n37948 );
buf ( n40254 , n36988 );
nand ( n40255 , n40253 , n40254 );
buf ( n40256 , n40255 );
buf ( n40257 , n40256 );
nand ( n40258 , n40252 , n40257 );
buf ( n40259 , n40258 );
and ( n40260 , n40235 , n40259 );
not ( n40261 , n40235 );
not ( n40262 , n40259 );
and ( n40263 , n40261 , n40262 );
nor ( n40264 , n40260 , n40263 );
buf ( n40265 , n38009 );
buf ( n40266 , n37875 );
and ( n40267 , n40265 , n40266 );
and ( n40268 , n36620 , n37882 );
not ( n40269 , n36620 );
and ( n40270 , n40269 , n37893 );
or ( n40271 , n40268 , n40270 );
buf ( n40272 , n40271 );
not ( n40273 , n40272 );
buf ( n40274 , n37922 );
not ( n40275 , n40274 );
buf ( n40276 , n40275 );
buf ( n40277 , n40276 );
nor ( n40278 , n40273 , n40277 );
buf ( n40279 , n40278 );
buf ( n40280 , n40279 );
nor ( n40281 , n40267 , n40280 );
buf ( n40282 , n40281 );
buf ( n40283 , n40282 );
not ( n40284 , n40283 );
buf ( n40285 , n40284 );
and ( n40286 , n40264 , n40285 );
not ( n40287 , n40264 );
and ( n40288 , n40287 , n40282 );
nor ( n40289 , n40286 , n40288 );
buf ( n40290 , n32972 );
not ( n40291 , n40290 );
buf ( n40292 , n33077 );
not ( n40293 , n40292 );
buf ( n40294 , n37971 );
not ( n40295 , n40294 );
or ( n40296 , n40293 , n40295 );
buf ( n40297 , n37977 );
buf ( n40298 , n33080 );
nand ( n40299 , n40297 , n40298 );
buf ( n40300 , n40299 );
buf ( n40301 , n40300 );
nand ( n40302 , n40296 , n40301 );
buf ( n40303 , n40302 );
buf ( n40304 , n40303 );
not ( n40305 , n40304 );
or ( n40306 , n40291 , n40305 );
buf ( n40307 , n38605 );
buf ( n40308 , n36107 );
nand ( n40309 , n40307 , n40308 );
buf ( n40310 , n40309 );
buf ( n40311 , n40310 );
nand ( n40312 , n40306 , n40311 );
buf ( n40313 , n40312 );
buf ( n40314 , n40313 );
not ( n40315 , n40314 );
buf ( n40316 , n36523 );
not ( n40317 , n40316 );
buf ( n40318 , n37278 );
not ( n40319 , n40318 );
buf ( n40320 , n40319 );
buf ( n40321 , n40320 );
not ( n40322 , n40321 );
or ( n40323 , n40317 , n40322 );
buf ( n40324 , n36533 );
not ( n40325 , n40324 );
buf ( n40326 , n38250 );
not ( n40327 , n40326 );
or ( n40328 , n40325 , n40327 );
buf ( n40329 , n38247 );
buf ( n40330 , n36578 );
nand ( n40331 , n40329 , n40330 );
buf ( n40332 , n40331 );
buf ( n40333 , n40332 );
nand ( n40334 , n40328 , n40333 );
buf ( n40335 , n40334 );
buf ( n40336 , n40335 );
buf ( n40337 , n36643 );
nand ( n40338 , n40336 , n40337 );
buf ( n40339 , n40338 );
buf ( n40340 , n40339 );
nand ( n40341 , n40323 , n40340 );
buf ( n40342 , n40341 );
buf ( n40343 , n40342 );
not ( n40344 , n40343 );
buf ( n40345 , n40344 );
buf ( n40346 , n40345 );
not ( n40347 , n40346 );
or ( n40348 , n40315 , n40347 );
buf ( n40349 , n40313 );
not ( n40350 , n40349 );
buf ( n40351 , n40350 );
buf ( n40352 , n40351 );
buf ( n40353 , n40342 );
nand ( n40354 , n40352 , n40353 );
buf ( n40355 , n40354 );
buf ( n40356 , n40355 );
nand ( n40357 , n40348 , n40356 );
buf ( n40358 , n40357 );
buf ( n40359 , n40358 );
buf ( n40360 , n37517 );
not ( n40361 , n40360 );
buf ( n40362 , n37483 );
not ( n40363 , n40362 );
or ( n40364 , n40361 , n40363 );
not ( n40365 , n37476 );
not ( n40366 , n35973 );
or ( n40367 , n40365 , n40366 );
buf ( n40368 , n35972 );
buf ( n40369 , n37545 );
nand ( n40370 , n40368 , n40369 );
buf ( n40371 , n40370 );
nand ( n40372 , n40367 , n40371 );
buf ( n40373 , n40372 );
buf ( n40374 , n37452 );
nand ( n40375 , n40373 , n40374 );
buf ( n40376 , n40375 );
buf ( n40377 , n40376 );
nand ( n40378 , n40364 , n40377 );
buf ( n40379 , n40378 );
buf ( n40380 , n40379 );
xor ( n40381 , n40359 , n40380 );
buf ( n40382 , n40381 );
xor ( n40383 , n40289 , n40382 );
buf ( n40384 , n38139 );
buf ( n40385 , n38016 );
or ( n40386 , n40384 , n40385 );
buf ( n40387 , n37991 );
nand ( n40388 , n40386 , n40387 );
buf ( n40389 , n40388 );
buf ( n40390 , n40389 );
buf ( n40391 , n38139 );
buf ( n40392 , n38016 );
nand ( n40393 , n40391 , n40392 );
buf ( n40394 , n40393 );
buf ( n40395 , n40394 );
nand ( n40396 , n40390 , n40395 );
buf ( n40397 , n40396 );
xnor ( n40398 , n40383 , n40397 );
buf ( n40399 , n40398 );
not ( n40400 , n40399 );
buf ( n40401 , n40400 );
buf ( n40402 , n40401 );
and ( n40403 , n40225 , n40402 );
not ( n40404 , n40225 );
buf ( n40405 , n40398 );
and ( n40406 , n40404 , n40405 );
nor ( n40407 , n40403 , n40406 );
buf ( n40408 , n40407 );
buf ( n40409 , n40408 );
buf ( n40410 , n37533 );
not ( n40411 , n40410 );
buf ( n40412 , n38142 );
not ( n40413 , n40412 );
or ( n40414 , n40411 , n40413 );
buf ( n40415 , n37933 );
nand ( n40416 , n40414 , n40415 );
buf ( n40417 , n40416 );
buf ( n40418 , n40417 );
nand ( n40419 , n38145 , n37532 );
buf ( n40420 , n40419 );
nand ( n40421 , n40418 , n40420 );
buf ( n40422 , n40421 );
not ( n40423 , n37526 );
not ( n40424 , n37303 );
or ( n40425 , n40423 , n40424 );
nand ( n40426 , n37521 , n37528 );
nand ( n40427 , n40425 , n40426 );
buf ( n40428 , n40427 );
buf ( n40429 , n38063 );
not ( n40430 , n40429 );
buf ( n40431 , n38074 );
not ( n40432 , n40431 );
buf ( n40433 , n36430 );
not ( n40434 , n40433 );
or ( n40435 , n40432 , n40434 );
buf ( n40436 , n36427 );
buf ( n40437 , n38083 );
nand ( n40438 , n40436 , n40437 );
buf ( n40439 , n40438 );
buf ( n40440 , n40439 );
nand ( n40441 , n40435 , n40440 );
buf ( n40442 , n40441 );
buf ( n40443 , n40442 );
not ( n40444 , n40443 );
or ( n40445 , n40430 , n40444 );
buf ( n40446 , n38089 );
buf ( n40447 , n38133 );
nand ( n40448 , n40446 , n40447 );
buf ( n40449 , n40448 );
buf ( n40450 , n40449 );
nand ( n40451 , n40445 , n40450 );
buf ( n40452 , n40451 );
buf ( n40453 , n40452 );
xor ( n40454 , n40428 , n40453 );
xor ( n40455 , n38616 , n38620 );
and ( n40456 , n40455 , n38632 );
and ( n40457 , n38616 , n38620 );
or ( n40458 , n40456 , n40457 );
buf ( n40459 , n40458 );
buf ( n40460 , n40459 );
xor ( n40461 , n40454 , n40460 );
buf ( n40462 , n40461 );
not ( n40463 , n40462 );
xor ( n40464 , n38585 , n38590 );
and ( n40465 , n40464 , n38634 );
and ( n40466 , n38585 , n38590 );
or ( n40467 , n40465 , n40466 );
buf ( n40468 , n40467 );
not ( n40469 , n40468 );
buf ( n40470 , n40469 );
not ( n40471 , n40470 );
or ( n40472 , n40463 , n40471 );
not ( n40473 , n40462 );
nand ( n40474 , n40473 , n40467 );
nand ( n40475 , n40472 , n40474 );
xnor ( n40476 , n40422 , n40475 );
buf ( n40477 , n40476 );
and ( n40478 , n40409 , n40477 );
not ( n40479 , n40409 );
buf ( n40480 , n40476 );
not ( n40481 , n40480 );
buf ( n40482 , n40481 );
buf ( n40483 , n40482 );
and ( n40484 , n40479 , n40483 );
nor ( n40485 , n40478 , n40484 );
buf ( n40486 , n40485 );
buf ( n40487 , n40486 );
xor ( n40488 , n38147 , n38718 );
and ( n40489 , n40488 , n39107 );
and ( n40490 , n38147 , n38718 );
or ( n40491 , n40489 , n40490 );
buf ( n40492 , n40491 );
buf ( n40493 , n40492 );
nand ( n40494 , n40487 , n40493 );
buf ( n40495 , n40494 );
buf ( n40496 , n40495 );
and ( n40497 , n40207 , n40496 );
buf ( n40498 , n40497 );
buf ( n40499 , n40498 );
buf ( n40500 , n32972 );
not ( n40501 , n40500 );
buf ( n40502 , n33083 );
not ( n40503 , n40502 );
buf ( n40504 , n36402 );
not ( n40505 , n40504 );
or ( n40506 , n40503 , n40505 );
buf ( n40507 , n36399 );
buf ( n40508 , n33080 );
nand ( n40509 , n40507 , n40508 );
buf ( n40510 , n40509 );
buf ( n40511 , n40510 );
nand ( n40512 , n40506 , n40511 );
buf ( n40513 , n40512 );
buf ( n40514 , n40513 );
not ( n40515 , n40514 );
or ( n40516 , n40501 , n40515 );
buf ( n40517 , n33083 );
not ( n40518 , n40517 );
buf ( n40519 , n37084 );
not ( n40520 , n40519 );
or ( n40521 , n40518 , n40520 );
buf ( n40522 , n37090 );
buf ( n40523 , n33080 );
nand ( n40524 , n40522 , n40523 );
buf ( n40525 , n40524 );
buf ( n40526 , n40525 );
nand ( n40527 , n40521 , n40526 );
buf ( n40528 , n40527 );
buf ( n40529 , n40528 );
buf ( n40530 , n36113 );
nand ( n40531 , n40529 , n40530 );
buf ( n40532 , n40531 );
buf ( n40533 , n40532 );
nand ( n40534 , n40516 , n40533 );
buf ( n40535 , n40534 );
buf ( n40536 , n40535 );
buf ( n40537 , n40276 );
not ( n40538 , n40537 );
buf ( n40539 , n37875 );
not ( n40540 , n40539 );
buf ( n40541 , n40540 );
buf ( n40542 , n40541 );
not ( n40543 , n40542 );
or ( n40544 , n40538 , n40543 );
buf ( n40545 , n37882 );
not ( n40546 , n40545 );
buf ( n40547 , n35973 );
not ( n40548 , n40547 );
or ( n40549 , n40546 , n40548 );
buf ( n40550 , n35972 );
buf ( n40551 , n37893 );
nand ( n40552 , n40550 , n40551 );
buf ( n40553 , n40552 );
buf ( n40554 , n40553 );
nand ( n40555 , n40549 , n40554 );
buf ( n40556 , n40555 );
buf ( n40557 , n40556 );
nand ( n40558 , n40544 , n40557 );
buf ( n40559 , n40558 );
buf ( n40560 , n40559 );
buf ( n40561 , n36456 );
not ( n40562 , n40561 );
buf ( n40563 , n36363 );
not ( n40564 , n40563 );
buf ( n40565 , n38221 );
not ( n40566 , n40565 );
or ( n40567 , n40564 , n40566 );
buf ( n40568 , n38227 );
buf ( n40569 , n36409 );
nand ( n40570 , n40568 , n40569 );
buf ( n40571 , n40570 );
buf ( n40572 , n40571 );
nand ( n40573 , n40567 , n40572 );
buf ( n40574 , n40573 );
buf ( n40575 , n40574 );
not ( n40576 , n40575 );
or ( n40577 , n40562 , n40576 );
and ( n40578 , n38250 , n36363 );
not ( n40579 , n38250 );
and ( n40580 , n40579 , n36409 );
or ( n40581 , n40578 , n40580 );
buf ( n40582 , C1 );
buf ( n40583 , n40582 );
nand ( n40584 , n40577 , n40583 );
buf ( n40585 , n40584 );
buf ( n40586 , n40585 );
xor ( n40587 , n40560 , n40586 );
buf ( n40588 , n38063 );
not ( n40589 , n40588 );
buf ( n40590 , n38074 );
not ( n40591 , n40590 );
buf ( n40592 , n36044 );
not ( n40593 , n40592 );
or ( n40594 , n40591 , n40593 );
buf ( n40595 , n38083 );
buf ( n40596 , n36057 );
nand ( n40597 , n40595 , n40596 );
buf ( n40598 , n40597 );
buf ( n40599 , n40598 );
nand ( n40600 , n40594 , n40599 );
buf ( n40601 , n40600 );
buf ( n40602 , n40601 );
not ( n40603 , n40602 );
or ( n40604 , n40589 , n40603 );
buf ( n40605 , n38074 );
not ( n40606 , n40605 );
buf ( n40607 , n36623 );
not ( n40608 , n40607 );
or ( n40609 , n40606 , n40608 );
buf ( n40610 , n36629 );
buf ( n40611 , n38083 );
nand ( n40612 , n40610 , n40611 );
buf ( n40613 , n40612 );
buf ( n40614 , n40613 );
nand ( n40615 , n40609 , n40614 );
buf ( n40616 , n40615 );
buf ( n40617 , n40616 );
buf ( n40618 , n38133 );
nand ( n40619 , n40617 , n40618 );
buf ( n40620 , n40619 );
buf ( n40621 , n40620 );
nand ( n40622 , n40604 , n40621 );
buf ( n40623 , n40622 );
buf ( n40624 , n40623 );
xor ( n40625 , n40587 , n40624 );
buf ( n40626 , n40625 );
buf ( n40627 , n40626 );
xor ( n40628 , n40536 , n40627 );
buf ( n40629 , n37875 );
not ( n40630 , n40629 );
buf ( n40631 , n37882 );
not ( n40632 , n40631 );
buf ( n40633 , n36041 );
not ( n40634 , n40633 );
or ( n40635 , n40632 , n40634 );
buf ( n40636 , n37481 );
buf ( n40637 , n37893 );
nand ( n40638 , n40636 , n40637 );
buf ( n40639 , n40638 );
buf ( n40640 , n40639 );
nand ( n40641 , n40635 , n40640 );
buf ( n40642 , n40641 );
buf ( n40643 , n40642 );
not ( n40644 , n40643 );
or ( n40645 , n40630 , n40644 );
buf ( n40646 , n40556 );
buf ( n40647 , n37922 );
nand ( n40648 , n40646 , n40647 );
buf ( n40649 , n40648 );
buf ( n40650 , n40649 );
nand ( n40651 , n40645 , n40650 );
buf ( n40652 , n40651 );
and ( n40653 , n37268 , n36363 );
not ( n40654 , n37268 );
and ( n40655 , n40654 , n36409 );
or ( n40656 , n40653 , n40655 );
buf ( n40657 , n40581 );
buf ( n40658 , n36456 );
nand ( n40659 , n40657 , n40658 );
buf ( n40660 , n40659 );
buf ( n40661 , n40660 );
nand ( n40662 , C1 , n40661 );
buf ( n40663 , n40662 );
xor ( n40664 , n40652 , n40663 );
buf ( n40665 , n33077 );
not ( n40666 , n40665 );
buf ( n40667 , n37149 );
not ( n40668 , n40667 );
or ( n40669 , n40666 , n40668 );
buf ( n40670 , n37153 );
buf ( n40671 , n33080 );
nand ( n40672 , n40670 , n40671 );
buf ( n40673 , n40672 );
buf ( n40674 , n40673 );
nand ( n40675 , n40669 , n40674 );
buf ( n40676 , n40675 );
buf ( n40677 , n40676 );
buf ( n40678 , n36113 );
nand ( n40679 , n40677 , n40678 );
buf ( n40680 , n40679 );
nand ( n40681 , n40528 , n32972 );
nand ( n40682 , n40680 , n40681 );
and ( n40683 , n40664 , n40682 );
and ( n40684 , n40652 , n40663 );
or ( n40685 , n40683 , n40684 );
buf ( n40686 , n40685 );
xnor ( n40687 , n40628 , n40686 );
buf ( n40688 , n40687 );
buf ( n40689 , n40688 );
not ( n40690 , n37514 );
not ( n40691 , n37449 );
or ( n40692 , n40690 , n40691 );
nand ( n40693 , n40692 , n40372 );
buf ( n40694 , n40693 );
not ( n40695 , n40694 );
buf ( n40696 , n37922 );
not ( n40697 , n40696 );
buf ( n40698 , n40642 );
not ( n40699 , n40698 );
or ( n40700 , n40697 , n40699 );
buf ( n40701 , n40271 );
buf ( n40702 , n37875 );
nand ( n40703 , n40701 , n40702 );
buf ( n40704 , n40703 );
buf ( n40705 , n40704 );
nand ( n40706 , n40700 , n40705 );
buf ( n40707 , n40706 );
buf ( n40708 , n40707 );
not ( n40709 , n40708 );
or ( n40710 , n40695 , n40709 );
buf ( n40711 , n40676 );
buf ( n40712 , n32972 );
and ( n40713 , n40711 , n40712 );
buf ( n40714 , n40303 );
not ( n40715 , n40714 );
buf ( n40716 , n36110 );
nor ( n40717 , n40715 , n40716 );
buf ( n40718 , n40717 );
buf ( n40719 , n40718 );
nor ( n40720 , n40713 , n40719 );
buf ( n40721 , n40720 );
buf ( n40722 , n40721 );
not ( n40723 , n40722 );
buf ( n40724 , n40707 );
not ( n40725 , n40724 );
buf ( n40726 , n40693 );
not ( n40727 , n40726 );
buf ( n40728 , n40727 );
buf ( n40729 , n40728 );
nand ( n40730 , n40725 , n40729 );
buf ( n40731 , n40730 );
buf ( n40732 , n40731 );
nand ( n40733 , n40723 , n40732 );
buf ( n40734 , n40733 );
buf ( n40735 , n40734 );
nand ( n40736 , n40710 , n40735 );
buf ( n40737 , n40736 );
not ( n40738 , n40737 );
xor ( n40739 , n40652 , n40663 );
xor ( n40740 , n40739 , n40682 );
not ( n40741 , n40740 );
nand ( n40742 , n40738 , n40741 );
buf ( n40743 , n40742 );
buf ( n40744 , n40234 );
buf ( n40745 , n36643 );
not ( n40746 , n40745 );
buf ( n40747 , n36578 );
buf ( n40748 , n38227 );
and ( n40749 , n40747 , n40748 );
not ( n40750 , n40747 );
buf ( n40751 , n38221 );
and ( n40752 , n40750 , n40751 );
nor ( n40753 , n40749 , n40752 );
buf ( n40754 , n40753 );
buf ( n40755 , n40754 );
not ( n40756 , n40755 );
buf ( n40757 , n40756 );
buf ( n40758 , n40757 );
not ( n40759 , n40758 );
or ( n40760 , n40746 , n40759 );
buf ( n40761 , n40335 );
buf ( n40762 , n36523 );
nand ( n40763 , n40761 , n40762 );
buf ( n40764 , n40763 );
buf ( n40765 , n40764 );
nand ( n40766 , n40760 , n40765 );
buf ( n40767 , n40766 );
buf ( n40768 , n40767 );
xor ( n40769 , n40744 , n40768 );
buf ( n40770 , n36456 );
not ( n40771 , n40770 );
buf ( n40772 , n40656 );
not ( n40773 , n40772 );
or ( n40774 , n40771 , n40773 );
buf ( n40775 , C1 );
buf ( n40776 , n40775 );
nand ( n40777 , n40774 , n40776 );
buf ( n40778 , n40777 );
buf ( n40779 , n40778 );
and ( n40780 , n40769 , n40779 );
and ( n40781 , n40744 , n40768 );
or ( n40782 , n40780 , n40781 );
buf ( n40783 , n40782 );
buf ( n40784 , n40783 );
and ( n40785 , n40743 , n40784 );
nor ( n40786 , n40741 , n40738 );
buf ( n40787 , n40786 );
nor ( n40788 , n40785 , n40787 );
buf ( n40789 , n40788 );
buf ( n40790 , n40789 );
not ( n40791 , n40790 );
buf ( n40792 , n36533 );
buf ( n40793 , n37977 );
and ( n40794 , n40792 , n40793 );
not ( n40795 , n40792 );
buf ( n40796 , n37971 );
and ( n40797 , n40795 , n40796 );
or ( n40798 , n40794 , n40797 );
buf ( n40799 , n40798 );
not ( n40800 , n40799 );
not ( n40801 , n36706 );
and ( n40802 , n40800 , n40801 );
buf ( n40803 , n40754 );
buf ( n40804 , n36688 );
nor ( n40805 , n40803 , n40804 );
buf ( n40806 , n40805 );
nor ( n40807 , n40802 , n40806 );
not ( n40808 , n40807 );
not ( n40809 , n40616 );
not ( n40810 , n38063 );
or ( n40811 , n40809 , n40810 );
buf ( n40812 , n36565 );
buf ( n40813 , n38074 );
and ( n40814 , n40812 , n40813 );
buf ( n40815 , n37543 );
buf ( n40816 , n38083 );
and ( n40817 , n40815 , n40816 );
nor ( n40818 , n40814 , n40817 );
buf ( n40819 , n40818 );
not ( n40820 , n40819 );
nand ( n40821 , n40820 , n38133 );
nand ( n40822 , n40811 , n40821 );
not ( n40823 , n40822 );
or ( n40824 , n40808 , n40823 );
or ( n40825 , n40822 , n40807 );
buf ( n40826 , n36988 );
not ( n40827 , n40826 );
and ( n40828 , n37887 , n36951 );
not ( n40829 , n37887 );
and ( n40830 , n40829 , n36935 );
nor ( n40831 , n40828 , n40830 );
buf ( n40832 , n40831 );
not ( n40833 , n40832 );
or ( n40834 , n40827 , n40833 );
and ( n40835 , n36430 , n36935 );
not ( n40836 , n36430 );
and ( n40837 , n40836 , n36951 );
or ( n40838 , n40835 , n40837 );
buf ( n40839 , n40838 );
buf ( n40840 , n36915 );
nand ( n40841 , n40839 , n40840 );
buf ( n40842 , n40841 );
buf ( n40843 , n40842 );
nand ( n40844 , n40834 , n40843 );
buf ( n40845 , n40844 );
not ( n40846 , n40845 );
not ( n40847 , n40846 );
nand ( n40848 , n40825 , n40847 );
nand ( n40849 , n40824 , n40848 );
not ( n40850 , n40849 );
buf ( n40851 , n36643 );
not ( n40852 , n40851 );
buf ( n40853 , n36533 );
not ( n40854 , n40853 );
buf ( n40855 , n37149 );
not ( n40856 , n40855 );
or ( n40857 , n40854 , n40856 );
buf ( n40858 , n37153 );
buf ( n40859 , n36578 );
nand ( n40860 , n40858 , n40859 );
buf ( n40861 , n40860 );
buf ( n40862 , n40861 );
nand ( n40863 , n40857 , n40862 );
buf ( n40864 , n40863 );
buf ( n40865 , n40864 );
not ( n40866 , n40865 );
or ( n40867 , n40852 , n40866 );
buf ( n40868 , n40799 );
not ( n40869 , n40868 );
buf ( n40870 , n36523 );
nand ( n40871 , n40869 , n40870 );
buf ( n40872 , n40871 );
buf ( n40873 , n40872 );
nand ( n40874 , n40867 , n40873 );
buf ( n40875 , n40874 );
xor ( n40876 , n40807 , n40875 );
buf ( n40877 , n36988 );
not ( n40878 , n40877 );
buf ( n40879 , n40838 );
not ( n40880 , n40879 );
or ( n40881 , n40878 , n40880 );
and ( n40882 , n36568 , n36935 );
not ( n40883 , n36568 );
and ( n40884 , n40883 , n36951 );
or ( n40885 , n40882 , n40884 );
buf ( n40886 , n40885 );
buf ( n40887 , n36915 );
nand ( n40888 , n40886 , n40887 );
buf ( n40889 , n40888 );
buf ( n40890 , n40889 );
nand ( n40891 , n40881 , n40890 );
buf ( n40892 , n40891 );
xor ( n40893 , n40876 , n40892 );
not ( n40894 , n40893 );
or ( n40895 , n40850 , n40894 );
or ( n40896 , n40893 , n40849 );
nand ( n40897 , n40895 , n40896 );
buf ( n40898 , n40897 );
not ( n40899 , n40898 );
and ( n40900 , n40791 , n40899 );
buf ( n40901 , n40789 );
buf ( n40902 , n40897 );
and ( n40903 , n40901 , n40902 );
nor ( n40904 , n40900 , n40903 );
buf ( n40905 , n40904 );
buf ( n40906 , n40905 );
xor ( n40907 , n40689 , n40906 );
buf ( n40908 , n40234 );
not ( n40909 , n40908 );
buf ( n40910 , n40282 );
not ( n40911 , n40910 );
or ( n40912 , n40909 , n40911 );
buf ( n40913 , n40259 );
nand ( n40914 , n40912 , n40913 );
buf ( n40915 , n40914 );
buf ( n40916 , n40915 );
buf ( n40917 , n40234 );
not ( n40918 , n40917 );
buf ( n40919 , n40285 );
nand ( n40920 , n40918 , n40919 );
buf ( n40921 , n40920 );
buf ( n40922 , n40921 );
and ( n40923 , n40916 , n40922 );
buf ( n40924 , n40923 );
not ( n40925 , n40924 );
xor ( n40926 , n40728 , n40707 );
xnor ( n40927 , n40926 , n40721 );
not ( n40928 , n40927 );
and ( n40929 , n40925 , n40928 );
buf ( n40930 , n40927 );
buf ( n40931 , n40924 );
nand ( n40932 , n40930 , n40931 );
buf ( n40933 , n40932 );
xor ( n40934 , n40744 , n40768 );
xor ( n40935 , n40934 , n40779 );
buf ( n40936 , n40935 );
and ( n40937 , n40933 , n40936 );
nor ( n40938 , n40929 , n40937 );
buf ( n40939 , n40938 );
not ( n40940 , n40939 );
buf ( n40941 , n40940 );
buf ( n40942 , n40819 );
not ( n40943 , n40942 );
buf ( n40944 , n38733 );
not ( n40945 , n40944 );
and ( n40946 , n40943 , n40945 );
buf ( n40947 , n40442 );
buf ( n40948 , n38133 );
and ( n40949 , n40947 , n40948 );
nor ( n40950 , n40946 , n40949 );
buf ( n40951 , n40950 );
buf ( n40952 , n40951 );
not ( n40953 , n40952 );
buf ( n40954 , n36915 );
not ( n40955 , n40954 );
buf ( n40956 , n40831 );
not ( n40957 , n40956 );
or ( n40958 , n40955 , n40957 );
buf ( n40959 , n40249 );
buf ( n40960 , n36988 );
nand ( n40961 , n40959 , n40960 );
buf ( n40962 , n40961 );
buf ( n40963 , n40962 );
nand ( n40964 , n40958 , n40963 );
buf ( n40965 , n40964 );
buf ( n40966 , n40965 );
not ( n40967 , n40966 );
buf ( n40968 , n40967 );
buf ( n40969 , n40968 );
not ( n40970 , n40969 );
or ( n40971 , n40953 , n40970 );
buf ( n40972 , n40345 );
buf ( n40973 , n40351 );
nand ( n40974 , n40972 , n40973 );
buf ( n40975 , n40974 );
not ( n40976 , n40975 );
not ( n40977 , n40379 );
or ( n40978 , n40976 , n40977 );
or ( n40979 , n40345 , n40351 );
nand ( n40980 , n40978 , n40979 );
buf ( n40981 , n40980 );
nand ( n40982 , n40971 , n40981 );
buf ( n40983 , n40982 );
buf ( n40984 , n40951 );
not ( n40985 , n40984 );
buf ( n40986 , n40965 );
nand ( n40987 , n40985 , n40986 );
buf ( n40988 , n40987 );
nand ( n40989 , n40983 , n40988 );
xor ( n40990 , n40807 , n40846 );
xnor ( n40991 , n40990 , n40822 );
or ( n40992 , n40989 , n40991 );
and ( n40993 , n40941 , n40992 );
and ( n40994 , n40991 , n40989 );
nor ( n40995 , n40993 , n40994 );
buf ( n40996 , n40995 );
xor ( n40997 , n40907 , n40996 );
buf ( n40998 , n40997 );
not ( n40999 , n40741 );
and ( n41000 , n40783 , n40738 );
not ( n41001 , n40783 );
and ( n41002 , n41001 , n40737 );
or ( n41003 , n41000 , n41002 );
not ( n41004 , n41003 );
or ( n41005 , n40999 , n41004 );
or ( n41006 , n41003 , n40741 );
nand ( n41007 , n41005 , n41006 );
not ( n41008 , n41007 );
not ( n41009 , n40938 );
xor ( n41010 , n40991 , n40989 );
not ( n41011 , n41010 );
or ( n41012 , n41009 , n41011 );
or ( n41013 , n40938 , n41010 );
nand ( n41014 , n41012 , n41013 );
not ( n41015 , n41014 );
and ( n41016 , n41008 , n41015 );
buf ( n41017 , n40397 );
buf ( n41018 , n40382 );
or ( n41019 , n41017 , n41018 );
buf ( n41020 , n40289 );
nand ( n41021 , n41019 , n41020 );
buf ( n41022 , n41021 );
buf ( n41023 , n41022 );
buf ( n41024 , n40397 );
buf ( n41025 , n40382 );
nand ( n41026 , n41024 , n41025 );
buf ( n41027 , n41026 );
buf ( n41028 , n41027 );
nand ( n41029 , n41023 , n41028 );
buf ( n41030 , n41029 );
not ( n41031 , n41030 );
xor ( n41032 , n40951 , n40965 );
xor ( n41033 , n41032 , n40980 );
nand ( n41034 , n41031 , n41033 );
buf ( n41035 , n41034 );
xor ( n41036 , n40428 , n40453 );
and ( n41037 , n41036 , n40460 );
and ( n41038 , n40428 , n40453 );
or ( n41039 , n41037 , n41038 );
buf ( n41040 , n41039 );
buf ( n41041 , n41040 );
buf ( n41042 , n41041 );
and ( n41043 , n41035 , n41042 );
not ( n41044 , n41030 );
nor ( n41045 , n41044 , n41033 );
buf ( n41046 , n41045 );
nor ( n41047 , n41043 , n41046 );
buf ( n41048 , n41047 );
nor ( n41049 , n41016 , n41048 );
and ( n41050 , n41007 , n41014 );
nor ( n41051 , n41049 , n41050 );
nand ( n41052 , n40998 , n41051 );
buf ( n41053 , n41052 );
not ( n41054 , n40849 );
nand ( n41055 , n41054 , n40893 );
buf ( n41056 , n41055 );
not ( n41057 , n41056 );
buf ( n41058 , n40789 );
not ( n41059 , n41058 );
buf ( n41060 , n41059 );
buf ( n41061 , n41060 );
not ( n41062 , n41061 );
or ( n41063 , n41057 , n41062 );
not ( n41064 , n40893 );
nand ( n41065 , n41064 , n40849 );
buf ( n41066 , n41065 );
nand ( n41067 , n41063 , n41066 );
buf ( n41068 , n41067 );
buf ( n41069 , n41068 );
buf ( n41070 , n40535 );
not ( n41071 , n41070 );
buf ( n41072 , n40685 );
not ( n41073 , n41072 );
or ( n41074 , n41071 , n41073 );
buf ( n41075 , n40535 );
buf ( n41076 , n40685 );
or ( n41077 , n41075 , n41076 );
buf ( n41078 , n40626 );
nand ( n41079 , n41077 , n41078 );
buf ( n41080 , n41079 );
buf ( n41081 , n41080 );
nand ( n41082 , n41074 , n41081 );
buf ( n41083 , n41082 );
buf ( n41084 , n41083 );
not ( n41085 , n41084 );
buf ( n41086 , n40807 );
not ( n41087 , n41086 );
buf ( n41088 , n40875 );
not ( n41089 , n41088 );
buf ( n41090 , n41089 );
buf ( n41091 , n41090 );
not ( n41092 , n41091 );
or ( n41093 , n41087 , n41092 );
buf ( n41094 , n40892 );
nand ( n41095 , n41093 , n41094 );
buf ( n41096 , n41095 );
buf ( n41097 , n41096 );
buf ( n41098 , n40807 );
not ( n41099 , n41098 );
buf ( n41100 , n40875 );
nand ( n41101 , n41099 , n41100 );
buf ( n41102 , n41101 );
buf ( n41103 , n41102 );
nand ( n41104 , n41097 , n41103 );
buf ( n41105 , n41104 );
buf ( n41106 , n41105 );
buf ( n41107 , n38133 );
not ( n41108 , n41107 );
buf ( n41109 , n40601 );
not ( n41110 , n41109 );
or ( n41111 , n41108 , n41110 );
buf ( n41112 , n38074 );
not ( n41113 , n41112 );
buf ( n41114 , n35973 );
not ( n41115 , n41114 );
or ( n41116 , n41113 , n41115 );
buf ( n41117 , n35979 );
buf ( n41118 , n38083 );
nand ( n41119 , n41117 , n41118 );
buf ( n41120 , n41119 );
buf ( n41121 , n41120 );
nand ( n41122 , n41116 , n41121 );
buf ( n41123 , n41122 );
buf ( n41124 , n41123 );
buf ( n41125 , n38063 );
nand ( n41126 , n41124 , n41125 );
buf ( n41127 , n41126 );
buf ( n41128 , n41127 );
nand ( n41129 , n41111 , n41128 );
buf ( n41130 , n41129 );
buf ( n41131 , n41130 );
and ( n41132 , n39280 , n36363 );
not ( n41133 , n39280 );
and ( n41134 , n41133 , n36409 );
or ( n41135 , n41132 , n41134 );
buf ( n41136 , n41135 );
buf ( n41137 , n36456 );
nand ( n41138 , n41136 , n41137 );
buf ( n41139 , n41138 );
buf ( n41140 , n41139 );
nand ( n41141 , C1 , n41140 );
buf ( n41142 , n41141 );
buf ( n41143 , n41142 );
not ( n41144 , n41143 );
buf ( n41145 , n41144 );
buf ( n41146 , n41145 );
xor ( n41147 , n41131 , n41146 );
buf ( n41148 , n36988 );
not ( n41149 , n41148 );
buf ( n41150 , n40885 );
not ( n41151 , n41150 );
or ( n41152 , n41149 , n41151 );
buf ( n41153 , n36935 );
not ( n41154 , n41153 );
buf ( n41155 , n36623 );
not ( n41156 , n41155 );
or ( n41157 , n41154 , n41156 );
buf ( n41158 , n36629 );
buf ( n41159 , n36951 );
nand ( n41160 , n41158 , n41159 );
buf ( n41161 , n41160 );
buf ( n41162 , n41161 );
nand ( n41163 , n41157 , n41162 );
buf ( n41164 , n41163 );
buf ( n41165 , n41164 );
buf ( n41166 , n36915 );
nand ( n41167 , n41165 , n41166 );
buf ( n41168 , n41167 );
buf ( n41169 , n41168 );
nand ( n41170 , n41152 , n41169 );
buf ( n41171 , n41170 );
buf ( n41172 , n41171 );
xor ( n41173 , n41147 , n41172 );
buf ( n41174 , n41173 );
buf ( n41175 , n41174 );
xor ( n41176 , n41106 , n41175 );
buf ( n41177 , n36643 );
not ( n41178 , n41177 );
buf ( n41179 , n36533 );
not ( n41180 , n41179 );
buf ( n41181 , n37084 );
not ( n41182 , n41181 );
or ( n41183 , n41180 , n41182 );
buf ( n41184 , n37090 );
buf ( n41185 , n36578 );
nand ( n41186 , n41184 , n41185 );
buf ( n41187 , n41186 );
buf ( n41188 , n41187 );
nand ( n41189 , n41183 , n41188 );
buf ( n41190 , n41189 );
buf ( n41191 , n41190 );
not ( n41192 , n41191 );
or ( n41193 , n41178 , n41192 );
buf ( n41194 , n40864 );
buf ( n41195 , n36523 );
nand ( n41196 , n41194 , n41195 );
buf ( n41197 , n41196 );
buf ( n41198 , n41197 );
nand ( n41199 , n41193 , n41198 );
buf ( n41200 , n41199 );
buf ( n41201 , n41200 );
xor ( n41202 , n40560 , n40586 );
and ( n41203 , n41202 , n40624 );
and ( n41204 , n40560 , n40586 );
or ( n41205 , n41203 , n41204 );
buf ( n41206 , n41205 );
buf ( n41207 , n41206 );
xor ( n41208 , n41201 , n41207 );
buf ( n41209 , n36113 );
not ( n41210 , n41209 );
buf ( n41211 , n40513 );
not ( n41212 , n41211 );
or ( n41213 , n41210 , n41212 );
and ( n41214 , n36430 , n33083 );
not ( n41215 , n36430 );
and ( n41216 , n41215 , n33080 );
or ( n41217 , n41214 , n41216 );
buf ( n41218 , n41217 );
buf ( n41219 , n32972 );
nand ( n41220 , n41218 , n41219 );
buf ( n41221 , n41220 );
buf ( n41222 , n41221 );
nand ( n41223 , n41213 , n41222 );
buf ( n41224 , n41223 );
buf ( n41225 , n41224 );
xor ( n41226 , n41208 , n41225 );
buf ( n41227 , n41226 );
buf ( n41228 , n41227 );
xor ( n41229 , n41176 , n41228 );
buf ( n41230 , n41229 );
buf ( n41231 , n41230 );
not ( n41232 , n41231 );
buf ( n41233 , n41232 );
buf ( n41234 , n41233 );
not ( n41235 , n41234 );
or ( n41236 , n41085 , n41235 );
buf ( n41237 , n41230 );
buf ( n41238 , n41083 );
not ( n41239 , n41238 );
buf ( n41240 , n41239 );
buf ( n41241 , n41240 );
nand ( n41242 , n41237 , n41241 );
buf ( n41243 , n41242 );
buf ( n41244 , n41243 );
nand ( n41245 , n41236 , n41244 );
buf ( n41246 , n41245 );
buf ( n41247 , n41246 );
not ( n41248 , n41247 );
xor ( n41249 , n41069 , n41248 );
buf ( n41250 , n41249 );
buf ( n41251 , n41250 );
xor ( n41252 , n40689 , n40906 );
and ( n41253 , n41252 , n40996 );
and ( n41254 , n40689 , n40906 );
or ( n41255 , n41253 , n41254 );
buf ( n41256 , n41255 );
buf ( n41257 , n41256 );
nand ( n41258 , n41251 , n41257 );
buf ( n41259 , n41258 );
buf ( n41260 , n41259 );
nand ( n41261 , n41053 , n41260 );
buf ( n41262 , n41261 );
buf ( n41263 , n41262 );
xor ( n41264 , n41007 , n41014 );
xnor ( n41265 , n41264 , n41048 );
buf ( n41266 , n41265 );
xor ( n41267 , n40924 , n40927 );
xor ( n41268 , n41267 , n40936 );
buf ( n41269 , n41268 );
and ( n41270 , n41033 , n41040 );
not ( n41271 , n41033 );
not ( n41272 , n41040 );
and ( n41273 , n41271 , n41272 );
nor ( n41274 , n41270 , n41273 );
xnor ( n41275 , n41030 , n41274 );
buf ( n41276 , n41275 );
xor ( n41277 , n41269 , n41276 );
buf ( n41278 , n40473 );
buf ( n41279 , n40470 );
nand ( n41280 , n41278 , n41279 );
buf ( n41281 , n41280 );
buf ( n41282 , n41281 );
not ( n41283 , n41282 );
buf ( n41284 , n40422 );
not ( n41285 , n41284 );
or ( n41286 , n41283 , n41285 );
buf ( n41287 , n40462 );
buf ( n41288 , n40467 );
nand ( n41289 , n41287 , n41288 );
buf ( n41290 , n41289 );
buf ( n41291 , n41290 );
nand ( n41292 , n41286 , n41291 );
buf ( n41293 , n41292 );
buf ( n41294 , n41293 );
and ( n41295 , n41277 , n41294 );
and ( n41296 , n41269 , n41276 );
or ( n41297 , n41295 , n41296 );
buf ( n41298 , n41297 );
buf ( n41299 , n41298 );
nor ( n41300 , n41266 , n41299 );
buf ( n41301 , n41300 );
not ( n41302 , n41301 );
not ( n41303 , n40401 );
not ( n41304 , n40482 );
or ( n41305 , n41303 , n41304 );
buf ( n41306 , n40398 );
not ( n41307 , n41306 );
buf ( n41308 , n40476 );
not ( n41309 , n41308 );
or ( n41310 , n41307 , n41309 );
buf ( n41311 , n40224 );
nand ( n41312 , n41310 , n41311 );
buf ( n41313 , n41312 );
nand ( n41314 , n41305 , n41313 );
xor ( n41315 , n41269 , n41276 );
xor ( n41316 , n41315 , n41294 );
buf ( n41317 , n41316 );
or ( n41318 , n41314 , n41317 );
nand ( n41319 , n41302 , n41318 );
buf ( n41320 , n41319 );
nor ( n41321 , n41263 , n41320 );
buf ( n41322 , n41321 );
buf ( n41323 , n41322 );
and ( n41324 , n40499 , n41323 );
buf ( n41325 , n41324 );
buf ( n41326 , n41240 );
not ( n41327 , n41326 );
buf ( n41328 , n41233 );
not ( n41329 , n41328 );
or ( n41330 , n41327 , n41329 );
buf ( n41331 , n41068 );
nand ( n41332 , n41330 , n41331 );
buf ( n41333 , n41332 );
buf ( n41334 , n41333 );
buf ( n41335 , n41230 );
buf ( n41336 , n41083 );
nand ( n41337 , n41335 , n41336 );
buf ( n41338 , n41337 );
buf ( n41339 , n41338 );
nand ( n41340 , n41334 , n41339 );
buf ( n41341 , n41340 );
buf ( n41342 , n41341 );
buf ( n41343 , n36456 );
not ( n41344 , n41343 );
buf ( n41345 , n37160 );
not ( n41346 , n41345 );
or ( n41347 , n41344 , n41346 );
buf ( n41348 , C1 );
buf ( n41349 , n41348 );
nand ( n41350 , n41347 , n41349 );
buf ( n41351 , n41350 );
buf ( n41352 , n41351 );
buf ( n41353 , n36113 );
not ( n41354 , n41353 );
buf ( n41355 , n41217 );
not ( n41356 , n41355 );
or ( n41357 , n41354 , n41356 );
buf ( n41358 , n37118 );
buf ( n41359 , n32972 );
nand ( n41360 , n41358 , n41359 );
buf ( n41361 , n41360 );
buf ( n41362 , n41361 );
nand ( n41363 , n41357 , n41362 );
buf ( n41364 , n41363 );
buf ( n41365 , n41364 );
xor ( n41366 , n41352 , n41365 );
buf ( n41367 , n36643 );
not ( n41368 , n41367 );
buf ( n41369 , n37189 );
not ( n41370 , n41369 );
or ( n41371 , n41368 , n41370 );
buf ( n41372 , n41190 );
buf ( n41373 , n36523 );
nand ( n41374 , n41372 , n41373 );
buf ( n41375 , n41374 );
buf ( n41376 , n41375 );
nand ( n41377 , n41371 , n41376 );
buf ( n41378 , n41377 );
buf ( n41379 , n41378 );
xor ( n41380 , n41366 , n41379 );
buf ( n41381 , n41380 );
buf ( n41382 , n41381 );
xor ( n41383 , n41131 , n41146 );
and ( n41384 , n41383 , n41172 );
and ( n41385 , n41131 , n41146 );
or ( n41386 , n41384 , n41385 );
buf ( n41387 , n41386 );
buf ( n41388 , n41387 );
buf ( n41389 , n38733 );
not ( n41390 , n41389 );
buf ( n41391 , n39633 );
not ( n41392 , n41391 );
or ( n41393 , n41390 , n41392 );
buf ( n41394 , n41123 );
nand ( n41395 , n41393 , n41394 );
buf ( n41396 , n41395 );
buf ( n41397 , n41396 );
buf ( n41398 , n36915 );
not ( n41399 , n41398 );
buf ( n41400 , n36957 );
not ( n41401 , n41400 );
or ( n41402 , n41399 , n41401 );
buf ( n41403 , n41164 );
buf ( n41404 , n36988 );
nand ( n41405 , n41403 , n41404 );
buf ( n41406 , n41405 );
buf ( n41407 , n41406 );
nand ( n41408 , n41402 , n41407 );
buf ( n41409 , n41408 );
buf ( n41410 , n41409 );
xor ( n41411 , n41397 , n41410 );
buf ( n41412 , n41142 );
xor ( n41413 , n41411 , n41412 );
buf ( n41414 , n41413 );
buf ( n41415 , n41414 );
xor ( n41416 , n41388 , n41415 );
xor ( n41417 , n41201 , n41207 );
and ( n41418 , n41417 , n41225 );
and ( n41419 , n41201 , n41207 );
or ( n41420 , n41418 , n41419 );
buf ( n41421 , n41420 );
buf ( n41422 , n41421 );
xor ( n41423 , n41416 , n41422 );
buf ( n41424 , n41423 );
buf ( n41425 , n41424 );
xor ( n41426 , n41382 , n41425 );
xor ( n41427 , n41106 , n41175 );
and ( n41428 , n41427 , n41228 );
and ( n41429 , n41106 , n41175 );
or ( n41430 , n41428 , n41429 );
buf ( n41431 , n41430 );
buf ( n41432 , n41431 );
xor ( n41433 , n41426 , n41432 );
buf ( n41434 , n41433 );
buf ( n41435 , n41434 );
or ( n41436 , n41342 , n41435 );
buf ( n41437 , n41436 );
buf ( n41438 , n41437 );
xor ( n41439 , n41352 , n41365 );
and ( n41440 , n41439 , n41379 );
and ( n41441 , n41352 , n41365 );
or ( n41442 , n41440 , n41441 );
buf ( n41443 , n41442 );
buf ( n41444 , n41443 );
xor ( n41445 , n41388 , n41415 );
and ( n41446 , n41445 , n41422 );
and ( n41447 , n41388 , n41415 );
or ( n41448 , n41446 , n41447 );
buf ( n41449 , n41448 );
buf ( n41450 , n41449 );
xor ( n41451 , n41444 , n41450 );
xor ( n41452 , n41397 , n41410 );
and ( n41453 , n41452 , n41412 );
and ( n41454 , n41397 , n41410 );
or ( n41455 , n41453 , n41454 );
buf ( n41456 , n41455 );
xor ( n41457 , n41456 , n36994 );
buf ( n41458 , n37123 );
not ( n41459 , n41458 );
buf ( n41460 , n37170 );
not ( n41461 , n41460 );
or ( n41462 , n41459 , n41461 );
buf ( n41463 , n37164 );
buf ( n41464 , n37120 );
nand ( n41465 , n41463 , n41464 );
buf ( n41466 , n41465 );
buf ( n41467 , n41466 );
nand ( n41468 , n41462 , n41467 );
buf ( n41469 , n41468 );
buf ( n41470 , n41469 );
buf ( n41471 , n37199 );
xnor ( n41472 , n41470 , n41471 );
buf ( n41473 , n41472 );
xor ( n41474 , n41457 , n41473 );
buf ( n41475 , n41474 );
xor ( n41476 , n41451 , n41475 );
buf ( n41477 , n41476 );
buf ( n41478 , n41477 );
xor ( n41479 , n41382 , n41425 );
and ( n41480 , n41479 , n41432 );
and ( n41481 , n41382 , n41425 );
or ( n41482 , n41480 , n41481 );
buf ( n41483 , n41482 );
buf ( n41484 , n41483 );
nor ( n41485 , n41478 , n41484 );
buf ( n41486 , n41485 );
buf ( n41487 , n41486 );
not ( n41488 , n41487 );
buf ( n41489 , n41488 );
buf ( n41490 , n41489 );
nand ( n41491 , n41438 , n41490 );
buf ( n41492 , n41491 );
xor ( n41493 , n41444 , n41450 );
and ( n41494 , n41493 , n41475 );
and ( n41495 , n41444 , n41450 );
or ( n41496 , n41494 , n41495 );
buf ( n41497 , n41496 );
buf ( n41498 , n41497 );
not ( n41499 , n41498 );
buf ( n41500 , n37011 );
not ( n41501 , n41500 );
buf ( n41502 , n36865 );
not ( n41503 , n41502 );
or ( n41504 , n41501 , n41503 );
buf ( n41505 , n36865 );
buf ( n41506 , n37011 );
or ( n41507 , n41505 , n41506 );
nand ( n41508 , n41504 , n41507 );
buf ( n41509 , n41508 );
xnor ( n41510 , n41509 , n36994 );
buf ( n41511 , n41510 );
buf ( n41512 , n37098 );
not ( n41513 , n41512 );
buf ( n41514 , n37061 );
not ( n41515 , n41514 );
and ( n41516 , n41513 , n41515 );
buf ( n41517 , n37061 );
buf ( n41518 , n37098 );
and ( n41519 , n41517 , n41518 );
nor ( n41520 , n41516 , n41519 );
buf ( n41521 , n41520 );
xor ( n41522 , n41521 , n37205 );
buf ( n41523 , n41522 );
xor ( n41524 , n41511 , n41523 );
buf ( n41525 , n41473 );
buf ( n41526 , n36994 );
nand ( n41527 , n41525 , n41526 );
buf ( n41528 , n41527 );
buf ( n41529 , n41528 );
buf ( n41530 , n41456 );
and ( n41531 , n41529 , n41530 );
buf ( n41532 , n41473 );
buf ( n41533 , n36994 );
nor ( n41534 , n41532 , n41533 );
buf ( n41535 , n41534 );
buf ( n41536 , n41535 );
nor ( n41537 , n41531 , n41536 );
buf ( n41538 , n41537 );
buf ( n41539 , n41538 );
xor ( n41540 , n41524 , n41539 );
buf ( n41541 , n41540 );
buf ( n41542 , n41541 );
nand ( n41543 , n41499 , n41542 );
buf ( n41544 , n41543 );
buf ( n41545 , n41544 );
xor ( n41546 , n37021 , n37036 );
xor ( n41547 , n41546 , n37217 );
buf ( n41548 , n41547 );
buf ( n41549 , n41548 );
not ( n41550 , n41549 );
xor ( n41551 , n41511 , n41523 );
and ( n41552 , n41551 , n41539 );
and ( n41553 , n41511 , n41523 );
or ( n41554 , n41552 , n41553 );
buf ( n41555 , n41554 );
buf ( n41556 , n41555 );
nand ( n41557 , n41550 , n41556 );
buf ( n41558 , n41557 );
buf ( n41559 , n41558 );
nand ( n41560 , n41545 , n41559 );
buf ( n41561 , n41560 );
nor ( n41562 , n41492 , n41561 );
nand ( n41563 , n41325 , n41562 );
buf ( n41564 , n41563 );
not ( n41565 , n41564 );
buf ( n41566 , n41565 );
not ( n41567 , n41566 );
buf ( n41568 , n25379 );
buf ( n41569 , n41568 );
buf ( n41570 , n41569 );
xnor ( n41571 , n41570 , n24978 );
buf ( n41572 , n41571 );
not ( n41573 , n41572 );
buf ( n41574 , n41573 );
buf ( n41575 , n41574 );
not ( n41576 , n41575 );
buf ( n41577 , n41576 );
buf ( n41578 , n41577 );
not ( n41579 , n41578 );
buf ( n41580 , n24978 );
not ( n41581 , n41580 );
buf ( n41582 , n41581 );
buf ( n41583 , n41582 );
buf ( n41584 , n25336 );
not ( n41585 , n41584 );
buf ( n41586 , n41585 );
buf ( n41587 , n41586 );
and ( n41588 , n41583 , n41587 );
not ( n41589 , n41583 );
buf ( n41590 , n25336 );
and ( n41591 , n41589 , n41590 );
nor ( n41592 , n41588 , n41591 );
buf ( n41593 , n41592 );
nand ( n41594 , n41593 , n41571 );
buf ( n41595 , n41594 );
not ( n41596 , n41595 );
buf ( n41597 , n41596 );
not ( n41598 , n41597 );
buf ( n41599 , n41598 );
buf ( n41600 , n41599 );
not ( n41601 , n41600 );
or ( n41602 , n41579 , n41601 );
nand ( n41603 , n25329 , n25332 );
and ( n41604 , n41603 , n25335 );
not ( n41605 , n41604 );
buf ( n41606 , n41605 );
buf ( n41607 , n41606 );
buf ( n41608 , n41607 );
buf ( n41609 , n41608 );
not ( n41610 , n41609 );
buf ( n41611 , n41610 );
buf ( n41612 , n41611 );
not ( n41613 , n41612 );
buf ( n41614 , n39005 );
not ( n41615 , n41614 );
or ( n41616 , n41613 , n41615 );
buf ( n41617 , n39005 );
not ( n41618 , n41617 );
buf ( n41619 , n41618 );
buf ( n41620 , n41619 );
buf ( n41621 , n41608 );
nand ( n41622 , n41620 , n41621 );
buf ( n41623 , n41622 );
buf ( n41624 , n41623 );
nand ( n41625 , n41616 , n41624 );
buf ( n41626 , n41625 );
buf ( n41627 , n41626 );
nand ( n41628 , n41602 , n41627 );
buf ( n41629 , n41628 );
buf ( n41630 , n41629 );
not ( n41631 , n24951 );
buf ( n41632 , n25009 );
not ( n41633 , n41632 );
buf ( n41634 , n41633 );
not ( n41635 , n41634 );
or ( n41636 , n41631 , n41635 );
not ( n41637 , n25008 );
nand ( n41638 , n25004 , n24994 );
not ( n41639 , n41638 );
or ( n41640 , n41637 , n41639 );
nand ( n41641 , n41640 , n24950 );
nand ( n41642 , n41636 , n41641 );
buf ( n41643 , n41642 );
not ( n41644 , n41643 );
buf ( n41645 , n41644 );
not ( n41646 , n41645 );
buf ( n41647 , n41646 );
buf ( n41648 , n41647 );
not ( n41649 , n41648 );
not ( n41650 , n24849 );
not ( n41651 , n24854 );
or ( n41652 , n41650 , n41651 );
not ( n41653 , n24849 );
nand ( n41654 , n41653 , n24855 );
nand ( n41655 , n41652 , n41654 );
not ( n41656 , n41655 );
buf ( n41657 , n41656 );
buf ( n41658 , n41657 );
buf ( n41659 , n41658 );
buf ( n41660 , n41659 );
buf ( n41661 , n41660 );
buf ( n41662 , n41661 );
buf ( n41663 , n41662 );
buf ( n41664 , n41663 );
not ( n41665 , n41664 );
buf ( n41666 , n41665 );
buf ( n41667 , n41666 );
not ( n41668 , n41667 );
buf ( n41669 , n37147 );
not ( n41670 , n41669 );
or ( n41671 , n41668 , n41670 );
buf ( n41672 , n37148 );
buf ( n41673 , n41663 );
nand ( n41674 , n41672 , n41673 );
buf ( n41675 , n41674 );
buf ( n41676 , n41675 );
nand ( n41677 , n41671 , n41676 );
buf ( n41678 , n41677 );
buf ( n41679 , n41678 );
not ( n41680 , n41679 );
or ( n41681 , n41649 , n41680 );
buf ( n41682 , n41666 );
not ( n41683 , n41682 );
buf ( n41684 , n37971 );
not ( n41685 , n41684 );
or ( n41686 , n41683 , n41685 );
buf ( n41687 , n39277 );
buf ( n41688 , n41663 );
nand ( n41689 , n41687 , n41688 );
buf ( n41690 , n41689 );
buf ( n41691 , n41690 );
nand ( n41692 , n41686 , n41691 );
buf ( n41693 , n41692 );
buf ( n41694 , n41693 );
not ( n41695 , n41642 );
buf ( n41696 , n41655 );
buf ( n41697 , n41696 );
buf ( n41698 , n41697 );
nand ( n41699 , n25010 , n41698 );
not ( n41700 , n24862 );
buf ( n41701 , n41634 );
nand ( n41702 , n41700 , n41701 );
nand ( n41703 , n41695 , n41699 , n41702 );
buf ( n41704 , n41703 );
not ( n41705 , n41704 );
buf ( n41706 , n41705 );
nand ( n41707 , n41694 , n41706 );
buf ( n41708 , n41707 );
buf ( n41709 , n41708 );
nand ( n41710 , n41681 , n41709 );
buf ( n41711 , n41710 );
buf ( n41712 , n41711 );
xor ( n41713 , n41630 , n41712 );
not ( n41714 , n13662 );
not ( n41715 , n39726 );
not ( n41716 , n41715 );
or ( n41717 , n41714 , n41716 );
not ( n41718 , n36527 );
buf ( n41719 , n13662 );
not ( n41720 , n41719 );
buf ( n41721 , n41720 );
nand ( n41722 , n41718 , n41721 );
nand ( n41723 , n41717 , n41722 );
not ( n41724 , n41723 );
buf ( n41725 , n41724 );
not ( n41726 , n41725 );
buf ( n41727 , n39806 );
not ( n41728 , n41727 );
or ( n41729 , n41726 , n41728 );
buf ( n41730 , n36643 );
buf ( n41731 , n28344 );
not ( n41732 , n41731 );
buf ( n41733 , n41732 );
buf ( n41734 , n41733 );
not ( n41735 , n41734 );
buf ( n41736 , n41735 );
buf ( n41737 , n41736 );
not ( n41738 , n41737 );
buf ( n41739 , n41715 );
not ( n41740 , n41739 );
buf ( n41741 , n41740 );
buf ( n41742 , n41741 );
not ( n41743 , n41742 );
or ( n41744 , n41738 , n41743 );
buf ( n41745 , n38471 );
buf ( n41746 , n41736 );
not ( n41747 , n41746 );
buf ( n41748 , n41747 );
buf ( n41749 , n41748 );
nand ( n41750 , n41745 , n41749 );
buf ( n41751 , n41750 );
buf ( n41752 , n41751 );
nand ( n41753 , n41744 , n41752 );
buf ( n41754 , n41753 );
buf ( n41755 , n41754 );
nand ( n41756 , n41730 , n41755 );
buf ( n41757 , n41756 );
buf ( n41758 , n41757 );
nand ( n41759 , n41729 , n41758 );
buf ( n41760 , n41759 );
buf ( n41761 , n41760 );
buf ( n41762 , n28720 );
not ( n41763 , n41762 );
not ( n41764 , n41763 );
buf ( n41765 , n41764 );
not ( n41766 , n41765 );
buf ( n41767 , n37336 );
buf ( n41768 , n41767 );
buf ( n41769 , n41768 );
buf ( n41770 , n41769 );
not ( n41771 , n41770 );
buf ( n41772 , n41771 );
buf ( n41773 , n41772 );
not ( n41774 , n41773 );
or ( n41775 , n41766 , n41774 );
buf ( n41776 , n37327 );
not ( n41777 , n41776 );
buf ( n41778 , n41777 );
not ( n41779 , n41778 );
buf ( n41780 , n41779 );
not ( n41781 , n28721 );
not ( n41782 , n41781 );
not ( n41783 , n41782 );
buf ( n41784 , n41783 );
nand ( n41785 , n41780 , n41784 );
buf ( n41786 , n41785 );
buf ( n41787 , n41786 );
nand ( n41788 , n41775 , n41787 );
buf ( n41789 , n41788 );
buf ( n41790 , n41789 );
not ( n41791 , n41790 );
buf ( n41792 , n37397 );
not ( n41793 , n41792 );
or ( n41794 , n41791 , n41793 );
not ( n41795 , n37329 );
not ( n41796 , n41795 );
buf ( n41797 , n29287 );
not ( n41798 , n41797 );
buf ( n41799 , n41798 );
not ( n41800 , n41799 );
or ( n41801 , n41796 , n41800 );
buf ( n41802 , n39653 );
buf ( n41803 , n41769 );
not ( n41804 , n41803 );
buf ( n41805 , n41804 );
buf ( n41806 , n41805 );
nand ( n41807 , n41802 , n41806 );
buf ( n41808 , n41807 );
nand ( n41809 , n41801 , n41808 );
nand ( n41810 , n41809 , n37413 );
buf ( n41811 , n41810 );
nand ( n41812 , n41794 , n41811 );
buf ( n41813 , n41812 );
buf ( n41814 , n41813 );
buf ( n41815 , n37514 );
not ( n41816 , n29323 );
not ( n41817 , n29319 );
not ( n41818 , n41817 );
or ( n41819 , n41816 , n41818 );
nand ( n41820 , n29319 , n29313 );
nand ( n41821 , n41819 , n41820 );
buf ( n41822 , n41821 );
buf ( n41823 , n41822 );
buf ( n41824 , n41823 );
buf ( n41825 , n37472 );
and ( n41826 , n41824 , n41825 );
not ( n41827 , n41824 );
not ( n41828 , n37472 );
buf ( n41829 , n41828 );
and ( n41830 , n41827 , n41829 );
nor ( n41831 , n41826 , n41830 );
buf ( n41832 , n41831 );
buf ( n41833 , n41832 );
or ( n41834 , n41815 , n41833 );
not ( n41835 , n28305 );
not ( n41836 , n41835 );
buf ( n41837 , n41836 );
buf ( n41838 , n41837 );
not ( n41839 , n41828 );
buf ( n41840 , n41839 );
and ( n41841 , n41838 , n41840 );
not ( n41842 , n41838 );
buf ( n41843 , n37501 );
buf ( n41844 , n41843 );
buf ( n41845 , n41844 );
and ( n41846 , n41842 , n41845 );
nor ( n41847 , n41841 , n41846 );
buf ( n41848 , n41847 );
buf ( n41849 , n41848 );
buf ( n41850 , n37440 );
buf ( n41851 , n41850 );
buf ( n41852 , n41851 );
buf ( n41853 , n41852 );
not ( n41854 , n41853 );
buf ( n41855 , n41854 );
buf ( n41856 , n41855 );
or ( n41857 , n41849 , n41856 );
nand ( n41858 , n41834 , n41857 );
buf ( n41859 , n41858 );
buf ( n41860 , n41859 );
xor ( n41861 , n41814 , n41860 );
buf ( n41862 , n37871 );
buf ( n41863 , n41862 );
not ( n41864 , n41863 );
buf ( n41865 , n41864 );
buf ( n41866 , n41865 );
and ( n41867 , n29371 , n29376 );
not ( n41868 , n29371 );
and ( n41869 , n41868 , n29375 );
nor ( n41870 , n41867 , n41869 );
buf ( n41871 , n41870 );
not ( n41872 , n41871 );
buf ( n41873 , n41872 );
buf ( n41874 , n41873 );
not ( n41875 , n41874 );
buf ( n41876 , n41875 );
buf ( n41877 , n41876 );
not ( n41878 , n41877 );
buf ( n41879 , n41878 );
buf ( n41880 , n41879 );
not ( n41881 , n41880 );
buf ( n41882 , n41881 );
buf ( n41883 , n41882 );
not ( n41884 , n41883 );
not ( n41885 , n37840 );
not ( n41886 , n37851 );
or ( n41887 , n41885 , n41886 );
nand ( n41888 , n41887 , n37857 );
buf ( n41889 , n41888 );
not ( n41890 , n41889 );
buf ( n41891 , n41890 );
not ( n41892 , n41891 );
or ( n41893 , n41884 , n41892 );
not ( n41894 , n41888 );
not ( n41895 , n41894 );
nand ( n41896 , n41895 , n41879 );
buf ( n41897 , n41896 );
nand ( n41898 , n41893 , n41897 );
buf ( n41899 , n41898 );
buf ( n41900 , n41899 );
not ( n41901 , n41900 );
buf ( n41902 , n41901 );
buf ( n41903 , n41902 );
or ( n41904 , n41866 , n41903 );
not ( n41905 , n37916 );
buf ( n41906 , n41905 );
not ( n41907 , n41906 );
buf ( n41908 , n41907 );
buf ( n41909 , n41908 );
buf ( n41910 , n29358 );
buf ( n41911 , n41910 );
buf ( n41912 , n41911 );
buf ( n41913 , n41912 );
not ( n41914 , n41913 );
buf ( n41915 , n41914 );
buf ( n41916 , n41915 );
buf ( n41917 , n41916 );
buf ( n41918 , n41917 );
buf ( n41919 , n41918 );
buf ( n41920 , n37881 );
and ( n41921 , n41919 , n41920 );
not ( n41922 , n41919 );
buf ( n41923 , n41889 );
not ( n41924 , n41923 );
buf ( n41925 , n41924 );
buf ( n41926 , n41925 );
and ( n41927 , n41922 , n41926 );
nor ( n41928 , n41921 , n41927 );
buf ( n41929 , n41928 );
buf ( n41930 , n41929 );
or ( n41931 , n41909 , n41930 );
nand ( n41932 , n41904 , n41931 );
buf ( n41933 , n41932 );
buf ( n41934 , n41933 );
and ( n41935 , n41861 , n41934 );
and ( n41936 , n41814 , n41860 );
or ( n41937 , n41935 , n41936 );
buf ( n41938 , n41937 );
buf ( n41939 , n41938 );
xor ( n41940 , n41761 , n41939 );
not ( n41941 , n37919 );
buf ( n41942 , n41823 );
not ( n41943 , n41942 );
buf ( n41944 , n41925 );
not ( n41945 , n41944 );
or ( n41946 , n41943 , n41945 );
buf ( n41947 , n41889 );
buf ( n41948 , n41947 );
buf ( n41949 , n41821 );
not ( n41950 , n41949 );
buf ( n41951 , n41950 );
buf ( n41952 , n41951 );
nand ( n41953 , n41948 , n41952 );
buf ( n41954 , n41953 );
buf ( n41955 , n41954 );
nand ( n41956 , n41946 , n41955 );
buf ( n41957 , n41956 );
not ( n41958 , n41957 );
or ( n41959 , n41941 , n41958 );
not ( n41960 , n41929 );
nand ( n41961 , n41960 , n37872 );
nand ( n41962 , n41959 , n41961 );
buf ( n41963 , n41962 );
buf ( n41964 , n37511 );
not ( n41965 , n41964 );
buf ( n41966 , n41965 );
buf ( n41967 , n41966 );
not ( n41968 , n41967 );
buf ( n41969 , n41968 );
buf ( n41970 , n41969 );
buf ( n41971 , n41848 );
or ( n41972 , n41970 , n41971 );
not ( n41973 , n37440 );
buf ( n41974 , n41973 );
not ( n41975 , n41762 );
not ( n41976 , n37472 );
not ( n41977 , n41976 );
not ( n41978 , n41977 );
and ( n41979 , n41975 , n41978 );
not ( n41980 , n41975 );
not ( n41981 , n37472 );
not ( n41982 , n41981 );
and ( n41983 , n41980 , n41982 );
nor ( n41984 , n41979 , n41983 );
buf ( n41985 , n41984 );
or ( n41986 , n41974 , n41985 );
nand ( n41987 , n41972 , n41986 );
buf ( n41988 , n41987 );
buf ( n41989 , n41988 );
xor ( n41990 , n41963 , n41989 );
buf ( n41991 , n41990 );
buf ( n41992 , n41991 );
buf ( n41993 , n28430 );
buf ( n41994 , n41993 );
buf ( n41995 , n37649 );
and ( n41996 , n41994 , n41995 );
not ( n41997 , n41994 );
buf ( n41998 , n38798 );
and ( n41999 , n41997 , n41998 );
nor ( n42000 , n41996 , n41999 );
buf ( n42001 , n42000 );
buf ( n42002 , n36444 );
not ( n42003 , n42002 );
buf ( n42004 , n42003 );
buf ( n42005 , n42004 );
buf ( n42006 , n29463 );
buf ( n42007 , n42006 );
buf ( n42008 , n42007 );
buf ( n42009 , n42008 );
not ( n42010 , n42009 );
buf ( n42011 , n37602 );
not ( n42012 , n42011 );
or ( n42013 , n42010 , n42012 );
buf ( n42014 , n36360 );
buf ( n42015 , n42008 );
not ( n42016 , n42015 );
buf ( n42017 , n42016 );
buf ( n42018 , n42017 );
nand ( n42019 , n42014 , n42018 );
buf ( n42020 , n42019 );
buf ( n42021 , n42020 );
nand ( n42022 , n42013 , n42021 );
buf ( n42023 , n42022 );
buf ( n42024 , n42023 );
not ( n42025 , n42024 );
buf ( n42026 , n42025 );
buf ( n42027 , n42026 );
or ( n42028 , n42005 , n42027 );
nand ( n42029 , C1 , n42028 );
buf ( n42030 , n42029 );
buf ( n42031 , n42030 );
xor ( n42032 , n41992 , n42031 );
buf ( n42033 , n42032 );
buf ( n42034 , n42033 );
and ( n42035 , n41940 , n42034 );
and ( n42036 , n41761 , n41939 );
or ( n42037 , n42035 , n42036 );
buf ( n42038 , n42037 );
buf ( n42039 , n42038 );
xor ( n42040 , n41713 , n42039 );
buf ( n42041 , n42040 );
buf ( n42042 , n42041 );
buf ( n42043 , n36973 );
buf ( n42044 , n42043 );
buf ( n42045 , n42044 );
buf ( n42046 , n42045 );
buf ( n42047 , n29754 );
buf ( n42048 , n42047 );
buf ( n42049 , n42048 );
buf ( n42050 , n42049 );
not ( n42051 , n42050 );
buf ( n42052 , n42051 );
buf ( n42053 , n42052 );
not ( n42054 , n42053 );
buf ( n42055 , n42054 );
buf ( n42056 , n42055 );
buf ( n42057 , n39139 );
and ( n42058 , n42056 , n42057 );
not ( n42059 , n42056 );
buf ( n42060 , n36920 );
buf ( n42061 , n42060 );
buf ( n42062 , n42061 );
buf ( n42063 , n42062 );
and ( n42064 , n42059 , n42063 );
nor ( n42065 , n42058 , n42064 );
buf ( n42066 , n42065 );
buf ( n42067 , n42066 );
or ( n42068 , n42046 , n42067 );
buf ( n42069 , n36909 );
buf ( n42070 , n28368 );
not ( n42071 , n42070 );
buf ( n42072 , n42071 );
buf ( n42073 , n42072 );
buf ( n42074 , n42073 );
buf ( n42075 , n42074 );
buf ( n42076 , n42075 );
buf ( n42077 , n42062 );
and ( n42078 , n42076 , n42077 );
not ( n42079 , n42076 );
buf ( n42080 , n36923 );
buf ( n42081 , n42080 );
buf ( n42082 , n42081 );
buf ( n42083 , n42082 );
and ( n42084 , n42079 , n42083 );
nor ( n42085 , n42078 , n42084 );
buf ( n42086 , n42085 );
buf ( n42087 , n42086 );
or ( n42088 , n42069 , n42087 );
nand ( n42089 , n42068 , n42088 );
buf ( n42090 , n42089 );
not ( n42091 , n42090 );
buf ( n42092 , n39803 );
not ( n42093 , n42092 );
buf ( n42094 , n42093 );
buf ( n42095 , n36527 );
not ( n42096 , n42095 );
buf ( n42097 , n42017 );
not ( n42098 , n42097 );
and ( n42099 , n42096 , n42098 );
buf ( n42100 , n36527 );
buf ( n42101 , n42017 );
and ( n42102 , n42100 , n42101 );
nor ( n42103 , n42099 , n42102 );
buf ( n42104 , n42103 );
or ( n42105 , n42094 , n42104 );
not ( n42106 , n36640 );
nand ( n42107 , n42106 , n41724 );
nand ( n42108 , n42105 , n42107 );
not ( n42109 , n42108 );
nand ( n42110 , n42091 , n42109 );
not ( n42111 , n42110 );
buf ( n42112 , n41805 );
not ( n42113 , n42112 );
buf ( n42114 , n42113 );
buf ( n42115 , n42114 );
buf ( n42116 , n28306 );
and ( n42117 , n42115 , n42116 );
not ( n42118 , n42115 );
not ( n42119 , n28305 );
buf ( n42120 , n42119 );
and ( n42121 , n42118 , n42120 );
nor ( n42122 , n42117 , n42121 );
buf ( n42123 , n42122 );
buf ( n42124 , n42123 );
not ( n42125 , n42124 );
buf ( n42126 , n37397 );
not ( n42127 , n42126 );
or ( n42128 , n42125 , n42127 );
buf ( n42129 , n41789 );
buf ( n42130 , n37410 );
not ( n42131 , n42130 );
buf ( n42132 , n42131 );
buf ( n42133 , n42132 );
not ( n42134 , n42133 );
buf ( n42135 , n42134 );
buf ( n42136 , n42135 );
nand ( n42137 , n42129 , n42136 );
buf ( n42138 , n42137 );
buf ( n42139 , n42138 );
nand ( n42140 , n42128 , n42139 );
buf ( n42141 , n42140 );
buf ( n42142 , n42141 );
and ( n42143 , n28390 , n28403 );
not ( n42144 , n28390 );
and ( n42145 , n42144 , n28408 );
nor ( n42146 , n42143 , n42145 );
buf ( n42147 , n42146 );
buf ( n42148 , n42147 );
buf ( n42149 , n42148 );
buf ( n42150 , n42149 );
buf ( n42151 , n42150 );
buf ( n42152 , n42151 );
buf ( n42153 , n42152 );
not ( n42154 , n42153 );
buf ( n42155 , n41925 );
not ( n42156 , n42155 );
or ( n42157 , n42154 , n42156 );
buf ( n42158 , n42152 );
not ( n42159 , n42158 );
buf ( n42160 , n42159 );
buf ( n42161 , n42160 );
buf ( n42162 , n41947 );
nand ( n42163 , n42161 , n42162 );
buf ( n42164 , n42163 );
buf ( n42165 , n42164 );
nand ( n42166 , n42157 , n42165 );
buf ( n42167 , n42166 );
buf ( n42168 , n42167 );
not ( n42169 , n42168 );
buf ( n42170 , n37872 );
not ( n42171 , n42170 );
or ( n42172 , n42169 , n42171 );
buf ( n42173 , n37916 );
not ( n42174 , n42173 );
buf ( n42175 , n42174 );
buf ( n42176 , n42175 );
buf ( n42177 , n41899 );
nand ( n42178 , n42176 , n42177 );
buf ( n42179 , n42178 );
buf ( n42180 , n42179 );
nand ( n42181 , n42172 , n42180 );
buf ( n42182 , n42181 );
buf ( n42183 , n42182 );
xor ( n42184 , n42142 , n42183 );
buf ( n42185 , n37514 );
buf ( n42186 , n41918 );
not ( n42187 , n42186 );
buf ( n42188 , n42187 );
buf ( n42189 , n42188 );
not ( n42190 , n42189 );
buf ( n42191 , n37472 );
not ( n42192 , n42191 );
or ( n42193 , n42190 , n42192 );
buf ( n42194 , n41981 );
buf ( n42195 , n29359 );
buf ( n42196 , n42195 );
buf ( n42197 , n42196 );
nand ( n42198 , n42194 , n42197 );
buf ( n42199 , n42198 );
buf ( n42200 , n42199 );
nand ( n42201 , n42193 , n42200 );
buf ( n42202 , n42201 );
buf ( n42203 , n42202 );
not ( n42204 , n42203 );
buf ( n42205 , n42204 );
buf ( n42206 , n42205 );
or ( n42207 , n42185 , n42206 );
buf ( n42208 , n37446 );
not ( n42209 , n42208 );
buf ( n42210 , n42209 );
buf ( n42211 , n42210 );
buf ( n42212 , n41832 );
or ( n42213 , n42211 , n42212 );
nand ( n42214 , n42207 , n42213 );
buf ( n42215 , n42214 );
buf ( n42216 , n42215 );
and ( n42217 , n42184 , n42216 );
and ( n42218 , n42142 , n42183 );
or ( n42219 , n42217 , n42218 );
buf ( n42220 , n42219 );
not ( n42221 , n42220 );
or ( n42222 , n42111 , n42221 );
nand ( n42223 , n42108 , n42090 );
nand ( n42224 , n42222 , n42223 );
buf ( n42225 , n42224 );
buf ( n42226 , n25336 );
buf ( n42227 , n42226 );
buf ( n42228 , n42227 );
xnor ( n42229 , n24883 , n42228 );
buf ( n42230 , n42229 );
buf ( n42231 , n25287 );
buf ( n42232 , n24883 );
nand ( n42233 , n42231 , n42232 );
buf ( n42234 , n42233 );
buf ( n42235 , n42234 );
buf ( n42236 , n25287 );
not ( n42237 , n42236 );
buf ( n42238 , n24884 );
nand ( n42239 , n42237 , n42238 );
buf ( n42240 , n42239 );
buf ( n42241 , n42240 );
nand ( n42242 , n42230 , n42235 , n42241 );
buf ( n42243 , n42242 );
buf ( n42244 , n42243 );
not ( n42245 , n42244 );
buf ( n42246 , n42245 );
buf ( n42247 , n42246 );
not ( n42248 , n42247 );
buf ( n42249 , n42248 );
buf ( n42250 , n42249 );
not ( n42251 , n42250 );
buf ( n42252 , n42251 );
buf ( n42253 , n42252 );
not ( n42254 , n42253 );
buf ( n42255 , n25287 );
not ( n42256 , n42255 );
buf ( n42257 , n42256 );
buf ( n42258 , n42257 );
buf ( n42259 , n42258 );
buf ( n42260 , n42259 );
buf ( n42261 , n42260 );
buf ( n42262 , n42261 );
buf ( n42263 , n42262 );
buf ( n42264 , n42263 );
not ( n42265 , n42264 );
buf ( n42266 , n42265 );
buf ( n42267 , n42266 );
not ( n42268 , n42267 );
buf ( n42269 , n36559 );
not ( n42270 , n42269 );
buf ( n42271 , n42270 );
buf ( n42272 , n42271 );
not ( n42273 , n42272 );
or ( n42274 , n42268 , n42273 );
buf ( n42275 , n36559 );
not ( n42276 , n42275 );
buf ( n42277 , n42276 );
buf ( n42278 , n42277 );
not ( n42279 , n42278 );
buf ( n42280 , n42279 );
buf ( n42281 , n42280 );
buf ( n42282 , n42263 );
nand ( n42283 , n42281 , n42282 );
buf ( n42284 , n42283 );
buf ( n42285 , n42284 );
nand ( n42286 , n42274 , n42285 );
buf ( n42287 , n42286 );
buf ( n42288 , n42287 );
not ( n42289 , n42288 );
or ( n42290 , n42254 , n42289 );
buf ( n42291 , n42266 );
not ( n42292 , n42291 );
buf ( n42293 , n39582 );
not ( n42294 , n42293 );
or ( n42295 , n42292 , n42294 );
buf ( n42296 , n36611 );
buf ( n42297 , n42263 );
nand ( n42298 , n42296 , n42297 );
buf ( n42299 , n42298 );
buf ( n42300 , n42299 );
nand ( n42301 , n42295 , n42300 );
buf ( n42302 , n42301 );
buf ( n42303 , n42302 );
buf ( n42304 , n42229 );
buf ( n42305 , n42304 );
buf ( n42306 , n42305 );
buf ( n42307 , n42306 );
not ( n42308 , n42307 );
buf ( n42309 , n42308 );
buf ( n42310 , n42309 );
not ( n42311 , n42310 );
buf ( n42312 , n42311 );
buf ( n42313 , n42312 );
not ( n42314 , n42313 );
buf ( n42315 , n42314 );
buf ( n42316 , n42315 );
nand ( n42317 , n42303 , n42316 );
buf ( n42318 , n42317 );
buf ( n42319 , n42318 );
nand ( n42320 , n42290 , n42319 );
buf ( n42321 , n42320 );
buf ( n42322 , n42321 );
xor ( n42323 , n42225 , n42322 );
not ( n42324 , n25225 );
not ( n42325 , n42324 );
not ( n42326 , n42325 );
not ( n42327 , n24923 );
not ( n42328 , n42327 );
or ( n42329 , n42326 , n42328 );
nand ( n42330 , n42324 , n24923 );
nand ( n42331 , n42329 , n42330 );
not ( n42332 , n42331 );
not ( n42333 , n42332 );
buf ( n42334 , n42333 );
not ( n42335 , n42334 );
buf ( n42336 , n42335 );
buf ( n42337 , n42336 );
buf ( n42338 , n42337 );
buf ( n42339 , n42338 );
buf ( n42340 , n42339 );
not ( n42341 , n42340 );
buf ( n42342 , n24950 );
not ( n42343 , n42342 );
buf ( n42344 , n42343 );
not ( n42345 , n42344 );
buf ( n42346 , n38098 );
not ( n42347 , n42346 );
or ( n42348 , n42345 , n42347 );
buf ( n42349 , n39340 );
not ( n42350 , n42343 );
buf ( n42351 , n42350 );
nand ( n42352 , n42349 , n42351 );
buf ( n42353 , n42352 );
buf ( n42354 , n42353 );
nand ( n42355 , n42348 , n42354 );
buf ( n42356 , n42355 );
buf ( n42357 , n42356 );
not ( n42358 , n42357 );
or ( n42359 , n42341 , n42358 );
not ( n42360 , n37146 );
and ( n42361 , n42343 , n42360 );
not ( n42362 , n42343 );
and ( n42363 , n42362 , n39860 );
or ( n42364 , n42361 , n42363 );
buf ( n42365 , n42364 );
not ( n42366 , n24950 );
nand ( n42367 , n42366 , n24926 );
buf ( n42368 , n24923 );
buf ( n42369 , n24950 );
nand ( n42370 , n42368 , n42369 );
buf ( n42371 , n42370 );
nand ( n42372 , n42331 , n42367 , n42371 );
buf ( n42373 , n42372 );
not ( n42374 , n42373 );
not ( n42375 , n42374 );
buf ( n42376 , n42375 );
not ( n42377 , n42376 );
buf ( n42378 , n42377 );
buf ( n42379 , n42378 );
nand ( n42380 , n42365 , n42379 );
buf ( n42381 , n42380 );
buf ( n42382 , n42381 );
nand ( n42383 , n42359 , n42382 );
buf ( n42384 , n42383 );
buf ( n42385 , n42384 );
and ( n42386 , n42323 , n42385 );
and ( n42387 , n42225 , n42322 );
or ( n42388 , n42386 , n42387 );
buf ( n42389 , n42388 );
buf ( n42390 , n42389 );
xor ( n42391 , n42042 , n42390 );
xor ( n42392 , n41761 , n41939 );
xor ( n42393 , n42392 , n42034 );
buf ( n42394 , n42393 );
buf ( n42395 , n42394 );
buf ( n42396 , n41799 );
not ( n42397 , n42396 );
buf ( n42398 , n42397 );
buf ( n42399 , n42398 );
not ( n42400 , n42399 );
buf ( n42401 , n38393 );
not ( n42402 , n42401 );
buf ( n42403 , n42402 );
buf ( n42404 , n42403 );
not ( n42405 , n42404 );
and ( n42406 , n42400 , n42405 );
buf ( n42407 , n39653 );
buf ( n42408 , n37381 );
buf ( n42409 , n42408 );
buf ( n42410 , n42409 );
buf ( n42411 , n42410 );
buf ( n42412 , n42411 );
not ( n42413 , n42412 );
buf ( n42414 , n42413 );
buf ( n42415 , n42414 );
and ( n42416 , n42407 , n42415 );
nor ( n42417 , n42406 , n42416 );
buf ( n42418 , n42417 );
not ( n42419 , n42418 );
not ( n42420 , n38407 );
and ( n42421 , n42419 , n42420 );
buf ( n42422 , n42414 );
buf ( n42423 , n29269 );
not ( n42424 , n42423 );
buf ( n42425 , n42424 );
buf ( n42426 , n42425 );
not ( n42427 , n42426 );
buf ( n42428 , n42427 );
buf ( n42429 , n42428 );
and ( n42430 , n42422 , n42429 );
not ( n42431 , n42422 );
buf ( n42432 , n29269 );
buf ( n42433 , n42432 );
buf ( n42434 , n42433 );
buf ( n42435 , n42434 );
not ( n42436 , n42435 );
buf ( n42437 , n42436 );
buf ( n42438 , n42437 );
and ( n42439 , n42431 , n42438 );
nor ( n42440 , n42430 , n42439 );
buf ( n42441 , n42440 );
buf ( n42442 , n42441 );
buf ( n42443 , n38383 );
nor ( n42444 , n42442 , n42443 );
buf ( n42445 , n42444 );
nor ( n42446 , n42421 , n42445 );
buf ( n42447 , n42446 );
not ( n42448 , n38973 );
buf ( n42449 , n42448 );
not ( n42450 , n42449 );
buf ( n42451 , n38979 );
not ( n42452 , n42451 );
buf ( n42453 , n38820 );
not ( n42454 , n42453 );
buf ( n42455 , n42454 );
buf ( n42456 , n42455 );
not ( n42457 , n42456 );
buf ( n42458 , n42457 );
buf ( n42459 , n42458 );
not ( n42460 , n42459 );
buf ( n42461 , n42460 );
buf ( n42462 , n42461 );
not ( n42463 , n42462 );
or ( n42464 , n42452 , n42463 );
buf ( n42465 , n38821 );
buf ( n42466 , n24638 );
buf ( n42467 , n42466 );
buf ( n42468 , n42467 );
buf ( n42469 , n42468 );
not ( n42470 , n42469 );
buf ( n42471 , n42470 );
buf ( n42472 , n42471 );
nand ( n42473 , n42465 , n42472 );
buf ( n42474 , n42473 );
buf ( n42475 , n42474 );
nand ( n42476 , n42464 , n42475 );
buf ( n42477 , n42476 );
buf ( n42478 , n42477 );
not ( n42479 , n42478 );
or ( n42480 , n42450 , n42479 );
buf ( n42481 , n38979 );
not ( n42482 , n42481 );
buf ( n42483 , n30187 );
not ( n42484 , n42483 );
buf ( n42485 , n42484 );
buf ( n42486 , n42485 );
not ( n42487 , n42486 );
or ( n42488 , n42482 , n42487 );
nand ( n42489 , n30187 , n42471 );
buf ( n42490 , n42489 );
nand ( n42491 , n42488 , n42490 );
buf ( n42492 , n42491 );
buf ( n42493 , n42492 );
buf ( n42494 , n38985 );
nand ( n42495 , n42493 , n42494 );
buf ( n42496 , n42495 );
buf ( n42497 , n42496 );
nand ( n42498 , n42480 , n42497 );
buf ( n42499 , n42498 );
buf ( n42500 , n42499 );
xor ( n42501 , n42447 , n42500 );
buf ( n42502 , n41721 );
not ( n42503 , n42502 );
buf ( n42504 , n42503 );
buf ( n42505 , n42504 );
not ( n42506 , n42505 );
buf ( n42507 , n39478 );
not ( n42508 , n42507 );
or ( n42509 , n42506 , n42508 );
buf ( n42510 , n33077 );
buf ( n42511 , n41721 );
nand ( n42512 , n42510 , n42511 );
buf ( n42513 , n42512 );
buf ( n42514 , n42513 );
nand ( n42515 , n42509 , n42514 );
buf ( n42516 , n42515 );
buf ( n42517 , n42516 );
not ( n42518 , n42517 );
buf ( n42519 , n36098 );
not ( n42520 , n42519 );
buf ( n42521 , n42520 );
buf ( n42522 , n42521 );
not ( n42523 , n42522 );
or ( n42524 , n42518 , n42523 );
buf ( n42525 , n32963 );
not ( n42526 , n42525 );
buf ( n42527 , n42526 );
buf ( n42528 , n42527 );
buf ( n42529 , n42528 );
buf ( n42530 , n42529 );
buf ( n42531 , n42530 );
buf ( n42532 , n41736 );
not ( n42533 , n42532 );
buf ( n42534 , n39478 );
not ( n42535 , n42534 );
or ( n42536 , n42533 , n42535 );
buf ( n42537 , n33077 );
buf ( n42538 , n41748 );
nand ( n42539 , n42537 , n42538 );
buf ( n42540 , n42539 );
buf ( n42541 , n42540 );
nand ( n42542 , n42536 , n42541 );
buf ( n42543 , n42542 );
buf ( n42544 , n42543 );
nand ( n42545 , n42531 , n42544 );
buf ( n42546 , n42545 );
buf ( n42547 , n42546 );
nand ( n42548 , n42524 , n42547 );
buf ( n42549 , n42548 );
buf ( n42550 , n42549 );
and ( n42551 , n42501 , n42550 );
and ( n42552 , n42447 , n42500 );
or ( n42553 , n42551 , n42552 );
buf ( n42554 , n42553 );
buf ( n42555 , n42554 );
not ( n42556 , n25179 );
and ( n42557 , n25070 , n42556 );
not ( n42558 , n25070 );
not ( n42559 , n25179 );
not ( n42560 , n42559 );
and ( n42561 , n42558 , n42560 );
nor ( n42562 , n42557 , n42561 );
buf ( n42563 , n42562 );
not ( n42564 , n42563 );
not ( n42565 , n42564 );
not ( n42566 , n42565 );
buf ( n42567 , n42566 );
not ( n42568 , n42567 );
buf ( n42569 , n25160 );
not ( n42570 , n42569 );
buf ( n42571 , n37705 );
not ( n42572 , n42571 );
buf ( n42573 , n42572 );
buf ( n42574 , n42573 );
not ( n42575 , n42574 );
or ( n42576 , n42570 , n42575 );
buf ( n42577 , n37692 );
buf ( n42578 , n25159 );
buf ( n42579 , n42578 );
not ( n42580 , n42579 );
buf ( n42581 , n42580 );
buf ( n42582 , n42581 );
nand ( n42583 , n42577 , n42582 );
buf ( n42584 , n42583 );
buf ( n42585 , n42584 );
nand ( n42586 , n42576 , n42585 );
buf ( n42587 , n42586 );
buf ( n42588 , n42587 );
not ( n42589 , n42588 );
or ( n42590 , n42568 , n42589 );
buf ( n42591 , n25160 );
not ( n42592 , n42591 );
not ( n42593 , n37729 );
not ( n42594 , n37737 );
or ( n42595 , n42593 , n42594 );
nand ( n42596 , n42595 , n37741 );
not ( n42597 , n42596 );
buf ( n42598 , n42597 );
not ( n42599 , n42598 );
or ( n42600 , n42592 , n42599 );
buf ( n42601 , n39522 );
buf ( n42602 , n42581 );
nand ( n42603 , n42601 , n42602 );
buf ( n42604 , n42603 );
buf ( n42605 , n42604 );
nand ( n42606 , n42600 , n42605 );
buf ( n42607 , n42606 );
buf ( n42608 , n42607 );
buf ( n42609 , n39973 );
not ( n42610 , n42609 );
buf ( n42611 , n25070 );
not ( n42612 , n42611 );
buf ( n42613 , n42612 );
buf ( n42614 , n42613 );
nand ( n42615 , n42610 , n42614 );
buf ( n42616 , n42615 );
buf ( n42617 , n42616 );
buf ( n42618 , n42562 );
nand ( n42619 , n25070 , n39973 );
buf ( n42620 , n42619 );
nand ( n42621 , n42617 , n42618 , n42620 );
buf ( n42622 , n42621 );
buf ( n42623 , n42622 );
buf ( n42624 , n42623 );
buf ( n42625 , n42624 );
buf ( n42626 , n42625 );
not ( n42627 , n42626 );
buf ( n42628 , n42627 );
buf ( n42629 , n42628 );
buf ( n42630 , n42629 );
buf ( n42631 , n42630 );
buf ( n42632 , n42631 );
nand ( n42633 , n42608 , n42632 );
buf ( n42634 , n42633 );
buf ( n42635 , n42634 );
nand ( n42636 , n42590 , n42635 );
buf ( n42637 , n42636 );
buf ( n42638 , n42637 );
xor ( n42639 , n42555 , n42638 );
xor ( n42640 , n41814 , n41860 );
xor ( n42641 , n42640 , n41934 );
buf ( n42642 , n42641 );
buf ( n42643 , n42642 );
and ( n42644 , n42639 , n42643 );
and ( n42645 , n42555 , n42638 );
or ( n42646 , n42644 , n42645 );
buf ( n42647 , n42646 );
buf ( n42648 , n42647 );
xor ( n42649 , n42395 , n42648 );
not ( n42650 , n42257 );
buf ( n42651 , n25242 );
buf ( n42652 , n25250 );
and ( n42653 , n42651 , n42652 );
not ( n42654 , n42651 );
buf ( n42655 , n25247 );
and ( n42656 , n42654 , n42655 );
nor ( n42657 , n42653 , n42656 );
buf ( n42658 , n42657 );
not ( n42659 , n42658 );
not ( n42660 , n42659 );
or ( n42661 , n42650 , n42660 );
not ( n42662 , n25303 );
nand ( n42663 , n42658 , n42662 );
nand ( n42664 , n42661 , n42663 );
not ( n42665 , n42664 );
buf ( n42666 , n42665 );
buf ( n42667 , n42666 );
buf ( n42668 , n42667 );
buf ( n42669 , n42668 );
not ( n42670 , n42669 );
buf ( n42671 , n25227 );
not ( n42672 , n42671 );
buf ( n42673 , n42672 );
not ( n42674 , n42673 );
buf ( n42675 , n40067 );
not ( n42676 , n42675 );
or ( n42677 , n42674 , n42676 );
buf ( n42678 , n36427 );
not ( n42679 , n42672 );
buf ( n42680 , n42679 );
nand ( n42681 , n42678 , n42680 );
buf ( n42682 , n42681 );
buf ( n42683 , n42682 );
nand ( n42684 , n42677 , n42683 );
buf ( n42685 , n42684 );
buf ( n42686 , n42685 );
not ( n42687 , n42686 );
or ( n42688 , n42670 , n42687 );
buf ( n42689 , n25228 );
not ( n42690 , n42689 );
buf ( n42691 , n39897 );
not ( n42692 , n42691 );
or ( n42693 , n42690 , n42692 );
buf ( n42694 , n36396 );
buf ( n42695 , n42679 );
nand ( n42696 , n42694 , n42695 );
buf ( n42697 , n42696 );
buf ( n42698 , n42697 );
nand ( n42699 , n42693 , n42698 );
buf ( n42700 , n42699 );
buf ( n42701 , n42700 );
buf ( n42702 , n25257 );
buf ( n42703 , n25225 );
nand ( n42704 , n42702 , n42703 );
buf ( n42705 , n42704 );
not ( n42706 , n25257 );
nand ( n42707 , n42706 , n42324 );
nand ( n42708 , n42705 , n42664 , n42707 );
not ( n42709 , n42708 );
not ( n42710 , n42709 );
buf ( n42711 , n42710 );
not ( n42712 , n42711 );
buf ( n42713 , n42712 );
nand ( n42714 , n42701 , n42713 );
buf ( n42715 , n42714 );
buf ( n42716 , n42715 );
nand ( n42717 , n42688 , n42716 );
buf ( n42718 , n42717 );
buf ( n42719 , n42718 );
and ( n42720 , n42649 , n42719 );
and ( n42721 , n42395 , n42648 );
or ( n42722 , n42720 , n42721 );
buf ( n42723 , n42722 );
buf ( n42724 , n42723 );
xor ( n42725 , n42391 , n42724 );
buf ( n42726 , n42725 );
buf ( n42727 , n42266 );
not ( n42728 , n42727 );
buf ( n42729 , n36430 );
not ( n42730 , n42729 );
or ( n42731 , n42728 , n42730 );
buf ( n42732 , n40067 );
not ( n42733 , n42732 );
buf ( n42734 , n42263 );
nand ( n42735 , n42733 , n42734 );
buf ( n42736 , n42735 );
buf ( n42737 , n42736 );
nand ( n42738 , n42731 , n42737 );
buf ( n42739 , n42738 );
buf ( n42740 , n42739 );
buf ( n42741 , n42252 );
and ( n42742 , n42740 , n42741 );
buf ( n42743 , n42287 );
not ( n42744 , n42743 );
buf ( n42745 , n42312 );
nor ( n42746 , n42744 , n42745 );
buf ( n42747 , n42746 );
buf ( n42748 , n42747 );
nor ( n42749 , n42742 , n42748 );
buf ( n42750 , n42749 );
buf ( n42751 , n42750 );
not ( n42752 , n42751 );
buf ( n42753 , n42752 );
buf ( n42754 , n42753 );
not ( n42755 , n42754 );
buf ( n42756 , n42668 );
not ( n42757 , n42756 );
buf ( n42758 , n42700 );
not ( n42759 , n42758 );
or ( n42760 , n42757 , n42759 );
buf ( n42761 , n42672 );
not ( n42762 , n42761 );
buf ( n42763 , n38098 );
not ( n42764 , n42763 );
or ( n42765 , n42762 , n42764 );
buf ( n42766 , n39340 );
buf ( n42767 , n42679 );
nand ( n42768 , n42766 , n42767 );
buf ( n42769 , n42768 );
buf ( n42770 , n42769 );
nand ( n42771 , n42765 , n42770 );
buf ( n42772 , n42771 );
buf ( n42773 , n42772 );
buf ( n42774 , n42712 );
nand ( n42775 , n42773 , n42774 );
buf ( n42776 , n42775 );
buf ( n42777 , n42776 );
nand ( n42778 , n42760 , n42777 );
buf ( n42779 , n42778 );
buf ( n42780 , n42779 );
not ( n42781 , n42780 );
or ( n42782 , n42755 , n42781 );
buf ( n42783 , n42779 );
buf ( n42784 , n42753 );
or ( n42785 , n42783 , n42784 );
buf ( n42786 , n42566 );
not ( n42787 , n42786 );
buf ( n42788 , n42607 );
not ( n42789 , n42788 );
or ( n42790 , n42787 , n42789 );
buf ( n42791 , n25160 );
not ( n42792 , n42791 );
buf ( n42793 , n38477 );
not ( n42794 , n42793 );
buf ( n42795 , n42794 );
buf ( n42796 , n42795 );
not ( n42797 , n42796 );
or ( n42798 , n42792 , n42797 );
buf ( n42799 , n37783 );
buf ( n42800 , n42581 );
nand ( n42801 , n42799 , n42800 );
buf ( n42802 , n42801 );
buf ( n42803 , n42802 );
nand ( n42804 , n42798 , n42803 );
buf ( n42805 , n42804 );
buf ( n42806 , n42805 );
buf ( n42807 , n42631 );
nand ( n42808 , n42806 , n42807 );
buf ( n42809 , n42808 );
buf ( n42810 , n42809 );
nand ( n42811 , n42790 , n42810 );
buf ( n42812 , n42811 );
buf ( n42813 , n42812 );
buf ( n42814 , n42008 );
not ( n42815 , n42814 );
buf ( n42816 , n39478 );
not ( n42817 , n42816 );
or ( n42818 , n42815 , n42817 );
buf ( n42819 , n33076 );
buf ( n42820 , n42017 );
nand ( n42821 , n42819 , n42820 );
buf ( n42822 , n42821 );
buf ( n42823 , n42822 );
nand ( n42824 , n42818 , n42823 );
buf ( n42825 , n42824 );
buf ( n42826 , n42825 );
not ( n42827 , n42826 );
buf ( n42828 , n36101 );
not ( n42829 , n42828 );
or ( n42830 , n42827 , n42829 );
buf ( n42831 , n42516 );
buf ( n42832 , n32966 );
not ( n42833 , n42832 );
buf ( n42834 , n42833 );
buf ( n42835 , n42834 );
nand ( n42836 , n42831 , n42835 );
buf ( n42837 , n42836 );
buf ( n42838 , n42837 );
nand ( n42839 , n42830 , n42838 );
buf ( n42840 , n42839 );
buf ( n42841 , n42840 );
buf ( n42842 , n26033 );
buf ( n42843 , n42842 );
buf ( n42844 , n42843 );
buf ( n42845 , n42844 );
buf ( n42846 , n42845 );
buf ( n42847 , n42846 );
and ( n42848 , n42847 , n37602 );
not ( n42849 , n42847 );
and ( n42850 , n42849 , n38834 );
or ( n42851 , n42848 , n42850 );
buf ( n42852 , n36444 );
not ( n42853 , n42852 );
buf ( n42854 , n42853 );
buf ( n42855 , n42854 );
buf ( n42856 , n29535 );
buf ( n42857 , n42856 );
not ( n42858 , n42857 );
buf ( n42859 , n42858 );
buf ( n42860 , n42859 );
buf ( n42861 , n42860 );
buf ( n42862 , n42861 );
buf ( n42863 , n42862 );
not ( n42864 , n42863 );
buf ( n42865 , n42864 );
buf ( n42866 , n42865 );
not ( n42867 , n42866 );
buf ( n42868 , n37602 );
not ( n42869 , n42868 );
or ( n42870 , n42867 , n42869 );
buf ( n42871 , n38798 );
buf ( n42872 , n42862 );
nand ( n42873 , n42871 , n42872 );
buf ( n42874 , n42873 );
buf ( n42875 , n42874 );
nand ( n42876 , n42870 , n42875 );
buf ( n42877 , n42876 );
not ( n42878 , n42877 );
buf ( n42879 , n42878 );
or ( n42880 , n42855 , n42879 );
nand ( n42881 , C1 , n42880 );
buf ( n42882 , n42881 );
buf ( n42883 , n42882 );
xor ( n42884 , n42841 , n42883 );
buf ( n42885 , n39986 );
not ( n42886 , n42885 );
buf ( n42887 , n39205 );
buf ( n42888 , n40009 );
nand ( n42889 , n42887 , n42888 );
buf ( n42890 , n42889 );
not ( n42891 , n39205 );
nand ( n42892 , n24092 , n42891 );
nand ( n42893 , n42890 , n42892 );
buf ( n42894 , n42893 );
not ( n42895 , n42894 );
or ( n42896 , n42886 , n42895 );
buf ( n42897 , n24092 );
not ( n42898 , n42897 );
not ( n42899 , n38821 );
buf ( n42900 , n42899 );
not ( n42901 , n42900 );
or ( n42902 , n42898 , n42901 );
not ( n42903 , n40010 );
nand ( n42904 , n42903 , n38830 );
buf ( n42905 , n42904 );
nand ( n42906 , n42902 , n42905 );
buf ( n42907 , n42906 );
buf ( n42908 , n42907 );
buf ( n42909 , n40002 );
nand ( n42910 , n42908 , n42909 );
buf ( n42911 , n42910 );
buf ( n42912 , n42911 );
nand ( n42913 , n42896 , n42912 );
buf ( n42914 , n42913 );
buf ( n42915 , n42914 );
and ( n42916 , n42884 , n42915 );
and ( n42917 , n42841 , n42883 );
or ( n42918 , n42916 , n42917 );
buf ( n42919 , n42918 );
buf ( n42920 , n42919 );
xor ( n42921 , n42813 , n42920 );
buf ( n42922 , n42339 );
not ( n42923 , n42922 );
buf ( n42924 , n37968 );
not ( n42925 , n42924 );
buf ( n42926 , n42925 );
buf ( n42927 , n42926 );
not ( n42928 , n42927 );
buf ( n42929 , n42928 );
xnor ( n42930 , n42929 , n42350 );
buf ( n42931 , n42930 );
not ( n42932 , n42931 );
or ( n42933 , n42923 , n42932 );
buf ( n42934 , n42343 );
not ( n42935 , n42934 );
buf ( n42936 , n38218 );
not ( n42937 , n42936 );
or ( n42938 , n42935 , n42937 );
buf ( n42939 , n39406 );
not ( n42940 , n42939 );
buf ( n42941 , n42940 );
buf ( n42942 , n42941 );
buf ( n42943 , n42350 );
nand ( n42944 , n42942 , n42943 );
buf ( n42945 , n42944 );
buf ( n42946 , n42945 );
nand ( n42947 , n42938 , n42946 );
buf ( n42948 , n42947 );
buf ( n42949 , n42948 );
buf ( n42950 , n42378 );
nand ( n42951 , n42949 , n42950 );
buf ( n42952 , n42951 );
buf ( n42953 , n42952 );
nand ( n42954 , n42933 , n42953 );
buf ( n42955 , n42954 );
buf ( n42956 , n42955 );
and ( n42957 , n42921 , n42956 );
and ( n42958 , n42813 , n42920 );
or ( n42959 , n42957 , n42958 );
buf ( n42960 , n42959 );
buf ( n42961 , n42960 );
nand ( n42962 , n42785 , n42961 );
buf ( n42963 , n42962 );
buf ( n42964 , n42963 );
nand ( n42965 , n42782 , n42964 );
buf ( n42966 , n42965 );
buf ( n42967 , n39986 );
not ( n42968 , n42967 );
buf ( n42969 , n24092 );
not ( n42970 , n42969 );
buf ( n42971 , n38477 );
not ( n42972 , n42971 );
buf ( n42973 , n42972 );
buf ( n42974 , n42973 );
not ( n42975 , n42974 );
or ( n42976 , n42970 , n42975 );
buf ( n42977 , n37783 );
buf ( n42978 , n40009 );
nand ( n42979 , n42977 , n42978 );
buf ( n42980 , n42979 );
buf ( n42981 , n42980 );
nand ( n42982 , n42976 , n42981 );
buf ( n42983 , n42982 );
buf ( n42984 , n42983 );
not ( n42985 , n42984 );
or ( n42986 , n42968 , n42985 );
buf ( n42987 , n40010 );
not ( n42988 , n42987 );
buf ( n42989 , n37598 );
not ( n42990 , n42989 );
buf ( n42991 , n42990 );
buf ( n42992 , n42991 );
not ( n42993 , n42992 );
or ( n42994 , n42988 , n42993 );
buf ( n42995 , n39489 );
buf ( n42996 , n40009 );
nand ( n42997 , n42995 , n42996 );
buf ( n42998 , n42997 );
buf ( n42999 , n42998 );
nand ( n43000 , n42994 , n42999 );
buf ( n43001 , n43000 );
buf ( n43002 , n43001 );
buf ( n43003 , n40002 );
nand ( n43004 , n43002 , n43003 );
buf ( n43005 , n43004 );
buf ( n43006 , n43005 );
nand ( n43007 , n42986 , n43006 );
buf ( n43008 , n43007 );
buf ( n43009 , n43008 );
buf ( n43010 , n41647 );
not ( n43011 , n43010 );
buf ( n43012 , n41666 );
not ( n43013 , n43012 );
buf ( n43014 , n39407 );
not ( n43015 , n43014 );
or ( n43016 , n43013 , n43015 );
buf ( n43017 , n42941 );
buf ( n43018 , n41663 );
nand ( n43019 , n43017 , n43018 );
buf ( n43020 , n43019 );
buf ( n43021 , n43020 );
nand ( n43022 , n43016 , n43021 );
buf ( n43023 , n43022 );
buf ( n43024 , n43023 );
not ( n43025 , n43024 );
or ( n43026 , n43011 , n43025 );
buf ( n43027 , n41666 );
not ( n43028 , n43027 );
buf ( n43029 , n38244 );
not ( n43030 , n43029 );
buf ( n43031 , n43030 );
buf ( n43032 , n43031 );
not ( n43033 , n43032 );
or ( n43034 , n43028 , n43033 );
buf ( n43035 , n38244 );
buf ( n43036 , n41663 );
nand ( n43037 , n43035 , n43036 );
buf ( n43038 , n43037 );
buf ( n43039 , n43038 );
nand ( n43040 , n43034 , n43039 );
buf ( n43041 , n43040 );
buf ( n43042 , n43041 );
buf ( n43043 , n41705 );
nand ( n43044 , n43042 , n43043 );
buf ( n43045 , n43044 );
buf ( n43046 , n43045 );
nand ( n43047 , n43026 , n43046 );
buf ( n43048 , n43047 );
buf ( n43049 , n43048 );
xor ( n43050 , n43009 , n43049 );
buf ( n43051 , n36444 );
buf ( n43052 , n43051 );
buf ( n43053 , n43052 );
buf ( n43054 , n43053 );
not ( n43055 , n29499 );
not ( n43056 , n43055 );
buf ( n43057 , n43056 );
not ( n43058 , n43057 );
buf ( n43059 , n37649 );
not ( n43060 , n43059 );
or ( n43061 , n43058 , n43060 );
buf ( n43062 , n36360 );
buf ( n43063 , n29500 );
not ( n43064 , n43063 );
buf ( n43065 , n43064 );
nand ( n43066 , n43062 , n43065 );
buf ( n43067 , n43066 );
buf ( n43068 , n43067 );
nand ( n43069 , n43061 , n43068 );
buf ( n43070 , n43069 );
buf ( n43071 , n43070 );
nand ( n43072 , n43054 , n43071 );
buf ( n43073 , n43072 );
buf ( n43074 , n43073 );
nand ( n43075 , C1 , n43074 );
buf ( n43076 , n43075 );
buf ( n43077 , n43076 );
buf ( n43078 , n39986 );
not ( n43079 , n43078 );
buf ( n43080 , n43001 );
not ( n43081 , n43080 );
or ( n43082 , n43079 , n43081 );
not ( n43083 , n42892 );
not ( n43084 , n42890 );
or ( n43085 , n43083 , n43084 );
nand ( n43086 , n43085 , n40002 );
buf ( n43087 , n43086 );
nand ( n43088 , n43082 , n43087 );
buf ( n43089 , n43088 );
buf ( n43090 , n43089 );
xor ( n43091 , n43077 , n43090 );
buf ( n43092 , n36982 );
buf ( n43093 , n42082 );
not ( n43094 , n43093 );
buf ( n43095 , n43094 );
buf ( n43096 , n43095 );
buf ( n43097 , n13653 );
not ( n43098 , n43097 );
buf ( n43099 , n43098 );
buf ( n43100 , n43099 );
and ( n43101 , n43096 , n43100 );
buf ( n43102 , n42062 );
not ( n43103 , n43102 );
buf ( n43104 , n43103 );
buf ( n43105 , n43104 );
buf ( n43106 , n43099 );
not ( n43107 , n43106 );
buf ( n43108 , n43107 );
buf ( n43109 , n43108 );
and ( n43110 , n43105 , n43109 );
nor ( n43111 , n43101 , n43110 );
buf ( n43112 , n43111 );
buf ( n43113 , n43112 );
or ( n43114 , n43092 , n43113 );
buf ( n43115 , n42066 );
buf ( n43116 , n36909 );
or ( n43117 , n43115 , n43116 );
nand ( n43118 , n43114 , n43117 );
buf ( n43119 , n43118 );
buf ( n43120 , n43119 );
and ( n43121 , n43091 , n43120 );
and ( n43122 , n43077 , n43090 );
or ( n43123 , n43121 , n43122 );
buf ( n43124 , n43123 );
buf ( n43125 , n43124 );
xor ( n43126 , n43050 , n43125 );
buf ( n43127 , n43126 );
not ( n43128 , n43127 );
xor ( n43129 , n42555 , n42638 );
xor ( n43130 , n43129 , n42643 );
buf ( n43131 , n43130 );
not ( n43132 , n43131 );
or ( n43133 , n43128 , n43132 );
or ( n43134 , n43127 , n43131 );
xor ( n43135 , n42447 , n42500 );
xor ( n43136 , n43135 , n42550 );
buf ( n43137 , n43136 );
buf ( n43138 , n43137 );
buf ( n43139 , n41705 );
not ( n43140 , n43139 );
not ( n43141 , n41666 );
buf ( n43142 , n37264 );
not ( n43143 , n43142 );
not ( n43144 , n43143 );
or ( n43145 , n43141 , n43144 );
buf ( n43146 , n37265 );
buf ( n43147 , n41663 );
nand ( n43148 , n43146 , n43147 );
buf ( n43149 , n43148 );
nand ( n43150 , n43145 , n43149 );
buf ( n43151 , n43150 );
not ( n43152 , n43151 );
or ( n43153 , n43140 , n43152 );
buf ( n43154 , n43041 );
buf ( n43155 , n41647 );
nand ( n43156 , n43154 , n43155 );
buf ( n43157 , n43156 );
buf ( n43158 , n43157 );
nand ( n43159 , n43153 , n43158 );
buf ( n43160 , n43159 );
buf ( n43161 , n43160 );
or ( n43162 , n43138 , n43161 );
xor ( n43163 , n43077 , n43090 );
xor ( n43164 , n43163 , n43120 );
buf ( n43165 , n43164 );
buf ( n43166 , n43165 );
nand ( n43167 , n43162 , n43166 );
buf ( n43168 , n43167 );
buf ( n43169 , n43168 );
buf ( n43170 , n43160 );
buf ( n43171 , n43137 );
nand ( n43172 , n43170 , n43171 );
buf ( n43173 , n43172 );
buf ( n43174 , n43173 );
nand ( n43175 , n43169 , n43174 );
buf ( n43176 , n43175 );
nand ( n43177 , n43134 , n43176 );
nand ( n43178 , n43133 , n43177 );
xor ( n43179 , n42966 , n43178 );
xor ( n43180 , n43009 , n43049 );
and ( n43181 , n43180 , n43125 );
and ( n43182 , n43009 , n43049 );
or ( n43183 , n43181 , n43182 );
buf ( n43184 , n43183 );
buf ( n43185 , n43184 );
buf ( n43186 , n40002 );
not ( n43187 , n43186 );
buf ( n43188 , n42983 );
not ( n43189 , n43188 );
or ( n43190 , n43187 , n43189 );
buf ( n43191 , n24092 );
not ( n43192 , n43191 );
buf ( n43193 , n37745 );
not ( n43194 , n43193 );
or ( n43195 , n43192 , n43194 );
buf ( n43196 , n37742 );
buf ( n43197 , n43196 );
buf ( n43198 , n43197 );
buf ( n43199 , n43198 );
buf ( n43200 , n40009 );
nand ( n43201 , n43199 , n43200 );
buf ( n43202 , n43201 );
buf ( n43203 , n43202 );
nand ( n43204 , n43195 , n43203 );
buf ( n43205 , n43204 );
buf ( n43206 , n43205 );
buf ( n43207 , n39986 );
nand ( n43208 , n43206 , n43207 );
buf ( n43209 , n43208 );
buf ( n43210 , n43209 );
nand ( n43211 , n43190 , n43210 );
buf ( n43212 , n43211 );
buf ( n43213 , n43212 );
buf ( n43214 , n42631 );
not ( n43215 , n43214 );
buf ( n43216 , n42587 );
not ( n43217 , n43216 );
or ( n43218 , n43215 , n43217 );
buf ( n43219 , n25160 );
not ( n43220 , n43219 );
buf ( n43221 , n37295 );
not ( n43222 , n43221 );
or ( n43223 , n43220 , n43222 );
not ( n43224 , n37293 );
buf ( n43225 , n43224 );
not ( n43226 , n43225 );
buf ( n43227 , n42581 );
nand ( n43228 , n43226 , n43227 );
buf ( n43229 , n43228 );
buf ( n43230 , n43229 );
nand ( n43231 , n43223 , n43230 );
buf ( n43232 , n43231 );
buf ( n43233 , n43232 );
buf ( n43234 , n42566 );
nand ( n43235 , n43233 , n43234 );
buf ( n43236 , n43235 );
buf ( n43237 , n43236 );
nand ( n43238 , n43218 , n43237 );
buf ( n43239 , n43238 );
buf ( n43240 , n43239 );
xor ( n43241 , n43213 , n43240 );
buf ( n43242 , n42446 );
not ( n43243 , n43242 );
buf ( n43244 , n43243 );
buf ( n43245 , n43244 );
buf ( n43246 , n42543 );
not ( n43247 , n43246 );
buf ( n43248 , n36095 );
not ( n43249 , n43248 );
buf ( n43250 , n43249 );
buf ( n43251 , n43250 );
not ( n43252 , n43251 );
or ( n43253 , n43247 , n43252 );
buf ( n43254 , n32969 );
buf ( n43255 , n43108 );
not ( n43256 , n43255 );
buf ( n43257 , n33076 );
not ( n43258 , n43257 );
buf ( n43259 , n43258 );
buf ( n43260 , n43259 );
not ( n43261 , n43260 );
or ( n43262 , n43256 , n43261 );
buf ( n43263 , n36500 );
not ( n43264 , n43263 );
buf ( n43265 , n43264 );
buf ( n43266 , n43265 );
buf ( n43267 , n43099 );
nand ( n43268 , n43266 , n43267 );
buf ( n43269 , n43268 );
buf ( n43270 , n43269 );
nand ( n43271 , n43262 , n43270 );
buf ( n43272 , n43271 );
buf ( n43273 , n43272 );
nand ( n43274 , n43254 , n43273 );
buf ( n43275 , n43274 );
buf ( n43276 , n43275 );
nand ( n43277 , n43253 , n43276 );
buf ( n43278 , n43277 );
buf ( n43279 , n43278 );
xor ( n43280 , n43245 , n43279 );
buf ( n43281 , n43053 );
not ( n43282 , n43281 );
buf ( n43283 , n43282 );
buf ( n43284 , n43283 );
buf ( n43285 , n42001 );
or ( n43286 , n43284 , n43285 );
nand ( n43287 , C1 , n43286 );
buf ( n43288 , n43287 );
buf ( n43289 , n43288 );
and ( n43290 , n43280 , n43289 );
and ( n43291 , n43245 , n43279 );
or ( n43292 , n43290 , n43291 );
buf ( n43293 , n43292 );
buf ( n43294 , n43293 );
xor ( n43295 , n43241 , n43294 );
buf ( n43296 , n43295 );
buf ( n43297 , n43296 );
xor ( n43298 , n43185 , n43297 );
buf ( n43299 , n38382 );
not ( n43300 , n43299 );
buf ( n43301 , n38413 );
not ( n43302 , n43301 );
buf ( n43303 , n38851 );
not ( n43304 , n43303 );
or ( n43305 , n43302 , n43304 );
buf ( n43306 , n30187 );
not ( n43307 , n43306 );
buf ( n43308 , n43307 );
buf ( n43309 , n43308 );
buf ( n43310 , n43309 );
buf ( n43311 , n43310 );
buf ( n43312 , n43311 );
not ( n43313 , n43312 );
buf ( n43314 , n43313 );
buf ( n43315 , n43314 );
buf ( n43316 , n38412 );
nand ( n43317 , n43315 , n43316 );
buf ( n43318 , n43317 );
buf ( n43319 , n43318 );
nand ( n43320 , n43305 , n43319 );
buf ( n43321 , n43320 );
buf ( n43322 , n43321 );
not ( n43323 , n43322 );
or ( n43324 , n43300 , n43323 );
buf ( n43325 , n42441 );
not ( n43326 , n43325 );
buf ( n43327 , n38775 );
nand ( n43328 , n43326 , n43327 );
buf ( n43329 , n43328 );
buf ( n43330 , n43329 );
nand ( n43331 , n43324 , n43330 );
buf ( n43332 , n43331 );
buf ( n43333 , n43332 );
buf ( n43334 , n42448 );
not ( n43335 , n43334 );
buf ( n43336 , n39000 );
not ( n43337 , n43336 );
buf ( n43338 , n37642 );
not ( n43339 , n43338 );
or ( n43340 , n43337 , n43339 );
buf ( n43341 , n39205 );
buf ( n43342 , n38997 );
nand ( n43343 , n43341 , n43342 );
buf ( n43344 , n43343 );
buf ( n43345 , n43344 );
nand ( n43346 , n43340 , n43345 );
buf ( n43347 , n43346 );
buf ( n43348 , n43347 );
not ( n43349 , n43348 );
or ( n43350 , n43335 , n43349 );
buf ( n43351 , n42477 );
buf ( n43352 , n38985 );
nand ( n43353 , n43351 , n43352 );
buf ( n43354 , n43353 );
buf ( n43355 , n43354 );
nand ( n43356 , n43350 , n43355 );
buf ( n43357 , n43356 );
buf ( n43358 , n43357 );
xor ( n43359 , n43333 , n43358 );
buf ( n43360 , n29407 );
not ( n43361 , n43360 );
buf ( n43362 , n43361 );
buf ( n43363 , n43362 );
buf ( n43364 , n43363 );
buf ( n43365 , n43364 );
buf ( n43366 , n43365 );
not ( n43367 , n43366 );
buf ( n43368 , n43367 );
buf ( n43369 , n43368 );
not ( n43370 , n43369 );
buf ( n43371 , n36878 );
buf ( n43372 , n43371 );
not ( n43373 , n43372 );
or ( n43374 , n43370 , n43373 );
buf ( n43375 , n38108 );
buf ( n43376 , n43365 );
nand ( n43377 , n43375 , n43376 );
buf ( n43378 , n43377 );
buf ( n43379 , n43378 );
nand ( n43380 , n43374 , n43379 );
buf ( n43381 , n43380 );
buf ( n43382 , n43381 );
not ( n43383 , n43382 );
buf ( n43384 , n38124 );
not ( n43385 , n43384 );
buf ( n43386 , n43385 );
buf ( n43387 , n43386 );
buf ( n43388 , n43387 );
buf ( n43389 , n43388 );
buf ( n43390 , n43389 );
not ( n43391 , n43390 );
or ( n43392 , n43383 , n43391 );
buf ( n43393 , n42152 );
not ( n43394 , n43393 );
buf ( n43395 , n38068 );
not ( n43396 , n43395 );
or ( n43397 , n43394 , n43396 );
buf ( n43398 , n36878 );
not ( n43399 , n43398 );
buf ( n43400 , n43399 );
buf ( n43401 , n43400 );
buf ( n43402 , n43401 );
buf ( n43403 , n43402 );
buf ( n43404 , n43403 );
buf ( n43405 , n42160 );
nand ( n43406 , n43404 , n43405 );
buf ( n43407 , n43406 );
buf ( n43408 , n43407 );
nand ( n43409 , n43397 , n43408 );
buf ( n43410 , n43409 );
buf ( n43411 , n43410 );
buf ( n43412 , n38057 );
not ( n43413 , n43412 );
buf ( n43414 , n43413 );
buf ( n43415 , n43414 );
nand ( n43416 , n43411 , n43415 );
buf ( n43417 , n43416 );
buf ( n43418 , n43417 );
nand ( n43419 , n43392 , n43418 );
buf ( n43420 , n43419 );
buf ( n43421 , n43420 );
and ( n43422 , n43359 , n43421 );
and ( n43423 , n43333 , n43358 );
or ( n43424 , n43422 , n43423 );
buf ( n43425 , n43424 );
buf ( n43426 , n43425 );
buf ( n43427 , n41809 );
not ( n43428 , n43427 );
buf ( n43429 , n37400 );
not ( n43430 , n43429 );
or ( n43431 , n43428 , n43430 );
buf ( n43432 , n37328 );
not ( n43433 , n43432 );
buf ( n43434 , n43433 );
buf ( n43435 , n43434 );
not ( n43436 , n43435 );
buf ( n43437 , n42425 );
not ( n43438 , n43437 );
or ( n43439 , n43436 , n43438 );
buf ( n43440 , n41769 );
not ( n43441 , n43440 );
buf ( n43442 , n43441 );
buf ( n43443 , n43442 );
buf ( n43444 , n39682 );
not ( n43445 , n43444 );
buf ( n43446 , n43445 );
buf ( n43447 , n43446 );
nand ( n43448 , n43443 , n43447 );
buf ( n43449 , n43448 );
buf ( n43450 , n43449 );
nand ( n43451 , n43439 , n43450 );
buf ( n43452 , n43451 );
buf ( n43453 , n43452 );
buf ( n43454 , n37413 );
nand ( n43455 , n43453 , n43454 );
buf ( n43456 , n43455 );
buf ( n43457 , n43456 );
nand ( n43458 , n43431 , n43457 );
buf ( n43459 , n43458 );
buf ( n43460 , n43459 );
buf ( n43461 , n43460 );
buf ( n43462 , n43461 );
buf ( n43463 , n43462 );
buf ( n43464 , n38412 );
buf ( n43465 , n38830 );
and ( n43466 , n43464 , n43465 );
not ( n43467 , n43464 );
buf ( n43468 , n42458 );
not ( n43469 , n43468 );
buf ( n43470 , n43469 );
buf ( n43471 , n43470 );
and ( n43472 , n43467 , n43471 );
nor ( n43473 , n43466 , n43472 );
buf ( n43474 , n43473 );
buf ( n43475 , n43474 );
not ( n43476 , n43475 );
buf ( n43477 , n38383 );
not ( n43478 , n43477 );
and ( n43479 , n43476 , n43478 );
buf ( n43480 , n43321 );
buf ( n43481 , n38775 );
and ( n43482 , n43480 , n43481 );
nor ( n43483 , n43479 , n43482 );
buf ( n43484 , n43483 );
buf ( n43485 , n43484 );
not ( n43486 , n43485 );
buf ( n43487 , n43486 );
buf ( n43488 , n43487 );
xor ( n43489 , n43463 , n43488 );
buf ( n43490 , n43272 );
not ( n43491 , n43490 );
buf ( n43492 , n36104 );
not ( n43493 , n43492 );
or ( n43494 , n43491 , n43493 );
buf ( n43495 , n39718 );
buf ( n43496 , n42055 );
not ( n43497 , n43496 );
buf ( n43498 , n39478 );
not ( n43499 , n43498 );
or ( n43500 , n43497 , n43499 );
buf ( n43501 , n39493 );
not ( n43502 , n43501 );
buf ( n43503 , n43502 );
buf ( n43504 , n43503 );
buf ( n43505 , n42052 );
nand ( n43506 , n43504 , n43505 );
buf ( n43507 , n43506 );
buf ( n43508 , n43507 );
nand ( n43509 , n43500 , n43508 );
buf ( n43510 , n43509 );
buf ( n43511 , n43510 );
nand ( n43512 , n43495 , n43511 );
buf ( n43513 , n43512 );
buf ( n43514 , n43513 );
nand ( n43515 , n43494 , n43514 );
buf ( n43516 , n43515 );
buf ( n43517 , n43516 );
xnor ( n43518 , n43489 , n43517 );
buf ( n43519 , n43518 );
buf ( n43520 , n43519 );
xor ( n43521 , n43426 , n43520 );
buf ( n43522 , n41705 );
not ( n43523 , n43522 );
buf ( n43524 , n43023 );
not ( n43525 , n43524 );
or ( n43526 , n43523 , n43525 );
buf ( n43527 , n41647 );
buf ( n43528 , n41693 );
nand ( n43529 , n43527 , n43528 );
buf ( n43530 , n43529 );
buf ( n43531 , n43530 );
nand ( n43532 , n43526 , n43531 );
buf ( n43533 , n43532 );
buf ( n43534 , n43533 );
xor ( n43535 , n43521 , n43534 );
buf ( n43536 , n43535 );
buf ( n43537 , n43536 );
xor ( n43538 , n43298 , n43537 );
buf ( n43539 , n43538 );
and ( n43540 , n43179 , n43539 );
and ( n43541 , n42966 , n43178 );
or ( n43542 , n43540 , n43541 );
xor ( n43543 , n42726 , n43542 );
buf ( n43544 , n43184 );
not ( n43545 , n43544 );
buf ( n43546 , n43296 );
not ( n43547 , n43546 );
or ( n43548 , n43545 , n43547 );
or ( n43549 , n43296 , n43184 );
nand ( n43550 , n43549 , n43536 );
buf ( n43551 , n43550 );
nand ( n43552 , n43548 , n43551 );
buf ( n43553 , n43552 );
buf ( n43554 , n43553 );
xor ( n43555 , n43213 , n43240 );
and ( n43556 , n43555 , n43294 );
and ( n43557 , n43213 , n43240 );
or ( n43558 , n43556 , n43557 );
buf ( n43559 , n43558 );
buf ( n43560 , n43559 );
buf ( n43561 , n42712 );
not ( n43562 , n43561 );
buf ( n43563 , n42685 );
not ( n43564 , n43563 );
or ( n43565 , n43562 , n43564 );
buf ( n43566 , n42672 );
not ( n43567 , n43566 );
buf ( n43568 , n39927 );
not ( n43569 , n43568 );
or ( n43570 , n43567 , n43569 );
buf ( n43571 , n39924 );
buf ( n43572 , n42671 );
nand ( n43573 , n43571 , n43572 );
buf ( n43574 , n43573 );
buf ( n43575 , n43574 );
nand ( n43576 , n43570 , n43575 );
buf ( n43577 , n43576 );
buf ( n43578 , n43577 );
buf ( n43579 , n42668 );
nand ( n43580 , n43578 , n43579 );
buf ( n43581 , n43580 );
buf ( n43582 , n43581 );
nand ( n43583 , n43565 , n43582 );
buf ( n43584 , n43583 );
buf ( n43585 , n43584 );
xor ( n43586 , n43560 , n43585 );
xor ( n43587 , n43426 , n43520 );
and ( n43588 , n43587 , n43534 );
and ( n43589 , n43426 , n43520 );
or ( n43590 , n43588 , n43589 );
buf ( n43591 , n43590 );
buf ( n43592 , n43591 );
xor ( n43593 , n43586 , n43592 );
buf ( n43594 , n43593 );
buf ( n43595 , n43594 );
xor ( n43596 , n43554 , n43595 );
not ( n43597 , n36395 );
xnor ( n43598 , n42343 , n43597 );
buf ( n43599 , n43598 );
buf ( n43600 , n42339 );
and ( n43601 , n43599 , n43600 );
buf ( n43602 , n42356 );
not ( n43603 , n43602 );
buf ( n43604 , n42375 );
nor ( n43605 , n43603 , n43604 );
buf ( n43606 , n43605 );
buf ( n43607 , n43606 );
nor ( n43608 , n43601 , n43607 );
buf ( n43609 , n43608 );
or ( n43610 , n41962 , n41988 );
nand ( n43611 , n42030 , n43610 );
and ( n43612 , n41963 , n41989 );
buf ( n43613 , n43612 );
not ( n43614 , n43613 );
nand ( n43615 , n43611 , n43614 );
buf ( n43616 , n43615 );
not ( n43617 , n43616 );
buf ( n43618 , n40010 );
not ( n43619 , n43618 );
buf ( n43620 , n42573 );
not ( n43621 , n43620 );
or ( n43622 , n43619 , n43621 );
buf ( n43623 , n37708 );
not ( n43624 , n43623 );
buf ( n43625 , n43624 );
buf ( n43626 , n43625 );
buf ( n43627 , n40009 );
nand ( n43628 , n43626 , n43627 );
buf ( n43629 , n43628 );
buf ( n43630 , n43629 );
nand ( n43631 , n43622 , n43630 );
buf ( n43632 , n43631 );
buf ( n43633 , n43632 );
buf ( n43634 , n39986 );
and ( n43635 , n43633 , n43634 );
buf ( n43636 , n43205 );
not ( n43637 , n43636 );
buf ( n43638 , n40005 );
nor ( n43639 , n43637 , n43638 );
buf ( n43640 , n43639 );
buf ( n43641 , n43640 );
nor ( n43642 , n43635 , n43641 );
buf ( n43643 , n43642 );
buf ( n43644 , n43643 );
buf ( n43645 , n43462 );
not ( n43646 , n43645 );
buf ( n43647 , n43484 );
not ( n43648 , n43647 );
or ( n43649 , n43646 , n43648 );
buf ( n43650 , n43516 );
nand ( n43651 , n43649 , n43650 );
buf ( n43652 , n43651 );
buf ( n43653 , n43652 );
buf ( n43654 , n43462 );
not ( n43655 , n43654 );
buf ( n43656 , n43487 );
nand ( n43657 , n43655 , n43656 );
buf ( n43658 , n43657 );
buf ( n43659 , n43658 );
nand ( n43660 , n43653 , n43659 );
buf ( n43661 , n43660 );
buf ( n43662 , n43661 );
xor ( n43663 , n43644 , n43662 );
buf ( n43664 , n43663 );
buf ( n43665 , n43664 );
not ( n43666 , n43665 );
or ( n43667 , n43617 , n43666 );
buf ( n43668 , n43664 );
buf ( n43669 , n43615 );
or ( n43670 , n43668 , n43669 );
nand ( n43671 , n43667 , n43670 );
buf ( n43672 , n43671 );
xor ( n43673 , n43609 , n43672 );
buf ( n43674 , n39000 );
not ( n43675 , n43674 );
buf ( n43676 , n38477 );
not ( n43677 , n43676 );
buf ( n43678 , n43677 );
buf ( n43679 , n43678 );
not ( n43680 , n43679 );
or ( n43681 , n43675 , n43680 );
buf ( n43682 , n42795 );
not ( n43683 , n43682 );
buf ( n43684 , n43683 );
buf ( n43685 , n43684 );
buf ( n43686 , n38997 );
nand ( n43687 , n43685 , n43686 );
buf ( n43688 , n43687 );
buf ( n43689 , n43688 );
nand ( n43690 , n43681 , n43689 );
buf ( n43691 , n43690 );
buf ( n43692 , n43691 );
buf ( n43693 , n39374 );
and ( n43694 , n43692 , n43693 );
buf ( n43695 , n39000 );
not ( n43696 , n43695 );
buf ( n43697 , n37595 );
not ( n43698 , n43697 );
or ( n43699 , n43696 , n43698 );
buf ( n43700 , n37586 );
buf ( n43701 , n38997 );
nand ( n43702 , n43700 , n43701 );
buf ( n43703 , n43702 );
buf ( n43704 , n43703 );
nand ( n43705 , n43699 , n43704 );
buf ( n43706 , n43705 );
buf ( n43707 , n43706 );
not ( n43708 , n43707 );
buf ( n43709 , n38988 );
nor ( n43710 , n43708 , n43709 );
buf ( n43711 , n43710 );
buf ( n43712 , n43711 );
nor ( n43713 , n43694 , n43712 );
buf ( n43714 , n43713 );
buf ( n43715 , n43714 );
not ( n43716 , n43715 );
buf ( n43717 , n39806 );
not ( n43718 , n43717 );
buf ( n43719 , n43718 );
buf ( n43720 , n43719 );
not ( n43721 , n43720 );
buf ( n43722 , n41754 );
not ( n43723 , n43722 );
buf ( n43724 , n43723 );
buf ( n43725 , n43724 );
not ( n43726 , n43725 );
and ( n43727 , n43721 , n43726 );
buf ( n43728 , n36640 );
buf ( n43729 , n43099 );
buf ( n43730 , n39729 );
and ( n43731 , n43729 , n43730 );
not ( n43732 , n43729 );
buf ( n43733 , n41741 );
and ( n43734 , n43732 , n43733 );
nor ( n43735 , n43731 , n43734 );
buf ( n43736 , n43735 );
buf ( n43737 , n43736 );
nor ( n43738 , n43728 , n43737 );
buf ( n43739 , n43738 );
buf ( n43740 , n43739 );
nor ( n43741 , n43727 , n43740 );
buf ( n43742 , n43741 );
buf ( n43743 , n43742 );
not ( n43744 , n43743 );
buf ( n43745 , n43744 );
buf ( n43746 , n43745 );
not ( n43747 , n43746 );
or ( n43748 , n43716 , n43747 );
buf ( n43749 , n43714 );
not ( n43750 , n43749 );
buf ( n43751 , n43750 );
buf ( n43752 , n43751 );
buf ( n43753 , n43742 );
nand ( n43754 , n43752 , n43753 );
buf ( n43755 , n43754 );
buf ( n43756 , n43755 );
nand ( n43757 , n43748 , n43756 );
buf ( n43758 , n43757 );
buf ( n43759 , n43758 );
buf ( n43760 , n43459 );
not ( n43761 , n41984 );
buf ( n43762 , n43761 );
not ( n43763 , n43762 );
buf ( n43764 , n37514 );
not ( n43765 , n43764 );
buf ( n43766 , n43765 );
buf ( n43767 , n43766 );
not ( n43768 , n43767 );
or ( n43769 , n43763 , n43768 );
buf ( n43770 , n41844 );
not ( n43771 , n43770 );
buf ( n43772 , n39656 );
not ( n43773 , n43772 );
or ( n43774 , n43771 , n43773 );
buf ( n43775 , n39656 );
buf ( n43776 , n43775 );
buf ( n43777 , n43776 );
buf ( n43778 , n43777 );
not ( n43779 , n43778 );
not ( n43780 , n41844 );
buf ( n43781 , n43780 );
nand ( n43782 , n43779 , n43781 );
buf ( n43783 , n43782 );
buf ( n43784 , n43783 );
nand ( n43785 , n43774 , n43784 );
buf ( n43786 , n43785 );
buf ( n43787 , n43786 );
buf ( n43788 , n41852 );
nand ( n43789 , n43787 , n43788 );
buf ( n43790 , n43789 );
buf ( n43791 , n43790 );
nand ( n43792 , n43769 , n43791 );
buf ( n43793 , n43792 );
buf ( n43794 , n43793 );
xor ( n43795 , n43760 , n43794 );
buf ( n43796 , n41862 );
not ( n43797 , n43796 );
buf ( n43798 , n43797 );
buf ( n43799 , n43798 );
buf ( n43800 , n41957 );
not ( n43801 , n43800 );
buf ( n43802 , n43801 );
buf ( n43803 , n43802 );
or ( n43804 , n43799 , n43803 );
buf ( n43805 , n41908 );
not ( n43806 , n41835 );
buf ( n43807 , n43806 );
buf ( n43808 , n41925 );
and ( n43809 , n43807 , n43808 );
not ( n43810 , n43807 );
buf ( n43811 , n41925 );
not ( n43812 , n43811 );
buf ( n43813 , n43812 );
buf ( n43814 , n43813 );
and ( n43815 , n43810 , n43814 );
nor ( n43816 , n43809 , n43815 );
buf ( n43817 , n43816 );
buf ( n43818 , n43817 );
or ( n43819 , n43805 , n43818 );
nand ( n43820 , n43804 , n43819 );
buf ( n43821 , n43820 );
buf ( n43822 , n43821 );
xor ( n43823 , n43795 , n43822 );
buf ( n43824 , n43823 );
buf ( n43825 , n43824 );
xnor ( n43826 , n43759 , n43825 );
buf ( n43827 , n43826 );
xor ( n43828 , n43673 , n43827 );
buf ( n43829 , n43828 );
xor ( n43830 , n43596 , n43829 );
buf ( n43831 , n43830 );
xor ( n43832 , n43543 , n43831 );
not ( n43833 , n43832 );
buf ( n43834 , n41611 );
buf ( n43835 , n36611 );
and ( n43836 , n43834 , n43835 );
not ( n43837 , n43834 );
buf ( n43838 , n36614 );
and ( n43839 , n43837 , n43838 );
nor ( n43840 , n43836 , n43839 );
buf ( n43841 , n43840 );
buf ( n43842 , n43841 );
not ( n43843 , n43842 );
buf ( n43844 , n41599 );
not ( n43845 , n43844 );
and ( n43846 , n43843 , n43845 );
buf ( n43847 , n41611 );
not ( n43848 , n43847 );
buf ( n43849 , n36032 );
not ( n43850 , n43849 );
buf ( n43851 , n43850 );
buf ( n43852 , n43851 );
not ( n43853 , n43852 );
or ( n43854 , n43848 , n43853 );
buf ( n43855 , n43851 );
not ( n43856 , n43855 );
buf ( n43857 , n43856 );
buf ( n43858 , n43857 );
buf ( n43859 , n41608 );
nand ( n43860 , n43858 , n43859 );
buf ( n43861 , n43860 );
buf ( n43862 , n43861 );
nand ( n43863 , n43854 , n43862 );
buf ( n43864 , n43863 );
buf ( n43865 , n43864 );
buf ( n43866 , n41577 );
not ( n43867 , n43866 );
buf ( n43868 , n43867 );
buf ( n43869 , n43868 );
and ( n43870 , n43865 , n43869 );
nor ( n43871 , n43846 , n43870 );
buf ( n43872 , n43871 );
buf ( n43873 , n43872 );
not ( n43874 , n43873 );
buf ( n43875 , n25184 );
not ( n43876 , n43875 );
buf ( n43877 , n37264 );
not ( n43878 , n43877 );
buf ( n43879 , n43878 );
buf ( n43880 , n43879 );
not ( n43881 , n43880 );
or ( n43882 , n43876 , n43881 );
buf ( n43883 , n43879 );
not ( n43884 , n43883 );
buf ( n43885 , n43884 );
buf ( n43886 , n43885 );
buf ( n43887 , n25183 );
nand ( n43888 , n43886 , n43887 );
buf ( n43889 , n43888 );
buf ( n43890 , n43889 );
nand ( n43891 , n43882 , n43890 );
buf ( n43892 , n43891 );
buf ( n43893 , n25028 );
not ( n43894 , n43893 );
buf ( n43895 , n43894 );
and ( n43896 , n41698 , n43895 );
not ( n43897 , n41698 );
buf ( n43898 , n25022 );
buf ( n43899 , n25025 );
xnor ( n43900 , n43898 , n43899 );
buf ( n43901 , n43900 );
and ( n43902 , n43897 , n43901 );
nor ( n43903 , n43896 , n43902 );
buf ( n43904 , n43903 );
not ( n43905 , n43904 );
not ( n43906 , n43905 );
buf ( n43907 , n43906 );
not ( n43908 , n43907 );
buf ( n43909 , n43908 );
and ( n43910 , n43892 , n43909 );
buf ( n43911 , n25184 );
not ( n43912 , n43911 );
buf ( n43913 , n38286 );
not ( n43914 , n43913 );
or ( n43915 , n43912 , n43914 );
buf ( n43916 , n37293 );
buf ( n43917 , n25183 );
nand ( n43918 , n43916 , n43917 );
buf ( n43919 , n43918 );
buf ( n43920 , n43919 );
nand ( n43921 , n43915 , n43920 );
buf ( n43922 , n43921 );
not ( n43923 , n43922 );
and ( n43924 , n25179 , n43901 );
not ( n43925 , n25179 );
buf ( n43926 , n43901 );
not ( n43927 , n43926 );
buf ( n43928 , n43927 );
and ( n43929 , n43925 , n43928 );
nor ( n43930 , n43924 , n43929 );
nand ( n43931 , n43930 , n43903 );
buf ( n43932 , n43931 );
buf ( n43933 , n43932 );
not ( n43934 , n43933 );
buf ( n43935 , n43934 );
buf ( n43936 , n43935 );
buf ( n43937 , n43936 );
buf ( n43938 , n43937 );
buf ( n43939 , n43938 );
not ( n43940 , n43939 );
buf ( n43941 , n43940 );
nor ( n43942 , n43923 , n43941 );
nor ( n43943 , n43910 , n43942 );
buf ( n43944 , n43943 );
not ( n43945 , n43944 );
buf ( n43946 , n43945 );
buf ( n43947 , n43946 );
not ( n43948 , n43947 );
or ( n43949 , n43874 , n43948 );
buf ( n43950 , n43946 );
buf ( n43951 , n43872 );
or ( n43952 , n43950 , n43951 );
nand ( n43953 , n43949 , n43952 );
buf ( n43954 , n43953 );
buf ( n43955 , n41993 );
not ( n43956 , n43955 );
buf ( n43957 , n36527 );
not ( n43958 , n43957 );
buf ( n43959 , n43958 );
buf ( n43960 , n43959 );
not ( n43961 , n43960 );
or ( n43962 , n43956 , n43961 );
buf ( n43963 , n36527 );
buf ( n43964 , n41993 );
not ( n43965 , n43964 );
buf ( n43966 , n43965 );
buf ( n43967 , n43966 );
nand ( n43968 , n43963 , n43967 );
buf ( n43969 , n43968 );
buf ( n43970 , n43969 );
nand ( n43971 , n43962 , n43970 );
buf ( n43972 , n43971 );
buf ( n43973 , n43972 );
not ( n43974 , n43973 );
buf ( n43975 , n36523 );
not ( n43976 , n43975 );
or ( n43977 , n43974 , n43976 );
buf ( n43978 , n42104 );
not ( n43979 , n43978 );
buf ( n43980 , n36640 );
not ( n43981 , n43980 );
buf ( n43982 , n43981 );
buf ( n43983 , n43982 );
nand ( n43984 , n43979 , n43983 );
buf ( n43985 , n43984 );
buf ( n43986 , n43985 );
nand ( n43987 , n43977 , n43986 );
buf ( n43988 , n43987 );
buf ( n43989 , n38127 );
not ( n43990 , n43989 );
buf ( n43991 , n43990 );
buf ( n43992 , n43991 );
not ( n43993 , n43992 );
buf ( n43994 , n42075 );
not ( n43995 , n43994 );
buf ( n43996 , n43995 );
buf ( n43997 , n43996 );
not ( n43998 , n43997 );
buf ( n43999 , n38068 );
not ( n44000 , n43999 );
or ( n44001 , n43998 , n44000 );
buf ( n44002 , n38068 );
not ( n44003 , n44002 );
buf ( n44004 , n44003 );
buf ( n44005 , n44004 );
buf ( n44006 , n42075 );
nand ( n44007 , n44005 , n44006 );
buf ( n44008 , n44007 );
buf ( n44009 , n44008 );
nand ( n44010 , n44001 , n44009 );
buf ( n44011 , n44010 );
buf ( n44012 , n44011 );
not ( n44013 , n44012 );
or ( n44014 , n43993 , n44013 );
buf ( n44015 , n43381 );
buf ( n44016 , n38060 );
nand ( n44017 , n44015 , n44016 );
buf ( n44018 , n44017 );
buf ( n44019 , n44018 );
nand ( n44020 , n44014 , n44019 );
buf ( n44021 , n44020 );
or ( n44022 , n43988 , n44021 );
buf ( n44023 , n42411 );
not ( n44024 , n44023 );
not ( n44025 , n28305 );
buf ( n44026 , n44025 );
not ( n44027 , n44026 );
or ( n44028 , n44024 , n44027 );
buf ( n44029 , n42119 );
not ( n44030 , n44029 );
buf ( n44031 , n42414 );
nand ( n44032 , n44030 , n44031 );
buf ( n44033 , n44032 );
buf ( n44034 , n44033 );
nand ( n44035 , n44028 , n44034 );
buf ( n44036 , n44035 );
buf ( n44037 , n44036 );
not ( n44038 , n44037 );
buf ( n44039 , n38403 );
buf ( n44040 , n44039 );
not ( n44041 , n44040 );
buf ( n44042 , n44041 );
buf ( n44043 , n44042 );
not ( n44044 , n44043 );
or ( n44045 , n44038 , n44044 );
buf ( n44046 , n42411 );
not ( n44047 , n44046 );
buf ( n44048 , n41783 );
not ( n44049 , n44048 );
or ( n44050 , n44047 , n44049 );
buf ( n44051 , n41764 );
buf ( n44052 , n42403 );
buf ( n44053 , n44052 );
buf ( n44054 , n44053 );
buf ( n44055 , n44054 );
nand ( n44056 , n44051 , n44055 );
buf ( n44057 , n44056 );
buf ( n44058 , n44057 );
nand ( n44059 , n44050 , n44058 );
buf ( n44060 , n44059 );
buf ( n44061 , n44060 );
buf ( n44062 , n38380 );
nand ( n44063 , n44061 , n44062 );
buf ( n44064 , n44063 );
buf ( n44065 , n44064 );
nand ( n44066 , n44045 , n44065 );
buf ( n44067 , n44066 );
buf ( n44068 , n44067 );
buf ( n44069 , n38382 );
not ( n44070 , n44069 );
buf ( n44071 , n42418 );
not ( n44072 , n44071 );
buf ( n44073 , n44072 );
buf ( n44074 , n44073 );
not ( n44075 , n44074 );
or ( n44076 , n44070 , n44075 );
buf ( n44077 , n38407 );
not ( n44078 , n44077 );
buf ( n44079 , n44060 );
nand ( n44080 , n44078 , n44079 );
buf ( n44081 , n44080 );
buf ( n44082 , n44081 );
nand ( n44083 , n44076 , n44082 );
buf ( n44084 , n44083 );
buf ( n44085 , n44084 );
xor ( n44086 , n44068 , n44085 );
buf ( n44087 , n41823 );
not ( n44088 , n44087 );
buf ( n44089 , n37328 );
not ( n44090 , n44089 );
or ( n44091 , n44088 , n44090 );
buf ( n44092 , n41769 );
buf ( n44093 , n41951 );
nand ( n44094 , n44092 , n44093 );
buf ( n44095 , n44094 );
buf ( n44096 , n44095 );
nand ( n44097 , n44091 , n44096 );
buf ( n44098 , n44097 );
buf ( n44099 , n44098 );
not ( n44100 , n44099 );
buf ( n44101 , n37400 );
not ( n44102 , n44101 );
or ( n44103 , n44100 , n44102 );
buf ( n44104 , n42123 );
buf ( n44105 , n37413 );
nand ( n44106 , n44104 , n44105 );
buf ( n44107 , n44106 );
buf ( n44108 , n44107 );
nand ( n44109 , n44103 , n44108 );
buf ( n44110 , n44109 );
buf ( n44111 , n44110 );
and ( n44112 , n44086 , n44111 );
and ( n44113 , n44068 , n44085 );
or ( n44114 , n44112 , n44113 );
buf ( n44115 , n44114 );
nand ( n44116 , n44022 , n44115 );
nand ( n44117 , n44021 , n43988 );
nand ( n44118 , n44116 , n44117 );
xor ( n44119 , n43954 , n44118 );
not ( n44120 , n44119 );
not ( n44121 , n43063 );
not ( n44122 , n41718 );
or ( n44123 , n44121 , n44122 );
buf ( n44124 , n36527 );
not ( n44125 , n43056 );
buf ( n44126 , n44125 );
nand ( n44127 , n44124 , n44126 );
buf ( n44128 , n44127 );
nand ( n44129 , n44123 , n44128 );
buf ( n44130 , n44129 );
not ( n44131 , n44130 );
buf ( n44132 , n36516 );
buf ( n44133 , n36497 );
and ( n44134 , n44132 , n44133 );
buf ( n44135 , n44134 );
buf ( n44136 , n44135 );
not ( n44137 , n44136 );
or ( n44138 , n44131 , n44137 );
buf ( n44139 , n36640 );
not ( n44140 , n44139 );
buf ( n44141 , n44140 );
buf ( n44142 , n44141 );
buf ( n44143 , n43972 );
nand ( n44144 , n44142 , n44143 );
buf ( n44145 , n44144 );
buf ( n44146 , n44145 );
nand ( n44147 , n44138 , n44146 );
buf ( n44148 , n44147 );
buf ( n44149 , n44148 );
not ( n44150 , n42566 );
not ( n44151 , n42805 );
or ( n44152 , n44150 , n44151 );
buf ( n44153 , n25160 );
not ( n44154 , n44153 );
buf ( n44155 , n37586 );
not ( n44156 , n44155 );
buf ( n44157 , n44156 );
buf ( n44158 , n44157 );
not ( n44159 , n44158 );
or ( n44160 , n44154 , n44159 );
buf ( n44161 , n37595 );
not ( n44162 , n44161 );
buf ( n44163 , n44162 );
buf ( n44164 , n44163 );
buf ( n44165 , n42581 );
nand ( n44166 , n44164 , n44165 );
buf ( n44167 , n44166 );
buf ( n44168 , n44167 );
nand ( n44169 , n44160 , n44168 );
buf ( n44170 , n44169 );
nand ( n44171 , n44170 , n42631 );
nand ( n44172 , n44152 , n44171 );
buf ( n44173 , n44172 );
xor ( n44174 , n44149 , n44173 );
not ( n44175 , n37397 );
not ( n44176 , n43442 );
buf ( n44177 , n42195 );
not ( n44178 , n44177 );
buf ( n44179 , n44178 );
not ( n44180 , n44179 );
or ( n44181 , n44176 , n44180 );
nand ( n44182 , n41779 , n42196 );
nand ( n44183 , n44181 , n44182 );
not ( n44184 , n44183 );
or ( n44185 , n44175 , n44184 );
buf ( n44186 , n44098 );
buf ( n44187 , n37413 );
nand ( n44188 , n44186 , n44187 );
buf ( n44189 , n44188 );
nand ( n44190 , n44185 , n44189 );
not ( n44191 , n42448 );
buf ( n44192 , n42468 );
not ( n44193 , n44192 );
buf ( n44194 , n42437 );
not ( n44195 , n44194 );
or ( n44196 , n44193 , n44195 );
buf ( n44197 , n29270 );
buf ( n44198 , n38994 );
nand ( n44199 , n44197 , n44198 );
buf ( n44200 , n44199 );
buf ( n44201 , n44200 );
nand ( n44202 , n44196 , n44201 );
buf ( n44203 , n44202 );
not ( n44204 , n44203 );
or ( n44205 , n44191 , n44204 );
buf ( n44206 , n42468 );
not ( n44207 , n44206 );
buf ( n44208 , n29287 );
not ( n44209 , n44208 );
buf ( n44210 , n44209 );
buf ( n44211 , n44210 );
not ( n44212 , n44211 );
or ( n44213 , n44207 , n44212 );
buf ( n44214 , n39653 );
buf ( n44215 , n42471 );
nand ( n44216 , n44214 , n44215 );
buf ( n44217 , n44216 );
buf ( n44218 , n44217 );
nand ( n44219 , n44213 , n44218 );
buf ( n44220 , n44219 );
not ( n44221 , n38982 );
nand ( n44222 , n44220 , n44221 );
nand ( n44223 , n44205 , n44222 );
xor ( n44224 , n44190 , n44223 );
buf ( n44225 , n42152 );
not ( n44226 , n44225 );
buf ( n44227 , n37472 );
not ( n44228 , n44227 );
or ( n44229 , n44226 , n44228 );
buf ( n44230 , n41843 );
buf ( n44231 , n42160 );
nand ( n44232 , n44230 , n44231 );
buf ( n44233 , n44232 );
buf ( n44234 , n44233 );
nand ( n44235 , n44229 , n44234 );
buf ( n44236 , n44235 );
not ( n44237 , n44236 );
not ( n44238 , n41966 );
or ( n44239 , n44237 , n44238 );
buf ( n44240 , n41876 );
not ( n44241 , n44240 );
buf ( n44242 , n41977 );
not ( n44243 , n44242 );
or ( n44244 , n44241 , n44243 );
buf ( n44245 , n41981 );
buf ( n44246 , n41879 );
nand ( n44247 , n44245 , n44246 );
buf ( n44248 , n44247 );
buf ( n44249 , n44248 );
nand ( n44250 , n44244 , n44249 );
buf ( n44251 , n44250 );
buf ( n44252 , n44251 );
buf ( n44253 , n37440 );
buf ( n44254 , n44253 );
nand ( n44255 , n44252 , n44254 );
buf ( n44256 , n44255 );
nand ( n44257 , n44239 , n44256 );
and ( n44258 , n44224 , n44257 );
and ( n44259 , n44190 , n44223 );
or ( n44260 , n44258 , n44259 );
buf ( n44261 , n44260 );
and ( n44262 , n44174 , n44261 );
and ( n44263 , n44149 , n44173 );
or ( n44264 , n44262 , n44263 );
buf ( n44265 , n44264 );
not ( n44266 , n44265 );
not ( n44267 , n41599 );
buf ( n44268 , n44267 );
not ( n44269 , n44268 );
buf ( n44270 , n41608 );
not ( n44271 , n44270 );
buf ( n44272 , n42277 );
not ( n44273 , n44272 );
or ( n44274 , n44271 , n44273 );
buf ( n44275 , n36562 );
buf ( n44276 , n41611 );
nand ( n44277 , n44275 , n44276 );
buf ( n44278 , n44277 );
buf ( n44279 , n44278 );
nand ( n44280 , n44274 , n44279 );
buf ( n44281 , n44280 );
buf ( n44282 , n44281 );
not ( n44283 , n44282 );
or ( n44284 , n44269 , n44283 );
buf ( n44285 , n43841 );
not ( n44286 , n44285 );
buf ( n44287 , n43868 );
nand ( n44288 , n44286 , n44287 );
buf ( n44289 , n44288 );
buf ( n44290 , n44289 );
nand ( n44291 , n44284 , n44290 );
buf ( n44292 , n44291 );
not ( n44293 , n44292 );
nand ( n44294 , n44266 , n44293 );
not ( n44295 , n44294 );
buf ( n44296 , n25184 );
not ( n44297 , n44296 );
buf ( n44298 , n37686 );
not ( n44299 , n44298 );
buf ( n44300 , n44299 );
buf ( n44301 , n44300 );
not ( n44302 , n44301 );
or ( n44303 , n44297 , n44302 );
buf ( n44304 , n37686 );
buf ( n44305 , n25183 );
nand ( n44306 , n44304 , n44305 );
buf ( n44307 , n44306 );
buf ( n44308 , n44307 );
nand ( n44309 , n44303 , n44308 );
buf ( n44310 , n44309 );
and ( n44311 , n44310 , n43909 );
buf ( n44312 , n25184 );
not ( n44313 , n44312 );
buf ( n44314 , n43198 );
not ( n44315 , n44314 );
buf ( n44316 , n44315 );
buf ( n44317 , n44316 );
not ( n44318 , n44317 );
or ( n44319 , n44313 , n44318 );
buf ( n44320 , n43198 );
buf ( n44321 , n25183 );
nand ( n44322 , n44320 , n44321 );
buf ( n44323 , n44322 );
buf ( n44324 , n44323 );
nand ( n44325 , n44319 , n44324 );
buf ( n44326 , n44325 );
not ( n44327 , n44326 );
nor ( n44328 , n44327 , n43941 );
nor ( n44329 , n44311 , n44328 );
buf ( n44330 , n44329 );
not ( n44331 , n44330 );
buf ( n44332 , n44331 );
not ( n44333 , n44332 );
buf ( n44334 , n44251 );
not ( n44335 , n44334 );
buf ( n44336 , n37511 );
not ( n44337 , n44336 );
buf ( n44338 , n44337 );
buf ( n44339 , n44338 );
not ( n44340 , n44339 );
or ( n44341 , n44335 , n44340 );
buf ( n44342 , n42202 );
buf ( n44343 , n41852 );
nand ( n44344 , n44342 , n44343 );
buf ( n44345 , n44344 );
buf ( n44346 , n44345 );
nand ( n44347 , n44341 , n44346 );
buf ( n44348 , n44347 );
buf ( n44349 , n44348 );
or ( n44350 , n30187 , n38994 );
nand ( n44351 , n44350 , n42489 );
not ( n44352 , n44351 );
not ( n44353 , n42448 );
or ( n44354 , n44352 , n44353 );
buf ( n44355 , n44203 );
buf ( n44356 , n44221 );
nand ( n44357 , n44355 , n44356 );
buf ( n44358 , n44357 );
nand ( n44359 , n44354 , n44358 );
not ( n44360 , n44359 );
buf ( n44361 , n44360 );
and ( n44362 , n44349 , n44361 );
not ( n44363 , n44349 );
buf ( n44364 , n42448 );
not ( n44365 , n44364 );
buf ( n44366 , n42492 );
not ( n44367 , n44366 );
or ( n44368 , n44365 , n44367 );
buf ( n44369 , n44358 );
nand ( n44370 , n44368 , n44369 );
buf ( n44371 , n44370 );
buf ( n44372 , n44371 );
and ( n44373 , n44363 , n44372 );
or ( n44374 , n44362 , n44373 );
buf ( n44375 , n44374 );
buf ( n44376 , n44375 );
buf ( n44377 , n43368 );
not ( n44378 , n44377 );
buf ( n44379 , n41889 );
not ( n44380 , n44379 );
buf ( n44381 , n44380 );
buf ( n44382 , n44381 );
not ( n44383 , n44382 );
or ( n44384 , n44378 , n44383 );
buf ( n44385 , n41947 );
buf ( n44386 , n43365 );
nand ( n44387 , n44385 , n44386 );
buf ( n44388 , n44387 );
buf ( n44389 , n44388 );
nand ( n44390 , n44384 , n44389 );
buf ( n44391 , n44390 );
buf ( n44392 , n44391 );
not ( n44393 , n44392 );
buf ( n44394 , n37872 );
not ( n44395 , n44394 );
or ( n44396 , n44393 , n44395 );
buf ( n44397 , n42167 );
buf ( n44398 , n42175 );
nand ( n44399 , n44397 , n44398 );
buf ( n44400 , n44399 );
buf ( n44401 , n44400 );
nand ( n44402 , n44396 , n44401 );
buf ( n44403 , n44402 );
buf ( n44404 , n44403 );
not ( n44405 , n44404 );
buf ( n44406 , n44405 );
buf ( n44407 , n44406 );
and ( n44408 , n44376 , n44407 );
not ( n44409 , n44376 );
buf ( n44410 , n44403 );
and ( n44411 , n44409 , n44410 );
nor ( n44412 , n44408 , n44411 );
buf ( n44413 , n44412 );
buf ( n44414 , n44413 );
not ( n44415 , n44414 );
buf ( n44416 , n44415 );
not ( n44417 , n44416 );
or ( n44418 , n44333 , n44417 );
buf ( n44419 , n44329 );
not ( n44420 , n44419 );
buf ( n44421 , n44413 );
not ( n44422 , n44421 );
or ( n44423 , n44420 , n44422 );
buf ( n44424 , n44067 );
not ( n44425 , n44424 );
buf ( n44426 , n44425 );
buf ( n44427 , n44426 );
buf ( n44428 , n43996 );
not ( n44429 , n44428 );
buf ( n44430 , n41890 );
not ( n44431 , n44430 );
or ( n44432 , n44429 , n44431 );
buf ( n44433 , n44381 );
not ( n44434 , n44433 );
buf ( n44435 , n44434 );
buf ( n44436 , n44435 );
buf ( n44437 , n42075 );
nand ( n44438 , n44436 , n44437 );
buf ( n44439 , n44438 );
buf ( n44440 , n44439 );
nand ( n44441 , n44432 , n44440 );
buf ( n44442 , n44441 );
buf ( n44443 , n44442 );
not ( n44444 , n44443 );
buf ( n44445 , n37872 );
not ( n44446 , n44445 );
or ( n44447 , n44444 , n44446 );
buf ( n44448 , n37919 );
buf ( n44449 , n44391 );
nand ( n44450 , n44448 , n44449 );
buf ( n44451 , n44450 );
buf ( n44452 , n44451 );
nand ( n44453 , n44447 , n44452 );
buf ( n44454 , n44453 );
buf ( n44455 , n44454 );
xor ( n44456 , n44427 , n44455 );
and ( n44457 , n41993 , n39493 );
not ( n44458 , n41993 );
and ( n44459 , n44458 , n33077 );
or ( n44460 , n44457 , n44459 );
buf ( n44461 , n44460 );
not ( n44462 , n44461 );
buf ( n44463 , n43250 );
not ( n44464 , n44463 );
or ( n44465 , n44462 , n44464 );
buf ( n44466 , n42530 );
buf ( n44467 , n42825 );
nand ( n44468 , n44466 , n44467 );
buf ( n44469 , n44468 );
buf ( n44470 , n44469 );
nand ( n44471 , n44465 , n44470 );
buf ( n44472 , n44471 );
buf ( n44473 , n44472 );
and ( n44474 , n44456 , n44473 );
and ( n44475 , n44427 , n44455 );
or ( n44476 , n44474 , n44475 );
buf ( n44477 , n44476 );
buf ( n44478 , n44477 );
nand ( n44479 , n44423 , n44478 );
buf ( n44480 , n44479 );
nand ( n44481 , n44418 , n44480 );
not ( n44482 , n44481 );
or ( n44483 , n44295 , n44482 );
nand ( n44484 , n44292 , n44265 );
nand ( n44485 , n44483 , n44484 );
not ( n44486 , n44485 );
or ( n44487 , n44120 , n44486 );
or ( n44488 , n44485 , n44119 );
buf ( n44489 , n24811 );
not ( n44490 , n44489 );
buf ( n44491 , n44490 );
buf ( n44492 , n44491 );
not ( n44493 , n44492 );
buf ( n44494 , n44493 );
xnor ( n44495 , n44494 , n24833 );
not ( n44496 , n44495 );
not ( n44497 , n44496 );
buf ( n44498 , n44497 );
not ( n44499 , n44498 );
not ( n44500 , n24835 );
buf ( n44501 , n25382 );
not ( n44502 , n44501 );
buf ( n44503 , n44502 );
not ( n44504 , n44503 );
or ( n44505 , n44500 , n44504 );
not ( n44506 , n24834 );
not ( n44507 , n25368 );
not ( n44508 , n25375 );
or ( n44509 , n44507 , n44508 );
nand ( n44510 , n44509 , n25378 );
not ( n44511 , n44510 );
not ( n44512 , n44511 );
or ( n44513 , n44506 , n44512 );
nand ( n44514 , n44513 , n44495 );
not ( n44515 , n44514 );
nand ( n44516 , n44505 , n44515 );
not ( n44517 , n44516 );
not ( n44518 , n44517 );
buf ( n44519 , n44518 );
not ( n44520 , n44519 );
or ( n44521 , n44499 , n44520 );
buf ( n44522 , n44503 );
buf ( n44523 , n44522 );
buf ( n44524 , n44523 );
buf ( n44525 , n44524 );
not ( n44526 , n44525 );
buf ( n44527 , n44526 );
buf ( n44528 , n44527 );
buf ( n44529 , n44528 );
buf ( n44530 , n44529 );
buf ( n44531 , n44530 );
not ( n44532 , n44531 );
buf ( n44533 , n44532 );
buf ( n44534 , n44533 );
not ( n44535 , n44534 );
buf ( n44536 , n35969 );
buf ( n44537 , n44536 );
buf ( n44538 , n44537 );
buf ( n44539 , n44538 );
not ( n44540 , n44539 );
or ( n44541 , n44535 , n44540 );
buf ( n44542 , n39005 );
buf ( n44543 , n44530 );
nand ( n44544 , n44542 , n44543 );
buf ( n44545 , n44544 );
buf ( n44546 , n44545 );
nand ( n44547 , n44541 , n44546 );
buf ( n44548 , n44547 );
buf ( n44549 , n44548 );
nand ( n44550 , n44521 , n44549 );
buf ( n44551 , n44550 );
buf ( n44552 , n44551 );
xor ( n44553 , n43245 , n43279 );
xor ( n44554 , n44553 , n43289 );
buf ( n44555 , n44554 );
buf ( n44556 , n44555 );
xor ( n44557 , n44552 , n44556 );
xor ( n44558 , n43333 , n43358 );
xor ( n44559 , n44558 , n43421 );
buf ( n44560 , n44559 );
buf ( n44561 , n44560 );
xor ( n44562 , n44557 , n44561 );
buf ( n44563 , n44562 );
nand ( n44564 , n44488 , n44563 );
nand ( n44565 , n44487 , n44564 );
buf ( n44566 , n44565 );
not ( n44567 , n43946 );
buf ( n44568 , n43872 );
not ( n44569 , n44568 );
buf ( n44570 , n44569 );
not ( n44571 , n44570 );
or ( n44572 , n44567 , n44571 );
not ( n44573 , n43872 );
not ( n44574 , n43943 );
or ( n44575 , n44573 , n44574 );
nand ( n44576 , n44575 , n44118 );
nand ( n44577 , n44572 , n44576 );
xor ( n44578 , n44552 , n44556 );
and ( n44579 , n44578 , n44561 );
and ( n44580 , n44552 , n44556 );
or ( n44581 , n44579 , n44580 );
buf ( n44582 , n44581 );
xor ( n44583 , n44577 , n44582 );
buf ( n44584 , n43941 );
not ( n44585 , n44584 );
buf ( n44586 , n44585 );
buf ( n44587 , n44586 );
not ( n44588 , n44587 );
buf ( n44589 , n43892 );
not ( n44590 , n44589 );
or ( n44591 , n44588 , n44590 );
buf ( n44592 , n43031 );
not ( n44593 , n44592 );
buf ( n44594 , n25184 );
not ( n44595 , n44594 );
or ( n44596 , n44593 , n44595 );
buf ( n44597 , n38244 );
buf ( n44598 , n25183 );
nand ( n44599 , n44597 , n44598 );
buf ( n44600 , n44599 );
buf ( n44601 , n44600 );
nand ( n44602 , n44596 , n44601 );
buf ( n44603 , n44602 );
buf ( n44604 , n44603 );
buf ( n44605 , n43909 );
nand ( n44606 , n44604 , n44605 );
buf ( n44607 , n44606 );
buf ( n44608 , n44607 );
nand ( n44609 , n44591 , n44608 );
buf ( n44610 , n44609 );
buf ( n44611 , n44610 );
buf ( n44612 , n44267 );
not ( n44613 , n44612 );
buf ( n44614 , n43864 );
not ( n44615 , n44614 );
or ( n44616 , n44613 , n44615 );
buf ( n44617 , n41626 );
buf ( n44618 , n43868 );
nand ( n44619 , n44617 , n44618 );
buf ( n44620 , n44619 );
buf ( n44621 , n44620 );
nand ( n44622 , n44616 , n44621 );
buf ( n44623 , n44622 );
buf ( n44624 , n44623 );
xor ( n44625 , n44611 , n44624 );
buf ( n44626 , n43410 );
not ( n44627 , n44626 );
buf ( n44628 , n38130 );
not ( n44629 , n44628 );
or ( n44630 , n44627 , n44629 );
buf ( n44631 , n41882 );
not ( n44632 , n44631 );
buf ( n44633 , n38108 );
not ( n44634 , n44633 );
buf ( n44635 , n44634 );
buf ( n44636 , n44635 );
not ( n44637 , n44636 );
or ( n44638 , n44632 , n44637 );
buf ( n44639 , n38108 );
buf ( n44640 , n41879 );
nand ( n44641 , n44639 , n44640 );
buf ( n44642 , n44641 );
buf ( n44643 , n44642 );
nand ( n44644 , n44638 , n44643 );
buf ( n44645 , n44644 );
buf ( n44646 , n44645 );
buf ( n44647 , n43414 );
nand ( n44648 , n44646 , n44647 );
buf ( n44649 , n44648 );
buf ( n44650 , n44649 );
nand ( n44651 , n44630 , n44650 );
buf ( n44652 , n44651 );
buf ( n44653 , n44652 );
buf ( n44654 , n42448 );
not ( n44655 , n44654 );
buf ( n44656 , n43706 );
not ( n44657 , n44656 );
or ( n44658 , n44655 , n44657 );
buf ( n44659 , n43347 );
buf ( n44660 , n38985 );
nand ( n44661 , n44659 , n44660 );
buf ( n44662 , n44661 );
buf ( n44663 , n44662 );
nand ( n44664 , n44658 , n44663 );
buf ( n44665 , n44664 );
buf ( n44666 , n44665 );
xor ( n44667 , n44653 , n44666 );
buf ( n44668 , n42045 );
buf ( n44669 , n44668 );
buf ( n44670 , n44669 );
buf ( n44671 , n44670 );
buf ( n44672 , n42086 );
or ( n44673 , n44671 , n44672 );
buf ( n44674 , n36906 );
not ( n44675 , n44674 );
buf ( n44676 , n44675 );
buf ( n44677 , n44676 );
buf ( n44678 , n44677 );
buf ( n44679 , n44678 );
buf ( n44680 , n44679 );
not ( n44681 , n44680 );
buf ( n44682 , n44681 );
buf ( n44683 , n44682 );
buf ( n44684 , n42062 );
buf ( n44685 , n43365 );
and ( n44686 , n44684 , n44685 );
buf ( n44687 , n43095 );
not ( n44688 , n44687 );
buf ( n44689 , n44688 );
buf ( n44690 , n44689 );
buf ( n44691 , n43368 );
and ( n44692 , n44690 , n44691 );
nor ( n44693 , n44686 , n44692 );
buf ( n44694 , n44693 );
buf ( n44695 , n44694 );
or ( n44696 , n44683 , n44695 );
nand ( n44697 , n44673 , n44696 );
buf ( n44698 , n44697 );
buf ( n44699 , n44698 );
xor ( n44700 , n44667 , n44699 );
buf ( n44701 , n44700 );
buf ( n44702 , n44701 );
xor ( n44703 , n44625 , n44702 );
buf ( n44704 , n44703 );
xor ( n44705 , n44583 , n44704 );
buf ( n44706 , n44705 );
xor ( n44707 , n44566 , n44706 );
not ( n44708 , n44518 );
buf ( n44709 , n44708 );
not ( n44710 , n44709 );
buf ( n44711 , n44533 );
not ( n44712 , n44711 );
buf ( n44713 , n36054 );
not ( n44714 , n44713 );
or ( n44715 , n44712 , n44714 );
buf ( n44716 , n36054 );
not ( n44717 , n44716 );
buf ( n44718 , n44717 );
buf ( n44719 , n44718 );
buf ( n44720 , n44530 );
nand ( n44721 , n44719 , n44720 );
buf ( n44722 , n44721 );
buf ( n44723 , n44722 );
nand ( n44724 , n44715 , n44723 );
buf ( n44725 , n44724 );
buf ( n44726 , n44725 );
not ( n44727 , n44726 );
or ( n44728 , n44710 , n44727 );
buf ( n44729 , n44548 );
buf ( n44730 , n44496 );
nand ( n44731 , n44729 , n44730 );
buf ( n44732 , n44731 );
buf ( n44733 , n44732 );
nand ( n44734 , n44728 , n44733 );
buf ( n44735 , n44734 );
buf ( n44736 , n42055 );
not ( n44737 , n44736 );
buf ( n44738 , n43371 );
not ( n44739 , n44738 );
or ( n44740 , n44737 , n44739 );
buf ( n44741 , n43403 );
buf ( n44742 , n42052 );
nand ( n44743 , n44741 , n44742 );
buf ( n44744 , n44743 );
buf ( n44745 , n44744 );
nand ( n44746 , n44740 , n44745 );
buf ( n44747 , n44746 );
buf ( n44748 , n44747 );
not ( n44749 , n44748 );
buf ( n44750 , n38130 );
not ( n44751 , n44750 );
or ( n44752 , n44749 , n44751 );
buf ( n44753 , n43414 );
buf ( n44754 , n44011 );
nand ( n44755 , n44753 , n44754 );
buf ( n44756 , n44755 );
buf ( n44757 , n44756 );
nand ( n44758 , n44752 , n44757 );
buf ( n44759 , n44758 );
buf ( n44760 , n44759 );
buf ( n44761 , n41748 );
buf ( n44762 , n36929 );
and ( n44763 , n44761 , n44762 );
not ( n44764 , n44761 );
buf ( n44765 , n42082 );
and ( n44766 , n44764 , n44765 );
nor ( n44767 , n44763 , n44766 );
buf ( n44768 , n44767 );
buf ( n44769 , n44768 );
not ( n44770 , n44769 );
buf ( n44771 , n44770 );
buf ( n44772 , n44771 );
not ( n44773 , n44772 );
buf ( n44774 , n42045 );
not ( n44775 , n44774 );
buf ( n44776 , n44775 );
buf ( n44777 , n44776 );
not ( n44778 , n44777 );
or ( n44779 , n44773 , n44778 );
buf ( n44780 , n43112 );
not ( n44781 , n44780 );
buf ( n44782 , n36912 );
nand ( n44783 , n44781 , n44782 );
buf ( n44784 , n44783 );
buf ( n44785 , n44784 );
nand ( n44786 , n44779 , n44785 );
buf ( n44787 , n44786 );
buf ( n44788 , n44787 );
xor ( n44789 , n44760 , n44788 );
xor ( n44790 , n44068 , n44085 );
xor ( n44791 , n44790 , n44111 );
buf ( n44792 , n44791 );
buf ( n44793 , n44792 );
and ( n44794 , n44789 , n44793 );
and ( n44795 , n44760 , n44788 );
or ( n44796 , n44794 , n44795 );
buf ( n44797 , n44796 );
xor ( n44798 , n44735 , n44797 );
buf ( n44799 , n42712 );
not ( n44800 , n44799 );
buf ( n44801 , n42672 );
not ( n44802 , n44801 );
buf ( n44803 , n38435 );
not ( n44804 , n44803 );
or ( n44805 , n44802 , n44804 );
buf ( n44806 , n37146 );
buf ( n44807 , n42679 );
nand ( n44808 , n44806 , n44807 );
buf ( n44809 , n44808 );
buf ( n44810 , n44809 );
nand ( n44811 , n44805 , n44810 );
buf ( n44812 , n44811 );
buf ( n44813 , n44812 );
not ( n44814 , n44813 );
or ( n44815 , n44800 , n44814 );
buf ( n44816 , n42772 );
buf ( n44817 , n42668 );
nand ( n44818 , n44816 , n44817 );
buf ( n44819 , n44818 );
buf ( n44820 , n44819 );
nand ( n44821 , n44815 , n44820 );
buf ( n44822 , n44821 );
and ( n44823 , n44798 , n44822 );
and ( n44824 , n44735 , n44797 );
or ( n44825 , n44823 , n44824 );
buf ( n44826 , n44825 );
xor ( n44827 , n42090 , n42108 );
xnor ( n44828 , n44827 , n42220 );
buf ( n44829 , n44828 );
buf ( n44830 , n44829 );
buf ( n44831 , n44830 );
buf ( n44832 , n44831 );
not ( n44833 , n44832 );
not ( n44834 , n42339 );
not ( n44835 , n42364 );
or ( n44836 , n44834 , n44835 );
nand ( n44837 , n42930 , n42374 );
nand ( n44838 , n44836 , n44837 );
not ( n44839 , n44838 );
buf ( n44840 , n43909 );
not ( n44841 , n44840 );
buf ( n44842 , n43922 );
not ( n44843 , n44842 );
or ( n44844 , n44841 , n44843 );
buf ( n44845 , n44310 );
buf ( n44846 , n44586 );
nand ( n44847 , n44845 , n44846 );
buf ( n44848 , n44847 );
buf ( n44849 , n44848 );
nand ( n44850 , n44844 , n44849 );
buf ( n44851 , n44850 );
buf ( n44852 , n44851 );
not ( n44853 , n44852 );
buf ( n44854 , n44853 );
buf ( n44855 , n44854 );
buf ( n44856 , n44403 );
not ( n44857 , n44856 );
buf ( n44858 , n44348 );
not ( n44859 , n44858 );
buf ( n44860 , n44360 );
nand ( n44861 , n44859 , n44860 );
buf ( n44862 , n44861 );
buf ( n44863 , n44862 );
not ( n44864 , n44863 );
or ( n44865 , n44857 , n44864 );
buf ( n44866 , n44371 );
buf ( n44867 , n44348 );
nand ( n44868 , n44866 , n44867 );
buf ( n44869 , n44868 );
buf ( n44870 , n44869 );
nand ( n44871 , n44865 , n44870 );
buf ( n44872 , n44871 );
buf ( n44873 , n44872 );
not ( n44874 , n44873 );
buf ( n44875 , n44874 );
buf ( n44876 , n44875 );
nand ( n44877 , n44855 , n44876 );
buf ( n44878 , n44877 );
buf ( n44879 , n44878 );
xor ( n44880 , n42142 , n42183 );
xor ( n44881 , n44880 , n42216 );
buf ( n44882 , n44881 );
buf ( n44883 , n44882 );
and ( n44884 , n44879 , n44883 );
and ( n44885 , n44851 , n44872 );
buf ( n44886 , n44885 );
nor ( n44887 , n44884 , n44886 );
buf ( n44888 , n44887 );
not ( n44889 , n44888 );
or ( n44890 , n44839 , n44889 );
or ( n44891 , n44888 , n44838 );
nand ( n44892 , n44890 , n44891 );
buf ( n44893 , n44892 );
not ( n44894 , n44893 );
or ( n44895 , n44833 , n44894 );
buf ( n44896 , n44892 );
buf ( n44897 , n44831 );
or ( n44898 , n44896 , n44897 );
nand ( n44899 , n44895 , n44898 );
buf ( n44900 , n44899 );
buf ( n44901 , n44900 );
xor ( n44902 , n44826 , n44901 );
buf ( n44903 , n44115 );
not ( n44904 , n44903 );
buf ( n44905 , n44904 );
and ( n44906 , n44021 , n44905 );
not ( n44907 , n44021 );
and ( n44908 , n44907 , n44115 );
or ( n44909 , n44906 , n44908 );
buf ( n44910 , n44909 );
buf ( n44911 , n43988 );
and ( n44912 , n44910 , n44911 );
not ( n44913 , n44910 );
buf ( n44914 , n43988 );
not ( n44915 , n44914 );
buf ( n44916 , n44915 );
buf ( n44917 , n44916 );
and ( n44918 , n44913 , n44917 );
nor ( n44919 , n44912 , n44918 );
buf ( n44920 , n44919 );
buf ( n44921 , n44920 );
buf ( n44922 , n42315 );
not ( n44923 , n44922 );
buf ( n44924 , n42739 );
not ( n44925 , n44924 );
or ( n44926 , n44923 , n44925 );
buf ( n44927 , n42266 );
buf ( n44928 , n36396 );
and ( n44929 , n44927 , n44928 );
not ( n44930 , n44927 );
buf ( n44931 , n43597 );
and ( n44932 , n44930 , n44931 );
nor ( n44933 , n44929 , n44932 );
buf ( n44934 , n44933 );
buf ( n44935 , n44934 );
buf ( n44936 , n42252 );
nand ( n44937 , n44935 , n44936 );
buf ( n44938 , n44937 );
buf ( n44939 , n44938 );
nand ( n44940 , n44926 , n44939 );
buf ( n44941 , n44940 );
buf ( n44942 , n44941 );
xor ( n44943 , n44921 , n44942 );
buf ( n44944 , n25997 );
not ( n44945 , n44944 );
buf ( n44946 , n44945 );
buf ( n44947 , n44946 );
buf ( n44948 , n44947 );
buf ( n44949 , n44948 );
buf ( n44950 , n44949 );
not ( n44951 , n44950 );
buf ( n44952 , n44951 );
buf ( n44953 , n44952 );
not ( n44954 , n44953 );
buf ( n44955 , n37649 );
not ( n44956 , n44955 );
or ( n44957 , n44954 , n44956 );
buf ( n44958 , n36360 );
buf ( n44959 , n44952 );
not ( n44960 , n44959 );
buf ( n44961 , n44960 );
buf ( n44962 , n44961 );
nand ( n44963 , n44958 , n44962 );
buf ( n44964 , n44963 );
buf ( n44965 , n44964 );
nand ( n44966 , n44957 , n44965 );
buf ( n44967 , n44966 );
buf ( n44968 , n43053 );
buf ( n44969 , n42851 );
nand ( n44970 , n44968 , n44969 );
buf ( n44971 , n44970 );
buf ( n44972 , n44971 );
nand ( n44973 , C1 , n44972 );
buf ( n44974 , n44973 );
buf ( n44975 , n44974 );
buf ( n44976 , n39986 );
not ( n44977 , n44976 );
buf ( n44978 , n42907 );
not ( n44979 , n44978 );
or ( n44980 , n44977 , n44979 );
buf ( n44981 , n24092 );
not ( n44982 , n44981 );
not ( n44983 , n30187 );
buf ( n44984 , n44983 );
not ( n44985 , n44984 );
or ( n44986 , n44982 , n44985 );
buf ( n44987 , n30187 );
not ( n44988 , n44987 );
buf ( n44989 , n44988 );
buf ( n44990 , n44989 );
not ( n44991 , n44990 );
buf ( n44992 , n44991 );
buf ( n44993 , n44992 );
buf ( n44994 , n40009 );
nand ( n44995 , n44993 , n44994 );
buf ( n44996 , n44995 );
buf ( n44997 , n44996 );
nand ( n44998 , n44986 , n44997 );
buf ( n44999 , n44998 );
buf ( n45000 , n44999 );
buf ( n45001 , n40002 );
nand ( n45002 , n45000 , n45001 );
buf ( n45003 , n45002 );
buf ( n45004 , n45003 );
nand ( n45005 , n44980 , n45004 );
buf ( n45006 , n45005 );
buf ( n45007 , n45006 );
or ( n45008 , n44975 , n45007 );
buf ( n45009 , n42631 );
not ( n45010 , n45009 );
buf ( n45011 , n25160 );
not ( n45012 , n45011 );
buf ( n45013 , n37642 );
not ( n45014 , n45013 );
or ( n45015 , n45012 , n45014 );
buf ( n45016 , n39205 );
buf ( n45017 , n42581 );
nand ( n45018 , n45016 , n45017 );
buf ( n45019 , n45018 );
buf ( n45020 , n45019 );
nand ( n45021 , n45015 , n45020 );
buf ( n45022 , n45021 );
buf ( n45023 , n45022 );
not ( n45024 , n45023 );
or ( n45025 , n45010 , n45024 );
buf ( n45026 , n44170 );
buf ( n45027 , n42566 );
nand ( n45028 , n45026 , n45027 );
buf ( n45029 , n45028 );
buf ( n45030 , n45029 );
nand ( n45031 , n45025 , n45030 );
buf ( n45032 , n45031 );
buf ( n45033 , n45032 );
nand ( n45034 , n45008 , n45033 );
buf ( n45035 , n45034 );
buf ( n45036 , n45035 );
buf ( n45037 , n45006 );
buf ( n45038 , n44974 );
nand ( n45039 , n45037 , n45038 );
buf ( n45040 , n45039 );
buf ( n45041 , n45040 );
nand ( n45042 , n45036 , n45041 );
buf ( n45043 , n45042 );
buf ( n45044 , n45043 );
xor ( n45045 , n42841 , n42883 );
xor ( n45046 , n45045 , n42915 );
buf ( n45047 , n45046 );
buf ( n45048 , n45047 );
xor ( n45049 , n45044 , n45048 );
not ( n45050 , n42448 );
not ( n45051 , n44220 );
or ( n45052 , n45050 , n45051 );
nand ( n45053 , n38972 , n38980 , n38981 );
buf ( n45054 , n45053 );
buf ( n45055 , n45054 );
buf ( n45056 , n45055 );
buf ( n45057 , n45056 );
not ( n45058 , n45057 );
buf ( n45059 , n45058 );
and ( n45060 , n38994 , n41762 );
not ( n45061 , n38994 );
and ( n45062 , n45061 , n28722 );
or ( n45063 , n45060 , n45062 );
nand ( n45064 , n45059 , n45063 );
nand ( n45065 , n45052 , n45064 );
buf ( n45066 , n45065 );
buf ( n45067 , n42408 );
not ( n45068 , n45067 );
buf ( n45069 , n45068 );
not ( n45070 , n45069 );
not ( n45071 , n41822 );
or ( n45072 , n45070 , n45071 );
buf ( n45073 , n29325 );
buf ( n45074 , n45073 );
buf ( n45075 , n45074 );
nand ( n45076 , n42411 , n45075 );
nand ( n45077 , n45072 , n45076 );
not ( n45078 , n45077 );
not ( n45079 , n38404 );
or ( n45080 , n45078 , n45079 );
buf ( n45081 , n44036 );
buf ( n45082 , n38380 );
nand ( n45083 , n45081 , n45082 );
buf ( n45084 , n45083 );
nand ( n45085 , n45080 , n45084 );
buf ( n45086 , n45085 );
xor ( n45087 , n45066 , n45086 );
buf ( n45088 , n43442 );
not ( n45089 , n45088 );
buf ( n45090 , n41876 );
not ( n45091 , n45090 );
or ( n45092 , n45089 , n45091 );
buf ( n45093 , n41779 );
buf ( n45094 , n41873 );
nand ( n45095 , n45093 , n45094 );
buf ( n45096 , n45095 );
buf ( n45097 , n45096 );
nand ( n45098 , n45092 , n45097 );
buf ( n45099 , n45098 );
buf ( n45100 , n45099 );
not ( n45101 , n45100 );
buf ( n45102 , n37397 );
not ( n45103 , n45102 );
or ( n45104 , n45101 , n45103 );
buf ( n45105 , n44183 );
buf ( n45106 , n37410 );
buf ( n45107 , n45106 );
buf ( n45108 , n45107 );
buf ( n45109 , n45108 );
nand ( n45110 , n45105 , n45109 );
buf ( n45111 , n45110 );
buf ( n45112 , n45111 );
nand ( n45113 , n45104 , n45112 );
buf ( n45114 , n45113 );
buf ( n45115 , n45114 );
and ( n45116 , n45087 , n45115 );
and ( n45117 , n45066 , n45086 );
or ( n45118 , n45116 , n45117 );
buf ( n45119 , n45118 );
buf ( n45120 , n45119 );
buf ( n45121 , n43108 );
not ( n45122 , n45121 );
buf ( n45123 , n44635 );
not ( n45124 , n45123 );
or ( n45125 , n45122 , n45124 );
buf ( n45126 , n43400 );
buf ( n45127 , n43099 );
nand ( n45128 , n45126 , n45127 );
buf ( n45129 , n45128 );
buf ( n45130 , n45129 );
nand ( n45131 , n45125 , n45130 );
buf ( n45132 , n45131 );
buf ( n45133 , n45132 );
not ( n45134 , n45133 );
buf ( n45135 , n43389 );
not ( n45136 , n45135 );
or ( n45137 , n45134 , n45136 );
buf ( n45138 , n44747 );
buf ( n45139 , n38054 );
not ( n45140 , n45139 );
buf ( n45141 , n45140 );
buf ( n45142 , n45141 );
not ( n45143 , n45142 );
buf ( n45144 , n45143 );
buf ( n45145 , n45144 );
nand ( n45146 , n45138 , n45145 );
buf ( n45147 , n45146 );
buf ( n45148 , n45147 );
nand ( n45149 , n45137 , n45148 );
buf ( n45150 , n45149 );
buf ( n45151 , n45150 );
xor ( n45152 , n45120 , n45151 );
buf ( n45153 , n36973 );
not ( n45154 , n45153 );
buf ( n45155 , n45154 );
buf ( n45156 , n45155 );
buf ( n45157 , n45156 );
buf ( n45158 , n45157 );
buf ( n45159 , n45158 );
not ( n45160 , n45159 );
buf ( n45161 , n45160 );
buf ( n45162 , n45161 );
buf ( n45163 , n42504 );
buf ( n45164 , n39139 );
and ( n45165 , n45163 , n45164 );
not ( n45166 , n45163 );
buf ( n45167 , n42062 );
and ( n45168 , n45166 , n45167 );
nor ( n45169 , n45165 , n45168 );
buf ( n45170 , n45169 );
buf ( n45171 , n45170 );
or ( n45172 , n45162 , n45171 );
buf ( n45173 , n44682 );
buf ( n45174 , n44768 );
or ( n45175 , n45173 , n45174 );
nand ( n45176 , n45172 , n45175 );
buf ( n45177 , n45176 );
buf ( n45178 , n45177 );
and ( n45179 , n45152 , n45178 );
and ( n45180 , n45120 , n45151 );
or ( n45181 , n45179 , n45180 );
buf ( n45182 , n45181 );
buf ( n45183 , n45182 );
and ( n45184 , n45049 , n45183 );
and ( n45185 , n45044 , n45048 );
or ( n45186 , n45184 , n45185 );
buf ( n45187 , n45186 );
buf ( n45188 , n45187 );
and ( n45189 , n44943 , n45188 );
and ( n45190 , n44921 , n44942 );
or ( n45191 , n45189 , n45190 );
buf ( n45192 , n45191 );
buf ( n45193 , n45192 );
and ( n45194 , n44902 , n45193 );
and ( n45195 , n44826 , n44901 );
or ( n45196 , n45194 , n45195 );
buf ( n45197 , n45196 );
buf ( n45198 , n45197 );
and ( n45199 , n44707 , n45198 );
and ( n45200 , n44566 , n44706 );
or ( n45201 , n45199 , n45200 );
buf ( n45202 , n45201 );
buf ( n45203 , n45202 );
not ( n45204 , n45203 );
buf ( n45205 , n45204 );
buf ( n45206 , n45205 );
not ( n45207 , n45206 );
xor ( n45208 , n44577 , n44582 );
and ( n45209 , n45208 , n44704 );
and ( n45210 , n44577 , n44582 );
or ( n45211 , n45209 , n45210 );
xor ( n45212 , n44611 , n44624 );
and ( n45213 , n45212 , n44702 );
and ( n45214 , n44611 , n44624 );
or ( n45215 , n45213 , n45214 );
buf ( n45216 , n45215 );
buf ( n45217 , n45216 );
buf ( n45218 , n43909 );
not ( n45219 , n45218 );
buf ( n45220 , n25184 );
not ( n45221 , n45220 );
buf ( n45222 , n39407 );
not ( n45223 , n45222 );
or ( n45224 , n45221 , n45223 );
buf ( n45225 , n38218 );
not ( n45226 , n45225 );
buf ( n45227 , n45226 );
buf ( n45228 , n45227 );
buf ( n45229 , n25183 );
nand ( n45230 , n45228 , n45229 );
buf ( n45231 , n45230 );
buf ( n45232 , n45231 );
nand ( n45233 , n45224 , n45232 );
buf ( n45234 , n45233 );
buf ( n45235 , n45234 );
not ( n45236 , n45235 );
or ( n45237 , n45219 , n45236 );
buf ( n45238 , n44586 );
buf ( n45239 , n44603 );
nand ( n45240 , n45238 , n45239 );
buf ( n45241 , n45240 );
buf ( n45242 , n45241 );
nand ( n45243 , n45237 , n45242 );
buf ( n45244 , n45243 );
buf ( n45245 , n45244 );
buf ( n45246 , n43053 );
buf ( n45247 , n42504 );
not ( n45248 , n45247 );
buf ( n45249 , n37602 );
not ( n45250 , n45249 );
or ( n45251 , n45248 , n45250 );
buf ( n45252 , n36360 );
buf ( n45253 , n41721 );
nand ( n45254 , n45252 , n45253 );
buf ( n45255 , n45254 );
buf ( n45256 , n45255 );
nand ( n45257 , n45251 , n45256 );
buf ( n45258 , n45257 );
buf ( n45259 , n45258 );
nand ( n45260 , n45246 , n45259 );
buf ( n45261 , n45260 );
buf ( n45262 , n45261 );
nand ( n45263 , C1 , n45262 );
buf ( n45264 , n45263 );
buf ( n45265 , n45264 );
buf ( n45266 , n38150 );
not ( n45267 , n45266 );
buf ( n45268 , n41779 );
not ( n45269 , n45268 );
buf ( n45270 , n45269 );
xor ( n45271 , n45270 , n43311 );
buf ( n45272 , n45271 );
not ( n45273 , n45272 );
or ( n45274 , n45267 , n45273 );
buf ( n45275 , n37400 );
buf ( n45276 , n43452 );
nand ( n45277 , n45275 , n45276 );
buf ( n45278 , n45277 );
buf ( n45279 , n45278 );
nand ( n45280 , n45274 , n45279 );
buf ( n45281 , n45280 );
buf ( n45282 , n45281 );
xor ( n45283 , n45265 , n45282 );
buf ( n45284 , n43510 );
not ( n45285 , n45284 );
buf ( n45286 , n36098 );
not ( n45287 , n45286 );
buf ( n45288 , n45287 );
buf ( n45289 , n45288 );
not ( n45290 , n45289 );
or ( n45291 , n45285 , n45290 );
buf ( n45292 , n42530 );
buf ( n45293 , n43996 );
not ( n45294 , n45293 );
buf ( n45295 , n39478 );
not ( n45296 , n45295 );
or ( n45297 , n45294 , n45296 );
buf ( n45298 , n39481 );
buf ( n45299 , n42075 );
nand ( n45300 , n45298 , n45299 );
buf ( n45301 , n45300 );
buf ( n45302 , n45301 );
nand ( n45303 , n45297 , n45302 );
buf ( n45304 , n45303 );
buf ( n45305 , n45304 );
nand ( n45306 , n45292 , n45305 );
buf ( n45307 , n45306 );
buf ( n45308 , n45307 );
nand ( n45309 , n45291 , n45308 );
buf ( n45310 , n45309 );
buf ( n45311 , n45310 );
xor ( n45312 , n45283 , n45311 );
buf ( n45313 , n45312 );
buf ( n45314 , n45313 );
xor ( n45315 , n45245 , n45314 );
xor ( n45316 , n44653 , n44666 );
and ( n45317 , n45316 , n44699 );
and ( n45318 , n44653 , n44666 );
or ( n45319 , n45317 , n45318 );
buf ( n45320 , n45319 );
buf ( n45321 , n45320 );
xor ( n45322 , n45315 , n45321 );
buf ( n45323 , n45322 );
buf ( n45324 , n45323 );
xor ( n45325 , n45217 , n45324 );
buf ( n45326 , n42315 );
not ( n45327 , n45326 );
buf ( n45328 , n42266 );
not ( n45329 , n45328 );
buf ( n45330 , n36054 );
not ( n45331 , n45330 );
or ( n45332 , n45329 , n45331 );
buf ( n45333 , n44718 );
buf ( n45334 , n42263 );
nand ( n45335 , n45333 , n45334 );
buf ( n45336 , n45335 );
buf ( n45337 , n45336 );
nand ( n45338 , n45332 , n45337 );
buf ( n45339 , n45338 );
buf ( n45340 , n45339 );
not ( n45341 , n45340 );
or ( n45342 , n45327 , n45341 );
buf ( n45343 , n42302 );
buf ( n45344 , n42252 );
nand ( n45345 , n45343 , n45344 );
buf ( n45346 , n45345 );
buf ( n45347 , n45346 );
nand ( n45348 , n45342 , n45347 );
buf ( n45349 , n45348 );
buf ( n45350 , n45349 );
not ( n45351 , n42566 );
and ( n45352 , n43142 , n42581 );
not ( n45353 , n43142 );
and ( n45354 , n45353 , n25160 );
or ( n45355 , n45352 , n45354 );
not ( n45356 , n45355 );
or ( n45357 , n45351 , n45356 );
buf ( n45358 , n43232 );
buf ( n45359 , n42631 );
nand ( n45360 , n45358 , n45359 );
buf ( n45361 , n45360 );
nand ( n45362 , n45357 , n45361 );
buf ( n45363 , n45362 );
xor ( n45364 , n45350 , n45363 );
buf ( n45365 , n44645 );
not ( n45366 , n45365 );
buf ( n45367 , n43389 );
not ( n45368 , n45367 );
or ( n45369 , n45366 , n45368 );
not ( n45370 , n42196 );
not ( n45371 , n45370 );
not ( n45372 , n38068 );
or ( n45373 , n45371 , n45372 );
buf ( n45374 , n38068 );
not ( n45375 , n45374 );
buf ( n45376 , n45375 );
buf ( n45377 , n45376 );
buf ( n45378 , n42196 );
nand ( n45379 , n45377 , n45378 );
buf ( n45380 , n45379 );
nand ( n45381 , n45373 , n45380 );
buf ( n45382 , n45381 );
buf ( n45383 , n43414 );
nand ( n45384 , n45382 , n45383 );
buf ( n45385 , n45384 );
buf ( n45386 , n45385 );
nand ( n45387 , n45369 , n45386 );
buf ( n45388 , n45387 );
buf ( n45389 , n45388 );
buf ( n45390 , n38758 );
not ( n45391 , n45390 );
buf ( n45392 , n38413 );
not ( n45393 , n45392 );
not ( n45394 , n37641 );
buf ( n45395 , n45394 );
not ( n45396 , n45395 );
or ( n45397 , n45393 , n45396 );
buf ( n45398 , n39205 );
buf ( n45399 , n38412 );
buf ( n45400 , n45399 );
buf ( n45401 , n45400 );
buf ( n45402 , n45401 );
nand ( n45403 , n45398 , n45402 );
buf ( n45404 , n45403 );
buf ( n45405 , n45404 );
nand ( n45406 , n45397 , n45405 );
buf ( n45407 , n45406 );
buf ( n45408 , n45407 );
not ( n45409 , n45408 );
or ( n45410 , n45391 , n45409 );
buf ( n45411 , n43474 );
not ( n45412 , n45411 );
buf ( n45413 , n38775 );
nand ( n45414 , n45412 , n45413 );
buf ( n45415 , n45414 );
buf ( n45416 , n45415 );
nand ( n45417 , n45410 , n45416 );
buf ( n45418 , n45417 );
buf ( n45419 , n45418 );
xor ( n45420 , n45389 , n45419 );
buf ( n45421 , n42045 );
not ( n45422 , n45421 );
buf ( n45423 , n45422 );
buf ( n45424 , n45423 );
not ( n45425 , n45424 );
buf ( n45426 , n45425 );
buf ( n45427 , n45426 );
buf ( n45428 , n44694 );
or ( n45429 , n45427 , n45428 );
buf ( n45430 , n44682 );
buf ( n45431 , n43095 );
buf ( n45432 , n42160 );
and ( n45433 , n45431 , n45432 );
buf ( n45434 , n44689 );
buf ( n45435 , n42152 );
and ( n45436 , n45434 , n45435 );
nor ( n45437 , n45433 , n45436 );
buf ( n45438 , n45437 );
buf ( n45439 , n45438 );
or ( n45440 , n45430 , n45439 );
nand ( n45441 , n45429 , n45440 );
buf ( n45442 , n45441 );
buf ( n45443 , n45442 );
xor ( n45444 , n45420 , n45443 );
buf ( n45445 , n45444 );
buf ( n45446 , n45445 );
xor ( n45447 , n45364 , n45446 );
buf ( n45448 , n45447 );
buf ( n45449 , n45448 );
xor ( n45450 , n45325 , n45449 );
buf ( n45451 , n45450 );
xor ( n45452 , n45211 , n45451 );
not ( n45453 , n44838 );
not ( n45454 , n45453 );
not ( n45455 , n44828 );
or ( n45456 , n45454 , n45455 );
buf ( n45457 , n44888 );
not ( n45458 , n45457 );
buf ( n45459 , n45458 );
nand ( n45460 , n45456 , n45459 );
buf ( n45461 , n45460 );
not ( n45462 , n44828 );
nand ( n45463 , n45462 , n44838 );
buf ( n45464 , n45463 );
nand ( n45465 , n45461 , n45464 );
buf ( n45466 , n45465 );
buf ( n45467 , n45466 );
xor ( n45468 , n42225 , n42322 );
xor ( n45469 , n45468 , n42385 );
buf ( n45470 , n45469 );
buf ( n45471 , n45470 );
xor ( n45472 , n45467 , n45471 );
xor ( n45473 , n42395 , n42648 );
xor ( n45474 , n45473 , n42719 );
buf ( n45475 , n45474 );
buf ( n45476 , n45475 );
and ( n45477 , n45472 , n45476 );
and ( n45478 , n45467 , n45471 );
or ( n45479 , n45477 , n45478 );
buf ( n45480 , n45479 );
xor ( n45481 , n45452 , n45480 );
buf ( n45482 , n45481 );
not ( n45483 , n45482 );
or ( n45484 , n45207 , n45483 );
xor ( n45485 , n45211 , n45451 );
xnor ( n45486 , n45485 , n45480 );
nand ( n45487 , n45486 , n45202 );
buf ( n45488 , n45487 );
nand ( n45489 , n45484 , n45488 );
buf ( n45490 , n45489 );
xor ( n45491 , n42750 , n42779 );
xor ( n45492 , n45491 , n42960 );
buf ( n45493 , n45492 );
not ( n45494 , n45493 );
buf ( n45495 , n43131 );
buf ( n45496 , n43176 );
xor ( n45497 , n45495 , n45496 );
buf ( n45498 , n43127 );
xnor ( n45499 , n45497 , n45498 );
buf ( n45500 , n45499 );
buf ( n45501 , n45500 );
not ( n45502 , n45501 );
or ( n45503 , n45494 , n45502 );
buf ( n45504 , n44872 );
buf ( n45505 , n44851 );
xor ( n45506 , n45504 , n45505 );
buf ( n45507 , n44882 );
xor ( n45508 , n45506 , n45507 );
buf ( n45509 , n45508 );
buf ( n45510 , n45509 );
xor ( n45511 , n42813 , n42920 );
xor ( n45512 , n45511 , n42956 );
buf ( n45513 , n45512 );
buf ( n45514 , n45513 );
xor ( n45515 , n45510 , n45514 );
buf ( n45516 , n41647 );
not ( n45517 , n45516 );
buf ( n45518 , n43150 );
not ( n45519 , n45518 );
or ( n45520 , n45517 , n45519 );
and ( n45521 , n37293 , n41663 );
not ( n45522 , n37293 );
and ( n45523 , n45522 , n41666 );
or ( n45524 , n45521 , n45523 );
buf ( n45525 , n45524 );
buf ( n45526 , n41705 );
nand ( n45527 , n45525 , n45526 );
buf ( n45528 , n45527 );
buf ( n45529 , n45528 );
nand ( n45530 , n45520 , n45529 );
buf ( n45531 , n45530 );
buf ( n45532 , n45531 );
buf ( n45533 , n42865 );
not ( n45534 , n45533 );
buf ( n45535 , n39726 );
not ( n45536 , n45535 );
or ( n45537 , n45534 , n45536 );
buf ( n45538 , n36527 );
buf ( n45539 , n42862 );
nand ( n45540 , n45538 , n45539 );
buf ( n45541 , n45540 );
buf ( n45542 , n45541 );
nand ( n45543 , n45537 , n45542 );
buf ( n45544 , n45543 );
buf ( n45545 , n45544 );
not ( n45546 , n45545 );
buf ( n45547 , n39803 );
not ( n45548 , n45547 );
or ( n45549 , n45546 , n45548 );
buf ( n45550 , n44141 );
buf ( n45551 , n44129 );
nand ( n45552 , n45550 , n45551 );
buf ( n45553 , n45552 );
buf ( n45554 , n45553 );
nand ( n45555 , n45549 , n45554 );
buf ( n45556 , n45555 );
buf ( n45557 , n45556 );
not ( n45558 , n42468 );
not ( n45559 , n44025 );
or ( n45560 , n45558 , n45559 );
buf ( n45561 , n28305 );
buf ( n45562 , n38994 );
nand ( n45563 , n45561 , n45562 );
buf ( n45564 , n45563 );
nand ( n45565 , n45560 , n45564 );
not ( n45566 , n45565 );
not ( n45567 , n44221 );
or ( n45568 , n45566 , n45567 );
nand ( n45569 , n42448 , n45063 );
nand ( n45570 , n45568 , n45569 );
buf ( n45571 , n45570 );
buf ( n45572 , n43368 );
not ( n45573 , n45572 );
buf ( n45574 , n41977 );
not ( n45575 , n45574 );
or ( n45576 , n45573 , n45575 );
buf ( n45577 , n41843 );
buf ( n45578 , n43365 );
nand ( n45579 , n45577 , n45578 );
buf ( n45580 , n45579 );
buf ( n45581 , n45580 );
nand ( n45582 , n45576 , n45581 );
buf ( n45583 , n45582 );
buf ( n45584 , n45583 );
not ( n45585 , n45584 );
buf ( n45586 , n44338 );
not ( n45587 , n45586 );
or ( n45588 , n45585 , n45587 );
buf ( n45589 , n41852 );
buf ( n45590 , n44236 );
nand ( n45591 , n45589 , n45590 );
buf ( n45592 , n45591 );
buf ( n45593 , n45592 );
nand ( n45594 , n45588 , n45593 );
buf ( n45595 , n45594 );
buf ( n45596 , n45595 );
xor ( n45597 , n45571 , n45596 );
buf ( n45598 , n42049 );
not ( n45599 , n45598 );
buf ( n45600 , n41890 );
not ( n45601 , n45600 );
or ( n45602 , n45599 , n45601 );
buf ( n45603 , n42052 );
buf ( n45604 , n41889 );
nand ( n45605 , n45603 , n45604 );
buf ( n45606 , n45605 );
buf ( n45607 , n45606 );
nand ( n45608 , n45602 , n45607 );
buf ( n45609 , n45608 );
buf ( n45610 , n45609 );
not ( n45611 , n45610 );
buf ( n45612 , n41862 );
not ( n45613 , n45612 );
or ( n45614 , n45611 , n45613 );
buf ( n45615 , n37916 );
not ( n45616 , n45615 );
buf ( n45617 , n45616 );
buf ( n45618 , n45617 );
buf ( n45619 , n44442 );
nand ( n45620 , n45618 , n45619 );
buf ( n45621 , n45620 );
buf ( n45622 , n45621 );
nand ( n45623 , n45614 , n45622 );
buf ( n45624 , n45623 );
buf ( n45625 , n45624 );
and ( n45626 , n45597 , n45625 );
and ( n45627 , n45571 , n45596 );
or ( n45628 , n45626 , n45627 );
buf ( n45629 , n45628 );
buf ( n45630 , n45629 );
xor ( n45631 , n45557 , n45630 );
xor ( n45632 , n44190 , n44223 );
xor ( n45633 , n45632 , n44257 );
buf ( n45634 , n45633 );
and ( n45635 , n45631 , n45634 );
and ( n45636 , n45557 , n45630 );
or ( n45637 , n45635 , n45636 );
buf ( n45638 , n45637 );
buf ( n45639 , n45638 );
xor ( n45640 , n45532 , n45639 );
buf ( n45641 , n44496 );
not ( n45642 , n45641 );
buf ( n45643 , n44725 );
not ( n45644 , n45643 );
or ( n45645 , n45642 , n45644 );
buf ( n45646 , n44533 );
not ( n45647 , n45646 );
buf ( n45648 , n36611 );
not ( n45649 , n45648 );
buf ( n45650 , n45649 );
buf ( n45651 , n45650 );
not ( n45652 , n45651 );
or ( n45653 , n45647 , n45652 );
buf ( n45654 , n36611 );
buf ( n45655 , n44530 );
nand ( n45656 , n45654 , n45655 );
buf ( n45657 , n45656 );
buf ( n45658 , n45657 );
nand ( n45659 , n45653 , n45658 );
buf ( n45660 , n45659 );
buf ( n45661 , n45660 );
buf ( n45662 , n44708 );
nand ( n45663 , n45661 , n45662 );
buf ( n45664 , n45663 );
buf ( n45665 , n45664 );
nand ( n45666 , n45645 , n45665 );
buf ( n45667 , n45666 );
buf ( n45668 , n45667 );
and ( n45669 , n45640 , n45668 );
and ( n45670 , n45532 , n45639 );
or ( n45671 , n45669 , n45670 );
buf ( n45672 , n45671 );
buf ( n45673 , n45672 );
and ( n45674 , n45515 , n45673 );
and ( n45675 , n45510 , n45514 );
or ( n45676 , n45674 , n45675 );
buf ( n45677 , n45676 );
buf ( n45678 , n45677 );
nand ( n45679 , n45503 , n45678 );
buf ( n45680 , n45679 );
buf ( n45681 , n45680 );
buf ( n45682 , n45500 );
not ( n45683 , n45682 );
buf ( n45684 , n45683 );
buf ( n45685 , n45684 );
buf ( n45686 , n45492 );
not ( n45687 , n45686 );
buf ( n45688 , n45687 );
buf ( n45689 , n45688 );
nand ( n45690 , n45685 , n45689 );
buf ( n45691 , n45690 );
buf ( n45692 , n45691 );
nand ( n45693 , n45681 , n45692 );
buf ( n45694 , n45693 );
xor ( n45695 , n45467 , n45471 );
xor ( n45696 , n45695 , n45476 );
buf ( n45697 , n45696 );
or ( n45698 , n45694 , n45697 );
xor ( n45699 , n42966 , n43178 );
xor ( n45700 , n45699 , n43539 );
nand ( n45701 , n45698 , n45700 );
nand ( n45702 , n45694 , n45697 );
nand ( n45703 , n45701 , n45702 );
and ( n45704 , n45490 , n45703 );
not ( n45705 , n45490 );
not ( n45706 , n45703 );
and ( n45707 , n45705 , n45706 );
nor ( n45708 , n45704 , n45707 );
not ( n45709 , n45708 );
xor ( n45710 , n43833 , n45709 );
not ( n45711 , n42339 );
not ( n45712 , n42948 );
or ( n45713 , n45711 , n45712 );
buf ( n45714 , n42378 );
xor ( n45715 , n42343 , n38244 );
buf ( n45716 , n45715 );
nand ( n45717 , n45714 , n45716 );
buf ( n45718 , n45717 );
nand ( n45719 , n45713 , n45718 );
buf ( n45720 , n45719 );
buf ( n45721 , n25431 );
buf ( n45722 , n45721 );
buf ( n45723 , n45722 );
buf ( n45724 , n45723 );
buf ( n45725 , n24784 );
xor ( n45726 , n45724 , n45725 );
buf ( n45727 , n45726 );
buf ( n45728 , n45727 );
not ( n45729 , n45728 );
buf ( n45730 , n45729 );
buf ( n45731 , n45730 );
not ( n45732 , n45731 );
and ( n45733 , n24811 , n24784 );
not ( n45734 , n24811 );
buf ( n45735 , n24784 );
not ( n45736 , n45735 );
buf ( n45737 , n45736 );
and ( n45738 , n45734 , n45737 );
nor ( n45739 , n45733 , n45738 );
nand ( n45740 , n45739 , n45730 );
not ( n45741 , n45740 );
not ( n45742 , n45741 );
buf ( n45743 , n45742 );
not ( n45744 , n45743 );
or ( n45745 , n45732 , n45744 );
buf ( n45746 , n24811 );
not ( n45747 , n45746 );
buf ( n45748 , n45747 );
buf ( n45749 , n45748 );
buf ( n45750 , n45749 );
buf ( n45751 , n45750 );
not ( n45752 , n45751 );
buf ( n45753 , n45752 );
buf ( n45754 , n45753 );
not ( n45755 , n45754 );
buf ( n45756 , n41619 );
not ( n45757 , n45756 );
or ( n45758 , n45755 , n45757 );
buf ( n45759 , n39005 );
buf ( n45760 , n45750 );
nand ( n45761 , n45759 , n45760 );
buf ( n45762 , n45761 );
buf ( n45763 , n45762 );
nand ( n45764 , n45758 , n45763 );
buf ( n45765 , n45764 );
buf ( n45766 , n45765 );
nand ( n45767 , n45745 , n45766 );
buf ( n45768 , n45767 );
buf ( n45769 , n45768 );
nor ( n45770 , n45720 , n45769 );
buf ( n45771 , n45770 );
buf ( n45772 , n45771 );
not ( n45773 , n45772 );
buf ( n45774 , n45773 );
buf ( n45775 , n45774 );
not ( n45776 , n45775 );
xor ( n45777 , n44760 , n44788 );
xor ( n45778 , n45777 , n44793 );
buf ( n45779 , n45778 );
buf ( n45780 , n45779 );
not ( n45781 , n45780 );
or ( n45782 , n45776 , n45781 );
nand ( n45783 , n45719 , n45768 );
buf ( n45784 , n45783 );
nand ( n45785 , n45782 , n45784 );
buf ( n45786 , n45785 );
not ( n45787 , n45786 );
buf ( n45788 , n43137 );
buf ( n45789 , n43160 );
xor ( n45790 , n45788 , n45789 );
buf ( n45791 , n43165 );
xnor ( n45792 , n45790 , n45791 );
buf ( n45793 , n45792 );
nand ( n45794 , n45787 , n45793 );
xor ( n45795 , n44735 , n44797 );
xor ( n45796 , n45795 , n44822 );
and ( n45797 , n45794 , n45796 );
nor ( n45798 , n45793 , n45787 );
nor ( n45799 , n45797 , n45798 );
buf ( n45800 , n45799 );
not ( n45801 , n45800 );
buf ( n45802 , n45801 );
buf ( n45803 , n45802 );
not ( n45804 , n45803 );
buf ( n45805 , n41608 );
not ( n45806 , n45805 );
buf ( n45807 , n40067 );
not ( n45808 , n45807 );
or ( n45809 , n45806 , n45808 );
buf ( n45810 , n36427 );
buf ( n45811 , n41611 );
nand ( n45812 , n45810 , n45811 );
buf ( n45813 , n45812 );
buf ( n45814 , n45813 );
nand ( n45815 , n45809 , n45814 );
buf ( n45816 , n45815 );
buf ( n45817 , n45816 );
buf ( n45818 , n44267 );
and ( n45819 , n45817 , n45818 );
not ( n45820 , n44281 );
nor ( n45821 , n45820 , n41577 );
buf ( n45822 , n45821 );
nor ( n45823 , n45819 , n45822 );
buf ( n45824 , n45823 );
buf ( n45825 , n45824 );
not ( n45826 , n45825 );
buf ( n45827 , n45826 );
buf ( n45828 , n45827 );
not ( n45829 , n45828 );
buf ( n45830 , n42315 );
not ( n45831 , n45830 );
buf ( n45832 , n44934 );
not ( n45833 , n45832 );
or ( n45834 , n45831 , n45833 );
buf ( n45835 , n42266 );
not ( n45836 , n45835 );
buf ( n45837 , n37078 );
not ( n45838 , n45837 );
buf ( n45839 , n45838 );
buf ( n45840 , n45839 );
not ( n45841 , n45840 );
or ( n45842 , n45836 , n45841 );
buf ( n45843 , n37078 );
buf ( n45844 , n42263 );
nand ( n45845 , n45843 , n45844 );
buf ( n45846 , n45845 );
buf ( n45847 , n45846 );
nand ( n45848 , n45842 , n45847 );
buf ( n45849 , n45848 );
buf ( n45850 , n45849 );
buf ( n45851 , n42252 );
nand ( n45852 , n45850 , n45851 );
buf ( n45853 , n45852 );
buf ( n45854 , n45853 );
nand ( n45855 , n45834 , n45854 );
buf ( n45856 , n45855 );
buf ( n45857 , n45856 );
not ( n45858 , n45857 );
or ( n45859 , n45829 , n45858 );
buf ( n45860 , n45827 );
buf ( n45861 , n45856 );
or ( n45862 , n45860 , n45861 );
xor ( n45863 , n44329 , n44477 );
xor ( n45864 , n45863 , n44413 );
buf ( n45865 , n45864 );
nand ( n45866 , n45862 , n45865 );
buf ( n45867 , n45866 );
buf ( n45868 , n45867 );
nand ( n45869 , n45859 , n45868 );
buf ( n45870 , n45869 );
buf ( n45871 , n45870 );
not ( n45872 , n45871 );
xor ( n45873 , n44265 , n44293 );
xnor ( n45874 , n45873 , n44481 );
buf ( n45875 , n45874 );
not ( n45876 , n45875 );
or ( n45877 , n45872 , n45876 );
buf ( n45878 , n45874 );
buf ( n45879 , n45870 );
or ( n45880 , n45878 , n45879 );
xor ( n45881 , n44149 , n44173 );
xor ( n45882 , n45881 , n44261 );
buf ( n45883 , n45882 );
buf ( n45884 , n45883 );
xor ( n45885 , n44427 , n44455 );
xor ( n45886 , n45885 , n44473 );
buf ( n45887 , n45886 );
not ( n45888 , n45887 );
buf ( n45889 , n41705 );
not ( n45890 , n45889 );
buf ( n45891 , n41663 );
buf ( n45892 , n42573 );
and ( n45893 , n45891 , n45892 );
not ( n45894 , n45891 );
buf ( n45895 , n37686 );
and ( n45896 , n45894 , n45895 );
nor ( n45897 , n45893 , n45896 );
buf ( n45898 , n45897 );
buf ( n45899 , n45898 );
not ( n45900 , n45899 );
or ( n45901 , n45890 , n45900 );
buf ( n45902 , n45524 );
buf ( n45903 , n41647 );
nand ( n45904 , n45902 , n45903 );
buf ( n45905 , n45904 );
buf ( n45906 , n45905 );
nand ( n45907 , n45901 , n45906 );
buf ( n45908 , n45907 );
buf ( n45909 , n44586 );
not ( n45910 , n45909 );
buf ( n45911 , n25184 );
not ( n45912 , n45911 );
buf ( n45913 , n42973 );
not ( n45914 , n45913 );
or ( n45915 , n45912 , n45914 );
not ( n45916 , n37782 );
buf ( n45917 , n45916 );
buf ( n45918 , n25183 );
nand ( n45919 , n45917 , n45918 );
buf ( n45920 , n45919 );
buf ( n45921 , n45920 );
nand ( n45922 , n45915 , n45921 );
buf ( n45923 , n45922 );
buf ( n45924 , n45923 );
not ( n45925 , n45924 );
or ( n45926 , n45910 , n45925 );
buf ( n45927 , n44326 );
buf ( n45928 , n43909 );
nand ( n45929 , n45927 , n45928 );
buf ( n45930 , n45929 );
buf ( n45931 , n45930 );
nand ( n45932 , n45926 , n45931 );
buf ( n45933 , n45932 );
or ( n45934 , n45908 , n45933 );
not ( n45935 , n45934 );
or ( n45936 , n45888 , n45935 );
nand ( n45937 , n45908 , n45933 );
nand ( n45938 , n45936 , n45937 );
buf ( n45939 , n45938 );
xor ( n45940 , n45884 , n45939 );
buf ( n45941 , n42668 );
not ( n45942 , n45941 );
buf ( n45943 , n44812 );
not ( n45944 , n45943 );
or ( n45945 , n45942 , n45944 );
buf ( n45946 , n42672 );
not ( n45947 , n45946 );
buf ( n45948 , n39280 );
not ( n45949 , n45948 );
or ( n45950 , n45947 , n45949 );
buf ( n45951 , n39277 );
buf ( n45952 , n42679 );
nand ( n45953 , n45951 , n45952 );
buf ( n45954 , n45953 );
buf ( n45955 , n45954 );
nand ( n45956 , n45950 , n45955 );
buf ( n45957 , n45956 );
buf ( n45958 , n45957 );
buf ( n45959 , n42712 );
nand ( n45960 , n45958 , n45959 );
buf ( n45961 , n45960 );
buf ( n45962 , n45961 );
nand ( n45963 , n45945 , n45962 );
buf ( n45964 , n45963 );
buf ( n45965 , n45964 );
and ( n45966 , n45940 , n45965 );
and ( n45967 , n45884 , n45939 );
or ( n45968 , n45966 , n45967 );
buf ( n45969 , n45968 );
buf ( n45970 , n45969 );
nand ( n45971 , n45880 , n45970 );
buf ( n45972 , n45971 );
buf ( n45973 , n45972 );
nand ( n45974 , n45877 , n45973 );
buf ( n45975 , n45974 );
buf ( n45976 , n45975 );
not ( n45977 , n45976 );
or ( n45978 , n45804 , n45977 );
buf ( n45979 , n45975 );
not ( n45980 , n45979 );
buf ( n45981 , n45980 );
buf ( n45982 , n45981 );
not ( n45983 , n45982 );
buf ( n45984 , n45799 );
not ( n45985 , n45984 );
or ( n45986 , n45983 , n45985 );
xor ( n45987 , n44485 , n44563 );
xor ( n45988 , n45987 , n44119 );
buf ( n45989 , n45988 );
nand ( n45990 , n45986 , n45989 );
buf ( n45991 , n45990 );
buf ( n45992 , n45991 );
nand ( n45993 , n45978 , n45992 );
buf ( n45994 , n45993 );
buf ( n45995 , n45994 );
not ( n45996 , n45995 );
xor ( n45997 , n44566 , n44706 );
xor ( n45998 , n45997 , n45198 );
buf ( n45999 , n45998 );
buf ( n46000 , n45999 );
not ( n46001 , n46000 );
buf ( n46002 , n46001 );
buf ( n46003 , n46002 );
nand ( n46004 , n45996 , n46003 );
buf ( n46005 , n46004 );
not ( n46006 , n46005 );
xor ( n46007 , n44826 , n44901 );
xor ( n46008 , n46007 , n45193 );
buf ( n46009 , n46008 );
buf ( n46010 , n46009 );
not ( n46011 , n46010 );
buf ( n46012 , n45677 );
buf ( n46013 , n45688 );
xor ( n46014 , n46012 , n46013 );
buf ( n46015 , n45684 );
xnor ( n46016 , n46014 , n46015 );
buf ( n46017 , n46016 );
buf ( n46018 , n46017 );
not ( n46019 , n46018 );
buf ( n46020 , n46019 );
buf ( n46021 , n46020 );
not ( n46022 , n46021 );
or ( n46023 , n46011 , n46022 );
buf ( n46024 , n46009 );
not ( n46025 , n46024 );
buf ( n46026 , n46025 );
buf ( n46027 , n46026 );
not ( n46028 , n46027 );
buf ( n46029 , n46017 );
not ( n46030 , n46029 );
or ( n46031 , n46028 , n46030 );
xor ( n46032 , n44921 , n44942 );
xor ( n46033 , n46032 , n45188 );
buf ( n46034 , n46033 );
buf ( n46035 , n46034 );
not ( n46036 , n42668 );
not ( n46037 , n45957 );
or ( n46038 , n46036 , n46037 );
not ( n46039 , n42672 );
not ( n46040 , n38218 );
or ( n46041 , n46039 , n46040 );
buf ( n46042 , n45227 );
buf ( n46043 , n42679 );
nand ( n46044 , n46042 , n46043 );
buf ( n46045 , n46044 );
nand ( n46046 , n46041 , n46045 );
not ( n46047 , n42710 );
nand ( n46048 , n46046 , n46047 );
nand ( n46049 , n46038 , n46048 );
not ( n46050 , n46049 );
buf ( n46051 , n45006 );
buf ( n46052 , n44974 );
xor ( n46053 , n46051 , n46052 );
buf ( n46054 , n45032 );
xnor ( n46055 , n46053 , n46054 );
buf ( n46056 , n46055 );
buf ( n46057 , n46056 );
not ( n46058 , n46057 );
buf ( n46059 , n46058 );
not ( n46060 , n46059 );
or ( n46061 , n46050 , n46060 );
not ( n46062 , n46056 );
buf ( n46063 , n46049 );
not ( n46064 , n46063 );
buf ( n46065 , n46064 );
not ( n46066 , n46065 );
or ( n46067 , n46062 , n46066 );
buf ( n46068 , n39986 );
not ( n46069 , n46068 );
buf ( n46070 , n44999 );
not ( n46071 , n46070 );
or ( n46072 , n46069 , n46071 );
not ( n46073 , n24092 );
and ( n46074 , n29269 , n46073 );
not ( n46075 , n29269 );
and ( n46076 , n46075 , n24092 );
or ( n46077 , n46074 , n46076 );
buf ( n46078 , n46077 );
buf ( n46079 , n40002 );
nand ( n46080 , n46078 , n46079 );
buf ( n46081 , n46080 );
buf ( n46082 , n46081 );
nand ( n46083 , n46072 , n46082 );
buf ( n46084 , n46083 );
buf ( n46085 , n46084 );
buf ( n46086 , n43063 );
not ( n46087 , n46086 );
buf ( n46088 , n39478 );
not ( n46089 , n46088 );
or ( n46090 , n46087 , n46089 );
buf ( n46091 , n43265 );
buf ( n46092 , n43064 );
nand ( n46093 , n46091 , n46092 );
buf ( n46094 , n46093 );
buf ( n46095 , n46094 );
nand ( n46096 , n46090 , n46095 );
buf ( n46097 , n46096 );
buf ( n46098 , n46097 );
not ( n46099 , n46098 );
buf ( n46100 , n42521 );
not ( n46101 , n46100 );
or ( n46102 , n46099 , n46101 );
buf ( n46103 , n39715 );
buf ( n46104 , n44460 );
nand ( n46105 , n46103 , n46104 );
buf ( n46106 , n46105 );
buf ( n46107 , n46106 );
nand ( n46108 , n46102 , n46107 );
buf ( n46109 , n46108 );
buf ( n46110 , n46109 );
xor ( n46111 , n46085 , n46110 );
buf ( n46112 , n25977 );
buf ( n46113 , n46112 );
buf ( n46114 , n46113 );
buf ( n46115 , n46114 );
buf ( n46116 , n46115 );
buf ( n46117 , n46116 );
buf ( n46118 , n46117 );
not ( n46119 , n46118 );
buf ( n46120 , n37602 );
not ( n46121 , n46120 );
or ( n46122 , n46119 , n46121 );
buf ( n46123 , n38798 );
buf ( n46124 , n46117 );
not ( n46125 , n46124 );
buf ( n46126 , n46125 );
buf ( n46127 , n46126 );
nand ( n46128 , n46123 , n46127 );
buf ( n46129 , n46128 );
buf ( n46130 , n46129 );
nand ( n46131 , n46122 , n46130 );
buf ( n46132 , n46131 );
buf ( n46133 , n39667 );
buf ( n46134 , n44967 );
not ( n46135 , n46134 );
buf ( n46136 , n46135 );
buf ( n46137 , n46136 );
or ( n46138 , n46133 , n46137 );
nand ( n46139 , C1 , n46138 );
buf ( n46140 , n46139 );
buf ( n46141 , n46140 );
and ( n46142 , n46111 , n46141 );
and ( n46143 , n46085 , n46110 );
or ( n46144 , n46142 , n46143 );
buf ( n46145 , n46144 );
nand ( n46146 , n46067 , n46145 );
nand ( n46147 , n46061 , n46146 );
buf ( n46148 , n46147 );
buf ( n46149 , n41736 );
not ( n46150 , n46149 );
buf ( n46151 , n44635 );
not ( n46152 , n46151 );
or ( n46153 , n46150 , n46152 );
buf ( n46154 , n43400 );
buf ( n46155 , n41748 );
nand ( n46156 , n46154 , n46155 );
buf ( n46157 , n46156 );
buf ( n46158 , n46157 );
nand ( n46159 , n46153 , n46158 );
buf ( n46160 , n46159 );
buf ( n46161 , n46160 );
not ( n46162 , n46161 );
buf ( n46163 , n38127 );
not ( n46164 , n46163 );
buf ( n46165 , n46164 );
buf ( n46166 , n46165 );
not ( n46167 , n46166 );
or ( n46168 , n46162 , n46167 );
buf ( n46169 , n45132 );
buf ( n46170 , n38054 );
buf ( n46171 , n46170 );
buf ( n46172 , n46171 );
buf ( n46173 , n46172 );
nand ( n46174 , n46169 , n46173 );
buf ( n46175 , n46174 );
buf ( n46176 , n46175 );
nand ( n46177 , n46168 , n46176 );
buf ( n46178 , n46177 );
buf ( n46179 , n46178 );
not ( n46180 , n46179 );
buf ( n46181 , n46180 );
buf ( n46182 , n46181 );
not ( n46183 , n46182 );
and ( n46184 , n45022 , n42566 );
and ( n46185 , n25160 , n42455 );
not ( n46186 , n25160 );
and ( n46187 , n46186 , n38821 );
or ( n46188 , n46185 , n46187 );
and ( n46189 , n46188 , n42631 );
nor ( n46190 , n46184 , n46189 );
buf ( n46191 , n46190 );
not ( n46192 , n46191 );
or ( n46193 , n46183 , n46192 );
buf ( n46194 , n36982 );
buf ( n46195 , n42008 );
buf ( n46196 , n36926 );
and ( n46197 , n46195 , n46196 );
not ( n46198 , n46195 );
buf ( n46199 , n42062 );
and ( n46200 , n46198 , n46199 );
nor ( n46201 , n46197 , n46200 );
buf ( n46202 , n46201 );
buf ( n46203 , n46202 );
or ( n46204 , n46194 , n46203 );
buf ( n46205 , n36909 );
buf ( n46206 , n45170 );
or ( n46207 , n46205 , n46206 );
nand ( n46208 , n46204 , n46207 );
buf ( n46209 , n46208 );
buf ( n46210 , n46209 );
nand ( n46211 , n46193 , n46210 );
buf ( n46212 , n46211 );
buf ( n46213 , n46212 );
buf ( n46214 , n46190 );
not ( n46215 , n46214 );
buf ( n46216 , n46215 );
buf ( n46217 , n46216 );
buf ( n46218 , n46178 );
nand ( n46219 , n46217 , n46218 );
buf ( n46220 , n46219 );
buf ( n46221 , n46220 );
nand ( n46222 , n46213 , n46221 );
buf ( n46223 , n46222 );
buf ( n46224 , n46223 );
buf ( n46225 , n45741 );
buf ( n46226 , n46225 );
not ( n46227 , n46226 );
buf ( n46228 , n45753 );
not ( n46229 , n46228 );
buf ( n46230 , n36054 );
not ( n46231 , n46230 );
or ( n46232 , n46229 , n46231 );
buf ( n46233 , n43851 );
buf ( n46234 , n45750 );
nand ( n46235 , n46233 , n46234 );
buf ( n46236 , n46235 );
buf ( n46237 , n46236 );
nand ( n46238 , n46232 , n46237 );
buf ( n46239 , n46238 );
buf ( n46240 , n46239 );
not ( n46241 , n46240 );
or ( n46242 , n46227 , n46241 );
buf ( n46243 , n45765 );
buf ( n46244 , n45730 );
not ( n46245 , n46244 );
buf ( n46246 , n46245 );
buf ( n46247 , n46246 );
nand ( n46248 , n46243 , n46247 );
buf ( n46249 , n46248 );
buf ( n46250 , n46249 );
nand ( n46251 , n46242 , n46250 );
buf ( n46252 , n46251 );
buf ( n46253 , n46252 );
xor ( n46254 , n46224 , n46253 );
xor ( n46255 , n45120 , n45151 );
xor ( n46256 , n46255 , n45178 );
buf ( n46257 , n46256 );
buf ( n46258 , n46257 );
and ( n46259 , n46254 , n46258 );
and ( n46260 , n46224 , n46253 );
or ( n46261 , n46259 , n46260 );
buf ( n46262 , n46261 );
buf ( n46263 , n46262 );
xor ( n46264 , n46148 , n46263 );
xor ( n46265 , n45044 , n45048 );
xor ( n46266 , n46265 , n45183 );
buf ( n46267 , n46266 );
buf ( n46268 , n46267 );
and ( n46269 , n46264 , n46268 );
and ( n46270 , n46148 , n46263 );
or ( n46271 , n46269 , n46270 );
buf ( n46272 , n46271 );
buf ( n46273 , n46272 );
xor ( n46274 , n46035 , n46273 );
buf ( n46275 , n42252 );
not ( n46276 , n46275 );
and ( n46277 , n37146 , n42263 );
not ( n46278 , n37146 );
and ( n46279 , n46278 , n42266 );
or ( n46280 , n46277 , n46279 );
buf ( n46281 , n46280 );
not ( n46282 , n46281 );
or ( n46283 , n46276 , n46282 );
buf ( n46284 , n45849 );
buf ( n46285 , n42315 );
nand ( n46286 , n46284 , n46285 );
buf ( n46287 , n46286 );
buf ( n46288 , n46287 );
nand ( n46289 , n46283 , n46288 );
buf ( n46290 , n46289 );
buf ( n46291 , n46290 );
buf ( n46292 , n43906 );
not ( n46293 , n46292 );
buf ( n46294 , n46293 );
buf ( n46295 , n46294 );
not ( n46296 , n46295 );
buf ( n46297 , n45923 );
not ( n46298 , n46297 );
or ( n46299 , n46296 , n46298 );
buf ( n46300 , n25184 );
not ( n46301 , n46300 );
buf ( n46302 , n37589 );
not ( n46303 , n46302 );
or ( n46304 , n46301 , n46303 );
buf ( n46305 , n37598 );
buf ( n46306 , n25183 );
nand ( n46307 , n46305 , n46306 );
buf ( n46308 , n46307 );
buf ( n46309 , n46308 );
nand ( n46310 , n46304 , n46309 );
buf ( n46311 , n46310 );
buf ( n46312 , n46311 );
buf ( n46313 , n44586 );
nand ( n46314 , n46312 , n46313 );
buf ( n46315 , n46314 );
buf ( n46316 , n46315 );
nand ( n46317 , n46299 , n46316 );
buf ( n46318 , n46317 );
buf ( n46319 , n46318 );
not ( n46320 , n46319 );
buf ( n46321 , n46320 );
not ( n46322 , n46321 );
buf ( n46323 , n42865 );
not ( n46324 , n46323 );
buf ( n46325 , n36500 );
not ( n46326 , n46325 );
or ( n46327 , n46324 , n46326 );
buf ( n46328 , n43265 );
buf ( n46329 , n42862 );
nand ( n46330 , n46328 , n46329 );
buf ( n46331 , n46330 );
buf ( n46332 , n46331 );
nand ( n46333 , n46327 , n46332 );
buf ( n46334 , n46333 );
buf ( n46335 , n46334 );
not ( n46336 , n46335 );
buf ( n46337 , n32963 );
buf ( n46338 , n36092 );
and ( n46339 , n46337 , n46338 );
buf ( n46340 , n46339 );
buf ( n46341 , n46340 );
not ( n46342 , n46341 );
or ( n46343 , n46336 , n46342 );
buf ( n46344 , n32963 );
not ( n46345 , n46344 );
buf ( n46346 , n46097 );
nand ( n46347 , n46345 , n46346 );
buf ( n46348 , n46347 );
buf ( n46349 , n46348 );
nand ( n46350 , n46343 , n46349 );
buf ( n46351 , n46350 );
buf ( n46352 , n46351 );
not ( n46353 , n46352 );
buf ( n46354 , n42631 );
not ( n46355 , n46354 );
not ( n46356 , n25159 );
buf ( n46357 , n46356 );
buf ( n46358 , n42485 );
and ( n46359 , n46357 , n46358 );
not ( n46360 , n46357 );
buf ( n46361 , n30187 );
and ( n46362 , n46360 , n46361 );
nor ( n46363 , n46359 , n46362 );
buf ( n46364 , n46363 );
buf ( n46365 , n46364 );
not ( n46366 , n46365 );
or ( n46367 , n46355 , n46366 );
buf ( n46368 , n46188 );
buf ( n46369 , n42566 );
nand ( n46370 , n46368 , n46369 );
buf ( n46371 , n46370 );
buf ( n46372 , n46371 );
nand ( n46373 , n46367 , n46372 );
buf ( n46374 , n46373 );
buf ( n46375 , n46374 );
not ( n46376 , n46375 );
buf ( n46377 , n46376 );
buf ( n46378 , n46377 );
nand ( n46379 , n46353 , n46378 );
buf ( n46380 , n46379 );
buf ( n46381 , n46380 );
buf ( n46382 , n25951 );
not ( n46383 , n46382 );
buf ( n46384 , n46383 );
buf ( n46385 , n46384 );
buf ( n46386 , n46385 );
buf ( n46387 , n46386 );
buf ( n46388 , n46387 );
not ( n46389 , n46388 );
buf ( n46390 , n46389 );
buf ( n46391 , n46390 );
not ( n46392 , n46391 );
buf ( n46393 , n46392 );
buf ( n46394 , n46393 );
buf ( n46395 , n38834 );
and ( n46396 , n46394 , n46395 );
not ( n46397 , n46394 );
buf ( n46398 , n37649 );
and ( n46399 , n46397 , n46398 );
nor ( n46400 , n46396 , n46399 );
buf ( n46401 , n46400 );
buf ( n46402 , n43053 );
buf ( n46403 , n46132 );
nand ( n46404 , n46402 , n46403 );
buf ( n46405 , n46404 );
buf ( n46406 , n46405 );
nand ( n46407 , C1 , n46406 );
buf ( n46408 , n46407 );
buf ( n46409 , n46408 );
and ( n46410 , n46381 , n46409 );
buf ( n46411 , n46351 );
buf ( n46412 , n46374 );
and ( n46413 , n46411 , n46412 );
buf ( n46414 , n46413 );
buf ( n46415 , n46414 );
nor ( n46416 , n46410 , n46415 );
buf ( n46417 , n46416 );
not ( n46418 , n46417 );
or ( n46419 , n46322 , n46418 );
buf ( n46420 , n45570 );
not ( n46421 , n46420 );
buf ( n46422 , n43108 );
not ( n46423 , n46422 );
buf ( n46424 , n44381 );
not ( n46425 , n46424 );
or ( n46426 , n46423 , n46425 );
buf ( n46427 , n37881 );
buf ( n46428 , n43099 );
nand ( n46429 , n46427 , n46428 );
buf ( n46430 , n46429 );
buf ( n46431 , n46430 );
nand ( n46432 , n46426 , n46431 );
buf ( n46433 , n46432 );
not ( n46434 , n46433 );
not ( n46435 , n41862 );
or ( n46436 , n46434 , n46435 );
nand ( n46437 , n45609 , n45617 );
nand ( n46438 , n46436 , n46437 );
buf ( n46439 , n46438 );
not ( n46440 , n46439 );
buf ( n46441 , n46440 );
buf ( n46442 , n46441 );
not ( n46443 , n46442 );
or ( n46444 , n46421 , n46443 );
buf ( n46445 , n41969 );
buf ( n46446 , n41981 );
not ( n46447 , n46446 );
buf ( n46448 , n42075 );
not ( n46449 , n46448 );
and ( n46450 , n46447 , n46449 );
buf ( n46451 , n41844 );
buf ( n46452 , n42075 );
and ( n46453 , n46451 , n46452 );
nor ( n46454 , n46450 , n46453 );
buf ( n46455 , n46454 );
buf ( n46456 , n46455 );
or ( n46457 , n46445 , n46456 );
buf ( n46458 , n45583 );
not ( n46459 , n46458 );
buf ( n46460 , n46459 );
buf ( n46461 , n46460 );
buf ( n46462 , n42210 );
or ( n46463 , n46461 , n46462 );
nand ( n46464 , n46457 , n46463 );
buf ( n46465 , n46464 );
buf ( n46466 , n46465 );
nand ( n46467 , n46444 , n46466 );
buf ( n46468 , n46467 );
buf ( n46469 , n46468 );
buf ( n46470 , n45570 );
not ( n46471 , n46470 );
buf ( n46472 , n46438 );
nand ( n46473 , n46471 , n46472 );
buf ( n46474 , n46473 );
buf ( n46475 , n46474 );
nand ( n46476 , n46469 , n46475 );
buf ( n46477 , n46476 );
not ( n46478 , n46477 );
not ( n46479 , n46478 );
nand ( n46480 , n46419 , n46479 );
buf ( n46481 , n46380 );
buf ( n46482 , n46408 );
and ( n46483 , n46481 , n46482 );
buf ( n46484 , n46414 );
nor ( n46485 , n46483 , n46484 );
buf ( n46486 , n46485 );
buf ( n46487 , n46486 );
not ( n46488 , n46487 );
buf ( n46489 , n46318 );
nand ( n46490 , n46488 , n46489 );
buf ( n46491 , n46490 );
nand ( n46492 , n46480 , n46491 );
buf ( n46493 , n46492 );
xor ( n46494 , n46291 , n46493 );
xor ( n46495 , n45557 , n45630 );
xor ( n46496 , n46495 , n45634 );
buf ( n46497 , n46496 );
buf ( n46498 , n46497 );
and ( n46499 , n46494 , n46498 );
and ( n46500 , n46291 , n46493 );
or ( n46501 , n46499 , n46500 );
buf ( n46502 , n46501 );
buf ( n46503 , n46502 );
buf ( n46504 , n45771 );
not ( n46505 , n46504 );
buf ( n46506 , n45783 );
nand ( n46507 , n46505 , n46506 );
buf ( n46508 , n46507 );
xnor ( n46509 , n46508 , n45779 );
buf ( n46510 , n46509 );
xor ( n46511 , n46503 , n46510 );
xor ( n46512 , n45532 , n45639 );
xor ( n46513 , n46512 , n45668 );
buf ( n46514 , n46513 );
buf ( n46515 , n46514 );
and ( n46516 , n46511 , n46515 );
and ( n46517 , n46503 , n46510 );
or ( n46518 , n46516 , n46517 );
buf ( n46519 , n46518 );
buf ( n46520 , n46519 );
and ( n46521 , n46274 , n46520 );
and ( n46522 , n46035 , n46273 );
or ( n46523 , n46521 , n46522 );
buf ( n46524 , n46523 );
buf ( n46525 , n46524 );
nand ( n46526 , n46031 , n46525 );
buf ( n46527 , n46526 );
buf ( n46528 , n46527 );
nand ( n46529 , n46023 , n46528 );
buf ( n46530 , n46529 );
not ( n46531 , n46530 );
or ( n46532 , n46006 , n46531 );
buf ( n46533 , n45999 );
buf ( n46534 , n45994 );
nand ( n46535 , n46533 , n46534 );
buf ( n46536 , n46535 );
nand ( n46537 , n46532 , n46536 );
xnor ( n46538 , n45710 , n46537 );
buf ( n46539 , n46538 );
buf ( n46540 , n45680 );
buf ( n46541 , n45691 );
nand ( n46542 , n46540 , n46541 );
buf ( n46543 , n46542 );
xor ( n46544 , n45697 , n46543 );
not ( n46545 , n45700 );
and ( n46546 , n46544 , n46545 );
not ( n46547 , n46544 );
and ( n46548 , n46547 , n45700 );
nor ( n46549 , n46546 , n46548 );
buf ( n46550 , n46549 );
buf ( n46551 , n45799 );
buf ( n46552 , n45981 );
and ( n46553 , n46551 , n46552 );
not ( n46554 , n46551 );
buf ( n46555 , n45975 );
and ( n46556 , n46554 , n46555 );
nor ( n46557 , n46553 , n46556 );
buf ( n46558 , n46557 );
buf ( n46559 , n45988 );
not ( n46560 , n46559 );
buf ( n46561 , n46560 );
and ( n46562 , n46558 , n46561 );
not ( n46563 , n46558 );
and ( n46564 , n46563 , n45988 );
nor ( n46565 , n46562 , n46564 );
xor ( n46566 , n45510 , n45514 );
xor ( n46567 , n46566 , n45673 );
buf ( n46568 , n46567 );
buf ( n46569 , n46568 );
buf ( n46570 , n45786 );
buf ( n46571 , n45793 );
xor ( n46572 , n46570 , n46571 );
buf ( n46573 , n45796 );
xnor ( n46574 , n46572 , n46573 );
buf ( n46575 , n46574 );
buf ( n46576 , n46575 );
xor ( n46577 , n46569 , n46576 );
buf ( n46578 , n42378 );
not ( n46579 , n46578 );
not ( n46580 , n42343 );
not ( n46581 , n38742 );
or ( n46582 , n46580 , n46581 );
or ( n46583 , n38742 , n42343 );
nand ( n46584 , n46582 , n46583 );
buf ( n46585 , n46584 );
not ( n46586 , n46585 );
or ( n46587 , n46579 , n46586 );
buf ( n46588 , n45715 );
buf ( n46589 , n42339 );
nand ( n46590 , n46588 , n46589 );
buf ( n46591 , n46590 );
buf ( n46592 , n46591 );
nand ( n46593 , n46587 , n46592 );
buf ( n46594 , n46593 );
buf ( n46595 , n46594 );
buf ( n46596 , n38374 );
buf ( n46597 , n24638 );
and ( n46598 , n46596 , n46597 );
not ( n46599 , n46596 );
buf ( n46600 , n38348 );
and ( n46601 , n46599 , n46600 );
nor ( n46602 , n46598 , n46601 );
buf ( n46603 , n46602 );
buf ( n46604 , n46603 );
not ( n46605 , n46604 );
buf ( n46606 , n46605 );
not ( n46607 , n46606 );
not ( n46608 , n45077 );
or ( n46609 , n46607 , n46608 );
nand ( n46610 , n46603 , n38397 );
not ( n46611 , n46610 );
buf ( n46612 , n42403 );
buf ( n46613 , n38371 );
not ( n46614 , n46613 );
buf ( n46615 , n46614 );
buf ( n46616 , n46615 );
nand ( n46617 , n46612 , n46616 );
buf ( n46618 , n46617 );
nand ( n46619 , n46611 , n46618 );
not ( n46620 , n46619 );
buf ( n46621 , n42403 );
not ( n46622 , n46621 );
buf ( n46623 , n46622 );
and ( n46624 , n46623 , n42195 );
not ( n46625 , n46623 );
and ( n46626 , n46625 , n29360 );
or ( n46627 , n46624 , n46626 );
nand ( n46628 , n46620 , n46627 );
nand ( n46629 , n46609 , n46628 );
not ( n46630 , n46629 );
buf ( n46631 , n39980 );
not ( n46632 , n46631 );
buf ( n46633 , n46632 );
not ( n46634 , n46633 );
not ( n46635 , n46077 );
or ( n46636 , n46634 , n46635 );
buf ( n46637 , n24092 );
not ( n46638 , n46637 );
buf ( n46639 , n29287 );
not ( n46640 , n46639 );
buf ( n46641 , n46640 );
buf ( n46642 , n46641 );
not ( n46643 , n46642 );
or ( n46644 , n46638 , n46643 );
buf ( n46645 , n39653 );
buf ( n46646 , n40009 );
nand ( n46647 , n46645 , n46646 );
buf ( n46648 , n46647 );
buf ( n46649 , n46648 );
nand ( n46650 , n46644 , n46649 );
buf ( n46651 , n46650 );
nand ( n46652 , n46651 , n40002 );
nand ( n46653 , n46636 , n46652 );
not ( n46654 , n46653 );
or ( n46655 , n46630 , n46654 );
or ( n46656 , n46653 , n46629 );
not ( n46657 , n28410 );
buf ( n46658 , n46657 );
not ( n46659 , n46658 );
buf ( n46660 , n46659 );
buf ( n46661 , n46660 );
not ( n46662 , n46661 );
buf ( n46663 , n41778 );
not ( n46664 , n46663 );
or ( n46665 , n46662 , n46664 );
not ( n46666 , n28411 );
nand ( n46667 , n46666 , n41769 );
buf ( n46668 , n46667 );
nand ( n46669 , n46665 , n46668 );
buf ( n46670 , n46669 );
not ( n46671 , n46670 );
not ( n46672 , n37397 );
or ( n46673 , n46671 , n46672 );
buf ( n46674 , n42132 );
not ( n46675 , n46674 );
buf ( n46676 , n45099 );
nand ( n46677 , n46675 , n46676 );
buf ( n46678 , n46677 );
nand ( n46679 , n46673 , n46678 );
nand ( n46680 , n46656 , n46679 );
nand ( n46681 , n46655 , n46680 );
not ( n46682 , n46681 );
buf ( n46683 , n42847 );
not ( n46684 , n46683 );
buf ( n46685 , n43959 );
not ( n46686 , n46685 );
or ( n46687 , n46684 , n46686 );
buf ( n46688 , n36527 );
buf ( n46689 , n42847 );
not ( n46690 , n46689 );
buf ( n46691 , n46690 );
buf ( n46692 , n46691 );
nand ( n46693 , n46688 , n46692 );
buf ( n46694 , n46693 );
buf ( n46695 , n46694 );
nand ( n46696 , n46687 , n46695 );
buf ( n46697 , n46696 );
not ( n46698 , n46697 );
not ( n46699 , n44135 );
or ( n46700 , n46698 , n46699 );
nand ( n46701 , n43982 , n45544 );
nand ( n46702 , n46700 , n46701 );
not ( n46703 , n46702 );
or ( n46704 , n46682 , n46703 );
buf ( n46705 , n46681 );
not ( n46706 , n46705 );
buf ( n46707 , n46706 );
buf ( n46708 , n46707 );
not ( n46709 , n46708 );
not ( n46710 , n46702 );
buf ( n46711 , n46710 );
not ( n46712 , n46711 );
or ( n46713 , n46709 , n46712 );
xor ( n46714 , n45066 , n45086 );
xor ( n46715 , n46714 , n45115 );
buf ( n46716 , n46715 );
buf ( n46717 , n46716 );
nand ( n46718 , n46713 , n46717 );
buf ( n46719 , n46718 );
nand ( n46720 , n46704 , n46719 );
buf ( n46721 , n46720 );
xor ( n46722 , n46595 , n46721 );
buf ( n46723 , n44708 );
not ( n46724 , n46723 );
buf ( n46725 , n44533 );
not ( n46726 , n46725 );
buf ( n46727 , n42271 );
not ( n46728 , n46727 );
or ( n46729 , n46726 , n46728 );
buf ( n46730 , n36559 );
buf ( n46731 , n44530 );
nand ( n46732 , n46730 , n46731 );
buf ( n46733 , n46732 );
buf ( n46734 , n46733 );
nand ( n46735 , n46729 , n46734 );
buf ( n46736 , n46735 );
buf ( n46737 , n46736 );
not ( n46738 , n46737 );
or ( n46739 , n46724 , n46738 );
buf ( n46740 , n45660 );
buf ( n46741 , n44496 );
nand ( n46742 , n46740 , n46741 );
buf ( n46743 , n46742 );
buf ( n46744 , n46743 );
nand ( n46745 , n46739 , n46744 );
buf ( n46746 , n46745 );
buf ( n46747 , n46746 );
and ( n46748 , n46722 , n46747 );
and ( n46749 , n46595 , n46721 );
or ( n46750 , n46748 , n46749 );
buf ( n46751 , n46750 );
buf ( n46752 , n46751 );
xor ( n46753 , n45884 , n45939 );
xor ( n46754 , n46753 , n45965 );
buf ( n46755 , n46754 );
buf ( n46756 , n46755 );
xor ( n46757 , n46752 , n46756 );
xor ( n46758 , n45571 , n45596 );
xor ( n46759 , n46758 , n45625 );
buf ( n46760 , n46759 );
not ( n46761 , n46760 );
buf ( n46762 , n41647 );
not ( n46763 , n46762 );
buf ( n46764 , n45898 );
not ( n46765 , n46764 );
or ( n46766 , n46763 , n46765 );
buf ( n46767 , n41666 );
not ( n46768 , n46767 );
buf ( n46769 , n44316 );
not ( n46770 , n46769 );
or ( n46771 , n46768 , n46770 );
buf ( n46772 , n43198 );
buf ( n46773 , n41663 );
nand ( n46774 , n46772 , n46773 );
buf ( n46775 , n46774 );
buf ( n46776 , n46775 );
nand ( n46777 , n46771 , n46776 );
buf ( n46778 , n46777 );
buf ( n46779 , n46778 );
buf ( n46780 , n41705 );
nand ( n46781 , n46779 , n46780 );
buf ( n46782 , n46781 );
buf ( n46783 , n46782 );
nand ( n46784 , n46766 , n46783 );
buf ( n46785 , n46784 );
not ( n46786 , n46785 );
nand ( n46787 , n46761 , n46786 );
not ( n46788 , n46787 );
xor ( n46789 , n46085 , n46110 );
xor ( n46790 , n46789 , n46141 );
buf ( n46791 , n46790 );
not ( n46792 , n46791 );
or ( n46793 , n46788 , n46792 );
nand ( n46794 , n46785 , n46760 );
nand ( n46795 , n46793 , n46794 );
xor ( n46796 , n45933 , n45908 );
xor ( n46797 , n46796 , n45887 );
xor ( n46798 , n46795 , n46797 );
not ( n46799 , n44267 );
buf ( n46800 , n41608 );
not ( n46801 , n46800 );
buf ( n46802 , n43597 );
not ( n46803 , n46802 );
or ( n46804 , n46801 , n46803 );
buf ( n46805 , n36396 );
buf ( n46806 , n41611 );
nand ( n46807 , n46805 , n46806 );
buf ( n46808 , n46807 );
buf ( n46809 , n46808 );
nand ( n46810 , n46804 , n46809 );
buf ( n46811 , n46810 );
not ( n46812 , n46811 );
or ( n46813 , n46799 , n46812 );
buf ( n46814 , n45816 );
buf ( n46815 , n43868 );
nand ( n46816 , n46814 , n46815 );
buf ( n46817 , n46816 );
nand ( n46818 , n46813 , n46817 );
and ( n46819 , n46798 , n46818 );
and ( n46820 , n46795 , n46797 );
or ( n46821 , n46819 , n46820 );
buf ( n46822 , n46821 );
and ( n46823 , n46757 , n46822 );
and ( n46824 , n46752 , n46756 );
or ( n46825 , n46823 , n46824 );
buf ( n46826 , n46825 );
buf ( n46827 , n46826 );
and ( n46828 , n46577 , n46827 );
and ( n46829 , n46569 , n46576 );
or ( n46830 , n46828 , n46829 );
buf ( n46831 , n46830 );
buf ( n46832 , n46831 );
not ( n46833 , n46832 );
buf ( n46834 , n46833 );
nand ( n46835 , n46565 , n46834 );
not ( n46836 , n46835 );
xor ( n46837 , n46035 , n46273 );
xor ( n46838 , n46837 , n46520 );
buf ( n46839 , n46838 );
not ( n46840 , n46839 );
xor ( n46841 , n45856 , n45824 );
xnor ( n46842 , n46841 , n45864 );
buf ( n46843 , n46842 );
buf ( n46844 , n42339 );
not ( n46845 , n46844 );
buf ( n46846 , n46584 );
not ( n46847 , n46846 );
or ( n46848 , n46845 , n46847 );
buf ( n46849 , n42343 );
not ( n46850 , n46849 );
not ( n46851 , n37293 );
buf ( n46852 , n46851 );
not ( n46853 , n46852 );
or ( n46854 , n46850 , n46853 );
buf ( n46855 , n42342 );
buf ( n46856 , n46855 );
buf ( n46857 , n37293 );
nand ( n46858 , n46856 , n46857 );
buf ( n46859 , n46858 );
buf ( n46860 , n46859 );
nand ( n46861 , n46854 , n46860 );
buf ( n46862 , n46861 );
buf ( n46863 , n46862 );
buf ( n46864 , n42378 );
nand ( n46865 , n46863 , n46864 );
buf ( n46866 , n46865 );
buf ( n46867 , n46866 );
nand ( n46868 , n46848 , n46867 );
buf ( n46869 , n46868 );
not ( n46870 , n46869 );
buf ( n46871 , n46870 );
not ( n46872 , n46871 );
buf ( n46873 , n45723 );
buf ( n46874 , n46873 );
buf ( n46875 , n46874 );
buf ( n46876 , n46875 );
not ( n46877 , n46876 );
buf ( n46878 , n35968 );
not ( n46879 , n46878 );
buf ( n46880 , n46879 );
buf ( n46881 , n46880 );
not ( n46882 , n46881 );
or ( n46883 , n46877 , n46882 );
buf ( n46884 , n35968 );
buf ( n46885 , n46875 );
not ( n46886 , n46885 );
buf ( n46887 , n46886 );
buf ( n46888 , n46887 );
buf ( n46889 , n46888 );
buf ( n46890 , n46889 );
buf ( n46891 , n46890 );
nand ( n46892 , n46884 , n46891 );
buf ( n46893 , n46892 );
buf ( n46894 , n46893 );
nand ( n46895 , n46883 , n46894 );
buf ( n46896 , n46895 );
buf ( n46897 , n46896 );
xor ( n46898 , n24750 , n25431 );
and ( n46899 , n24750 , n24714 );
not ( n46900 , n24750 );
buf ( n46901 , n24714 );
not ( n46902 , n46901 );
buf ( n46903 , n46902 );
and ( n46904 , n46900 , n46903 );
or ( n46905 , n46899 , n46904 );
nand ( n46906 , n46898 , n46905 );
not ( n46907 , n46906 );
buf ( n46908 , n46907 );
not ( n46909 , n46908 );
buf ( n46910 , n46909 );
buf ( n46911 , n46910 );
not ( n46912 , n46905 );
buf ( n46913 , n46912 );
not ( n46914 , n46913 );
buf ( n46915 , n46914 );
buf ( n46916 , n46915 );
nand ( n46917 , n46911 , n46916 );
buf ( n46918 , n46917 );
buf ( n46919 , n46918 );
nand ( n46920 , n46897 , n46919 );
buf ( n46921 , n46920 );
buf ( n46922 , n46921 );
not ( n46923 , n46922 );
buf ( n46924 , n46923 );
buf ( n46925 , n46924 );
not ( n46926 , n46925 );
or ( n46927 , n46872 , n46926 );
buf ( n46928 , n46246 );
not ( n46929 , n46928 );
buf ( n46930 , n46239 );
not ( n46931 , n46930 );
or ( n46932 , n46929 , n46931 );
buf ( n46933 , n45753 );
not ( n46934 , n46933 );
buf ( n46935 , n45650 );
not ( n46936 , n46935 );
or ( n46937 , n46934 , n46936 );
buf ( n46938 , n36611 );
buf ( n46939 , n45750 );
nand ( n46940 , n46938 , n46939 );
buf ( n46941 , n46940 );
buf ( n46942 , n46941 );
nand ( n46943 , n46937 , n46942 );
buf ( n46944 , n46943 );
buf ( n46945 , n46944 );
buf ( n46946 , n46225 );
nand ( n46947 , n46945 , n46946 );
buf ( n46948 , n46947 );
buf ( n46949 , n46948 );
nand ( n46950 , n46932 , n46949 );
buf ( n46951 , n46950 );
buf ( n46952 , n46951 );
nand ( n46953 , n46927 , n46952 );
buf ( n46954 , n46953 );
buf ( n46955 , n46954 );
buf ( n46956 , n46921 );
buf ( n46957 , n46869 );
nand ( n46958 , n46956 , n46957 );
buf ( n46959 , n46958 );
buf ( n46960 , n46959 );
nand ( n46961 , n46955 , n46960 );
buf ( n46962 , n46961 );
buf ( n46963 , n46962 );
not ( n46964 , n46963 );
buf ( n46965 , n46145 );
buf ( n46966 , n46049 );
xor ( n46967 , n46965 , n46966 );
buf ( n46968 , n46059 );
xnor ( n46969 , n46967 , n46968 );
buf ( n46970 , n46969 );
buf ( n46971 , n46970 );
not ( n46972 , n46971 );
buf ( n46973 , n46972 );
buf ( n46974 , n46973 );
not ( n46975 , n46974 );
or ( n46976 , n46964 , n46975 );
buf ( n46977 , n46962 );
not ( n46978 , n46977 );
buf ( n46979 , n46978 );
not ( n46980 , n46979 );
not ( n46981 , n46970 );
or ( n46982 , n46980 , n46981 );
not ( n46983 , n42668 );
not ( n46984 , n46046 );
or ( n46985 , n46983 , n46984 );
and ( n46986 , n38244 , n42679 );
not ( n46987 , n38244 );
and ( n46988 , n46987 , n42672 );
or ( n46989 , n46986 , n46988 );
buf ( n46990 , n46989 );
buf ( n46991 , n42712 );
nand ( n46992 , n46990 , n46991 );
buf ( n46993 , n46992 );
nand ( n46994 , n46985 , n46993 );
buf ( n46995 , n38979 );
not ( n46996 , n46995 );
not ( n46997 , n29344 );
not ( n46998 , n29351 );
or ( n46999 , n46997 , n46998 );
nand ( n47000 , n46999 , n29357 );
not ( n47001 , n47000 );
buf ( n47002 , n47001 );
not ( n47003 , n47002 );
or ( n47004 , n46996 , n47003 );
buf ( n47005 , n29360 );
buf ( n47006 , n42471 );
nand ( n47007 , n47005 , n47006 );
buf ( n47008 , n47007 );
buf ( n47009 , n47008 );
nand ( n47010 , n47004 , n47009 );
buf ( n47011 , n47010 );
buf ( n47012 , n47011 );
not ( n47013 , n47012 );
and ( n47014 , n38972 , n38980 , n38981 );
buf ( n47015 , n47014 );
not ( n47016 , n47015 );
or ( n47017 , n47013 , n47016 );
not ( n47018 , n38972 );
not ( n47019 , n47018 );
buf ( n47020 , n47019 );
buf ( n47021 , n47020 );
not ( n47022 , n47021 );
buf ( n47023 , n38979 );
not ( n47024 , n47023 );
buf ( n47025 , n41951 );
not ( n47026 , n47025 );
or ( n47027 , n47024 , n47026 );
buf ( n47028 , n41821 );
buf ( n47029 , n38979 );
not ( n47030 , n47029 );
buf ( n47031 , n47030 );
buf ( n47032 , n47031 );
nand ( n47033 , n47028 , n47032 );
buf ( n47034 , n47033 );
buf ( n47035 , n47034 );
nand ( n47036 , n47027 , n47035 );
buf ( n47037 , n47036 );
buf ( n47038 , n47037 );
nand ( n47039 , n47022 , n47038 );
buf ( n47040 , n47039 );
buf ( n47041 , n47040 );
nand ( n47042 , n47017 , n47041 );
buf ( n47043 , n47042 );
buf ( n47044 , n47043 );
not ( n47045 , n45565 );
not ( n47046 , n42448 );
or ( n47047 , n47045 , n47046 );
buf ( n47048 , n45053 );
not ( n47049 , n47048 );
buf ( n47050 , n47049 );
buf ( n47051 , n47050 );
buf ( n47052 , n47037 );
nand ( n47053 , n47051 , n47052 );
buf ( n47054 , n47053 );
nand ( n47055 , n47047 , n47054 );
buf ( n47056 , n47055 );
xor ( n47057 , n47044 , n47056 );
not ( n47058 , n46627 );
not ( n47059 , n38380 );
or ( n47060 , n47058 , n47059 );
buf ( n47061 , n41873 );
not ( n47062 , n47061 );
buf ( n47063 , n47062 );
buf ( n47064 , n47063 );
not ( n47065 , n47064 );
buf ( n47066 , n38411 );
not ( n47067 , n47066 );
buf ( n47068 , n47067 );
buf ( n47069 , n47068 );
nor ( n47070 , n47065 , n47069 );
buf ( n47071 , n47070 );
not ( n47072 , n29380 );
and ( n47073 , n46623 , n47072 );
nor ( n47074 , n47071 , n47073 );
or ( n47075 , n47074 , n44039 );
nand ( n47076 , n47060 , n47075 );
buf ( n47077 , n47076 );
and ( n47078 , n47057 , n47077 );
and ( n47079 , n47044 , n47056 );
or ( n47080 , n47078 , n47079 );
buf ( n47081 , n47080 );
buf ( n47082 , n42504 );
not ( n47083 , n47082 );
buf ( n47084 , n43371 );
not ( n47085 , n47084 );
or ( n47086 , n47083 , n47085 );
buf ( n47087 , n45376 );
buf ( n47088 , n41721 );
nand ( n47089 , n47087 , n47088 );
buf ( n47090 , n47089 );
buf ( n47091 , n47090 );
nand ( n47092 , n47086 , n47091 );
buf ( n47093 , n47092 );
buf ( n47094 , n47093 );
not ( n47095 , n47094 );
buf ( n47096 , n43386 );
not ( n47097 , n47096 );
buf ( n47098 , n47097 );
buf ( n47099 , n47098 );
not ( n47100 , n47099 );
buf ( n47101 , n47100 );
buf ( n47102 , n47101 );
not ( n47103 , n47102 );
or ( n47104 , n47095 , n47103 );
buf ( n47105 , n46160 );
buf ( n47106 , n45141 );
not ( n47107 , n47106 );
buf ( n47108 , n47107 );
buf ( n47109 , n47108 );
nand ( n47110 , n47105 , n47109 );
buf ( n47111 , n47110 );
buf ( n47112 , n47111 );
nand ( n47113 , n47104 , n47112 );
buf ( n47114 , n47113 );
xor ( n47115 , n47081 , n47114 );
not ( n47116 , n44586 );
buf ( n47117 , n25184 );
not ( n47118 , n47117 );
not ( n47119 , n37641 );
buf ( n47120 , n47119 );
not ( n47121 , n47120 );
or ( n47122 , n47118 , n47121 );
buf ( n47123 , n39205 );
buf ( n47124 , n25183 );
nand ( n47125 , n47123 , n47124 );
buf ( n47126 , n47125 );
buf ( n47127 , n47126 );
nand ( n47128 , n47122 , n47127 );
buf ( n47129 , n47128 );
not ( n47130 , n47129 );
or ( n47131 , n47116 , n47130 );
nand ( n47132 , n43909 , n46311 );
nand ( n47133 , n47131 , n47132 );
and ( n47134 , n47115 , n47133 );
and ( n47135 , n47081 , n47114 );
or ( n47136 , n47134 , n47135 );
xor ( n47137 , n46994 , n47136 );
buf ( n47138 , n46209 );
buf ( n47139 , n46178 );
not ( n47140 , n47139 );
buf ( n47141 , n46190 );
not ( n47142 , n47141 );
or ( n47143 , n47140 , n47142 );
buf ( n47144 , n46216 );
buf ( n47145 , n46181 );
nand ( n47146 , n47144 , n47145 );
buf ( n47147 , n47146 );
buf ( n47148 , n47147 );
nand ( n47149 , n47143 , n47148 );
buf ( n47150 , n47149 );
buf ( n47151 , n47150 );
xor ( n47152 , n47138 , n47151 );
buf ( n47153 , n47152 );
and ( n47154 , n47137 , n47153 );
and ( n47155 , n46994 , n47136 );
or ( n47156 , n47154 , n47155 );
buf ( n47157 , n47156 );
nand ( n47158 , n46982 , n47157 );
buf ( n47159 , n47158 );
nand ( n47160 , n46976 , n47159 );
buf ( n47161 , n47160 );
buf ( n47162 , n47161 );
xor ( n47163 , n46843 , n47162 );
xor ( n47164 , n46148 , n46263 );
xor ( n47165 , n47164 , n46268 );
buf ( n47166 , n47165 );
buf ( n47167 , n47166 );
and ( n47168 , n47163 , n47167 );
and ( n47169 , n46843 , n47162 );
or ( n47170 , n47168 , n47169 );
buf ( n47171 , n47170 );
buf ( n47172 , n47171 );
not ( n47173 , n47172 );
buf ( n47174 , n47173 );
buf ( n47175 , n47174 );
and ( n47176 , n45969 , n45870 );
not ( n47177 , n45969 );
buf ( n47178 , n45870 );
not ( n47179 , n47178 );
buf ( n47180 , n47179 );
and ( n47181 , n47177 , n47180 );
or ( n47182 , n47176 , n47181 );
buf ( n47183 , n45874 );
xor ( n47184 , n47182 , n47183 );
buf ( n47185 , n47184 );
nand ( n47186 , n47175 , n47185 );
buf ( n47187 , n47186 );
not ( n47188 , n47187 );
or ( n47189 , n46840 , n47188 );
buf ( n47190 , n47171 );
buf ( n47191 , n47184 );
not ( n47192 , n47191 );
buf ( n47193 , n47192 );
buf ( n47194 , n47193 );
nand ( n47195 , n47190 , n47194 );
buf ( n47196 , n47195 );
nand ( n47197 , n47189 , n47196 );
not ( n47198 , n47197 );
or ( n47199 , n46836 , n47198 );
not ( n47200 , n46565 );
nand ( n47201 , n47200 , n46831 );
nand ( n47202 , n47199 , n47201 );
buf ( n47203 , n47202 );
not ( n47204 , n47203 );
buf ( n47205 , n47204 );
buf ( n47206 , n47205 );
xor ( n47207 , n46550 , n47206 );
buf ( n47208 , n45994 );
buf ( n47209 , n46002 );
and ( n47210 , n47208 , n47209 );
not ( n47211 , n47208 );
buf ( n47212 , n45999 );
and ( n47213 , n47211 , n47212 );
nor ( n47214 , n47210 , n47213 );
buf ( n47215 , n47214 );
xor ( n47216 , n47215 , n46530 );
buf ( n47217 , n47216 );
and ( n47218 , n47207 , n47217 );
and ( n47219 , n46550 , n47206 );
or ( n47220 , n47218 , n47219 );
buf ( n47221 , n47220 );
buf ( n47222 , n47221 );
nand ( n47223 , n46539 , n47222 );
buf ( n47224 , n47223 );
buf ( n47225 , n47224 );
xor ( n47226 , n46550 , n47206 );
xor ( n47227 , n47226 , n47217 );
buf ( n47228 , n47227 );
buf ( n47229 , n47228 );
buf ( n47230 , n46009 );
buf ( n47231 , n46524 );
xor ( n47232 , n47230 , n47231 );
buf ( n47233 , n46020 );
xnor ( n47234 , n47232 , n47233 );
buf ( n47235 , n47234 );
xor ( n47236 , n46752 , n46756 );
xor ( n47237 , n47236 , n46822 );
buf ( n47238 , n47237 );
buf ( n47239 , n47238 );
not ( n47240 , n47239 );
xor ( n47241 , n46843 , n47162 );
xor ( n47242 , n47241 , n47167 );
buf ( n47243 , n47242 );
buf ( n47244 , n47243 );
not ( n47245 , n47244 );
or ( n47246 , n47240 , n47245 );
buf ( n47247 , n47243 );
buf ( n47248 , n47238 );
or ( n47249 , n47247 , n47248 );
xor ( n47250 , n46795 , n46797 );
xor ( n47251 , n47250 , n46818 );
buf ( n47252 , n47251 );
not ( n47253 , n47252 );
xor ( n47254 , n46962 , n47156 );
xnor ( n47255 , n47254 , n46970 );
buf ( n47256 , n47255 );
not ( n47257 , n47256 );
or ( n47258 , n47253 , n47257 );
not ( n47259 , n47251 );
not ( n47260 , n47259 );
or ( n47261 , n47260 , n47255 );
xor ( n47262 , n46994 , n47136 );
xor ( n47263 , n47262 , n47153 );
not ( n47264 , n47263 );
buf ( n47265 , n46408 );
buf ( n47266 , n46351 );
buf ( n47267 , n46374 );
and ( n47268 , n47266 , n47267 );
not ( n47269 , n47266 );
buf ( n47270 , n46377 );
and ( n47271 , n47269 , n47270 );
nor ( n47272 , n47268 , n47271 );
buf ( n47273 , n47272 );
buf ( n47274 , n47273 );
xor ( n47275 , n47265 , n47274 );
buf ( n47276 , n47275 );
buf ( n47277 , n47276 );
buf ( n47278 , n45570 );
buf ( n47279 , n46438 );
xor ( n47280 , n47278 , n47279 );
buf ( n47281 , n46465 );
xnor ( n47282 , n47280 , n47281 );
buf ( n47283 , n47282 );
buf ( n47284 , n47283 );
xor ( n47285 , n47277 , n47284 );
buf ( n47286 , n42339 );
not ( n47287 , n47286 );
buf ( n47288 , n46862 );
not ( n47289 , n47288 );
or ( n47290 , n47287 , n47289 );
buf ( n47291 , n42343 );
not ( n47292 , n47291 );
buf ( n47293 , n42573 );
not ( n47294 , n47293 );
or ( n47295 , n47292 , n47294 );
buf ( n47296 , n37683 );
buf ( n47297 , n46855 );
nand ( n47298 , n47296 , n47297 );
buf ( n47299 , n47298 );
buf ( n47300 , n47299 );
nand ( n47301 , n47295 , n47300 );
buf ( n47302 , n47301 );
buf ( n47303 , n47302 );
buf ( n47304 , n42378 );
nand ( n47305 , n47303 , n47304 );
buf ( n47306 , n47305 );
buf ( n47307 , n47306 );
nand ( n47308 , n47290 , n47307 );
buf ( n47309 , n47308 );
buf ( n47310 , n47309 );
and ( n47311 , n47285 , n47310 );
and ( n47312 , n47277 , n47284 );
or ( n47313 , n47311 , n47312 );
buf ( n47314 , n47313 );
not ( n47315 , n47314 );
or ( n47316 , n47264 , n47315 );
or ( n47317 , n47263 , n47314 );
not ( n47318 , n42672 );
not ( n47319 , n38743 );
not ( n47320 , n47319 );
or ( n47321 , n47318 , n47320 );
nand ( n47322 , n42679 , n38743 );
nand ( n47323 , n47321 , n47322 );
and ( n47324 , n47323 , n42712 );
and ( n47325 , n46989 , n42668 );
nor ( n47326 , n47324 , n47325 );
not ( n47327 , n47326 );
not ( n47328 , n47327 );
buf ( n47329 , n46910 );
not ( n47330 , n47329 );
buf ( n47331 , n47330 );
buf ( n47332 , n47331 );
not ( n47333 , n47332 );
buf ( n47334 , n46875 );
not ( n47335 , n47334 );
buf ( n47336 , n36032 );
not ( n47337 , n47336 );
or ( n47338 , n47335 , n47337 );
buf ( n47339 , n43851 );
buf ( n47340 , n46890 );
nand ( n47341 , n47339 , n47340 );
buf ( n47342 , n47341 );
buf ( n47343 , n47342 );
nand ( n47344 , n47338 , n47343 );
buf ( n47345 , n47344 );
buf ( n47346 , n47345 );
not ( n47347 , n47346 );
or ( n47348 , n47333 , n47347 );
buf ( n47349 , n46896 );
buf ( n47350 , n46912 );
nand ( n47351 , n47349 , n47350 );
buf ( n47352 , n47351 );
buf ( n47353 , n47352 );
nand ( n47354 , n47348 , n47353 );
buf ( n47355 , n47354 );
not ( n47356 , n47355 );
or ( n47357 , n47328 , n47356 );
or ( n47358 , n47355 , n47327 );
xor ( n47359 , n47081 , n47114 );
xor ( n47360 , n47359 , n47133 );
buf ( n47361 , n47360 );
nand ( n47362 , n47358 , n47361 );
nand ( n47363 , n47357 , n47362 );
nand ( n47364 , n47317 , n47363 );
nand ( n47365 , n47316 , n47364 );
buf ( n47366 , n47365 );
nand ( n47367 , n47261 , n47366 );
buf ( n47368 , n47367 );
nand ( n47369 , n47258 , n47368 );
buf ( n47370 , n47369 );
buf ( n47371 , n47370 );
nand ( n47372 , n47249 , n47371 );
buf ( n47373 , n47372 );
buf ( n47374 , n47373 );
nand ( n47375 , n47246 , n47374 );
buf ( n47376 , n47375 );
not ( n47377 , n47376 );
xor ( n47378 , n46569 , n46576 );
xor ( n47379 , n47378 , n46827 );
buf ( n47380 , n47379 );
buf ( n47381 , n47380 );
not ( n47382 , n47381 );
buf ( n47383 , n47382 );
buf ( n47384 , n47383 );
xor ( n47385 , n46595 , n46721 );
xor ( n47386 , n47385 , n46747 );
buf ( n47387 , n47386 );
buf ( n47388 , n47387 );
buf ( n47389 , n41993 );
buf ( n47390 , n36926 );
and ( n47391 , n47389 , n47390 );
not ( n47392 , n47389 );
buf ( n47393 , n42062 );
and ( n47394 , n47392 , n47393 );
nor ( n47395 , n47391 , n47394 );
buf ( n47396 , n47395 );
buf ( n47397 , n47396 );
not ( n47398 , n47397 );
buf ( n47399 , n47398 );
buf ( n47400 , n47399 );
not ( n47401 , n47400 );
buf ( n47402 , n44776 );
not ( n47403 , n47402 );
or ( n47404 , n47401 , n47403 );
buf ( n47405 , n46202 );
not ( n47406 , n47405 );
buf ( n47407 , n36909 );
not ( n47408 , n47407 );
buf ( n47409 , n47408 );
buf ( n47410 , n47409 );
nand ( n47411 , n47406 , n47410 );
buf ( n47412 , n47411 );
buf ( n47413 , n47412 );
nand ( n47414 , n47404 , n47413 );
buf ( n47415 , n47414 );
buf ( n47416 , n47415 );
xor ( n47417 , n46629 , n46653 );
and ( n47418 , n47417 , n46679 );
not ( n47419 , n47417 );
not ( n47420 , n46679 );
and ( n47421 , n47419 , n47420 );
nor ( n47422 , n47418 , n47421 );
buf ( n47423 , n47422 );
or ( n47424 , n47416 , n47423 );
buf ( n47425 , n47424 );
buf ( n47426 , n47425 );
buf ( n47427 , n41778 );
not ( n47428 , n47427 );
buf ( n47429 , n47428 );
not ( n47430 , n47429 );
not ( n47431 , n29399 );
nand ( n47432 , n47431 , n29394 );
not ( n47433 , n29394 );
nand ( n47434 , n47433 , n29399 );
nand ( n47435 , n47432 , n47434 );
not ( n47436 , n47435 );
not ( n47437 , n47436 );
or ( n47438 , n47430 , n47437 );
buf ( n47439 , n29407 );
nand ( n47440 , n47439 , n37328 );
nand ( n47441 , n47438 , n47440 );
buf ( n47442 , n47441 );
not ( n47443 , n47442 );
buf ( n47444 , n37394 );
not ( n47445 , n47444 );
or ( n47446 , n47443 , n47445 );
buf ( n47447 , n46670 );
buf ( n47448 , n37410 );
nand ( n47449 , n47447 , n47448 );
buf ( n47450 , n47449 );
buf ( n47451 , n47450 );
nand ( n47452 , n47446 , n47451 );
buf ( n47453 , n47452 );
buf ( n47454 , n47453 );
not ( n47455 , n47454 );
buf ( n47456 , n47455 );
not ( n47457 , n47456 );
buf ( n47458 , n39983 );
not ( n47459 , n47458 );
buf ( n47460 , n46651 );
not ( n47461 , n47460 );
or ( n47462 , n47459 , n47461 );
buf ( n47463 , n28721 );
not ( n47464 , n47463 );
buf ( n47465 , n40009 );
not ( n47466 , n47465 );
and ( n47467 , n47464 , n47466 );
buf ( n47468 , n41782 );
not ( n47469 , n24092 );
buf ( n47470 , n47469 );
and ( n47471 , n47468 , n47470 );
nor ( n47472 , n47467 , n47471 );
buf ( n47473 , n47472 );
buf ( n47474 , n47473 );
not ( n47475 , n47474 );
buf ( n47476 , n40002 );
nand ( n47477 , n47475 , n47476 );
buf ( n47478 , n47477 );
buf ( n47479 , n47478 );
nand ( n47480 , n47462 , n47479 );
buf ( n47481 , n47480 );
buf ( n47482 , n47481 );
buf ( n47483 , n47482 );
buf ( n47484 , n47483 );
nor ( n47485 , n47457 , n47484 );
not ( n47486 , n37499 );
not ( n47487 , n37502 );
or ( n47488 , n47486 , n47487 );
nand ( n47489 , n47488 , n37505 );
nand ( n47490 , n47489 , n37509 );
buf ( n47491 , n47490 );
not ( n47492 , n47491 );
buf ( n47493 , n42052 );
buf ( n47494 , n41981 );
and ( n47495 , n47493 , n47494 );
not ( n47496 , n47493 );
buf ( n47497 , n41977 );
and ( n47498 , n47496 , n47497 );
nor ( n47499 , n47495 , n47498 );
buf ( n47500 , n47499 );
buf ( n47501 , n47500 );
not ( n47502 , n47501 );
and ( n47503 , n47492 , n47502 );
buf ( n47504 , n46455 );
buf ( n47505 , n37443 );
nor ( n47506 , n47504 , n47505 );
buf ( n47507 , n47506 );
buf ( n47508 , n47507 );
nor ( n47509 , n47503 , n47508 );
buf ( n47510 , n47509 );
or ( n47511 , n47485 , n47510 );
buf ( n47512 , n47453 );
buf ( n47513 , n47484 );
nand ( n47514 , n47512 , n47513 );
buf ( n47515 , n47514 );
nand ( n47516 , n47511 , n47515 );
buf ( n47517 , n47516 );
and ( n47518 , n47426 , n47517 );
buf ( n47519 , n47422 );
buf ( n47520 , n47415 );
and ( n47521 , n47519 , n47520 );
buf ( n47522 , n47521 );
buf ( n47523 , n47522 );
nor ( n47524 , n47518 , n47523 );
buf ( n47525 , n47524 );
buf ( n47526 , n47525 );
not ( n47527 , n47526 );
buf ( n47528 , n42315 );
not ( n47529 , n47528 );
buf ( n47530 , n46280 );
not ( n47531 , n47530 );
or ( n47532 , n47529 , n47531 );
buf ( n47533 , n42266 );
not ( n47534 , n47533 );
buf ( n47535 , n42926 );
not ( n47536 , n47535 );
or ( n47537 , n47534 , n47536 );
buf ( n47538 , n39277 );
buf ( n47539 , n42263 );
nand ( n47540 , n47538 , n47539 );
buf ( n47541 , n47540 );
buf ( n47542 , n47541 );
nand ( n47543 , n47537 , n47542 );
buf ( n47544 , n47543 );
buf ( n47545 , n47544 );
buf ( n47546 , n42252 );
nand ( n47547 , n47545 , n47546 );
buf ( n47548 , n47547 );
buf ( n47549 , n47548 );
nand ( n47550 , n47532 , n47549 );
buf ( n47551 , n47550 );
buf ( n47552 , n47551 );
not ( n47553 , n47552 );
buf ( n47554 , n47553 );
buf ( n47555 , n47554 );
not ( n47556 , n47555 );
or ( n47557 , n47527 , n47556 );
not ( n47558 , n46702 );
not ( n47559 , n46681 );
or ( n47560 , n47558 , n47559 );
nand ( n47561 , n46707 , n46710 );
nand ( n47562 , n47560 , n47561 );
not ( n47563 , n46716 );
and ( n47564 , n47562 , n47563 );
not ( n47565 , n47562 );
and ( n47566 , n47565 , n46716 );
nor ( n47567 , n47564 , n47566 );
buf ( n47568 , n47567 );
nand ( n47569 , n47557 , n47568 );
buf ( n47570 , n47569 );
buf ( n47571 , n47570 );
buf ( n47572 , n47525 );
not ( n47573 , n47572 );
buf ( n47574 , n47551 );
nand ( n47575 , n47573 , n47574 );
buf ( n47576 , n47575 );
buf ( n47577 , n47576 );
nand ( n47578 , n47571 , n47577 );
buf ( n47579 , n47578 );
buf ( n47580 , n47579 );
xor ( n47581 , n47388 , n47580 );
xor ( n47582 , n46224 , n46253 );
xor ( n47583 , n47582 , n46258 );
buf ( n47584 , n47583 );
buf ( n47585 , n47584 );
and ( n47586 , n47581 , n47585 );
and ( n47587 , n47388 , n47580 );
or ( n47588 , n47586 , n47587 );
buf ( n47589 , n47588 );
not ( n47590 , n47589 );
xor ( n47591 , n46503 , n46510 );
xor ( n47592 , n47591 , n46515 );
buf ( n47593 , n47592 );
not ( n47594 , n47593 );
xor ( n47595 , n46291 , n46493 );
xor ( n47596 , n47595 , n46498 );
buf ( n47597 , n47596 );
buf ( n47598 , n47597 );
buf ( n47599 , n44952 );
not ( n47600 , n47599 );
buf ( n47601 , n41718 );
not ( n47602 , n47601 );
or ( n47603 , n47600 , n47602 );
buf ( n47604 , n39726 );
not ( n47605 , n47604 );
buf ( n47606 , n44961 );
nand ( n47607 , n47605 , n47606 );
buf ( n47608 , n47607 );
buf ( n47609 , n47608 );
nand ( n47610 , n47603 , n47609 );
buf ( n47611 , n47610 );
not ( n47612 , n47611 );
not ( n47613 , n39803 );
or ( n47614 , n47612 , n47613 );
buf ( n47615 , n43982 );
buf ( n47616 , n46697 );
nand ( n47617 , n47615 , n47616 );
buf ( n47618 , n47617 );
nand ( n47619 , n47614 , n47618 );
buf ( n47620 , n47619 );
buf ( n47621 , n41705 );
not ( n47622 , n47621 );
buf ( n47623 , n41660 );
buf ( n47624 , n38477 );
not ( n47625 , n47624 );
buf ( n47626 , n47625 );
buf ( n47627 , n47626 );
and ( n47628 , n47623 , n47627 );
not ( n47629 , n47623 );
buf ( n47630 , n45916 );
and ( n47631 , n47629 , n47630 );
nor ( n47632 , n47628 , n47631 );
buf ( n47633 , n47632 );
buf ( n47634 , n47633 );
not ( n47635 , n47634 );
or ( n47636 , n47622 , n47635 );
buf ( n47637 , n46778 );
buf ( n47638 , n41644 );
not ( n47639 , n47638 );
buf ( n47640 , n47639 );
buf ( n47641 , n47640 );
nand ( n47642 , n47637 , n47641 );
buf ( n47643 , n47642 );
buf ( n47644 , n47643 );
nand ( n47645 , n47636 , n47644 );
buf ( n47646 , n47645 );
buf ( n47647 , n47646 );
xor ( n47648 , n47620 , n47647 );
buf ( n47649 , n42566 );
not ( n47650 , n47649 );
buf ( n47651 , n46364 );
not ( n47652 , n47651 );
or ( n47653 , n47650 , n47652 );
not ( n47654 , n25159 );
and ( n47655 , n29263 , n47654 );
not ( n47656 , n29263 );
not ( n47657 , n46356 );
and ( n47658 , n47656 , n47657 );
or ( n47659 , n47655 , n47658 );
and ( n47660 , n29018 , n47659 );
not ( n47661 , n29018 );
not ( n47662 , n25159 );
and ( n47663 , n29266 , n47662 );
not ( n47664 , n29266 );
not ( n47665 , n46356 );
and ( n47666 , n47664 , n47665 );
or ( n47667 , n47663 , n47666 );
and ( n47668 , n47661 , n47667 );
or ( n47669 , n47660 , n47668 );
buf ( n47670 , n47669 );
not ( n47671 , n47670 );
buf ( n47672 , n42631 );
nand ( n47673 , n47671 , n47672 );
buf ( n47674 , n47673 );
buf ( n47675 , n47674 );
nand ( n47676 , n47653 , n47675 );
buf ( n47677 , n47676 );
buf ( n47678 , n47677 );
not ( n47679 , n47678 );
buf ( n47680 , n41736 );
not ( n47681 , n47680 );
buf ( n47682 , n41890 );
not ( n47683 , n47682 );
or ( n47684 , n47681 , n47683 );
buf ( n47685 , n41889 );
buf ( n47686 , n41748 );
nand ( n47687 , n47685 , n47686 );
buf ( n47688 , n47687 );
buf ( n47689 , n47688 );
nand ( n47690 , n47684 , n47689 );
buf ( n47691 , n47690 );
buf ( n47692 , n47691 );
not ( n47693 , n47692 );
buf ( n47694 , n41862 );
not ( n47695 , n47694 );
or ( n47696 , n47693 , n47695 );
buf ( n47697 , n37919 );
buf ( n47698 , n46433 );
nand ( n47699 , n47697 , n47698 );
buf ( n47700 , n47699 );
buf ( n47701 , n47700 );
nand ( n47702 , n47696 , n47701 );
buf ( n47703 , n47702 );
buf ( n47704 , n47703 );
not ( n47705 , n47704 );
buf ( n47706 , n47705 );
buf ( n47707 , n47706 );
nand ( n47708 , n47679 , n47707 );
buf ( n47709 , n47708 );
not ( n47710 , n47709 );
buf ( n47711 , n25938 );
not ( n47712 , n47711 );
buf ( n47713 , n47712 );
buf ( n47714 , n47713 );
not ( n47715 , n47714 );
buf ( n47716 , n47715 );
buf ( n47717 , n47716 );
not ( n47718 , n47717 );
buf ( n47719 , n37649 );
not ( n47720 , n47719 );
or ( n47721 , n47718 , n47720 );
buf ( n47722 , n38834 );
buf ( n47723 , n47716 );
not ( n47724 , n47723 );
buf ( n47725 , n47724 );
buf ( n47726 , n47725 );
nand ( n47727 , n47722 , n47726 );
buf ( n47728 , n47727 );
buf ( n47729 , n47728 );
nand ( n47730 , n47721 , n47729 );
buf ( n47731 , n47730 );
or ( n47732 , n36447 , n46401 );
nand ( n47733 , C1 , n47732 );
not ( n47734 , n47733 );
or ( n47735 , n47710 , n47734 );
buf ( n47736 , n47703 );
buf ( n47737 , n47677 );
nand ( n47738 , n47736 , n47737 );
buf ( n47739 , n47738 );
nand ( n47740 , n47735 , n47739 );
buf ( n47741 , n47740 );
and ( n47742 , n47648 , n47741 );
and ( n47743 , n47620 , n47647 );
or ( n47744 , n47742 , n47743 );
buf ( n47745 , n47744 );
buf ( n47746 , n47745 );
not ( n47747 , n46417 );
not ( n47748 , n47747 );
and ( n47749 , n46318 , n46478 );
not ( n47750 , n46318 );
and ( n47751 , n47750 , n46477 );
nor ( n47752 , n47749 , n47751 );
not ( n47753 , n47752 );
or ( n47754 , n47748 , n47753 );
or ( n47755 , n47752 , n47747 );
nand ( n47756 , n47754 , n47755 );
buf ( n47757 , n47756 );
xor ( n47758 , n47746 , n47757 );
not ( n47759 , n46785 );
not ( n47760 , n46761 );
or ( n47761 , n47759 , n47760 );
nand ( n47762 , n46760 , n46786 );
nand ( n47763 , n47761 , n47762 );
and ( n47764 , n47763 , n46791 );
not ( n47765 , n47763 );
not ( n47766 , n46791 );
and ( n47767 , n47765 , n47766 );
nor ( n47768 , n47764 , n47767 );
buf ( n47769 , n47768 );
and ( n47770 , n47758 , n47769 );
and ( n47771 , n47746 , n47757 );
or ( n47772 , n47770 , n47771 );
buf ( n47773 , n47772 );
buf ( n47774 , n47773 );
xor ( n47775 , n47598 , n47774 );
buf ( n47776 , n44708 );
not ( n47777 , n47776 );
buf ( n47778 , n44533 );
not ( n47779 , n47778 );
buf ( n47780 , n40067 );
not ( n47781 , n47780 );
or ( n47782 , n47779 , n47781 );
buf ( n47783 , n36427 );
buf ( n47784 , n44530 );
nand ( n47785 , n47783 , n47784 );
buf ( n47786 , n47785 );
buf ( n47787 , n47786 );
nand ( n47788 , n47782 , n47787 );
buf ( n47789 , n47788 );
buf ( n47790 , n47789 );
not ( n47791 , n47790 );
or ( n47792 , n47777 , n47791 );
buf ( n47793 , n46736 );
buf ( n47794 , n44496 );
nand ( n47795 , n47793 , n47794 );
buf ( n47796 , n47795 );
buf ( n47797 , n47796 );
nand ( n47798 , n47792 , n47797 );
buf ( n47799 , n47798 );
buf ( n47800 , n47799 );
buf ( n47801 , n43868 );
not ( n47802 , n47801 );
buf ( n47803 , n46811 );
not ( n47804 , n47803 );
or ( n47805 , n47802 , n47804 );
buf ( n47806 , n41608 );
not ( n47807 , n47806 );
buf ( n47808 , n38098 );
not ( n47809 , n47808 );
or ( n47810 , n47807 , n47809 );
buf ( n47811 , n37078 );
not ( n47812 , n47811 );
buf ( n47813 , n47812 );
buf ( n47814 , n47813 );
not ( n47815 , n47814 );
buf ( n47816 , n41611 );
nand ( n47817 , n47815 , n47816 );
buf ( n47818 , n47817 );
buf ( n47819 , n47818 );
nand ( n47820 , n47810 , n47819 );
buf ( n47821 , n47820 );
buf ( n47822 , n47821 );
buf ( n47823 , n44267 );
nand ( n47824 , n47822 , n47823 );
buf ( n47825 , n47824 );
buf ( n47826 , n47825 );
nand ( n47827 , n47805 , n47826 );
buf ( n47828 , n47827 );
buf ( n47829 , n47828 );
xor ( n47830 , n47800 , n47829 );
not ( n47831 , n47074 );
not ( n47832 , n38379 );
and ( n47833 , n47831 , n47832 );
buf ( n47834 , n46660 );
not ( n47835 , n47834 );
buf ( n47836 , n47835 );
buf ( n47837 , n47836 );
buf ( n47838 , n44054 );
and ( n47839 , n47837 , n47838 );
not ( n47840 , n47837 );
buf ( n47841 , n46623 );
and ( n47842 , n47840 , n47841 );
or ( n47843 , n47839 , n47842 );
buf ( n47844 , n47843 );
not ( n47845 , n47844 );
and ( n47846 , n44042 , n47845 );
nor ( n47847 , n47833 , n47846 );
not ( n47848 , n47847 );
not ( n47849 , n47848 );
or ( n47850 , n47473 , n39980 );
buf ( n47851 , n24092 );
not ( n47852 , n47851 );
buf ( n47853 , n44025 );
not ( n47854 , n47853 );
or ( n47855 , n47852 , n47854 );
buf ( n47856 , n28305 );
not ( n47857 , n24092 );
buf ( n47858 , n47857 );
nand ( n47859 , n47856 , n47858 );
buf ( n47860 , n47859 );
buf ( n47861 , n47860 );
nand ( n47862 , n47855 , n47861 );
buf ( n47863 , n47862 );
nand ( n47864 , n47863 , n39999 );
nand ( n47865 , n47850 , n47864 );
not ( n47866 , n47865 );
or ( n47867 , n47849 , n47866 );
not ( n47868 , n47865 );
not ( n47869 , n47868 );
not ( n47870 , n47847 );
or ( n47871 , n47869 , n47870 );
not ( n47872 , n42563 );
not ( n47873 , n47872 );
not ( n47874 , n47669 );
not ( n47875 , n47874 );
or ( n47876 , n47873 , n47875 );
buf ( n47877 , n25160 );
not ( n47878 , n47877 );
buf ( n47879 , n46641 );
not ( n47880 , n47879 );
or ( n47881 , n47878 , n47880 );
buf ( n47882 , n29287 );
buf ( n47883 , n46356 );
nand ( n47884 , n47882 , n47883 );
buf ( n47885 , n47884 );
buf ( n47886 , n47885 );
nand ( n47887 , n47881 , n47886 );
buf ( n47888 , n47887 );
nand ( n47889 , n47888 , n42628 );
nand ( n47890 , n47876 , n47889 );
nand ( n47891 , n47871 , n47890 );
nand ( n47892 , n47867 , n47891 );
buf ( n47893 , n47892 );
buf ( n47894 , n42008 );
not ( n47895 , n47894 );
buf ( n47896 , n43400 );
not ( n47897 , n47896 );
buf ( n47898 , n47897 );
buf ( n47899 , n47898 );
not ( n47900 , n47899 );
or ( n47901 , n47895 , n47900 );
buf ( n47902 , n45376 );
buf ( n47903 , n42017 );
nand ( n47904 , n47902 , n47903 );
buf ( n47905 , n47904 );
buf ( n47906 , n47905 );
nand ( n47907 , n47901 , n47906 );
buf ( n47908 , n47907 );
buf ( n47909 , n47908 );
not ( n47910 , n47909 );
buf ( n47911 , n43386 );
not ( n47912 , n47911 );
or ( n47913 , n47910 , n47912 );
buf ( n47914 , n45144 );
buf ( n47915 , n47093 );
nand ( n47916 , n47914 , n47915 );
buf ( n47917 , n47916 );
buf ( n47918 , n47917 );
nand ( n47919 , n47913 , n47918 );
buf ( n47920 , n47919 );
buf ( n47921 , n47920 );
xor ( n47922 , n47893 , n47921 );
buf ( n47923 , n46294 );
not ( n47924 , n47923 );
buf ( n47925 , n47129 );
not ( n47926 , n47925 );
or ( n47927 , n47924 , n47926 );
buf ( n47928 , n25182 );
not ( n47929 , n47928 );
buf ( n47930 , n38821 );
not ( n47931 , n47930 );
buf ( n47932 , n47931 );
buf ( n47933 , n47932 );
not ( n47934 , n47933 );
or ( n47935 , n47929 , n47934 );
buf ( n47936 , n42458 );
buf ( n47937 , n25181 );
nand ( n47938 , n47936 , n47937 );
buf ( n47939 , n47938 );
buf ( n47940 , n47939 );
nand ( n47941 , n47935 , n47940 );
buf ( n47942 , n47941 );
buf ( n47943 , n47942 );
buf ( n47944 , n44586 );
nand ( n47945 , n47943 , n47944 );
buf ( n47946 , n47945 );
buf ( n47947 , n47946 );
nand ( n47948 , n47927 , n47947 );
buf ( n47949 , n47948 );
buf ( n47950 , n47949 );
and ( n47951 , n47922 , n47950 );
and ( n47952 , n47893 , n47921 );
or ( n47953 , n47951 , n47952 );
buf ( n47954 , n47953 );
buf ( n47955 , n47954 );
buf ( n47956 , n47955 );
buf ( n47957 , n47956 );
buf ( n47958 , n47957 );
not ( n47959 , n47958 );
buf ( n47960 , n42252 );
not ( n47961 , n47960 );
buf ( n47962 , n42266 );
not ( n47963 , n47962 );
buf ( n47964 , n38218 );
not ( n47965 , n47964 );
or ( n47966 , n47963 , n47965 );
buf ( n47967 , n39406 );
not ( n47968 , n47967 );
buf ( n47969 , n47968 );
buf ( n47970 , n47969 );
buf ( n47971 , n42263 );
nand ( n47972 , n47970 , n47971 );
buf ( n47973 , n47972 );
buf ( n47974 , n47973 );
nand ( n47975 , n47966 , n47974 );
buf ( n47976 , n47975 );
buf ( n47977 , n47976 );
not ( n47978 , n47977 );
or ( n47979 , n47961 , n47978 );
buf ( n47980 , n47544 );
buf ( n47981 , n42315 );
nand ( n47982 , n47980 , n47981 );
buf ( n47983 , n47982 );
buf ( n47984 , n47983 );
nand ( n47985 , n47979 , n47984 );
buf ( n47986 , n47985 );
buf ( n47987 , n47986 );
not ( n47988 , n47987 );
or ( n47989 , n47959 , n47988 );
buf ( n47990 , n47957 );
buf ( n47991 , n47986 );
or ( n47992 , n47990 , n47991 );
buf ( n47993 , n42847 );
not ( n47994 , n47993 );
buf ( n47995 , n43259 );
not ( n47996 , n47995 );
or ( n47997 , n47994 , n47996 );
buf ( n47998 , n43503 );
buf ( n47999 , n46691 );
nand ( n48000 , n47998 , n47999 );
buf ( n48001 , n48000 );
buf ( n48002 , n48001 );
nand ( n48003 , n47997 , n48002 );
buf ( n48004 , n48003 );
buf ( n48005 , n48004 );
not ( n48006 , n48005 );
buf ( n48007 , n42521 );
not ( n48008 , n48007 );
or ( n48009 , n48006 , n48008 );
buf ( n48010 , n42530 );
buf ( n48011 , n46334 );
nand ( n48012 , n48010 , n48011 );
buf ( n48013 , n48012 );
buf ( n48014 , n48013 );
nand ( n48015 , n48009 , n48014 );
buf ( n48016 , n48015 );
buf ( n48017 , n48016 );
xor ( n48018 , n47044 , n47056 );
xor ( n48019 , n48018 , n47077 );
buf ( n48020 , n48019 );
buf ( n48021 , n48020 );
xor ( n48022 , n48017 , n48021 );
buf ( n48023 , n43063 );
not ( n48024 , n48023 );
buf ( n48025 , n42082 );
not ( n48026 , n48025 );
or ( n48027 , n48024 , n48026 );
buf ( n48028 , n42062 );
buf ( n48029 , n44125 );
nand ( n48030 , n48028 , n48029 );
buf ( n48031 , n48030 );
buf ( n48032 , n48031 );
nand ( n48033 , n48027 , n48032 );
buf ( n48034 , n48033 );
buf ( n48035 , n48034 );
not ( n48036 , n48035 );
buf ( n48037 , n45158 );
not ( n48038 , n48037 );
or ( n48039 , n48036 , n48038 );
buf ( n48040 , n47396 );
not ( n48041 , n48040 );
buf ( n48042 , n36912 );
nand ( n48043 , n48041 , n48042 );
buf ( n48044 , n48043 );
buf ( n48045 , n48044 );
nand ( n48046 , n48039 , n48045 );
buf ( n48047 , n48046 );
buf ( n48048 , n48047 );
and ( n48049 , n48022 , n48048 );
and ( n48050 , n48017 , n48021 );
or ( n48051 , n48049 , n48050 );
buf ( n48052 , n48051 );
buf ( n48053 , n48052 );
nand ( n48054 , n47992 , n48053 );
buf ( n48055 , n48054 );
buf ( n48056 , n48055 );
nand ( n48057 , n47989 , n48056 );
buf ( n48058 , n48057 );
buf ( n48059 , n48058 );
and ( n48060 , n47830 , n48059 );
and ( n48061 , n47800 , n47829 );
or ( n48062 , n48060 , n48061 );
buf ( n48063 , n48062 );
buf ( n48064 , n48063 );
and ( n48065 , n47775 , n48064 );
and ( n48066 , n47598 , n47774 );
or ( n48067 , n48065 , n48066 );
buf ( n48068 , n48067 );
buf ( n48069 , n48068 );
not ( n48070 , n48069 );
buf ( n48071 , n48070 );
nand ( n48072 , n47594 , n48071 );
not ( n48073 , n48072 );
or ( n48074 , n47590 , n48073 );
buf ( n48075 , n48068 );
buf ( n48076 , n47593 );
nand ( n48077 , n48075 , n48076 );
buf ( n48078 , n48077 );
nand ( n48079 , n48074 , n48078 );
buf ( n48080 , n48079 );
not ( n48081 , n48080 );
buf ( n48082 , n48081 );
buf ( n48083 , n48082 );
nand ( n48084 , n47384 , n48083 );
buf ( n48085 , n48084 );
not ( n48086 , n48085 );
or ( n48087 , n47377 , n48086 );
buf ( n48088 , n47383 );
buf ( n48089 , n48082 );
or ( n48090 , n48088 , n48089 );
buf ( n48091 , n48090 );
nand ( n48092 , n48087 , n48091 );
not ( n48093 , n48092 );
xor ( n48094 , n47235 , n48093 );
xor ( n48095 , n46831 , n46565 );
xor ( n48096 , n48095 , n47197 );
and ( n48097 , n48094 , n48096 );
and ( n48098 , n47235 , n48093 );
or ( n48099 , n48097 , n48098 );
buf ( n48100 , n48099 );
nand ( n48101 , n47229 , n48100 );
buf ( n48102 , n48101 );
buf ( n48103 , n48102 );
xor ( n48104 , n47235 , n48093 );
xor ( n48105 , n48104 , n48096 );
buf ( n48106 , n47171 );
buf ( n48107 , n47193 );
and ( n48108 , n48106 , n48107 );
not ( n48109 , n48106 );
buf ( n48110 , n47184 );
and ( n48111 , n48109 , n48110 );
nor ( n48112 , n48108 , n48111 );
buf ( n48113 , n48112 );
buf ( n48114 , n48113 );
buf ( n48115 , n46839 );
not ( n48116 , n48115 );
buf ( n48117 , n48116 );
buf ( n48118 , n48117 );
and ( n48119 , n48114 , n48118 );
not ( n48120 , n48114 );
buf ( n48121 , n46839 );
and ( n48122 , n48120 , n48121 );
nor ( n48123 , n48119 , n48122 );
buf ( n48124 , n48123 );
buf ( n48125 , n48124 );
and ( n48126 , n47380 , n48079 );
not ( n48127 , n47380 );
and ( n48128 , n48127 , n48082 );
nor ( n48129 , n48126 , n48128 );
not ( n48130 , n47376 );
and ( n48131 , n48129 , n48130 );
not ( n48132 , n48129 );
and ( n48133 , n48132 , n47376 );
nor ( n48134 , n48131 , n48133 );
buf ( n48135 , n48134 );
xor ( n48136 , n48125 , n48135 );
buf ( n48137 , n47589 );
buf ( n48138 , n47593 );
xor ( n48139 , n48137 , n48138 );
buf ( n48140 , n48068 );
xnor ( n48141 , n48139 , n48140 );
buf ( n48142 , n48141 );
buf ( n48143 , n48142 );
xor ( n48144 , n47388 , n47580 );
xor ( n48145 , n48144 , n47585 );
buf ( n48146 , n48145 );
buf ( n48147 , n48146 );
not ( n48148 , n48147 );
buf ( n48149 , n48148 );
buf ( n48150 , n48149 );
buf ( n48151 , n48150 );
buf ( n48152 , n48151 );
not ( n48153 , n48152 );
xor ( n48154 , n47598 , n47774 );
xor ( n48155 , n48154 , n48064 );
buf ( n48156 , n48155 );
buf ( n48157 , n48156 );
not ( n48158 , n48157 );
buf ( n48159 , n48158 );
not ( n48160 , n48159 );
or ( n48161 , n48153 , n48160 );
or ( n48162 , n48152 , n48159 );
buf ( n48163 , n37394 );
not ( n48164 , n48163 );
buf ( n48165 , n48164 );
not ( n48166 , n48165 );
buf ( n48167 , n28368 );
not ( n48168 , n48167 );
buf ( n48169 , n48168 );
buf ( n48170 , n48169 );
not ( n48171 , n48170 );
buf ( n48172 , n48171 );
buf ( n48173 , n48172 );
buf ( n48174 , n41778 );
and ( n48175 , n48173 , n48174 );
not ( n48176 , n48173 );
buf ( n48177 , n47429 );
and ( n48178 , n48176 , n48177 );
nor ( n48179 , n48175 , n48178 );
buf ( n48180 , n48179 );
not ( n48181 , n48180 );
and ( n48182 , n48166 , n48181 );
not ( n48183 , n42132 );
buf ( n48184 , n41769 );
not ( n48185 , n48184 );
buf ( n48186 , n43362 );
not ( n48187 , n48186 );
and ( n48188 , n48185 , n48187 );
buf ( n48189 , n47429 );
buf ( n48190 , n47436 );
and ( n48191 , n48189 , n48190 );
nor ( n48192 , n48188 , n48191 );
buf ( n48193 , n48192 );
not ( n48194 , n48193 );
and ( n48195 , n48183 , n48194 );
nor ( n48196 , n48182 , n48195 );
buf ( n48197 , n48196 );
not ( n48198 , n48197 );
buf ( n48199 , n47043 );
not ( n48200 , n48199 );
or ( n48201 , n48198 , n48200 );
buf ( n48202 , n47490 );
buf ( n48203 , n43099 );
buf ( n48204 , n41828 );
and ( n48205 , n48203 , n48204 );
not ( n48206 , n48203 );
not ( n48207 , n41843 );
buf ( n48208 , n48207 );
and ( n48209 , n48206 , n48208 );
nor ( n48210 , n48205 , n48209 );
buf ( n48211 , n48210 );
buf ( n48212 , n48211 );
or ( n48213 , n48202 , n48212 );
buf ( n48214 , n37443 );
buf ( n48215 , n47500 );
or ( n48216 , n48214 , n48215 );
nand ( n48217 , n48213 , n48216 );
buf ( n48218 , n48217 );
buf ( n48219 , n48218 );
nand ( n48220 , n48201 , n48219 );
buf ( n48221 , n48220 );
buf ( n48222 , n48221 );
buf ( n48223 , n47043 );
not ( n48224 , n48223 );
buf ( n48225 , n48196 );
not ( n48226 , n48225 );
buf ( n48227 , n48226 );
buf ( n48228 , n48227 );
nand ( n48229 , n48224 , n48228 );
buf ( n48230 , n48229 );
buf ( n48231 , n48230 );
nand ( n48232 , n48222 , n48231 );
buf ( n48233 , n48232 );
buf ( n48234 , n48233 );
buf ( n48235 , n46117 );
not ( n48236 , n48235 );
buf ( n48237 , n43959 );
not ( n48238 , n48237 );
or ( n48239 , n48236 , n48238 );
buf ( n48240 , n39726 );
not ( n48241 , n48240 );
buf ( n48242 , n46126 );
nand ( n48243 , n48241 , n48242 );
buf ( n48244 , n48243 );
buf ( n48245 , n48244 );
nand ( n48246 , n48239 , n48245 );
buf ( n48247 , n48246 );
buf ( n48248 , n48247 );
not ( n48249 , n48248 );
buf ( n48250 , n44135 );
not ( n48251 , n48250 );
or ( n48252 , n48249 , n48251 );
buf ( n48253 , n36640 );
not ( n48254 , n48253 );
buf ( n48255 , n47611 );
nand ( n48256 , n48254 , n48255 );
buf ( n48257 , n48256 );
buf ( n48258 , n48257 );
nand ( n48259 , n48252 , n48258 );
buf ( n48260 , n48259 );
buf ( n48261 , n48260 );
xor ( n48262 , n48234 , n48261 );
buf ( n48263 , n47510 );
not ( n48264 , n48263 );
buf ( n48265 , n47456 );
not ( n48266 , n48265 );
buf ( n48267 , n47481 );
not ( n48268 , n48267 );
or ( n48269 , n48266 , n48268 );
buf ( n48270 , n47456 );
buf ( n48271 , n47481 );
or ( n48272 , n48270 , n48271 );
nand ( n48273 , n48269 , n48272 );
buf ( n48274 , n48273 );
buf ( n48275 , n48274 );
not ( n48276 , n48275 );
or ( n48277 , n48264 , n48276 );
buf ( n48278 , n47510 );
buf ( n48279 , n48274 );
or ( n48280 , n48278 , n48279 );
nand ( n48281 , n48277 , n48280 );
buf ( n48282 , n48281 );
buf ( n48283 , n48282 );
and ( n48284 , n48262 , n48283 );
and ( n48285 , n48234 , n48261 );
or ( n48286 , n48284 , n48285 );
buf ( n48287 , n48286 );
buf ( n48288 , n48287 );
not ( n48289 , n48288 );
buf ( n48290 , n48289 );
buf ( n48291 , n48290 );
not ( n48292 , n48291 );
buf ( n48293 , n41862 );
not ( n48294 , n48293 );
buf ( n48295 , n42504 );
not ( n48296 , n48295 );
buf ( n48297 , n41890 );
not ( n48298 , n48297 );
or ( n48299 , n48296 , n48298 );
buf ( n48300 , n41947 );
buf ( n48301 , n41721 );
nand ( n48302 , n48300 , n48301 );
buf ( n48303 , n48302 );
buf ( n48304 , n48303 );
nand ( n48305 , n48299 , n48304 );
buf ( n48306 , n48305 );
buf ( n48307 , n48306 );
not ( n48308 , n48307 );
or ( n48309 , n48294 , n48308 );
buf ( n48310 , n45617 );
buf ( n48311 , n47691 );
nand ( n48312 , n48310 , n48311 );
buf ( n48313 , n48312 );
buf ( n48314 , n48313 );
nand ( n48315 , n48309 , n48314 );
buf ( n48316 , n48315 );
not ( n48317 , n48316 );
buf ( n48318 , n25925 );
not ( n48319 , n48318 );
buf ( n48320 , n48319 );
buf ( n48321 , n48320 );
not ( n48322 , n48321 );
buf ( n48323 , n48322 );
buf ( n48324 , n48323 );
not ( n48325 , n48324 );
buf ( n48326 , n37649 );
not ( n48327 , n48326 );
or ( n48328 , n48325 , n48327 );
buf ( n48329 , n38834 );
buf ( n48330 , n48320 );
nand ( n48331 , n48329 , n48330 );
buf ( n48332 , n48331 );
buf ( n48333 , n48332 );
nand ( n48334 , n48328 , n48333 );
buf ( n48335 , n48334 );
buf ( n48336 , n36444 );
buf ( n48337 , n47731 );
nand ( n48338 , n48336 , n48337 );
buf ( n48339 , n48338 );
buf ( n48340 , n48339 );
nand ( n48341 , C1 , n48340 );
buf ( n48342 , n48341 );
not ( n48343 , n48342 );
or ( n48344 , n48317 , n48343 );
buf ( n48345 , n48342 );
buf ( n48346 , n48316 );
nor ( n48347 , n48345 , n48346 );
buf ( n48348 , n48347 );
buf ( n48349 , n44586 );
not ( n48350 , n48349 );
buf ( n48351 , n25182 );
not ( n48352 , n48351 );
buf ( n48353 , n44989 );
not ( n48354 , n48353 );
or ( n48355 , n48352 , n48354 );
buf ( n48356 , n25180 );
buf ( n48357 , n48356 );
buf ( n48358 , n48357 );
not ( n48359 , n48358 );
buf ( n48360 , n30187 );
nand ( n48361 , n48359 , n48360 );
buf ( n48362 , n48361 );
buf ( n48363 , n48362 );
nand ( n48364 , n48355 , n48363 );
buf ( n48365 , n48364 );
buf ( n48366 , n48365 );
not ( n48367 , n48366 );
or ( n48368 , n48350 , n48367 );
buf ( n48369 , n47942 );
buf ( n48370 , n46294 );
nand ( n48371 , n48369 , n48370 );
buf ( n48372 , n48371 );
buf ( n48373 , n48372 );
nand ( n48374 , n48368 , n48373 );
buf ( n48375 , n48374 );
buf ( n48376 , n48375 );
not ( n48377 , n48376 );
buf ( n48378 , n48377 );
or ( n48379 , n48348 , n48378 );
nand ( n48380 , n48344 , n48379 );
buf ( n48381 , n48380 );
not ( n48382 , n48381 );
buf ( n48383 , n41647 );
not ( n48384 , n48383 );
buf ( n48385 , n47633 );
not ( n48386 , n48385 );
or ( n48387 , n48384 , n48386 );
buf ( n48388 , n41660 );
not ( n48389 , n48388 );
buf ( n48390 , n48389 );
buf ( n48391 , n48390 );
not ( n48392 , n48391 );
buf ( n48393 , n37595 );
not ( n48394 , n48393 );
or ( n48395 , n48392 , n48394 );
buf ( n48396 , n37586 );
buf ( n48397 , n41660 );
nand ( n48398 , n48396 , n48397 );
buf ( n48399 , n48398 );
buf ( n48400 , n48399 );
nand ( n48401 , n48395 , n48400 );
buf ( n48402 , n48401 );
buf ( n48403 , n48402 );
buf ( n48404 , n41705 );
nand ( n48405 , n48403 , n48404 );
buf ( n48406 , n48405 );
buf ( n48407 , n48406 );
nand ( n48408 , n48387 , n48407 );
buf ( n48409 , n48408 );
buf ( n48410 , n48409 );
not ( n48411 , n48410 );
buf ( n48412 , n42343 );
buf ( n48413 , n37745 );
and ( n48414 , n48412 , n48413 );
not ( n48415 , n48412 );
buf ( n48416 , n42596 );
and ( n48417 , n48415 , n48416 );
nor ( n48418 , n48414 , n48417 );
buf ( n48419 , n48418 );
buf ( n48420 , n48419 );
not ( n48421 , n48420 );
buf ( n48422 , n42375 );
not ( n48423 , n48422 );
and ( n48424 , n48421 , n48423 );
buf ( n48425 , n47302 );
buf ( n48426 , n42339 );
and ( n48427 , n48425 , n48426 );
nor ( n48428 , n48424 , n48427 );
buf ( n48429 , n48428 );
buf ( n48430 , n48429 );
nand ( n48431 , n48411 , n48430 );
buf ( n48432 , n48431 );
buf ( n48433 , n48432 );
not ( n48434 , n48433 );
or ( n48435 , n48382 , n48434 );
buf ( n48436 , n48429 );
not ( n48437 , n48436 );
buf ( n48438 , n48409 );
buf ( n48439 , n48438 );
buf ( n48440 , n48439 );
buf ( n48441 , n48440 );
nand ( n48442 , n48437 , n48441 );
buf ( n48443 , n48442 );
buf ( n48444 , n48443 );
nand ( n48445 , n48435 , n48444 );
buf ( n48446 , n48445 );
buf ( n48447 , n48446 );
not ( n48448 , n48447 );
buf ( n48449 , n48448 );
buf ( n48450 , n48449 );
not ( n48451 , n48450 );
or ( n48452 , n48292 , n48451 );
xor ( n48453 , n47519 , n47520 );
buf ( n48454 , n48453 );
xor ( n48455 , n47516 , n48454 );
buf ( n48456 , n48455 );
nand ( n48457 , n48452 , n48456 );
buf ( n48458 , n48457 );
buf ( n48459 , n48458 );
buf ( n48460 , n48446 );
buf ( n48461 , n48287 );
nand ( n48462 , n48460 , n48461 );
buf ( n48463 , n48462 );
buf ( n48464 , n48463 );
nand ( n48465 , n48459 , n48464 );
buf ( n48466 , n48465 );
buf ( n48467 , n48466 );
not ( n48468 , n48467 );
buf ( n48469 , n48468 );
buf ( n48470 , n48469 );
not ( n48471 , n48470 );
buf ( n48472 , n46921 );
buf ( n48473 , n46869 );
and ( n48474 , n48472 , n48473 );
not ( n48475 , n48472 );
buf ( n48476 , n46870 );
and ( n48477 , n48475 , n48476 );
nor ( n48478 , n48474 , n48477 );
buf ( n48479 , n48478 );
buf ( n48480 , n48479 );
buf ( n48481 , n46951 );
xnor ( n48482 , n48480 , n48481 );
buf ( n48483 , n48482 );
buf ( n48484 , n48483 );
not ( n48485 , n48484 );
or ( n48486 , n48471 , n48485 );
buf ( n48487 , n46225 );
not ( n48488 , n48487 );
buf ( n48489 , n45753 );
not ( n48490 , n48489 );
buf ( n48491 , n39927 );
not ( n48492 , n48491 );
or ( n48493 , n48490 , n48492 );
buf ( n48494 , n36562 );
buf ( n48495 , n45750 );
nand ( n48496 , n48494 , n48495 );
buf ( n48497 , n48496 );
buf ( n48498 , n48497 );
nand ( n48499 , n48493 , n48498 );
buf ( n48500 , n48499 );
buf ( n48501 , n48500 );
not ( n48502 , n48501 );
or ( n48503 , n48488 , n48502 );
buf ( n48504 , n46944 );
buf ( n48505 , n46246 );
nand ( n48506 , n48504 , n48505 );
buf ( n48507 , n48506 );
buf ( n48508 , n48507 );
nand ( n48509 , n48503 , n48508 );
buf ( n48510 , n48509 );
buf ( n48511 , n48510 );
not ( n48512 , n48511 );
buf ( n48513 , n37146 );
not ( n48514 , n48513 );
buf ( n48515 , n41611 );
not ( n48516 , n48515 );
and ( n48517 , n48514 , n48516 );
buf ( n48518 , n39860 );
buf ( n48519 , n41611 );
and ( n48520 , n48518 , n48519 );
nor ( n48521 , n48517 , n48520 );
buf ( n48522 , n48521 );
buf ( n48523 , n48522 );
not ( n48524 , n48523 );
buf ( n48525 , n41599 );
not ( n48526 , n48525 );
and ( n48527 , n48524 , n48526 );
buf ( n48528 , n47821 );
buf ( n48529 , n43868 );
and ( n48530 , n48528 , n48529 );
nor ( n48531 , n48527 , n48530 );
buf ( n48532 , n48531 );
buf ( n48533 , n48532 );
not ( n48534 , n48533 );
buf ( n48535 , n48534 );
buf ( n48536 , n48535 );
not ( n48537 , n48536 );
or ( n48538 , n48512 , n48537 );
buf ( n48539 , n48535 );
buf ( n48540 , n48510 );
or ( n48541 , n48539 , n48540 );
xor ( n48542 , n47277 , n47284 );
xor ( n48543 , n48542 , n47310 );
buf ( n48544 , n48543 );
buf ( n48545 , n48544 );
nand ( n48546 , n48541 , n48545 );
buf ( n48547 , n48546 );
buf ( n48548 , n48547 );
nand ( n48549 , n48538 , n48548 );
buf ( n48550 , n48549 );
buf ( n48551 , n48550 );
nand ( n48552 , n48486 , n48551 );
buf ( n48553 , n48552 );
buf ( n48554 , n48553 );
buf ( n48555 , n48483 );
not ( n48556 , n48555 );
buf ( n48557 , n48466 );
nand ( n48558 , n48556 , n48557 );
buf ( n48559 , n48558 );
buf ( n48560 , n48559 );
nand ( n48561 , n48554 , n48560 );
buf ( n48562 , n48561 );
not ( n48563 , n48562 );
nand ( n48564 , n48162 , n48563 );
nand ( n48565 , n48161 , n48564 );
buf ( n48566 , n48565 );
xor ( n48567 , n48143 , n48566 );
not ( n48568 , n47567 );
not ( n48569 , n47554 );
or ( n48570 , n48568 , n48569 );
not ( n48571 , n47567 );
nand ( n48572 , n48571 , n47551 );
nand ( n48573 , n48570 , n48572 );
buf ( n48574 , n48573 );
buf ( n48575 , n47525 );
buf ( n48576 , n48575 );
buf ( n48577 , n48576 );
buf ( n48578 , n48577 );
not ( n48579 , n48578 );
buf ( n48580 , n48579 );
buf ( n48581 , n48580 );
and ( n48582 , n48574 , n48581 );
not ( n48583 , n48574 );
buf ( n48584 , n48577 );
and ( n48585 , n48583 , n48584 );
nor ( n48586 , n48582 , n48585 );
buf ( n48587 , n48586 );
buf ( n48588 , n48587 );
xor ( n48589 , n47620 , n47647 );
xor ( n48590 , n48589 , n47741 );
buf ( n48591 , n48590 );
buf ( n48592 , n48591 );
not ( n48593 , n48592 );
buf ( n48594 , n44708 );
not ( n48595 , n48594 );
buf ( n48596 , n44533 );
not ( n48597 , n48596 );
buf ( n48598 , n43597 );
not ( n48599 , n48598 );
or ( n48600 , n48597 , n48599 );
buf ( n48601 , n36396 );
buf ( n48602 , n44530 );
nand ( n48603 , n48601 , n48602 );
buf ( n48604 , n48603 );
buf ( n48605 , n48604 );
nand ( n48606 , n48600 , n48605 );
buf ( n48607 , n48606 );
buf ( n48608 , n48607 );
not ( n48609 , n48608 );
or ( n48610 , n48595 , n48609 );
buf ( n48611 , n47789 );
buf ( n48612 , n44496 );
nand ( n48613 , n48611 , n48612 );
buf ( n48614 , n48613 );
buf ( n48615 , n48614 );
nand ( n48616 , n48610 , n48615 );
buf ( n48617 , n48616 );
buf ( n48618 , n48617 );
not ( n48619 , n48618 );
or ( n48620 , n48593 , n48619 );
buf ( n48621 , n48617 );
buf ( n48622 , n48591 );
or ( n48623 , n48621 , n48622 );
xor ( n48624 , n47677 , n47706 );
xnor ( n48625 , n48624 , n47733 );
buf ( n48626 , n48625 );
buf ( n48627 , n41993 );
not ( n48628 , n48627 );
buf ( n48629 , n47898 );
not ( n48630 , n48629 );
or ( n48631 , n48628 , n48630 );
buf ( n48632 , n44004 );
buf ( n48633 , n43966 );
nand ( n48634 , n48632 , n48633 );
buf ( n48635 , n48634 );
buf ( n48636 , n48635 );
nand ( n48637 , n48631 , n48636 );
buf ( n48638 , n48637 );
buf ( n48639 , n48638 );
not ( n48640 , n48639 );
buf ( n48641 , n43386 );
not ( n48642 , n48641 );
or ( n48643 , n48640 , n48642 );
buf ( n48644 , n47908 );
buf ( n48645 , n46172 );
nand ( n48646 , n48644 , n48645 );
buf ( n48647 , n48646 );
buf ( n48648 , n48647 );
nand ( n48649 , n48643 , n48648 );
buf ( n48650 , n48649 );
buf ( n48651 , n48650 );
not ( n48652 , n48651 );
buf ( n48653 , n41705 );
not ( n48654 , n48653 );
buf ( n48655 , n48390 );
not ( n48656 , n48655 );
buf ( n48657 , n39701 );
not ( n48658 , n48657 );
or ( n48659 , n48656 , n48658 );
buf ( n48660 , n37641 );
buf ( n48661 , n41660 );
nand ( n48662 , n48660 , n48661 );
buf ( n48663 , n48662 );
buf ( n48664 , n48663 );
nand ( n48665 , n48659 , n48664 );
buf ( n48666 , n48665 );
buf ( n48667 , n48666 );
not ( n48668 , n48667 );
or ( n48669 , n48654 , n48668 );
buf ( n48670 , n48402 );
buf ( n48671 , n41643 );
buf ( n48672 , n48671 );
nand ( n48673 , n48670 , n48672 );
buf ( n48674 , n48673 );
buf ( n48675 , n48674 );
nand ( n48676 , n48669 , n48675 );
buf ( n48677 , n48676 );
buf ( n48678 , n48677 );
not ( n48679 , n48678 );
or ( n48680 , n48652 , n48679 );
buf ( n48681 , n48677 );
buf ( n48682 , n48650 );
or ( n48683 , n48681 , n48682 );
not ( n48684 , n39999 );
buf ( n48685 , n24092 );
not ( n48686 , n48685 );
buf ( n48687 , n41915 );
not ( n48688 , n48687 );
or ( n48689 , n48686 , n48688 );
buf ( n48690 , n41912 );
buf ( n48691 , n47857 );
nand ( n48692 , n48690 , n48691 );
buf ( n48693 , n48692 );
buf ( n48694 , n48693 );
nand ( n48695 , n48689 , n48694 );
buf ( n48696 , n48695 );
not ( n48697 , n48696 );
or ( n48698 , n48684 , n48697 );
not ( n48699 , n24092 );
or ( n48700 , n45075 , n48699 );
not ( n48701 , n29328 );
nand ( n48702 , n48701 , n48699 );
buf ( n48703 , n39980 );
not ( n48704 , n48703 );
buf ( n48705 , n48704 );
nand ( n48706 , n48700 , n48702 , n48705 );
nand ( n48707 , n48698 , n48706 );
buf ( n48708 , n48707 );
buf ( n48709 , n42566 );
not ( n48710 , n48709 );
buf ( n48711 , n47888 );
not ( n48712 , n48711 );
or ( n48713 , n48710 , n48712 );
buf ( n48714 , n41762 );
not ( n48715 , n48714 );
buf ( n48716 , n46356 );
not ( n48717 , n48716 );
and ( n48718 , n48715 , n48717 );
buf ( n48719 , n28723 );
buf ( n48720 , n46356 );
and ( n48721 , n48719 , n48720 );
nor ( n48722 , n48718 , n48721 );
buf ( n48723 , n48722 );
buf ( n48724 , n48723 );
not ( n48725 , n48724 );
buf ( n48726 , n42631 );
nand ( n48727 , n48725 , n48726 );
buf ( n48728 , n48727 );
buf ( n48729 , n48728 );
nand ( n48730 , n48713 , n48729 );
buf ( n48731 , n48730 );
buf ( n48732 , n48731 );
xor ( n48733 , n48708 , n48732 );
not ( n48734 , n42052 );
not ( n48735 , n42114 );
or ( n48736 , n48734 , n48735 );
nand ( n48737 , n41772 , n42049 );
nand ( n48738 , n48736 , n48737 );
buf ( n48739 , n48738 );
not ( n48740 , n48739 );
buf ( n48741 , n37397 );
not ( n48742 , n48741 );
or ( n48743 , n48740 , n48742 );
buf ( n48744 , n48180 );
not ( n48745 , n48744 );
buf ( n48746 , n37413 );
nand ( n48747 , n48745 , n48746 );
buf ( n48748 , n48747 );
buf ( n48749 , n48748 );
nand ( n48750 , n48743 , n48749 );
buf ( n48751 , n48750 );
buf ( n48752 , n48751 );
and ( n48753 , n48733 , n48752 );
and ( n48754 , n48708 , n48732 );
or ( n48755 , n48753 , n48754 );
buf ( n48756 , n48755 );
buf ( n48757 , n48756 );
nand ( n48758 , n48683 , n48757 );
buf ( n48759 , n48758 );
buf ( n48760 , n48759 );
nand ( n48761 , n48680 , n48760 );
buf ( n48762 , n48761 );
buf ( n48763 , n48762 );
xor ( n48764 , n48626 , n48763 );
buf ( n48765 , n42315 );
not ( n48766 , n48765 );
buf ( n48767 , n47976 );
not ( n48768 , n48767 );
or ( n48769 , n48766 , n48768 );
buf ( n48770 , n42266 );
not ( n48771 , n48770 );
buf ( n48772 , n43031 );
not ( n48773 , n48772 );
or ( n48774 , n48771 , n48773 );
buf ( n48775 , n38244 );
buf ( n48776 , n42263 );
nand ( n48777 , n48775 , n48776 );
buf ( n48778 , n48777 );
buf ( n48779 , n48778 );
nand ( n48780 , n48774 , n48779 );
buf ( n48781 , n48780 );
buf ( n48782 , n48781 );
buf ( n48783 , n42252 );
nand ( n48784 , n48782 , n48783 );
buf ( n48785 , n48784 );
buf ( n48786 , n48785 );
nand ( n48787 , n48769 , n48786 );
buf ( n48788 , n48787 );
buf ( n48789 , n48788 );
and ( n48790 , n48764 , n48789 );
and ( n48791 , n48626 , n48763 );
or ( n48792 , n48790 , n48791 );
buf ( n48793 , n48792 );
buf ( n48794 , n48793 );
nand ( n48795 , n48623 , n48794 );
buf ( n48796 , n48795 );
buf ( n48797 , n48796 );
nand ( n48798 , n48620 , n48797 );
buf ( n48799 , n48798 );
buf ( n48800 , n48799 );
xor ( n48801 , n48588 , n48800 );
xor ( n48802 , n47954 , n47986 );
xnor ( n48803 , n48802 , n48052 );
buf ( n48804 , n48803 );
not ( n48805 , n48804 );
buf ( n48806 , n48805 );
not ( n48807 , n48806 );
not ( n48808 , n24713 );
buf ( n48809 , n48808 );
not ( n48810 , n48809 );
buf ( n48811 , n35969 );
not ( n48812 , n48811 );
or ( n48813 , n48810 , n48812 );
buf ( n48814 , n46880 );
not ( n48815 , n48814 );
buf ( n48816 , n48808 );
not ( n48817 , n48816 );
buf ( n48818 , n48817 );
buf ( n48819 , n48818 );
buf ( n48820 , n48819 );
buf ( n48821 , n48820 );
buf ( n48822 , n48821 );
nand ( n48823 , n48815 , n48822 );
buf ( n48824 , n48823 );
buf ( n48825 , n48824 );
nand ( n48826 , n48813 , n48825 );
buf ( n48827 , n48826 );
buf ( n48828 , n48827 );
buf ( n48829 , n24689 );
not ( n48830 , n48829 );
buf ( n48831 , n48830 );
buf ( n48832 , n48831 );
not ( n48833 , n48832 );
buf ( n48834 , n48833 );
nand ( n48835 , n24714 , n48834 );
buf ( n48836 , n24661 );
buf ( n48837 , n48836 );
not ( n48838 , n48837 );
buf ( n48839 , n48838 );
buf ( n48840 , n48839 );
buf ( n48841 , n24689 );
xor ( n48842 , n48840 , n48841 );
buf ( n48843 , n48842 );
buf ( n48844 , n24713 );
buf ( n48845 , n48831 );
nand ( n48846 , n48844 , n48845 );
buf ( n48847 , n48846 );
and ( n48848 , n48835 , n48843 , n48847 );
not ( n48849 , n48848 );
buf ( n48850 , n48849 );
not ( n48851 , n48850 );
buf ( n48852 , n48851 );
buf ( n48853 , n48852 );
buf ( n48854 , n48853 );
buf ( n48855 , n48854 );
buf ( n48856 , n48855 );
not ( n48857 , n48856 );
buf ( n48858 , n48857 );
buf ( n48859 , n48858 );
buf ( n48860 , n48843 );
not ( n48861 , n48860 );
buf ( n48862 , n48861 );
buf ( n48863 , n48862 );
buf ( n48864 , n48863 );
buf ( n48865 , n48864 );
buf ( n48866 , n48865 );
buf ( n48867 , n48866 );
buf ( n48868 , n48867 );
buf ( n48869 , n48868 );
not ( n48870 , n48869 );
buf ( n48871 , n48870 );
buf ( n48872 , n48871 );
nand ( n48873 , n48859 , n48872 );
buf ( n48874 , n48873 );
buf ( n48875 , n48874 );
nand ( n48876 , n48828 , n48875 );
buf ( n48877 , n48876 );
buf ( n48878 , n48877 );
buf ( n48879 , n46912 );
not ( n48880 , n48879 );
buf ( n48881 , n47345 );
not ( n48882 , n48881 );
or ( n48883 , n48880 , n48882 );
buf ( n48884 , n46875 );
not ( n48885 , n48884 );
buf ( n48886 , n45650 );
not ( n48887 , n48886 );
or ( n48888 , n48885 , n48887 );
buf ( n48889 , n36611 );
buf ( n48890 , n46887 );
nand ( n48891 , n48889 , n48890 );
buf ( n48892 , n48891 );
buf ( n48893 , n48892 );
nand ( n48894 , n48888 , n48893 );
buf ( n48895 , n48894 );
buf ( n48896 , n48895 );
buf ( n48897 , n47331 );
nand ( n48898 , n48896 , n48897 );
buf ( n48899 , n48898 );
buf ( n48900 , n48899 );
nand ( n48901 , n48883 , n48900 );
buf ( n48902 , n48901 );
buf ( n48903 , n48902 );
xor ( n48904 , n48878 , n48903 );
not ( n48905 , n42668 );
not ( n48906 , n47323 );
or ( n48907 , n48905 , n48906 );
buf ( n48908 , n42672 );
not ( n48909 , n48908 );
buf ( n48910 , n43224 );
not ( n48911 , n48910 );
or ( n48912 , n48909 , n48911 );
buf ( n48913 , n37294 );
buf ( n48914 , n42671 );
nand ( n48915 , n48913 , n48914 );
buf ( n48916 , n48915 );
buf ( n48917 , n48916 );
nand ( n48918 , n48912 , n48917 );
buf ( n48919 , n48918 );
buf ( n48920 , n48919 );
buf ( n48921 , n42712 );
nand ( n48922 , n48920 , n48921 );
buf ( n48923 , n48922 );
nand ( n48924 , n48907 , n48923 );
buf ( n48925 , n48924 );
and ( n48926 , n48904 , n48925 );
and ( n48927 , n48878 , n48903 );
or ( n48928 , n48926 , n48927 );
buf ( n48929 , n48928 );
not ( n48930 , n48929 );
or ( n48931 , n48807 , n48930 );
buf ( n48932 , n48929 );
not ( n48933 , n48932 );
buf ( n48934 , n48933 );
not ( n48935 , n48934 );
not ( n48936 , n48803 );
or ( n48937 , n48935 , n48936 );
buf ( n48938 , n42448 );
not ( n48939 , n48938 );
buf ( n48940 , n47011 );
not ( n48941 , n48940 );
or ( n48942 , n48939 , n48941 );
buf ( n48943 , n47014 );
buf ( n48944 , n47063 );
not ( n48945 , n48944 );
buf ( n48946 , n47031 );
not ( n48947 , n48946 );
or ( n48948 , n48945 , n48947 );
buf ( n48949 , n38979 );
buf ( n48950 , n41873 );
nand ( n48951 , n48949 , n48950 );
buf ( n48952 , n48951 );
buf ( n48953 , n48952 );
nand ( n48954 , n48948 , n48953 );
buf ( n48955 , n48954 );
buf ( n48956 , n48955 );
nand ( n48957 , n48943 , n48956 );
buf ( n48958 , n48957 );
buf ( n48959 , n48958 );
nand ( n48960 , n48942 , n48959 );
buf ( n48961 , n48960 );
buf ( n48962 , n48961 );
not ( n48963 , n48962 );
buf ( n48964 , n48963 );
buf ( n48965 , n48964 );
not ( n48966 , n48965 );
or ( n48967 , n45075 , n48699 );
nand ( n48968 , n48967 , n48702 );
not ( n48969 , n48968 );
buf ( n48970 , n39998 );
not ( n48971 , n48970 );
and ( n48972 , n48969 , n48971 );
buf ( n48973 , n39980 );
not ( n48974 , n48973 );
buf ( n48975 , n48974 );
and ( n48976 , n47863 , n48975 );
nor ( n48977 , n48972 , n48976 );
buf ( n48978 , n48977 );
not ( n48979 , n48978 );
or ( n48980 , n48966 , n48979 );
buf ( n48981 , n44039 );
buf ( n48982 , n45069 );
not ( n48983 , n48982 );
buf ( n48984 , n48983 );
buf ( n48985 , n48984 );
not ( n48986 , n48985 );
buf ( n48987 , n47436 );
not ( n48988 , n48987 );
and ( n48989 , n48986 , n48988 );
buf ( n48990 , n47068 );
buf ( n48991 , n47436 );
and ( n48992 , n48990 , n48991 );
nor ( n48993 , n48989 , n48992 );
buf ( n48994 , n48993 );
buf ( n48995 , n48994 );
or ( n48996 , n48981 , n48995 );
buf ( n48997 , n47844 );
buf ( n48998 , n38381 );
or ( n48999 , n48997 , n48998 );
nand ( n49000 , n48996 , n48999 );
buf ( n49001 , n49000 );
buf ( n49002 , n49001 );
nand ( n49003 , n48980 , n49002 );
buf ( n49004 , n49003 );
buf ( n49005 , n49004 );
buf ( n49006 , n48977 );
not ( n49007 , n49006 );
buf ( n49008 , n48961 );
nand ( n49009 , n49007 , n49008 );
buf ( n49010 , n49009 );
buf ( n49011 , n49010 );
nand ( n49012 , n49005 , n49011 );
buf ( n49013 , n49012 );
buf ( n49014 , n44952 );
not ( n49015 , n49014 );
buf ( n49016 , n43259 );
not ( n49017 , n49016 );
or ( n49018 , n49015 , n49017 );
buf ( n49019 , n43503 );
buf ( n49020 , n44961 );
nand ( n49021 , n49019 , n49020 );
buf ( n49022 , n49021 );
buf ( n49023 , n49022 );
nand ( n49024 , n49018 , n49023 );
buf ( n49025 , n49024 );
not ( n49026 , n49025 );
not ( n49027 , n42521 );
or ( n49028 , n49026 , n49027 );
buf ( n49029 , n48004 );
buf ( n49030 , n42834 );
nand ( n49031 , n49029 , n49030 );
buf ( n49032 , n49031 );
nand ( n49033 , n49028 , n49032 );
xor ( n49034 , n49013 , n49033 );
not ( n49035 , n47868 );
not ( n49036 , n47890 );
and ( n49037 , n49035 , n49036 );
and ( n49038 , n47868 , n47890 );
nor ( n49039 , n49037 , n49038 );
buf ( n49040 , n47847 );
and ( n49041 , n49039 , n49040 );
not ( n49042 , n49039 );
not ( n49043 , n49040 );
and ( n49044 , n49042 , n49043 );
nor ( n49045 , n49041 , n49044 );
and ( n49046 , n49034 , n49045 );
and ( n49047 , n49013 , n49033 );
or ( n49048 , n49046 , n49047 );
not ( n49049 , n49048 );
not ( n49050 , n49049 );
xor ( n49051 , n47893 , n47921 );
xor ( n49052 , n49051 , n47950 );
buf ( n49053 , n49052 );
not ( n49054 , n49053 );
not ( n49055 , n49054 );
or ( n49056 , n49050 , n49055 );
xor ( n49057 , n48017 , n48021 );
xor ( n49058 , n49057 , n48048 );
buf ( n49059 , n49058 );
nand ( n49060 , n49056 , n49059 );
not ( n49061 , n49054 );
nand ( n49062 , n49061 , n49048 );
nand ( n49063 , n49060 , n49062 );
nand ( n49064 , n48937 , n49063 );
nand ( n49065 , n48931 , n49064 );
buf ( n49066 , n49065 );
and ( n49067 , n48801 , n49066 );
and ( n49068 , n48588 , n48800 );
or ( n49069 , n49067 , n49068 );
buf ( n49070 , n49069 );
not ( n49071 , n49070 );
buf ( n49072 , n47365 );
buf ( n49073 , n47251 );
and ( n49074 , n49072 , n49073 );
not ( n49075 , n49072 );
buf ( n49076 , n47259 );
and ( n49077 , n49075 , n49076 );
nor ( n49078 , n49074 , n49077 );
buf ( n49079 , n49078 );
not ( n49080 , n47255 );
and ( n49081 , n49079 , n49080 );
not ( n49082 , n49079 );
and ( n49083 , n49082 , n47255 );
nor ( n49084 , n49081 , n49083 );
nand ( n49085 , n49071 , n49084 );
buf ( n49086 , n49085 );
xor ( n49087 , n47800 , n47829 );
xor ( n49088 , n49087 , n48059 );
buf ( n49089 , n49088 );
buf ( n49090 , n49089 );
not ( n49091 , n49090 );
xor ( n49092 , n47746 , n47757 );
xor ( n49093 , n49092 , n47769 );
buf ( n49094 , n49093 );
not ( n49095 , n49094 );
nand ( n49096 , n49091 , n49095 );
not ( n49097 , n49096 );
not ( n49098 , n47263 );
not ( n49099 , n49098 );
xor ( n49100 , n47314 , n47363 );
not ( n49101 , n49100 );
or ( n49102 , n49099 , n49101 );
or ( n49103 , n49100 , n49098 );
nand ( n49104 , n49102 , n49103 );
not ( n49105 , n49104 );
or ( n49106 , n49097 , n49105 );
nand ( n49107 , n49090 , n49094 );
nand ( n49108 , n49106 , n49107 );
buf ( n49109 , n49108 );
and ( n49110 , n49086 , n49109 );
buf ( n49111 , n49070 );
not ( n49112 , n49111 );
buf ( n49113 , n49084 );
nor ( n49114 , n49112 , n49113 );
buf ( n49115 , n49114 );
buf ( n49116 , n49115 );
nor ( n49117 , n49110 , n49116 );
buf ( n49118 , n49117 );
buf ( n49119 , n49118 );
and ( n49120 , n48567 , n49119 );
and ( n49121 , n48143 , n48566 );
or ( n49122 , n49120 , n49121 );
buf ( n49123 , n49122 );
buf ( n49124 , n49123 );
and ( n49125 , n48136 , n49124 );
and ( n49126 , n48125 , n48135 );
or ( n49127 , n49125 , n49126 );
buf ( n49128 , n49127 );
nand ( n49129 , n48105 , n49128 );
buf ( n49130 , n49129 );
nand ( n49131 , n43833 , n45709 );
not ( n49132 , n49131 );
not ( n49133 , n46537 );
or ( n49134 , n49132 , n49133 );
nand ( n49135 , n43832 , n45708 );
nand ( n49136 , n49134 , n49135 );
buf ( n49137 , n49136 );
not ( n49138 , n49137 );
xor ( n49139 , n42726 , n43542 );
and ( n49140 , n49139 , n43831 );
and ( n49141 , n42726 , n43542 );
or ( n49142 , n49140 , n49141 );
buf ( n49143 , n49142 );
not ( n49144 , n45481 );
not ( n49145 , n45202 );
or ( n49146 , n49144 , n49145 );
not ( n49147 , n45481 );
not ( n49148 , n49147 );
not ( n49149 , n45205 );
or ( n49150 , n49148 , n49149 );
nand ( n49151 , n49150 , n45703 );
nand ( n49152 , n49146 , n49151 );
buf ( n49153 , n49152 );
xor ( n49154 , n49143 , n49153 );
xor ( n49155 , n45211 , n45451 );
and ( n49156 , n49155 , n45480 );
and ( n49157 , n45211 , n45451 );
or ( n49158 , n49156 , n49157 );
xor ( n49159 , n45217 , n45324 );
and ( n49160 , n49159 , n45449 );
and ( n49161 , n45217 , n45324 );
or ( n49162 , n49160 , n49161 );
buf ( n49163 , n49162 );
buf ( n49164 , n49163 );
xor ( n49165 , n45350 , n45363 );
and ( n49166 , n49165 , n45446 );
and ( n49167 , n45350 , n45363 );
or ( n49168 , n49166 , n49167 );
buf ( n49169 , n49168 );
buf ( n49170 , n49169 );
buf ( n49171 , n39986 );
not ( n49172 , n49171 );
buf ( n49173 , n40010 );
not ( n49174 , n49173 );
buf ( n49175 , n38286 );
not ( n49176 , n49175 );
or ( n49177 , n49174 , n49176 );
not ( n49178 , n37293 );
not ( n49179 , n49178 );
buf ( n49180 , n49179 );
buf ( n49181 , n40009 );
nand ( n49182 , n49180 , n49181 );
buf ( n49183 , n49182 );
buf ( n49184 , n49183 );
nand ( n49185 , n49177 , n49184 );
buf ( n49186 , n49185 );
buf ( n49187 , n49186 );
not ( n49188 , n49187 );
or ( n49189 , n49172 , n49188 );
buf ( n49190 , n43632 );
buf ( n49191 , n40002 );
nand ( n49192 , n49190 , n49191 );
buf ( n49193 , n49192 );
buf ( n49194 , n49193 );
nand ( n49195 , n49189 , n49194 );
buf ( n49196 , n49195 );
buf ( n49197 , n49196 );
xor ( n49198 , n45389 , n45419 );
and ( n49199 , n49198 , n45443 );
and ( n49200 , n45389 , n45419 );
or ( n49201 , n49199 , n49200 );
buf ( n49202 , n49201 );
buf ( n49203 , n49202 );
xor ( n49204 , n49197 , n49203 );
not ( n49205 , n42004 );
buf ( n49206 , n38834 );
not ( n49207 , n49206 );
buf ( n49208 , n41748 );
not ( n49209 , n49208 );
and ( n49210 , n49207 , n49209 );
buf ( n49211 , n38798 );
buf ( n49212 , n41748 );
and ( n49213 , n49211 , n49212 );
nor ( n49214 , n49210 , n49213 );
buf ( n49215 , n49214 );
not ( n49216 , n49215 );
and ( n49217 , n49205 , n49216 );
nor ( n49218 , n49217 , C0 );
buf ( n49219 , n43798 );
not ( n49220 , n49219 );
buf ( n49221 , n43817 );
not ( n49222 , n49221 );
and ( n49223 , n49220 , n49222 );
buf ( n49224 , n37916 );
buf ( n49225 , n41975 );
buf ( n49226 , n37880 );
not ( n49227 , n49226 );
buf ( n49228 , n49227 );
buf ( n49229 , n49228 );
and ( n49230 , n49225 , n49229 );
not ( n49231 , n49225 );
buf ( n49232 , n41894 );
and ( n49233 , n49231 , n49232 );
nor ( n49234 , n49230 , n49233 );
buf ( n49235 , n49234 );
buf ( n49236 , n49235 );
nor ( n49237 , n49224 , n49236 );
buf ( n49238 , n49237 );
buf ( n49239 , n49238 );
nor ( n49240 , n49223 , n49239 );
buf ( n49241 , n49240 );
buf ( n49242 , n49241 );
not ( n49243 , n49242 );
buf ( n49244 , n49243 );
buf ( n49245 , n49244 );
buf ( n49246 , n45304 );
not ( n49247 , n49246 );
buf ( n49248 , n36104 );
not ( n49249 , n49248 );
or ( n49250 , n49247 , n49249 );
buf ( n49251 , n39718 );
buf ( n49252 , n43368 );
not ( n49253 , n49252 );
buf ( n49254 , n39493 );
not ( n49255 , n49254 );
or ( n49256 , n49253 , n49255 );
buf ( n49257 , n43503 );
buf ( n49258 , n43365 );
nand ( n49259 , n49257 , n49258 );
buf ( n49260 , n49259 );
buf ( n49261 , n49260 );
nand ( n49262 , n49256 , n49261 );
buf ( n49263 , n49262 );
buf ( n49264 , n49263 );
nand ( n49265 , n49251 , n49264 );
buf ( n49266 , n49265 );
buf ( n49267 , n49266 );
nand ( n49268 , n49250 , n49267 );
buf ( n49269 , n49268 );
buf ( n49270 , n49269 );
xor ( n49271 , n49245 , n49270 );
buf ( n49272 , n49271 );
not ( n49273 , n49272 );
xor ( n49274 , n49218 , n49273 );
buf ( n49275 , n49274 );
xor ( n49276 , n49204 , n49275 );
buf ( n49277 , n49276 );
buf ( n49278 , n49277 );
xor ( n49279 , n49170 , n49278 );
buf ( n49280 , n38150 );
not ( n49281 , n49280 );
buf ( n49282 , n43434 );
not ( n49283 , n49282 );
buf ( n49284 , n42899 );
not ( n49285 , n49284 );
or ( n49286 , n49283 , n49285 );
buf ( n49287 , n38830 );
buf ( n49288 , n37328 );
nand ( n49289 , n49287 , n49288 );
buf ( n49290 , n49289 );
buf ( n49291 , n49290 );
nand ( n49292 , n49286 , n49291 );
buf ( n49293 , n49292 );
buf ( n49294 , n49293 );
not ( n49295 , n49294 );
or ( n49296 , n49281 , n49295 );
buf ( n49297 , n37400 );
buf ( n49298 , n45271 );
nand ( n49299 , n49297 , n49298 );
buf ( n49300 , n49299 );
buf ( n49301 , n49300 );
nand ( n49302 , n49296 , n49301 );
buf ( n49303 , n49302 );
buf ( n49304 , n49303 );
buf ( n49305 , n43786 );
not ( n49306 , n49305 );
buf ( n49307 , n43766 );
not ( n49308 , n49307 );
or ( n49309 , n49306 , n49308 );
and ( n49310 , n42434 , n43780 );
not ( n49311 , n42434 );
and ( n49312 , n49311 , n41844 );
nor ( n49313 , n49310 , n49312 );
buf ( n49314 , n49313 );
not ( n49315 , n49314 );
buf ( n49316 , n44253 );
nand ( n49317 , n49315 , n49316 );
buf ( n49318 , n49317 );
buf ( n49319 , n49318 );
nand ( n49320 , n49309 , n49319 );
buf ( n49321 , n49320 );
buf ( n49322 , n49321 );
not ( n49323 , n49322 );
buf ( n49324 , n49323 );
buf ( n49325 , n49324 );
xor ( n49326 , n49304 , n49325 );
buf ( n49327 , n38775 );
not ( n49328 , n49327 );
buf ( n49329 , n45407 );
not ( n49330 , n49329 );
or ( n49331 , n49328 , n49330 );
buf ( n49332 , n38413 );
not ( n49333 , n49332 );
buf ( n49334 , n39489 );
not ( n49335 , n49334 );
buf ( n49336 , n49335 );
buf ( n49337 , n49336 );
not ( n49338 , n49337 );
or ( n49339 , n49333 , n49338 );
buf ( n49340 , n39489 );
buf ( n49341 , n45401 );
nand ( n49342 , n49340 , n49341 );
buf ( n49343 , n49342 );
buf ( n49344 , n49343 );
nand ( n49345 , n49339 , n49344 );
buf ( n49346 , n49345 );
buf ( n49347 , n49346 );
buf ( n49348 , n38758 );
nand ( n49349 , n49347 , n49348 );
buf ( n49350 , n49349 );
buf ( n49351 , n49350 );
nand ( n49352 , n49331 , n49351 );
buf ( n49353 , n49352 );
buf ( n49354 , n49353 );
xor ( n49355 , n49326 , n49354 );
buf ( n49356 , n49355 );
buf ( n49357 , n49356 );
buf ( n49358 , n42712 );
not ( n49359 , n49358 );
buf ( n49360 , n43577 );
not ( n49361 , n49360 );
or ( n49362 , n49359 , n49361 );
and ( n49363 , n39582 , n25228 );
not ( n49364 , n39582 );
and ( n49365 , n49364 , n42671 );
or ( n49366 , n49363 , n49365 );
buf ( n49367 , n49366 );
buf ( n49368 , n42668 );
nand ( n49369 , n49367 , n49368 );
buf ( n49370 , n49369 );
buf ( n49371 , n49370 );
nand ( n49372 , n49362 , n49371 );
buf ( n49373 , n49372 );
buf ( n49374 , n49373 );
xor ( n49375 , n49357 , n49374 );
buf ( n49376 , n38127 );
buf ( n49377 , n45381 );
not ( n49378 , n49377 );
buf ( n49379 , n49378 );
buf ( n49380 , n49379 );
or ( n49381 , n49376 , n49380 );
buf ( n49382 , n41823 );
buf ( n49383 , n43403 );
not ( n49384 , n49383 );
buf ( n49385 , n49384 );
buf ( n49386 , n49385 );
and ( n49387 , n49382 , n49386 );
not ( n49388 , n49382 );
buf ( n49389 , n43371 );
not ( n49390 , n49389 );
buf ( n49391 , n49390 );
buf ( n49392 , n49391 );
and ( n49393 , n49388 , n49392 );
nor ( n49394 , n49387 , n49393 );
buf ( n49395 , n49394 );
buf ( n49396 , n49395 );
buf ( n49397 , n38057 );
or ( n49398 , n49396 , n49397 );
nand ( n49399 , n49381 , n49398 );
buf ( n49400 , n49399 );
buf ( n49401 , n49400 );
buf ( n49402 , n43736 );
not ( n49403 , n49402 );
buf ( n49404 , n49403 );
not ( n49405 , n49404 );
not ( n49406 , n36523 );
or ( n49407 , n49405 , n49406 );
not ( n49408 , n36533 );
not ( n49409 , n42052 );
or ( n49410 , n49408 , n49409 );
nand ( n49411 , n36530 , n42055 );
nand ( n49412 , n49410 , n49411 );
nand ( n49413 , n49412 , n44141 );
nand ( n49414 , n49407 , n49413 );
buf ( n49415 , n49414 );
xor ( n49416 , n49401 , n49415 );
buf ( n49417 , n44670 );
buf ( n49418 , n45438 );
or ( n49419 , n49417 , n49418 );
buf ( n49420 , n37005 );
buf ( n49421 , n41882 );
not ( n49422 , n49421 );
buf ( n49423 , n39136 );
not ( n49424 , n49423 );
buf ( n49425 , n49424 );
buf ( n49426 , n49425 );
not ( n49427 , n49426 );
or ( n49428 , n49422 , n49427 );
buf ( n49429 , n43095 );
buf ( n49430 , n41879 );
nand ( n49431 , n49429 , n49430 );
buf ( n49432 , n49431 );
buf ( n49433 , n49432 );
nand ( n49434 , n49428 , n49433 );
buf ( n49435 , n49434 );
buf ( n49436 , n49435 );
not ( n49437 , n49436 );
buf ( n49438 , n49437 );
buf ( n49439 , n49438 );
or ( n49440 , n49420 , n49439 );
nand ( n49441 , n49419 , n49440 );
buf ( n49442 , n49441 );
buf ( n49443 , n49442 );
xor ( n49444 , n49416 , n49443 );
buf ( n49445 , n49444 );
buf ( n49446 , n49445 );
xor ( n49447 , n49375 , n49446 );
buf ( n49448 , n49447 );
buf ( n49449 , n49448 );
xor ( n49450 , n49279 , n49449 );
buf ( n49451 , n49450 );
buf ( n49452 , n49451 );
xor ( n49453 , n49164 , n49452 );
xor ( n49454 , n41630 , n41712 );
and ( n49455 , n49454 , n42039 );
and ( n49456 , n41630 , n41712 );
or ( n49457 , n49455 , n49456 );
buf ( n49458 , n49457 );
buf ( n49459 , n49458 );
not ( n49460 , n42315 );
buf ( n49461 , n39008 );
not ( n49462 , n49461 );
buf ( n49463 , n42263 );
nand ( n49464 , n49462 , n49463 );
buf ( n49465 , n49464 );
nand ( n49466 , n42266 , n41619 );
nand ( n49467 , n49465 , n49466 );
not ( n49468 , n49467 );
or ( n49469 , n49460 , n49468 );
buf ( n49470 , n45339 );
buf ( n49471 , n42252 );
nand ( n49472 , n49470 , n49471 );
buf ( n49473 , n49472 );
nand ( n49474 , n49469 , n49473 );
not ( n49475 , n45355 );
not ( n49476 , n42631 );
or ( n49477 , n49475 , n49476 );
buf ( n49478 , n25160 );
not ( n49479 , n49478 );
buf ( n49480 , n43031 );
not ( n49481 , n49480 );
or ( n49482 , n49479 , n49481 );
buf ( n49483 , n38247 );
buf ( n49484 , n42581 );
nand ( n49485 , n49483 , n49484 );
buf ( n49486 , n49485 );
buf ( n49487 , n49486 );
nand ( n49488 , n49482 , n49487 );
buf ( n49489 , n49488 );
buf ( n49490 , n49489 );
buf ( n49491 , n42566 );
nand ( n49492 , n49490 , n49491 );
buf ( n49493 , n49492 );
nand ( n49494 , n49477 , n49493 );
xor ( n49495 , n49474 , n49494 );
not ( n49496 , n44586 );
not ( n49497 , n45234 );
or ( n49498 , n49496 , n49497 );
not ( n49499 , n43906 );
buf ( n49500 , n25184 );
not ( n49501 , n49500 );
buf ( n49502 , n39280 );
not ( n49503 , n49502 );
or ( n49504 , n49501 , n49503 );
buf ( n49505 , n39277 );
buf ( n49506 , n25183 );
nand ( n49507 , n49505 , n49506 );
buf ( n49508 , n49507 );
buf ( n49509 , n49508 );
nand ( n49510 , n49504 , n49509 );
buf ( n49511 , n49510 );
nand ( n49512 , n49499 , n49511 );
nand ( n49513 , n49498 , n49512 );
xor ( n49514 , n49495 , n49513 );
buf ( n49515 , n49514 );
xor ( n49516 , n49459 , n49515 );
xor ( n49517 , n43560 , n43585 );
and ( n49518 , n49517 , n43592 );
and ( n49519 , n43560 , n43585 );
or ( n49520 , n49518 , n49519 );
buf ( n49521 , n49520 );
buf ( n49522 , n49521 );
xor ( n49523 , n49516 , n49522 );
buf ( n49524 , n49523 );
buf ( n49525 , n49524 );
xor ( n49526 , n49453 , n49525 );
buf ( n49527 , n49526 );
not ( n49528 , n49527 );
xor ( n49529 , n49158 , n49528 );
xor ( n49530 , n42042 , n42390 );
and ( n49531 , n49530 , n42724 );
and ( n49532 , n42042 , n42390 );
or ( n49533 , n49531 , n49532 );
buf ( n49534 , n49533 );
buf ( n49535 , n49534 );
xor ( n49536 , n43554 , n43595 );
and ( n49537 , n49536 , n43829 );
and ( n49538 , n43554 , n43595 );
or ( n49539 , n49537 , n49538 );
buf ( n49540 , n49539 );
buf ( n49541 , n49540 );
xor ( n49542 , n49535 , n49541 );
buf ( n49543 , n43745 );
not ( n49544 , n49543 );
buf ( n49545 , n43751 );
not ( n49546 , n49545 );
or ( n49547 , n49544 , n49546 );
buf ( n49548 , n43742 );
not ( n49549 , n49548 );
buf ( n49550 , n43714 );
not ( n49551 , n49550 );
or ( n49552 , n49549 , n49551 );
buf ( n49553 , n43824 );
nand ( n49554 , n49552 , n49553 );
buf ( n49555 , n49554 );
buf ( n49556 , n49555 );
nand ( n49557 , n49547 , n49556 );
buf ( n49558 , n49557 );
buf ( n49559 , n49558 );
nand ( n49560 , n43643 , n43611 , n43614 );
not ( n49561 , n49560 );
not ( n49562 , n43661 );
or ( n49563 , n49561 , n49562 );
not ( n49564 , n43614 );
not ( n49565 , n43611 );
or ( n49566 , n49564 , n49565 );
not ( n49567 , n43643 );
nand ( n49568 , n49566 , n49567 );
nand ( n49569 , n49563 , n49568 );
buf ( n49570 , n49569 );
xor ( n49571 , n49559 , n49570 );
buf ( n49572 , n41647 );
not ( n49573 , n49572 );
buf ( n49574 , n41666 );
not ( n49575 , n49574 );
buf ( n49576 , n37081 );
not ( n49577 , n49576 );
or ( n49578 , n49575 , n49577 );
nand ( n49579 , n40089 , n41663 );
buf ( n49580 , n49579 );
nand ( n49581 , n49578 , n49580 );
buf ( n49582 , n49581 );
buf ( n49583 , n49582 );
not ( n49584 , n49583 );
or ( n49585 , n49573 , n49584 );
buf ( n49586 , n41678 );
buf ( n49587 , n41705 );
nand ( n49588 , n49586 , n49587 );
buf ( n49589 , n49588 );
buf ( n49590 , n49589 );
nand ( n49591 , n49585 , n49590 );
buf ( n49592 , n49591 );
buf ( n49593 , n49592 );
xor ( n49594 , n49571 , n49593 );
buf ( n49595 , n49594 );
buf ( n49596 , n49595 );
buf ( n49597 , n43609 );
not ( n49598 , n49597 );
buf ( n49599 , n43827 );
not ( n49600 , n49599 );
or ( n49601 , n49598 , n49600 );
buf ( n49602 , n43672 );
nand ( n49603 , n49601 , n49602 );
buf ( n49604 , n49603 );
buf ( n49605 , n49604 );
buf ( n49606 , n43827 );
buf ( n49607 , n43609 );
or ( n49608 , n49606 , n49607 );
buf ( n49609 , n49608 );
buf ( n49610 , n49609 );
nand ( n49611 , n49605 , n49610 );
buf ( n49612 , n49611 );
buf ( n49613 , n49612 );
xor ( n49614 , n49596 , n49613 );
xor ( n49615 , n43760 , n43794 );
and ( n49616 , n49615 , n43822 );
and ( n49617 , n43760 , n43794 );
or ( n49618 , n49616 , n49617 );
buf ( n49619 , n49618 );
buf ( n49620 , n49619 );
buf ( n49621 , n38985 );
not ( n49622 , n49621 );
buf ( n49623 , n43691 );
not ( n49624 , n49623 );
or ( n49625 , n49622 , n49624 );
buf ( n49626 , n39000 );
not ( n49627 , n49626 );
buf ( n49628 , n39518 );
not ( n49629 , n49628 );
or ( n49630 , n49627 , n49629 );
buf ( n49631 , n39522 );
buf ( n49632 , n38997 );
nand ( n49633 , n49631 , n49632 );
buf ( n49634 , n49633 );
buf ( n49635 , n49634 );
nand ( n49636 , n49630 , n49635 );
buf ( n49637 , n49636 );
buf ( n49638 , n49637 );
buf ( n49639 , n42448 );
nand ( n49640 , n49638 , n49639 );
buf ( n49641 , n49640 );
buf ( n49642 , n49641 );
nand ( n49643 , n49625 , n49642 );
buf ( n49644 , n49643 );
buf ( n49645 , n49644 );
xor ( n49646 , n49620 , n49645 );
xor ( n49647 , n45265 , n45282 );
and ( n49648 , n49647 , n45311 );
and ( n49649 , n45265 , n45282 );
or ( n49650 , n49648 , n49649 );
buf ( n49651 , n49650 );
buf ( n49652 , n49651 );
xor ( n49653 , n49646 , n49652 );
buf ( n49654 , n49653 );
buf ( n49655 , n42339 );
not ( n49656 , n49655 );
and ( n49657 , n42343 , n36430 );
not ( n49658 , n42343 );
and ( n49659 , n49658 , n36427 );
or ( n49660 , n49657 , n49659 );
buf ( n49661 , n49660 );
not ( n49662 , n49661 );
or ( n49663 , n49656 , n49662 );
buf ( n49664 , n43598 );
buf ( n49665 , n42378 );
nand ( n49666 , n49664 , n49665 );
buf ( n49667 , n49666 );
buf ( n49668 , n49667 );
nand ( n49669 , n49663 , n49668 );
buf ( n49670 , n49669 );
xor ( n49671 , n49654 , n49670 );
xor ( n49672 , n45245 , n45314 );
and ( n49673 , n49672 , n45321 );
and ( n49674 , n45245 , n45314 );
or ( n49675 , n49673 , n49674 );
buf ( n49676 , n49675 );
xor ( n49677 , n49671 , n49676 );
buf ( n49678 , n49677 );
xor ( n49679 , n49614 , n49678 );
buf ( n49680 , n49679 );
buf ( n49681 , n49680 );
xor ( n49682 , n49542 , n49681 );
buf ( n49683 , n49682 );
xnor ( n49684 , n49529 , n49683 );
buf ( n49685 , n49684 );
xnor ( n49686 , n49154 , n49685 );
buf ( n49687 , n49686 );
buf ( n49688 , n49687 );
nand ( n49689 , n49138 , n49688 );
buf ( n49690 , n49689 );
buf ( n49691 , n49690 );
and ( n49692 , n47225 , n48103 , n49130 , n49691 );
buf ( n49693 , n49692 );
xor ( n49694 , n49071 , n49108 );
buf ( n49695 , n49084 );
xnor ( n49696 , n49694 , n49695 );
buf ( n49697 , n48562 );
not ( n49698 , n49697 );
buf ( n49699 , n48149 );
not ( n49700 , n49699 );
or ( n49701 , n49698 , n49700 );
buf ( n49702 , n48146 );
buf ( n49703 , n48562 );
not ( n49704 , n49703 );
buf ( n49705 , n49704 );
buf ( n49706 , n49705 );
nand ( n49707 , n49702 , n49706 );
buf ( n49708 , n49707 );
buf ( n49709 , n49708 );
nand ( n49710 , n49701 , n49709 );
buf ( n49711 , n49710 );
and ( n49712 , n49711 , n48156 );
not ( n49713 , n49711 );
and ( n49714 , n49713 , n48159 );
nor ( n49715 , n49712 , n49714 );
not ( n49716 , n47360 );
not ( n49717 , n47355 );
not ( n49718 , n47326 );
or ( n49719 , n49717 , n49718 );
not ( n49720 , n47355 );
nand ( n49721 , n49720 , n47327 );
nand ( n49722 , n49719 , n49721 );
xor ( n49723 , n49716 , n49722 );
buf ( n49724 , n49723 );
not ( n49725 , n49724 );
buf ( n49726 , n49725 );
not ( n49727 , n49726 );
buf ( n49728 , n46390 );
not ( n49729 , n49728 );
buf ( n49730 , n38468 );
not ( n49731 , n49730 );
or ( n49732 , n49729 , n49731 );
buf ( n49733 , n36527 );
buf ( n49734 , n46393 );
nand ( n49735 , n49733 , n49734 );
buf ( n49736 , n49735 );
buf ( n49737 , n49736 );
nand ( n49738 , n49732 , n49737 );
buf ( n49739 , n49738 );
buf ( n49740 , n49739 );
not ( n49741 , n49740 );
buf ( n49742 , n44135 );
not ( n49743 , n49742 );
or ( n49744 , n49741 , n49743 );
buf ( n49745 , n36640 );
not ( n49746 , n49745 );
buf ( n49747 , n48247 );
nand ( n49748 , n49746 , n49747 );
buf ( n49749 , n49748 );
buf ( n49750 , n49749 );
nand ( n49751 , n49744 , n49750 );
buf ( n49752 , n49751 );
buf ( n49753 , n49752 );
not ( n49754 , n49753 );
buf ( n49755 , n42865 );
not ( n49756 , n49755 );
buf ( n49757 , n42082 );
not ( n49758 , n49757 );
or ( n49759 , n49756 , n49758 );
buf ( n49760 , n42062 );
buf ( n49761 , n42862 );
nand ( n49762 , n49760 , n49761 );
buf ( n49763 , n49762 );
buf ( n49764 , n49763 );
nand ( n49765 , n49759 , n49764 );
buf ( n49766 , n49765 );
buf ( n49767 , n49766 );
not ( n49768 , n49767 );
buf ( n49769 , n45155 );
not ( n49770 , n49769 );
or ( n49771 , n49768 , n49770 );
not ( n49772 , n36909 );
nand ( n49773 , n49772 , n48034 );
buf ( n49774 , n49773 );
nand ( n49775 , n49771 , n49774 );
buf ( n49776 , n49775 );
buf ( n49777 , n49776 );
not ( n49778 , n49777 );
or ( n49779 , n49754 , n49778 );
buf ( n49780 , n49776 );
buf ( n49781 , n49752 );
or ( n49782 , n49780 , n49781 );
xor ( n49783 , n47043 , n48227 );
xnor ( n49784 , n49783 , n48218 );
buf ( n49785 , n49784 );
nand ( n49786 , n49782 , n49785 );
buf ( n49787 , n49786 );
buf ( n49788 , n49787 );
nand ( n49789 , n49779 , n49788 );
buf ( n49790 , n49789 );
buf ( n49791 , n49790 );
xor ( n49792 , n48234 , n48261 );
xor ( n49793 , n49792 , n48283 );
buf ( n49794 , n49793 );
buf ( n49795 , n49794 );
xor ( n49796 , n49791 , n49795 );
buf ( n49797 , n41608 );
not ( n49798 , n49797 );
buf ( n49799 , n42926 );
not ( n49800 , n49799 );
or ( n49801 , n49798 , n49800 );
buf ( n49802 , n37968 );
buf ( n49803 , n49802 );
buf ( n49804 , n49803 );
buf ( n49805 , n49804 );
buf ( n49806 , n41611 );
nand ( n49807 , n49805 , n49806 );
buf ( n49808 , n49807 );
buf ( n49809 , n49808 );
nand ( n49810 , n49801 , n49809 );
buf ( n49811 , n49810 );
not ( n49812 , n49811 );
not ( n49813 , n44267 );
or ( n49814 , n49812 , n49813 );
or ( n49815 , n48522 , n41577 );
nand ( n49816 , n49814 , n49815 );
buf ( n49817 , n49816 );
and ( n49818 , n49796 , n49817 );
and ( n49819 , n49791 , n49795 );
or ( n49820 , n49818 , n49819 );
buf ( n49821 , n49820 );
not ( n49822 , n49821 );
or ( n49823 , n49727 , n49822 );
buf ( n49824 , n49723 );
not ( n49825 , n49824 );
buf ( n49826 , n49821 );
not ( n49827 , n49826 );
buf ( n49828 , n49827 );
buf ( n49829 , n49828 );
not ( n49830 , n49829 );
or ( n49831 , n49825 , n49830 );
buf ( n49832 , n48409 );
buf ( n49833 , n48429 );
xor ( n49834 , n49832 , n49833 );
buf ( n49835 , n48380 );
xor ( n49836 , n49834 , n49835 );
buf ( n49837 , n49836 );
buf ( n49838 , n49837 );
not ( n49839 , n49838 );
buf ( n49840 , n49839 );
buf ( n49841 , n49840 );
not ( n49842 , n49841 );
buf ( n49843 , n42378 );
not ( n49844 , n49843 );
buf ( n49845 , n42343 );
not ( n49846 , n49845 );
buf ( n49847 , n42795 );
not ( n49848 , n49847 );
or ( n49849 , n49846 , n49848 );
buf ( n49850 , n37783 );
buf ( n49851 , n46855 );
nand ( n49852 , n49850 , n49851 );
buf ( n49853 , n49852 );
buf ( n49854 , n49853 );
nand ( n49855 , n49849 , n49854 );
buf ( n49856 , n49855 );
buf ( n49857 , n49856 );
not ( n49858 , n49857 );
or ( n49859 , n49844 , n49858 );
buf ( n49860 , n48419 );
not ( n49861 , n49860 );
buf ( n49862 , n42339 );
nand ( n49863 , n49861 , n49862 );
buf ( n49864 , n49863 );
buf ( n49865 , n49864 );
nand ( n49866 , n49859 , n49865 );
buf ( n49867 , n49866 );
buf ( n49868 , n49867 );
buf ( n49869 , n41905 );
buf ( n49870 , n48306 );
nand ( n49871 , n49869 , n49870 );
buf ( n49872 , n49871 );
buf ( n49873 , n42017 );
buf ( n49874 , n41889 );
and ( n49875 , n49873 , n49874 );
not ( n49876 , n49873 );
buf ( n49877 , n37881 );
not ( n49878 , n49877 );
buf ( n49879 , n49878 );
buf ( n49880 , n49879 );
and ( n49881 , n49876 , n49880 );
nor ( n49882 , n49875 , n49881 );
buf ( n49883 , n49882 );
not ( n49884 , n49883 );
nand ( n49885 , n49884 , n41862 );
nand ( n49886 , n49872 , n49885 );
buf ( n49887 , n49886 );
buf ( n49888 , n41736 );
not ( n49889 , n49888 );
buf ( n49890 , n48207 );
not ( n49891 , n49890 );
or ( n49892 , n49889 , n49891 );
buf ( n49893 , n41748 );
buf ( n49894 , n37473 );
nand ( n49895 , n49893 , n49894 );
buf ( n49896 , n49895 );
buf ( n49897 , n49896 );
nand ( n49898 , n49892 , n49897 );
buf ( n49899 , n49898 );
not ( n49900 , n49899 );
not ( n49901 , n44338 );
or ( n49902 , n49900 , n49901 );
buf ( n49903 , n48211 );
not ( n49904 , n49903 );
buf ( n49905 , n41852 );
nand ( n49906 , n49904 , n49905 );
buf ( n49907 , n49906 );
nand ( n49908 , n49902 , n49907 );
buf ( n49909 , n49908 );
or ( n49910 , n49887 , n49909 );
buf ( n49911 , n43250 );
not ( n49912 , n49911 );
buf ( n49913 , n46117 );
not ( n49914 , n49913 );
buf ( n49915 , n43259 );
not ( n49916 , n49915 );
or ( n49917 , n49914 , n49916 );
buf ( n49918 , n43503 );
buf ( n49919 , n46126 );
nand ( n49920 , n49918 , n49919 );
buf ( n49921 , n49920 );
buf ( n49922 , n49921 );
nand ( n49923 , n49917 , n49922 );
buf ( n49924 , n49923 );
buf ( n49925 , n49924 );
not ( n49926 , n49925 );
or ( n49927 , n49912 , n49926 );
buf ( n49928 , n42834 );
buf ( n49929 , n49025 );
nand ( n49930 , n49928 , n49929 );
buf ( n49931 , n49930 );
buf ( n49932 , n49931 );
nand ( n49933 , n49927 , n49932 );
buf ( n49934 , n49933 );
buf ( n49935 , n49934 );
nand ( n49936 , n49910 , n49935 );
buf ( n49937 , n49936 );
buf ( n49938 , n49937 );
not ( n49939 , n49885 );
not ( n49940 , n49872 );
or ( n49941 , n49939 , n49940 );
not ( n49942 , n49899 );
not ( n49943 , n44338 );
or ( n49944 , n49942 , n49943 );
nand ( n49945 , n49944 , n49907 );
nand ( n49946 , n49941 , n49945 );
buf ( n49947 , n49946 );
nand ( n49948 , n49938 , n49947 );
buf ( n49949 , n49948 );
buf ( n49950 , n49949 );
xor ( n49951 , n49868 , n49950 );
buf ( n49952 , n42668 );
not ( n49953 , n49952 );
buf ( n49954 , n48919 );
not ( n49955 , n49954 );
or ( n49956 , n49953 , n49955 );
buf ( n49957 , n42672 );
not ( n49958 , n49957 );
buf ( n49959 , n37714 );
not ( n49960 , n49959 );
or ( n49961 , n49958 , n49960 );
buf ( n49962 , n43625 );
buf ( n49963 , n42671 );
nand ( n49964 , n49962 , n49963 );
buf ( n49965 , n49964 );
buf ( n49966 , n49965 );
nand ( n49967 , n49961 , n49966 );
buf ( n49968 , n49967 );
buf ( n49969 , n49968 );
buf ( n49970 , n42712 );
nand ( n49971 , n49969 , n49970 );
buf ( n49972 , n49971 );
buf ( n49973 , n49972 );
nand ( n49974 , n49956 , n49973 );
buf ( n49975 , n49974 );
buf ( n49976 , n49975 );
and ( n49977 , n49951 , n49976 );
and ( n49978 , n49868 , n49950 );
or ( n49979 , n49977 , n49978 );
buf ( n49980 , n49979 );
buf ( n49981 , n49980 );
not ( n49982 , n49981 );
or ( n49983 , n49842 , n49982 );
buf ( n49984 , n49837 );
not ( n49985 , n49984 );
buf ( n49986 , n49980 );
not ( n49987 , n49986 );
buf ( n49988 , n49987 );
buf ( n49989 , n49988 );
not ( n49990 , n49989 );
or ( n49991 , n49985 , n49990 );
xor ( n49992 , n48375 , n48316 );
xor ( n49993 , n49992 , n48342 );
buf ( n49994 , n49993 );
not ( n49995 , n49994 );
buf ( n49996 , n44267 );
not ( n49997 , n49996 );
buf ( n49998 , n41611 );
not ( n49999 , n49998 );
buf ( n50000 , n42941 );
not ( n50001 , n50000 );
or ( n50002 , n49999 , n50001 );
buf ( n50003 , n47969 );
not ( n50004 , n50003 );
buf ( n50005 , n41608 );
nand ( n50006 , n50004 , n50005 );
buf ( n50007 , n50006 );
buf ( n50008 , n50007 );
nand ( n50009 , n50002 , n50008 );
buf ( n50010 , n50009 );
buf ( n50011 , n50010 );
not ( n50012 , n50011 );
or ( n50013 , n49997 , n50012 );
buf ( n50014 , n49811 );
buf ( n50015 , n43868 );
nand ( n50016 , n50014 , n50015 );
buf ( n50017 , n50016 );
buf ( n50018 , n50017 );
nand ( n50019 , n50013 , n50018 );
buf ( n50020 , n50019 );
buf ( n50021 , n50020 );
not ( n50022 , n50021 );
or ( n50023 , n49995 , n50022 );
buf ( n50024 , n50020 );
buf ( n50025 , n49993 );
or ( n50026 , n50024 , n50025 );
buf ( n50027 , n46294 );
not ( n50028 , n50027 );
buf ( n50029 , n48365 );
not ( n50030 , n50029 );
or ( n50031 , n50028 , n50030 );
buf ( n50032 , n43938 );
buf ( n50033 , n25182 );
not ( n50034 , n50033 );
buf ( n50035 , n39671 );
not ( n50036 , n50035 );
or ( n50037 , n50034 , n50036 );
buf ( n50038 , n29269 );
not ( n50039 , n50038 );
buf ( n50040 , n50039 );
buf ( n50041 , n50040 );
not ( n50042 , n50041 );
buf ( n50043 , n50042 );
buf ( n50044 , n50043 );
not ( n50045 , n48357 );
buf ( n50046 , n50045 );
nand ( n50047 , n50044 , n50046 );
buf ( n50048 , n50047 );
buf ( n50049 , n50048 );
nand ( n50050 , n50037 , n50049 );
buf ( n50051 , n50050 );
buf ( n50052 , n50051 );
nand ( n50053 , n50032 , n50052 );
buf ( n50054 , n50053 );
buf ( n50055 , n50054 );
nand ( n50056 , n50031 , n50055 );
buf ( n50057 , n50056 );
buf ( n50058 , n50057 );
and ( n50059 , n25893 , n25895 , n25898 , n25899 );
not ( n50060 , n50059 );
buf ( n50061 , n50060 );
not ( n50062 , n50061 );
buf ( n50063 , n37602 );
not ( n50064 , n50063 );
or ( n50065 , n50062 , n50064 );
buf ( n50066 , n38834 );
not ( n50067 , n50060 );
buf ( n50068 , n50067 );
nand ( n50069 , n50066 , n50068 );
buf ( n50070 , n50069 );
buf ( n50071 , n50070 );
nand ( n50072 , n50065 , n50071 );
buf ( n50073 , n50072 );
buf ( n50074 , n36444 );
buf ( n50075 , n48335 );
nand ( n50076 , n50074 , n50075 );
buf ( n50077 , n50076 );
buf ( n50078 , n50077 );
nand ( n50079 , C1 , n50078 );
buf ( n50080 , n50079 );
buf ( n50081 , n50080 );
xor ( n50082 , n50058 , n50081 );
buf ( n50083 , n42152 );
not ( n50084 , n50083 );
buf ( n50085 , n38994 );
not ( n50086 , n50085 );
or ( n50087 , n50084 , n50086 );
buf ( n50088 , n38979 );
buf ( n50089 , n42149 );
not ( n50090 , n50089 );
buf ( n50091 , n50090 );
buf ( n50092 , n50091 );
nand ( n50093 , n50088 , n50092 );
buf ( n50094 , n50093 );
buf ( n50095 , n50094 );
nand ( n50096 , n50087 , n50095 );
buf ( n50097 , n50096 );
buf ( n50098 , n50097 );
not ( n50099 , n50098 );
buf ( n50100 , n47050 );
not ( n50101 , n50100 );
or ( n50102 , n50099 , n50101 );
buf ( n50103 , n48955 );
not ( n50104 , n38973 );
buf ( n50105 , n50104 );
nand ( n50106 , n50103 , n50105 );
buf ( n50107 , n50106 );
buf ( n50108 , n50107 );
nand ( n50109 , n50102 , n50108 );
buf ( n50110 , n50109 );
buf ( n50111 , n50110 );
not ( n50112 , n50111 );
buf ( n50113 , n42578 );
not ( n50114 , n50113 );
buf ( n50115 , n41835 );
not ( n50116 , n50115 );
or ( n50117 , n50114 , n50116 );
buf ( n50118 , n28306 );
buf ( n50119 , n46356 );
nand ( n50120 , n50118 , n50119 );
buf ( n50121 , n50120 );
buf ( n50122 , n50121 );
nand ( n50123 , n50117 , n50122 );
buf ( n50124 , n50123 );
buf ( n50125 , n50124 );
buf ( n50126 , n42622 );
not ( n50127 , n50126 );
buf ( n50128 , n50127 );
buf ( n50129 , n50128 );
and ( n50130 , n50125 , n50129 );
buf ( n50131 , n48723 );
buf ( n50132 , n42565 );
nor ( n50133 , n50131 , n50132 );
buf ( n50134 , n50133 );
buf ( n50135 , n50134 );
nor ( n50136 , n50130 , n50135 );
buf ( n50137 , n50136 );
buf ( n50138 , n50137 );
not ( n50139 , n50138 );
buf ( n50140 , n50139 );
buf ( n50141 , n50140 );
not ( n50142 , n50141 );
or ( n50143 , n50112 , n50142 );
buf ( n50144 , n50110 );
not ( n50145 , n50144 );
buf ( n50146 , n50145 );
buf ( n50147 , n50146 );
not ( n50148 , n50147 );
buf ( n50149 , n50137 );
not ( n50150 , n50149 );
or ( n50151 , n50148 , n50150 );
not ( n50152 , n38404 );
buf ( n50153 , n42411 );
not ( n50154 , n50153 );
buf ( n50155 , n42072 );
not ( n50156 , n50155 );
and ( n50157 , n50154 , n50156 );
buf ( n50158 , n48984 );
buf ( n50159 , n42072 );
and ( n50160 , n50158 , n50159 );
nor ( n50161 , n50157 , n50160 );
buf ( n50162 , n50161 );
not ( n50163 , n50162 );
not ( n50164 , n50163 );
or ( n50165 , n50152 , n50164 );
buf ( n50166 , n48994 );
not ( n50167 , n50166 );
buf ( n50168 , n38382 );
nand ( n50169 , n50167 , n50168 );
buf ( n50170 , n50169 );
nand ( n50171 , n50165 , n50170 );
buf ( n50172 , n50171 );
nand ( n50173 , n50151 , n50172 );
buf ( n50174 , n50173 );
buf ( n50175 , n50174 );
nand ( n50176 , n50143 , n50175 );
buf ( n50177 , n50176 );
buf ( n50178 , n50177 );
and ( n50179 , n50082 , n50178 );
and ( n50180 , n50058 , n50081 );
or ( n50181 , n50179 , n50180 );
buf ( n50182 , n50181 );
buf ( n50183 , n50182 );
nand ( n50184 , n50026 , n50183 );
buf ( n50185 , n50184 );
buf ( n50186 , n50185 );
nand ( n50187 , n50023 , n50186 );
buf ( n50188 , n50187 );
buf ( n50189 , n50188 );
nand ( n50190 , n49991 , n50189 );
buf ( n50191 , n50190 );
buf ( n50192 , n50191 );
nand ( n50193 , n49983 , n50192 );
buf ( n50194 , n50193 );
buf ( n50195 , n50194 );
nand ( n50196 , n49831 , n50195 );
buf ( n50197 , n50196 );
nand ( n50198 , n49823 , n50197 );
not ( n50199 , n50198 );
not ( n50200 , n48550 );
not ( n50201 , n48483 );
not ( n50202 , n48466 );
or ( n50203 , n50201 , n50202 );
or ( n50204 , n48483 , n48466 );
nand ( n50205 , n50203 , n50204 );
not ( n50206 , n50205 );
or ( n50207 , n50200 , n50206 );
or ( n50208 , n48550 , n50205 );
nand ( n50209 , n50207 , n50208 );
nand ( n50210 , n50199 , n50209 );
not ( n50211 , n50210 );
xor ( n50212 , n48588 , n48800 );
xor ( n50213 , n50212 , n49066 );
buf ( n50214 , n50213 );
not ( n50215 , n50214 );
or ( n50216 , n50211 , n50215 );
not ( n50217 , n50209 );
nand ( n50218 , n50217 , n50198 );
nand ( n50219 , n50216 , n50218 );
and ( n50220 , n49715 , n50219 );
not ( n50221 , n49715 );
buf ( n50222 , n50219 );
not ( n50223 , n50222 );
buf ( n50224 , n50223 );
and ( n50225 , n50221 , n50224 );
nor ( n50226 , n50220 , n50225 );
xor ( n50227 , n48510 , n48532 );
xnor ( n50228 , n50227 , n48544 );
not ( n50229 , n50228 );
xor ( n50230 , n48287 , n48449 );
xnor ( n50231 , n50230 , n48455 );
buf ( n50232 , n50231 );
buf ( n50233 , n50232 );
buf ( n50234 , n50233 );
not ( n50235 , n50234 );
or ( n50236 , n50229 , n50235 );
buf ( n50237 , n50234 );
buf ( n50238 , n50228 );
or ( n50239 , n50237 , n50238 );
xor ( n50240 , n48626 , n48763 );
xor ( n50241 , n50240 , n48789 );
buf ( n50242 , n50241 );
not ( n50243 , n50242 );
buf ( n50244 , n46225 );
not ( n50245 , n50244 );
buf ( n50246 , n45753 );
not ( n50247 , n50246 );
buf ( n50248 , n40067 );
not ( n50249 , n50248 );
or ( n50250 , n50247 , n50249 );
buf ( n50251 , n36427 );
buf ( n50252 , n45750 );
nand ( n50253 , n50251 , n50252 );
buf ( n50254 , n50253 );
buf ( n50255 , n50254 );
nand ( n50256 , n50250 , n50255 );
buf ( n50257 , n50256 );
buf ( n50258 , n50257 );
not ( n50259 , n50258 );
or ( n50260 , n50245 , n50259 );
buf ( n50261 , n45730 );
not ( n50262 , n50261 );
buf ( n50263 , n48500 );
nand ( n50264 , n50262 , n50263 );
buf ( n50265 , n50264 );
buf ( n50266 , n50265 );
nand ( n50267 , n50260 , n50266 );
buf ( n50268 , n50267 );
buf ( n50269 , n44496 );
not ( n50270 , n50269 );
buf ( n50271 , n48607 );
not ( n50272 , n50271 );
or ( n50273 , n50270 , n50272 );
buf ( n50274 , n44533 );
not ( n50275 , n50274 );
buf ( n50276 , n38098 );
not ( n50277 , n50276 );
or ( n50278 , n50275 , n50277 );
buf ( n50279 , n37081 );
not ( n50280 , n50279 );
buf ( n50281 , n44530 );
nand ( n50282 , n50280 , n50281 );
buf ( n50283 , n50282 );
buf ( n50284 , n50283 );
nand ( n50285 , n50278 , n50284 );
buf ( n50286 , n50285 );
buf ( n50287 , n50286 );
buf ( n50288 , n44708 );
nand ( n50289 , n50287 , n50288 );
buf ( n50290 , n50289 );
buf ( n50291 , n50290 );
nand ( n50292 , n50273 , n50291 );
buf ( n50293 , n50292 );
or ( n50294 , n50268 , n50293 );
not ( n50295 , n50294 );
or ( n50296 , n50243 , n50295 );
buf ( n50297 , n50268 );
buf ( n50298 , n50293 );
nand ( n50299 , n50297 , n50298 );
buf ( n50300 , n50299 );
nand ( n50301 , n50296 , n50300 );
buf ( n50302 , n50301 );
nand ( n50303 , n50239 , n50302 );
buf ( n50304 , n50303 );
nand ( n50305 , n50236 , n50304 );
not ( n50306 , n50305 );
not ( n50307 , n49094 );
not ( n50308 , n49089 );
not ( n50309 , n50308 );
or ( n50310 , n50307 , n50309 );
nand ( n50311 , n49089 , n49095 );
nand ( n50312 , n50310 , n50311 );
xor ( n50313 , n49098 , n49100 );
and ( n50314 , n50312 , n50313 );
not ( n50315 , n50312 );
and ( n50316 , n50315 , n49104 );
nor ( n50317 , n50314 , n50316 );
not ( n50318 , n50317 );
not ( n50319 , n50318 );
or ( n50320 , n50306 , n50319 );
not ( n50321 , n50305 );
not ( n50322 , n50321 );
not ( n50323 , n50317 );
or ( n50324 , n50322 , n50323 );
buf ( n50325 , n48591 );
buf ( n50326 , n48617 );
xor ( n50327 , n50325 , n50326 );
buf ( n50328 , n48793 );
xor ( n50329 , n50327 , n50328 );
buf ( n50330 , n50329 );
buf ( n50331 , n50330 );
buf ( n50332 , n47331 );
not ( n50333 , n50332 );
buf ( n50334 , n46875 );
not ( n50335 , n50334 );
buf ( n50336 , n42277 );
not ( n50337 , n50336 );
or ( n50338 , n50335 , n50337 );
buf ( n50339 , n39924 );
buf ( n50340 , n46887 );
nand ( n50341 , n50339 , n50340 );
buf ( n50342 , n50341 );
buf ( n50343 , n50342 );
nand ( n50344 , n50338 , n50343 );
buf ( n50345 , n50344 );
buf ( n50346 , n50345 );
not ( n50347 , n50346 );
or ( n50348 , n50333 , n50347 );
buf ( n50349 , n48895 );
buf ( n50350 , n46912 );
nand ( n50351 , n50349 , n50350 );
buf ( n50352 , n50351 );
buf ( n50353 , n50352 );
nand ( n50354 , n50348 , n50353 );
buf ( n50355 , n50354 );
buf ( n50356 , n50355 );
not ( n50357 , n50356 );
xor ( n50358 , n48708 , n48732 );
xor ( n50359 , n50358 , n48752 );
buf ( n50360 , n50359 );
buf ( n50361 , n50360 );
not ( n50362 , n47716 );
not ( n50363 , n41741 );
or ( n50364 , n50362 , n50363 );
buf ( n50365 , n36527 );
buf ( n50366 , n47725 );
nand ( n50367 , n50365 , n50366 );
buf ( n50368 , n50367 );
nand ( n50369 , n50364 , n50368 );
buf ( n50370 , n50369 );
not ( n50371 , n50370 );
buf ( n50372 , n36520 );
not ( n50373 , n50372 );
buf ( n50374 , n50373 );
buf ( n50375 , n50374 );
not ( n50376 , n50375 );
or ( n50377 , n50371 , n50376 );
buf ( n50378 , n43982 );
buf ( n50379 , n49739 );
nand ( n50380 , n50378 , n50379 );
buf ( n50381 , n50380 );
buf ( n50382 , n50381 );
nand ( n50383 , n50377 , n50382 );
buf ( n50384 , n50383 );
buf ( n50385 , n50384 );
xor ( n50386 , n50361 , n50385 );
buf ( n50387 , n42339 );
not ( n50388 , n50387 );
buf ( n50389 , n49856 );
not ( n50390 , n50389 );
or ( n50391 , n50388 , n50390 );
buf ( n50392 , n42343 );
not ( n50393 , n50392 );
buf ( n50394 , n42991 );
not ( n50395 , n50394 );
or ( n50396 , n50393 , n50395 );
buf ( n50397 , n44163 );
buf ( n50398 , n46855 );
nand ( n50399 , n50397 , n50398 );
buf ( n50400 , n50399 );
buf ( n50401 , n50400 );
nand ( n50402 , n50396 , n50401 );
buf ( n50403 , n50402 );
buf ( n50404 , n50403 );
buf ( n50405 , n42378 );
nand ( n50406 , n50404 , n50405 );
buf ( n50407 , n50406 );
buf ( n50408 , n50407 );
nand ( n50409 , n50391 , n50408 );
buf ( n50410 , n50409 );
buf ( n50411 , n50410 );
and ( n50412 , n50386 , n50411 );
and ( n50413 , n50361 , n50385 );
or ( n50414 , n50412 , n50413 );
buf ( n50415 , n50414 );
buf ( n50416 , n50415 );
not ( n50417 , n50416 );
or ( n50418 , n50357 , n50417 );
buf ( n50419 , n50355 );
buf ( n50420 , n50415 );
or ( n50421 , n50419 , n50420 );
xor ( n50422 , n49784 , n49752 );
xor ( n50423 , n50422 , n49776 );
buf ( n50424 , n50423 );
nand ( n50425 , n50421 , n50424 );
buf ( n50426 , n50425 );
buf ( n50427 , n50426 );
nand ( n50428 , n50418 , n50427 );
buf ( n50429 , n50428 );
not ( n50430 , n50429 );
buf ( n50431 , n48868 );
not ( n50432 , n50431 );
buf ( n50433 , n48827 );
not ( n50434 , n50433 );
or ( n50435 , n50432 , n50434 );
buf ( n50436 , n48808 );
not ( n50437 , n50436 );
buf ( n50438 , n43857 );
not ( n50439 , n50438 );
or ( n50440 , n50437 , n50439 );
buf ( n50441 , n36051 );
buf ( n50442 , n48818 );
nand ( n50443 , n50441 , n50442 );
buf ( n50444 , n50443 );
buf ( n50445 , n50444 );
nand ( n50446 , n50440 , n50445 );
buf ( n50447 , n50446 );
buf ( n50448 , n50447 );
buf ( n50449 , n48855 );
nand ( n50450 , n50448 , n50449 );
buf ( n50451 , n50450 );
buf ( n50452 , n50451 );
nand ( n50453 , n50435 , n50452 );
buf ( n50454 , n50453 );
not ( n50455 , n50454 );
buf ( n50456 , n42252 );
not ( n50457 , n50456 );
buf ( n50458 , n42266 );
not ( n50459 , n50458 );
buf ( n50460 , n43879 );
not ( n50461 , n50460 );
or ( n50462 , n50459 , n50461 );
not ( n50463 , n38742 );
buf ( n50464 , n50463 );
buf ( n50465 , n42263 );
nand ( n50466 , n50464 , n50465 );
buf ( n50467 , n50466 );
buf ( n50468 , n50467 );
nand ( n50469 , n50462 , n50468 );
buf ( n50470 , n50469 );
buf ( n50471 , n50470 );
not ( n50472 , n50471 );
or ( n50473 , n50457 , n50472 );
buf ( n50474 , n48781 );
buf ( n50475 , n42315 );
nand ( n50476 , n50474 , n50475 );
buf ( n50477 , n50476 );
buf ( n50478 , n50477 );
nand ( n50479 , n50473 , n50478 );
buf ( n50480 , n50479 );
buf ( n50481 , n50480 );
not ( n50482 , n50481 );
buf ( n50483 , n50482 );
nand ( n50484 , n50455 , n50483 );
not ( n50485 , n50484 );
buf ( n50486 , n42847 );
buf ( n50487 , n42062 );
and ( n50488 , n50486 , n50487 );
not ( n50489 , n50486 );
buf ( n50490 , n42082 );
and ( n50491 , n50489 , n50490 );
nor ( n50492 , n50488 , n50491 );
buf ( n50493 , n50492 );
buf ( n50494 , n50493 );
not ( n50495 , n50494 );
buf ( n50496 , n44776 );
not ( n50497 , n50496 );
or ( n50498 , n50495 , n50497 );
buf ( n50499 , n44676 );
buf ( n50500 , n49766 );
nand ( n50501 , n50499 , n50500 );
buf ( n50502 , n50501 );
buf ( n50503 , n50502 );
nand ( n50504 , n50498 , n50503 );
buf ( n50505 , n50504 );
not ( n50506 , n50505 );
not ( n50507 , n50506 );
buf ( n50508 , n50507 );
not ( n50509 , n50508 );
buf ( n50510 , n43063 );
not ( n50511 , n50510 );
buf ( n50512 , n47898 );
not ( n50513 , n50512 );
or ( n50514 , n50511 , n50513 );
buf ( n50515 , n38108 );
buf ( n50516 , n43064 );
nand ( n50517 , n50515 , n50516 );
buf ( n50518 , n50517 );
buf ( n50519 , n50518 );
nand ( n50520 , n50514 , n50519 );
buf ( n50521 , n50520 );
buf ( n50522 , n50521 );
not ( n50523 , n50522 );
buf ( n50524 , n43386 );
not ( n50525 , n50524 );
or ( n50526 , n50523 , n50525 );
buf ( n50527 , n48638 );
buf ( n50528 , n45144 );
nand ( n50529 , n50527 , n50528 );
buf ( n50530 , n50529 );
buf ( n50531 , n50530 );
nand ( n50532 , n50526 , n50531 );
buf ( n50533 , n50532 );
buf ( n50534 , n50533 );
not ( n50535 , n50534 );
or ( n50536 , n50509 , n50535 );
buf ( n50537 , n50533 );
not ( n50538 , n50537 );
buf ( n50539 , n50538 );
buf ( n50540 , n50539 );
not ( n50541 , n50540 );
buf ( n50542 , n50506 );
not ( n50543 , n50542 );
or ( n50544 , n50541 , n50543 );
buf ( n50545 , n41993 );
not ( n50546 , n50545 );
buf ( n50547 , n41894 );
not ( n50548 , n50547 );
or ( n50549 , n50546 , n50548 );
buf ( n50550 , n41889 );
buf ( n50551 , n43966 );
nand ( n50552 , n50550 , n50551 );
buf ( n50553 , n50552 );
buf ( n50554 , n50553 );
nand ( n50555 , n50549 , n50554 );
buf ( n50556 , n50555 );
buf ( n50557 , n50556 );
not ( n50558 , n50557 );
buf ( n50559 , n37872 );
not ( n50560 , n50559 );
or ( n50561 , n50558 , n50560 );
buf ( n50562 , n49883 );
not ( n50563 , n50562 );
buf ( n50564 , n45617 );
nand ( n50565 , n50563 , n50564 );
buf ( n50566 , n50565 );
buf ( n50567 , n50566 );
nand ( n50568 , n50561 , n50567 );
buf ( n50569 , n50568 );
not ( n50570 , n50569 );
not ( n50571 , n48705 );
not ( n50572 , n24092 );
buf ( n50573 , n41870 );
buf ( n50574 , n50573 );
buf ( n50575 , n50574 );
buf ( n50576 , n50575 );
not ( n50577 , n50576 );
buf ( n50578 , n50577 );
not ( n50579 , n50578 );
or ( n50580 , n50572 , n50579 );
buf ( n50581 , n47072 );
not ( n50582 , n50581 );
buf ( n50583 , n50582 );
buf ( n50584 , n50583 );
buf ( n50585 , n46073 );
nand ( n50586 , n50584 , n50585 );
buf ( n50587 , n50586 );
nand ( n50588 , n50580 , n50587 );
not ( n50589 , n50588 );
or ( n50590 , n50571 , n50589 );
buf ( n50591 , n38963 );
buf ( n50592 , n50591 );
not ( n50593 , n50592 );
buf ( n50594 , n46657 );
not ( n50595 , n50594 );
or ( n50596 , n50593 , n50595 );
buf ( n50597 , n42149 );
buf ( n50598 , n38963 );
not ( n50599 , n50598 );
buf ( n50600 , n50599 );
nand ( n50601 , n50597 , n50600 );
buf ( n50602 , n50601 );
buf ( n50603 , n50602 );
nand ( n50604 , n50596 , n50603 );
buf ( n50605 , n50604 );
buf ( n50606 , n39998 );
not ( n50607 , n50606 );
buf ( n50608 , n50607 );
nand ( n50609 , n50605 , n50608 );
nand ( n50610 , n50590 , n50609 );
buf ( n50611 , n50610 );
buf ( n50612 , n39983 );
not ( n50613 , n50612 );
buf ( n50614 , n48696 );
not ( n50615 , n50614 );
or ( n50616 , n50613 , n50615 );
nand ( n50617 , n50588 , n39999 );
buf ( n50618 , n50617 );
nand ( n50619 , n50616 , n50618 );
buf ( n50620 , n50619 );
buf ( n50621 , n50620 );
xor ( n50622 , n50611 , n50621 );
buf ( n50623 , n45056 );
not ( n50624 , n29406 );
buf ( n50625 , n50624 );
not ( n50626 , n50625 );
buf ( n50627 , n47031 );
not ( n50628 , n50627 );
or ( n50629 , n50626 , n50628 );
buf ( n50630 , n42468 );
buf ( n50631 , n43362 );
nand ( n50632 , n50630 , n50631 );
buf ( n50633 , n50632 );
buf ( n50634 , n50633 );
nand ( n50635 , n50629 , n50634 );
buf ( n50636 , n50635 );
buf ( n50637 , n50636 );
not ( n50638 , n50637 );
buf ( n50639 , n50638 );
buf ( n50640 , n50639 );
or ( n50641 , n50623 , n50640 );
buf ( n50642 , n50097 );
not ( n50643 , n50642 );
buf ( n50644 , n50643 );
buf ( n50645 , n50644 );
buf ( n50646 , n47020 );
or ( n50647 , n50645 , n50646 );
nand ( n50648 , n50641 , n50647 );
buf ( n50649 , n50648 );
buf ( n50650 , n50649 );
and ( n50651 , n50622 , n50650 );
and ( n50652 , n50611 , n50621 );
or ( n50653 , n50651 , n50652 );
buf ( n50654 , n50653 );
buf ( n50655 , n42504 );
not ( n50656 , n50655 );
buf ( n50657 , n37472 );
not ( n50658 , n50657 );
or ( n50659 , n50656 , n50658 );
buf ( n50660 , n37473 );
buf ( n50661 , n41721 );
nand ( n50662 , n50660 , n50661 );
buf ( n50663 , n50662 );
buf ( n50664 , n50663 );
nand ( n50665 , n50659 , n50664 );
buf ( n50666 , n50665 );
buf ( n50667 , n50666 );
not ( n50668 , n50667 );
buf ( n50669 , n47490 );
not ( n50670 , n50669 );
buf ( n50671 , n50670 );
buf ( n50672 , n50671 );
not ( n50673 , n50672 );
or ( n50674 , n50668 , n50673 );
buf ( n50675 , n41852 );
buf ( n50676 , n49899 );
nand ( n50677 , n50675 , n50676 );
buf ( n50678 , n50677 );
buf ( n50679 , n50678 );
nand ( n50680 , n50674 , n50679 );
buf ( n50681 , n50680 );
or ( n50682 , n50654 , n50681 );
not ( n50683 , n50682 );
or ( n50684 , n50570 , n50683 );
nand ( n50685 , n50654 , n50681 );
nand ( n50686 , n50684 , n50685 );
buf ( n50687 , n50686 );
nand ( n50688 , n50544 , n50687 );
buf ( n50689 , n50688 );
buf ( n50690 , n50689 );
nand ( n50691 , n50536 , n50690 );
buf ( n50692 , n50691 );
not ( n50693 , n50692 );
or ( n50694 , n50485 , n50693 );
buf ( n50695 , n50454 );
buf ( n50696 , n50480 );
nand ( n50697 , n50695 , n50696 );
buf ( n50698 , n50697 );
nand ( n50699 , n50694 , n50698 );
not ( n50700 , n50699 );
buf ( n50701 , n48666 );
buf ( n50702 , n48671 );
and ( n50703 , n50701 , n50702 );
not ( n50704 , n48390 );
not ( n50705 , n47932 );
or ( n50706 , n50704 , n50705 );
buf ( n50707 , n38821 );
buf ( n50708 , n41660 );
nand ( n50709 , n50707 , n50708 );
buf ( n50710 , n50709 );
nand ( n50711 , n50706 , n50710 );
and ( n50712 , n50711 , n41705 );
buf ( n50713 , n50712 );
nor ( n50714 , n50703 , n50713 );
buf ( n50715 , n50714 );
buf ( n50716 , n50715 );
not ( n50717 , n50716 );
buf ( n50718 , n50717 );
not ( n50719 , n50718 );
buf ( n50720 , n48977 );
buf ( n50721 , n48964 );
and ( n50722 , n50720 , n50721 );
not ( n50723 , n50720 );
buf ( n50724 , n48961 );
and ( n50725 , n50723 , n50724 );
nor ( n50726 , n50722 , n50725 );
buf ( n50727 , n50726 );
buf ( n50728 , n50727 );
buf ( n50729 , n49001 );
not ( n50730 , n50729 );
buf ( n50731 , n50730 );
buf ( n50732 , n50731 );
and ( n50733 , n50728 , n50732 );
not ( n50734 , n50728 );
buf ( n50735 , n49001 );
and ( n50736 , n50734 , n50735 );
nor ( n50737 , n50733 , n50736 );
buf ( n50738 , n50737 );
buf ( n50739 , n50738 );
not ( n50740 , n50739 );
buf ( n50741 , n50740 );
not ( n50742 , n50741 );
or ( n50743 , n50719 , n50742 );
not ( n50744 , n50715 );
not ( n50745 , n50738 );
or ( n50746 , n50744 , n50745 );
buf ( n50747 , n48707 );
not ( n50748 , n50747 );
buf ( n50749 , n50748 );
buf ( n50750 , n50749 );
buf ( n50751 , n43108 );
not ( n50752 , n50751 );
buf ( n50753 , n37328 );
not ( n50754 , n50753 );
or ( n50755 , n50752 , n50754 );
buf ( n50756 , n41779 );
buf ( n50757 , n43099 );
nand ( n50758 , n50756 , n50757 );
buf ( n50759 , n50758 );
buf ( n50760 , n50759 );
nand ( n50761 , n50755 , n50760 );
buf ( n50762 , n50761 );
buf ( n50763 , n50762 );
not ( n50764 , n50763 );
buf ( n50765 , n37397 );
not ( n50766 , n50765 );
or ( n50767 , n50764 , n50766 );
nand ( n50768 , n45108 , n48738 );
buf ( n50769 , n50768 );
nand ( n50770 , n50767 , n50769 );
buf ( n50771 , n50770 );
buf ( n50772 , n50771 );
xor ( n50773 , n50750 , n50772 );
buf ( n50774 , n43938 );
not ( n50775 , n50774 );
buf ( n50776 , n48357 );
not ( n50777 , n50776 );
buf ( n50778 , n41799 );
not ( n50779 , n50778 );
or ( n50780 , n50777 , n50779 );
buf ( n50781 , n44210 );
not ( n50782 , n50781 );
buf ( n50783 , n50782 );
buf ( n50784 , n50783 );
buf ( n50785 , n50045 );
nand ( n50786 , n50784 , n50785 );
buf ( n50787 , n50786 );
buf ( n50788 , n50787 );
nand ( n50789 , n50780 , n50788 );
buf ( n50790 , n50789 );
buf ( n50791 , n50790 );
not ( n50792 , n50791 );
or ( n50793 , n50775 , n50792 );
buf ( n50794 , n50051 );
buf ( n50795 , n46294 );
nand ( n50796 , n50794 , n50795 );
buf ( n50797 , n50796 );
buf ( n50798 , n50797 );
nand ( n50799 , n50793 , n50798 );
buf ( n50800 , n50799 );
buf ( n50801 , n50800 );
and ( n50802 , n50773 , n50801 );
and ( n50803 , n50750 , n50772 );
or ( n50804 , n50802 , n50803 );
buf ( n50805 , n50804 );
nand ( n50806 , n50746 , n50805 );
nand ( n50807 , n50743 , n50806 );
buf ( n50808 , n50807 );
xor ( n50809 , n49013 , n49033 );
xor ( n50810 , n50809 , n49045 );
buf ( n50811 , n50810 );
xor ( n50812 , n50808 , n50811 );
xor ( n50813 , n48650 , n48677 );
xor ( n50814 , n50813 , n48756 );
buf ( n50815 , n50814 );
and ( n50816 , n50812 , n50815 );
and ( n50817 , n50808 , n50811 );
or ( n50818 , n50816 , n50817 );
buf ( n50819 , n50818 );
buf ( n50820 , n50819 );
not ( n50821 , n50820 );
buf ( n50822 , n50821 );
nand ( n50823 , n50700 , n50822 );
not ( n50824 , n50823 );
or ( n50825 , n50430 , n50824 );
not ( n50826 , n50822 );
nand ( n50827 , n50826 , n50699 );
nand ( n50828 , n50825 , n50827 );
buf ( n50829 , n50828 );
xor ( n50830 , n50331 , n50829 );
not ( n50831 , n48934 );
not ( n50832 , n49063 );
not ( n50833 , n50832 );
or ( n50834 , n50831 , n50833 );
or ( n50835 , n48934 , n50832 );
nand ( n50836 , n50834 , n50835 );
not ( n50837 , n50836 );
xor ( n50838 , n48806 , n50837 );
buf ( n50839 , n50838 );
and ( n50840 , n50830 , n50839 );
and ( n50841 , n50331 , n50829 );
or ( n50842 , n50840 , n50841 );
buf ( n50843 , n50842 );
nand ( n50844 , n50324 , n50843 );
nand ( n50845 , n50320 , n50844 );
not ( n50846 , n50845 );
and ( n50847 , n50226 , n50846 );
not ( n50848 , n50226 );
and ( n50849 , n50848 , n50845 );
nor ( n50850 , n50847 , n50849 );
xor ( n50851 , n49696 , n50850 );
buf ( n50852 , n50198 );
buf ( n50853 , n50217 );
xor ( n50854 , n50852 , n50853 );
buf ( n50855 , n50214 );
xnor ( n50856 , n50854 , n50855 );
buf ( n50857 , n50856 );
buf ( n50858 , n50857 );
xor ( n50859 , n49053 , n49049 );
xor ( n50860 , n50859 , n49059 );
xor ( n50861 , n48878 , n48903 );
xor ( n50862 , n50861 , n48925 );
buf ( n50863 , n50862 );
not ( n50864 , n50863 );
nand ( n50865 , n50860 , n50864 );
buf ( n50866 , n50865 );
not ( n50867 , n50866 );
buf ( n50868 , n44708 );
not ( n50869 , n50868 );
not ( n50870 , n44533 );
not ( n50871 , n37148 );
not ( n50872 , n50871 );
or ( n50873 , n50870 , n50872 );
buf ( n50874 , n44533 );
not ( n50875 , n50874 );
not ( n50876 , n42360 );
buf ( n50877 , n50876 );
nand ( n50878 , n50875 , n50877 );
buf ( n50879 , n50878 );
nand ( n50880 , n50873 , n50879 );
buf ( n50881 , n50880 );
not ( n50882 , n50881 );
or ( n50883 , n50869 , n50882 );
buf ( n50884 , n50286 );
buf ( n50885 , n44496 );
nand ( n50886 , n50884 , n50885 );
buf ( n50887 , n50886 );
buf ( n50888 , n50887 );
nand ( n50889 , n50883 , n50888 );
buf ( n50890 , n50889 );
buf ( n50891 , n50890 );
not ( n50892 , n50891 );
buf ( n50893 , n50892 );
buf ( n50894 , n50893 );
not ( n50895 , n50894 );
buf ( n50896 , n46225 );
not ( n50897 , n50896 );
and ( n50898 , n45753 , n39897 );
not ( n50899 , n45753 );
and ( n50900 , n50899 , n36396 );
or ( n50901 , n50898 , n50900 );
buf ( n50902 , n50901 );
not ( n50903 , n50902 );
or ( n50904 , n50897 , n50903 );
buf ( n50905 , n50257 );
buf ( n50906 , n46246 );
nand ( n50907 , n50905 , n50906 );
buf ( n50908 , n50907 );
buf ( n50909 , n50908 );
nand ( n50910 , n50904 , n50909 );
buf ( n50911 , n50910 );
not ( n50912 , n50911 );
buf ( n50913 , n50912 );
not ( n50914 , n50913 );
or ( n50915 , n50895 , n50914 );
buf ( n50916 , n42668 );
not ( n50917 , n50916 );
buf ( n50918 , n49968 );
not ( n50919 , n50918 );
or ( n50920 , n50917 , n50919 );
buf ( n50921 , n42672 );
not ( n50922 , n50921 );
buf ( n50923 , n43198 );
not ( n50924 , n50923 );
buf ( n50925 , n50924 );
buf ( n50926 , n50925 );
not ( n50927 , n50926 );
or ( n50928 , n50922 , n50927 );
buf ( n50929 , n43198 );
buf ( n50930 , n42671 );
nand ( n50931 , n50929 , n50930 );
buf ( n50932 , n50931 );
buf ( n50933 , n50932 );
nand ( n50934 , n50928 , n50933 );
buf ( n50935 , n50934 );
buf ( n50936 , n50935 );
buf ( n50937 , n42712 );
nand ( n50938 , n50936 , n50937 );
buf ( n50939 , n50938 );
buf ( n50940 , n50939 );
nand ( n50941 , n50920 , n50940 );
buf ( n50942 , n50941 );
not ( n50943 , n50942 );
buf ( n50944 , n49908 );
buf ( n50945 , n49886 );
xor ( n50946 , n50944 , n50945 );
buf ( n50947 , n49934 );
xnor ( n50948 , n50946 , n50947 );
buf ( n50949 , n50948 );
buf ( n50950 , n50949 );
not ( n50951 , n50950 );
buf ( n50952 , n50951 );
not ( n50953 , n50952 );
or ( n50954 , n50943 , n50953 );
buf ( n50955 , n50942 );
not ( n50956 , n50955 );
buf ( n50957 , n50956 );
not ( n50958 , n50957 );
not ( n50959 , n50949 );
or ( n50960 , n50958 , n50959 );
buf ( n50961 , n48671 );
not ( n50962 , n50961 );
buf ( n50963 , n50711 );
not ( n50964 , n50963 );
or ( n50965 , n50962 , n50964 );
buf ( n50966 , n48390 );
not ( n50967 , n50966 );
buf ( n50968 , n44989 );
not ( n50969 , n50968 );
or ( n50970 , n50967 , n50969 );
buf ( n50971 , n30187 );
buf ( n50972 , n41660 );
nand ( n50973 , n50971 , n50972 );
buf ( n50974 , n50973 );
buf ( n50975 , n50974 );
nand ( n50976 , n50970 , n50975 );
buf ( n50977 , n50976 );
buf ( n50978 , n50977 );
buf ( n50979 , n41703 );
buf ( n50980 , n50979 );
not ( n50981 , n50980 );
buf ( n50982 , n50981 );
buf ( n50983 , n50982 );
nand ( n50984 , n50978 , n50983 );
buf ( n50985 , n50984 );
buf ( n50986 , n50985 );
nand ( n50987 , n50965 , n50986 );
buf ( n50988 , n50987 );
buf ( n50989 , n50988 );
buf ( n50990 , n25879 );
not ( n50991 , n50990 );
buf ( n50992 , n50991 );
buf ( n50993 , n50992 );
not ( n50994 , n50993 );
buf ( n50995 , n50994 );
buf ( n50996 , n50995 );
not ( n50997 , n50996 );
buf ( n50998 , n50997 );
buf ( n50999 , n50998 );
buf ( n51000 , n50999 );
buf ( n51001 , n51000 );
buf ( n51002 , n51001 );
not ( n51003 , n51002 );
buf ( n51004 , n51003 );
buf ( n51005 , n51004 );
not ( n51006 , n51005 );
buf ( n51007 , n37649 );
not ( n51008 , n51007 );
or ( n51009 , n51006 , n51008 );
buf ( n51010 , n36360 );
buf ( n51011 , n51001 );
nand ( n51012 , n51010 , n51011 );
buf ( n51013 , n51012 );
buf ( n51014 , n51013 );
nand ( n51015 , n51009 , n51014 );
buf ( n51016 , n51015 );
buf ( n51017 , n43053 );
buf ( n51018 , n50073 );
nand ( n51019 , n51017 , n51018 );
buf ( n51020 , n51019 );
buf ( n51021 , n51020 );
nand ( n51022 , C1 , n51021 );
buf ( n51023 , n51022 );
buf ( n51024 , n51023 );
xor ( n51025 , n50989 , n51024 );
and ( n51026 , n46390 , n43259 );
not ( n51027 , n46390 );
buf ( n51028 , n39478 );
not ( n51029 , n51028 );
buf ( n51030 , n51029 );
and ( n51031 , n51027 , n51030 );
or ( n51032 , n51026 , n51031 );
buf ( n51033 , n51032 );
not ( n51034 , n51033 );
buf ( n51035 , n36101 );
not ( n51036 , n51035 );
or ( n51037 , n51034 , n51036 );
buf ( n51038 , n42530 );
buf ( n51039 , n49924 );
nand ( n51040 , n51038 , n51039 );
buf ( n51041 , n51040 );
buf ( n51042 , n51041 );
nand ( n51043 , n51037 , n51042 );
buf ( n51044 , n51043 );
buf ( n51045 , n51044 );
and ( n51046 , n51025 , n51045 );
and ( n51047 , n50989 , n51024 );
or ( n51048 , n51046 , n51047 );
buf ( n51049 , n51048 );
nand ( n51050 , n50960 , n51049 );
nand ( n51051 , n50954 , n51050 );
buf ( n51052 , n51051 );
buf ( n51053 , n51052 );
buf ( n51054 , n51053 );
buf ( n51055 , n51054 );
nand ( n51056 , n50915 , n51055 );
buf ( n51057 , n51056 );
buf ( n51058 , n51057 );
buf ( n51059 , n50890 );
buf ( n51060 , n50911 );
nand ( n51061 , n51059 , n51060 );
buf ( n51062 , n51061 );
buf ( n51063 , n51062 );
nand ( n51064 , n51058 , n51063 );
buf ( n51065 , n51064 );
buf ( n51066 , n51065 );
not ( n51067 , n51066 );
or ( n51068 , n50867 , n51067 );
not ( n51069 , n50860 );
nand ( n51070 , n51069 , n50863 );
buf ( n51071 , n51070 );
nand ( n51072 , n51068 , n51071 );
buf ( n51073 , n51072 );
not ( n51074 , n51073 );
buf ( n51075 , n50231 );
buf ( n51076 , n50301 );
xor ( n51077 , n51075 , n51076 );
buf ( n51078 , n50228 );
xnor ( n51079 , n51077 , n51078 );
buf ( n51080 , n51079 );
not ( n51081 , n51080 );
not ( n51082 , n51081 );
or ( n51083 , n51074 , n51082 );
buf ( n51084 , n51073 );
not ( n51085 , n51084 );
buf ( n51086 , n51085 );
buf ( n51087 , n51086 );
not ( n51088 , n51087 );
buf ( n51089 , n51080 );
not ( n51090 , n51089 );
or ( n51091 , n51088 , n51090 );
xor ( n51092 , n49723 , n49821 );
xor ( n51093 , n51092 , n50194 );
buf ( n51094 , n51093 );
not ( n51095 , n51094 );
buf ( n51096 , n51095 );
buf ( n51097 , n51096 );
nand ( n51098 , n51091 , n51097 );
buf ( n51099 , n51098 );
nand ( n51100 , n51083 , n51099 );
not ( n51101 , n51100 );
buf ( n51102 , n51101 );
xor ( n51103 , n50858 , n51102 );
xor ( n51104 , n49791 , n49795 );
xor ( n51105 , n51104 , n49817 );
buf ( n51106 , n51105 );
not ( n51107 , n51106 );
buf ( n51108 , n50293 );
buf ( n51109 , n50268 );
xor ( n51110 , n51108 , n51109 );
buf ( n51111 , n50242 );
xnor ( n51112 , n51110 , n51111 );
buf ( n51113 , n51112 );
nand ( n51114 , n51107 , n51113 );
not ( n51115 , n51114 );
xor ( n51116 , n49868 , n49950 );
xor ( n51117 , n51116 , n49976 );
buf ( n51118 , n51117 );
buf ( n51119 , n51118 );
not ( n51120 , n51119 );
xor ( n51121 , n50058 , n50081 );
xor ( n51122 , n51121 , n50178 );
buf ( n51123 , n51122 );
buf ( n51124 , n51123 );
not ( n51125 , n51124 );
buf ( n51126 , n51125 );
buf ( n51127 , n51126 );
not ( n51128 , n51127 );
buf ( n51129 , n50010 );
buf ( n51130 , n43868 );
and ( n51131 , n51129 , n51130 );
and ( n51132 , n38244 , n41611 );
not ( n51133 , n38244 );
and ( n51134 , n51133 , n41608 );
or ( n51135 , n51132 , n51134 );
buf ( n51136 , n51135 );
buf ( n51137 , n44267 );
and ( n51138 , n51136 , n51137 );
buf ( n51139 , n51138 );
buf ( n51140 , n51139 );
nor ( n51141 , n51131 , n51140 );
buf ( n51142 , n51141 );
buf ( n51143 , n51142 );
not ( n51144 , n51143 );
or ( n51145 , n51128 , n51144 );
buf ( n51146 , n47098 );
buf ( n51147 , n42862 );
buf ( n51148 , n38108 );
and ( n51149 , n51147 , n51148 );
not ( n51150 , n51147 );
buf ( n51151 , n49385 );
and ( n51152 , n51150 , n51151 );
nor ( n51153 , n51149 , n51152 );
buf ( n51154 , n51153 );
buf ( n51155 , n51154 );
or ( n51156 , n51146 , n51155 );
buf ( n51157 , n46172 );
not ( n51158 , n51157 );
buf ( n51159 , n51158 );
buf ( n51160 , n51159 );
buf ( n51161 , n50521 );
not ( n51162 , n51161 );
buf ( n51163 , n51162 );
buf ( n51164 , n51163 );
or ( n51165 , n51160 , n51164 );
nand ( n51166 , n51156 , n51165 );
buf ( n51167 , n51166 );
buf ( n51168 , n51167 );
buf ( n51169 , n50110 );
buf ( n51170 , n50140 );
xor ( n51171 , n51169 , n51170 );
buf ( n51172 , n50171 );
xor ( n51173 , n51171 , n51172 );
buf ( n51174 , n51173 );
buf ( n51175 , n51174 );
xor ( n51176 , n51168 , n51175 );
buf ( n51177 , n44670 );
and ( n51178 , n44952 , n44689 );
not ( n51179 , n44952 );
and ( n51180 , n51179 , n39235 );
nor ( n51181 , n51178 , n51180 );
buf ( n51182 , n51181 );
or ( n51183 , n51177 , n51182 );
buf ( n51184 , n44682 );
buf ( n51185 , n50493 );
not ( n51186 , n51185 );
buf ( n51187 , n51186 );
buf ( n51188 , n51187 );
or ( n51189 , n51184 , n51188 );
nand ( n51190 , n51183 , n51189 );
buf ( n51191 , n51190 );
buf ( n51192 , n51191 );
and ( n51193 , n51176 , n51192 );
and ( n51194 , n51168 , n51175 );
or ( n51195 , n51193 , n51194 );
buf ( n51196 , n51195 );
buf ( n51197 , n51196 );
nand ( n51198 , n51145 , n51197 );
buf ( n51199 , n51198 );
buf ( n51200 , n51199 );
buf ( n51201 , n51142 );
not ( n51202 , n51201 );
buf ( n51203 , n51202 );
buf ( n51204 , n51203 );
buf ( n51205 , n51123 );
nand ( n51206 , n51204 , n51205 );
buf ( n51207 , n51206 );
buf ( n51208 , n51207 );
nand ( n51209 , n51200 , n51208 );
buf ( n51210 , n51209 );
buf ( n51211 , n51210 );
not ( n51212 , n51211 );
or ( n51213 , n51120 , n51212 );
buf ( n51214 , n51118 );
not ( n51215 , n51214 );
buf ( n51216 , n51215 );
buf ( n51217 , n51216 );
not ( n51218 , n51217 );
not ( n51219 , n51210 );
buf ( n51220 , n51219 );
not ( n51221 , n51220 );
or ( n51222 , n51218 , n51221 );
buf ( n51223 , n50539 );
not ( n51224 , n51223 );
buf ( n51225 , n50505 );
not ( n51226 , n51225 );
or ( n51227 , n51224 , n51226 );
buf ( n51228 , n50505 );
buf ( n51229 , n50539 );
or ( n51230 , n51228 , n51229 );
nand ( n51231 , n51227 , n51230 );
buf ( n51232 , n51231 );
buf ( n51233 , n51232 );
buf ( n51234 , n50686 );
not ( n51235 , n51234 );
buf ( n51236 , n51235 );
buf ( n51237 , n51236 );
and ( n51238 , n51233 , n51237 );
not ( n51239 , n51233 );
buf ( n51240 , n50686 );
and ( n51241 , n51239 , n51240 );
nor ( n51242 , n51238 , n51241 );
buf ( n51243 , n51242 );
not ( n51244 , n51243 );
not ( n51245 , n47872 );
not ( n51246 , n50124 );
or ( n51247 , n51245 , n51246 );
buf ( n51248 , n25160 );
not ( n51249 , n51248 );
not ( n51250 , n41821 );
buf ( n51251 , n51250 );
not ( n51252 , n51251 );
or ( n51253 , n51249 , n51252 );
buf ( n51254 , n41822 );
buf ( n51255 , n46356 );
nand ( n51256 , n51254 , n51255 );
buf ( n51257 , n51256 );
buf ( n51258 , n51257 );
nand ( n51259 , n51253 , n51258 );
buf ( n51260 , n51259 );
buf ( n51261 , n51260 );
buf ( n51262 , n50128 );
nand ( n51263 , n51261 , n51262 );
buf ( n51264 , n51263 );
nand ( n51265 , n51247 , n51264 );
not ( n51266 , n51265 );
not ( n51267 , n51266 );
not ( n51268 , n38404 );
buf ( n51269 , n42049 );
not ( n51270 , n51269 );
buf ( n51271 , n42403 );
not ( n51272 , n51271 );
or ( n51273 , n51270 , n51272 );
buf ( n51274 , n48984 );
buf ( n51275 , n42052 );
nand ( n51276 , n51274 , n51275 );
buf ( n51277 , n51276 );
buf ( n51278 , n51277 );
nand ( n51279 , n51273 , n51278 );
buf ( n51280 , n51279 );
not ( n51281 , n51280 );
or ( n51282 , n51268 , n51281 );
nand ( n51283 , n50163 , n38380 );
nand ( n51284 , n51282 , n51283 );
buf ( n51285 , n51284 );
not ( n51286 , n51285 );
buf ( n51287 , n51286 );
not ( n51288 , n51287 );
or ( n51289 , n51267 , n51288 );
not ( n51290 , n37400 );
buf ( n51291 , n41736 );
not ( n51292 , n51291 );
buf ( n51293 , n43442 );
not ( n51294 , n51293 );
or ( n51295 , n51292 , n51294 );
buf ( n51296 , n41778 );
not ( n51297 , n51296 );
buf ( n51298 , n41748 );
nand ( n51299 , n51297 , n51298 );
buf ( n51300 , n51299 );
buf ( n51301 , n51300 );
nand ( n51302 , n51295 , n51301 );
buf ( n51303 , n51302 );
not ( n51304 , n51303 );
or ( n51305 , n51290 , n51304 );
buf ( n51306 , n50762 );
buf ( n51307 , n37413 );
nand ( n51308 , n51306 , n51307 );
buf ( n51309 , n51308 );
nand ( n51310 , n51305 , n51309 );
nand ( n51311 , n51289 , n51310 );
buf ( n51312 , n51265 );
buf ( n51313 , n51284 );
nand ( n51314 , n51312 , n51313 );
buf ( n51315 , n51314 );
and ( n51316 , n51311 , n51315 );
buf ( n51317 , n50403 );
buf ( n51318 , n42339 );
and ( n51319 , n51317 , n51318 );
not ( n51320 , n45394 );
not ( n51321 , n42343 );
or ( n51322 , n51320 , n51321 );
buf ( n51323 , n37641 );
buf ( n51324 , n46855 );
nand ( n51325 , n51323 , n51324 );
buf ( n51326 , n51325 );
nand ( n51327 , n51322 , n51326 );
not ( n51328 , n51327 );
nor ( n51329 , n51328 , n42375 );
buf ( n51330 , n51329 );
nor ( n51331 , n51319 , n51330 );
buf ( n51332 , n51331 );
xor ( n51333 , n51316 , n51332 );
buf ( n51334 , n48323 );
not ( n51335 , n51334 );
buf ( n51336 , n41741 );
not ( n51337 , n51336 );
or ( n51338 , n51335 , n51337 );
buf ( n51339 , n38471 );
buf ( n51340 , n48320 );
nand ( n51341 , n51339 , n51340 );
buf ( n51342 , n51341 );
buf ( n51343 , n51342 );
nand ( n51344 , n51338 , n51343 );
buf ( n51345 , n51344 );
buf ( n51346 , n51345 );
not ( n51347 , n51346 );
buf ( n51348 , n51347 );
buf ( n51349 , n51348 );
not ( n51350 , n51349 );
buf ( n51351 , n36520 );
not ( n51352 , n51351 );
and ( n51353 , n51350 , n51352 );
not ( n51354 , n50369 );
nor ( n51355 , n51354 , n39813 );
buf ( n51356 , n51355 );
nor ( n51357 , n51353 , n51356 );
buf ( n51358 , n51357 );
and ( n51359 , n51333 , n51358 );
and ( n51360 , n51316 , n51332 );
or ( n51361 , n51359 , n51360 );
not ( n51362 , n51361 );
and ( n51363 , n51244 , n51362 );
buf ( n51364 , n51361 );
buf ( n51365 , n51243 );
nand ( n51366 , n51364 , n51365 );
buf ( n51367 , n51366 );
not ( n51368 , n50715 );
not ( n51369 , n50741 );
or ( n51370 , n51368 , n51369 );
buf ( n51371 , n50718 );
buf ( n51372 , n50738 );
nand ( n51373 , n51371 , n51372 );
buf ( n51374 , n51373 );
nand ( n51375 , n51370 , n51374 );
xor ( n51376 , n51375 , n50805 );
and ( n51377 , n51367 , n51376 );
nor ( n51378 , n51363 , n51377 );
buf ( n51379 , n51378 );
not ( n51380 , n51379 );
buf ( n51381 , n51380 );
buf ( n51382 , n51381 );
nand ( n51383 , n51222 , n51382 );
buf ( n51384 , n51383 );
buf ( n51385 , n51384 );
nand ( n51386 , n51213 , n51385 );
buf ( n51387 , n51386 );
not ( n51388 , n51387 );
or ( n51389 , n51115 , n51388 );
buf ( n51390 , n51113 );
not ( n51391 , n51390 );
buf ( n51392 , n51106 );
nand ( n51393 , n51391 , n51392 );
buf ( n51394 , n51393 );
nand ( n51395 , n51389 , n51394 );
buf ( n51396 , n51395 );
not ( n51397 , n51396 );
buf ( n51398 , n49980 );
buf ( n51399 , n49840 );
xor ( n51400 , n51398 , n51399 );
buf ( n51401 , n50188 );
xnor ( n51402 , n51400 , n51401 );
buf ( n51403 , n51402 );
buf ( n51404 , n51403 );
not ( n51405 , n51404 );
and ( n51406 , n50699 , n50822 );
not ( n51407 , n50699 );
and ( n51408 , n51407 , n50819 );
nor ( n51409 , n51406 , n51408 );
xor ( n51410 , n50429 , n51409 );
buf ( n51411 , n51410 );
not ( n51412 , n51411 );
or ( n51413 , n51405 , n51412 );
buf ( n51414 , n48868 );
not ( n51415 , n51414 );
buf ( n51416 , n50447 );
not ( n51417 , n51416 );
or ( n51418 , n51415 , n51417 );
buf ( n51419 , n48808 );
buf ( n51420 , n36611 );
and ( n51421 , n51419 , n51420 );
not ( n51422 , n51419 );
buf ( n51423 , n45650 );
and ( n51424 , n51422 , n51423 );
nor ( n51425 , n51421 , n51424 );
buf ( n51426 , n51425 );
buf ( n51427 , n51426 );
buf ( n51428 , n48855 );
nand ( n51429 , n51427 , n51428 );
buf ( n51430 , n51429 );
buf ( n51431 , n51430 );
nand ( n51432 , n51418 , n51431 );
buf ( n51433 , n51432 );
not ( n51434 , n51433 );
buf ( n51435 , n50470 );
buf ( n51436 , n42315 );
and ( n51437 , n51435 , n51436 );
buf ( n51438 , n42266 );
not ( n51439 , n51438 );
buf ( n51440 , n46851 );
not ( n51441 , n51440 );
or ( n51442 , n51439 , n51441 );
buf ( n51443 , n37293 );
buf ( n51444 , n42263 );
nand ( n51445 , n51443 , n51444 );
buf ( n51446 , n51445 );
buf ( n51447 , n51446 );
nand ( n51448 , n51442 , n51447 );
buf ( n51449 , n51448 );
buf ( n51450 , n51449 );
not ( n51451 , n51450 );
buf ( n51452 , n42249 );
nor ( n51453 , n51451 , n51452 );
buf ( n51454 , n51453 );
buf ( n51455 , n51454 );
nor ( n51456 , n51437 , n51455 );
buf ( n51457 , n51456 );
nand ( n51458 , n51434 , n51457 );
not ( n51459 , n51458 );
buf ( n51460 , n23565 );
nand ( n51461 , C1 , n51460 );
buf ( n51462 , n51461 );
not ( n51463 , n51462 );
not ( n51464 , n23615 );
and ( n51465 , n51464 , C1 );
or ( n51466 , n51465 , C0 );
and ( n51467 , n51463 , n51466 );
not ( n51468 , n51463 );
and ( n51469 , n23615 , C1 );
or ( n51470 , n51469 , C0 );
and ( n51471 , n51468 , n51470 );
or ( n51472 , n51467 , n51471 );
not ( n51473 , n51472 );
buf ( n51474 , n51473 );
not ( n51475 , n51474 );
not ( n51476 , n51473 );
not ( n51477 , n23615 );
not ( n51478 , n51463 );
or ( n51479 , n51477 , n51478 );
nand ( n51480 , n51462 , n51464 );
nand ( n51481 , n51479 , n51480 );
not ( n51482 , n51481 );
and ( n51483 , n24661 , n51482 );
not ( n51484 , n24661 );
and ( n51485 , n51484 , n51481 );
or ( n51486 , n51483 , n51485 );
nor ( n51487 , n51476 , n51486 );
buf ( n51488 , n51487 );
not ( n51489 , n51488 );
buf ( n51490 , n51489 );
not ( n51491 , n51490 );
or ( n51492 , n51475 , n51491 );
not ( n51493 , n48836 );
buf ( n51494 , n51493 );
not ( n51495 , n51494 );
buf ( n51496 , n51495 );
buf ( n51497 , n51496 );
not ( n51498 , n51497 );
buf ( n51499 , n41619 );
not ( n51500 , n51499 );
or ( n51501 , n51498 , n51500 );
buf ( n51502 , n39005 );
buf ( n51503 , n51493 );
nand ( n51504 , n51502 , n51503 );
buf ( n51505 , n51504 );
buf ( n51506 , n51505 );
nand ( n51507 , n51501 , n51506 );
buf ( n51508 , n51507 );
buf ( n51509 , n51508 );
nand ( n51510 , n51492 , n51509 );
buf ( n51511 , n51510 );
not ( n51512 , n51511 );
or ( n51513 , n51459 , n51512 );
buf ( n51514 , n51457 );
not ( n51515 , n51514 );
buf ( n51516 , n51433 );
nand ( n51517 , n51515 , n51516 );
buf ( n51518 , n51517 );
nand ( n51519 , n51513 , n51518 );
buf ( n51520 , n51519 );
not ( n51521 , n51520 );
buf ( n51522 , n50182 );
buf ( n51523 , n49993 );
xor ( n51524 , n51522 , n51523 );
buf ( n51525 , n50020 );
xnor ( n51526 , n51524 , n51525 );
buf ( n51527 , n51526 );
buf ( n51528 , n51527 );
not ( n51529 , n51528 );
buf ( n51530 , n51529 );
buf ( n51531 , n51530 );
not ( n51532 , n51531 );
or ( n51533 , n51521 , n51532 );
buf ( n51534 , n51519 );
not ( n51535 , n51534 );
buf ( n51536 , n51535 );
buf ( n51537 , n51536 );
not ( n51538 , n51537 );
buf ( n51539 , n51527 );
not ( n51540 , n51539 );
or ( n51541 , n51538 , n51540 );
xor ( n51542 , n50808 , n50811 );
xor ( n51543 , n51542 , n50815 );
buf ( n51544 , n51543 );
buf ( n51545 , n51544 );
nand ( n51546 , n51541 , n51545 );
buf ( n51547 , n51546 );
buf ( n51548 , n51547 );
nand ( n51549 , n51533 , n51548 );
buf ( n51550 , n51549 );
buf ( n51551 , n51550 );
nand ( n51552 , n51413 , n51551 );
buf ( n51553 , n51552 );
not ( n51554 , n51403 );
buf ( n51555 , n51410 );
not ( n51556 , n51555 );
buf ( n51557 , n51556 );
nand ( n51558 , n51554 , n51557 );
nand ( n51559 , n51553 , n51558 );
buf ( n51560 , n51559 );
not ( n51561 , n51560 );
buf ( n51562 , n51561 );
buf ( n51563 , n51562 );
nand ( n51564 , n51397 , n51563 );
buf ( n51565 , n51564 );
buf ( n51566 , n51565 );
xor ( n51567 , n50331 , n50829 );
xor ( n51568 , n51567 , n50839 );
buf ( n51569 , n51568 );
buf ( n51570 , n51569 );
and ( n51571 , n51566 , n51570 );
buf ( n51572 , n51395 );
buf ( n51573 , n51559 );
and ( n51574 , n51572 , n51573 );
buf ( n51575 , n51574 );
buf ( n51576 , n51575 );
nor ( n51577 , n51571 , n51576 );
buf ( n51578 , n51577 );
buf ( n51579 , n51578 );
and ( n51580 , n51103 , n51579 );
and ( n51581 , n50858 , n51102 );
or ( n51582 , n51580 , n51581 );
buf ( n51583 , n51582 );
xor ( n51584 , n50851 , n51583 );
buf ( n51585 , n50305 );
buf ( n51586 , n50843 );
xor ( n51587 , n51585 , n51586 );
buf ( n51588 , n50318 );
xor ( n51589 , n51587 , n51588 );
buf ( n51590 , n51589 );
not ( n51591 , n51590 );
xor ( n51592 , n50858 , n51102 );
xor ( n51593 , n51592 , n51579 );
buf ( n51594 , n51593 );
not ( n51595 , n51594 );
not ( n51596 , n51595 );
or ( n51597 , n51591 , n51596 );
not ( n51598 , n51590 );
not ( n51599 , n51598 );
not ( n51600 , n51594 );
or ( n51601 , n51599 , n51600 );
buf ( n51602 , n51073 );
buf ( n51603 , n51093 );
xor ( n51604 , n51602 , n51603 );
buf ( n51605 , n51080 );
xnor ( n51606 , n51604 , n51605 );
buf ( n51607 , n51606 );
not ( n51608 , n51607 );
xor ( n51609 , n50454 , n50483 );
xnor ( n51610 , n51609 , n50692 );
buf ( n51611 , n51610 );
buf ( n51612 , n50345 );
not ( n51613 , n51612 );
buf ( n51614 , n51613 );
buf ( n51615 , n51614 );
not ( n51616 , n51615 );
buf ( n51617 , n46915 );
not ( n51618 , n51617 );
and ( n51619 , n51616 , n51618 );
buf ( n51620 , n46890 );
not ( n51621 , n51620 );
buf ( n51622 , n51621 );
buf ( n51623 , n51622 );
not ( n51624 , n51623 );
buf ( n51625 , n40067 );
not ( n51626 , n51625 );
or ( n51627 , n51624 , n51626 );
buf ( n51628 , n36427 );
buf ( n51629 , n46887 );
nand ( n51630 , n51628 , n51629 );
buf ( n51631 , n51630 );
buf ( n51632 , n51631 );
nand ( n51633 , n51627 , n51632 );
buf ( n51634 , n51633 );
buf ( n51635 , n51634 );
buf ( n51636 , n47331 );
and ( n51637 , n51635 , n51636 );
nor ( n51638 , n51619 , n51637 );
buf ( n51639 , n51638 );
buf ( n51640 , n51639 );
not ( n51641 , n51640 );
buf ( n51642 , n44533 );
not ( n51643 , n51642 );
buf ( n51644 , n39280 );
not ( n51645 , n51644 );
or ( n51646 , n51643 , n51645 );
buf ( n51647 , n42929 );
buf ( n51648 , n44530 );
nand ( n51649 , n51647 , n51648 );
buf ( n51650 , n51649 );
buf ( n51651 , n51650 );
nand ( n51652 , n51646 , n51651 );
buf ( n51653 , n51652 );
buf ( n51654 , n51653 );
not ( n51655 , n51654 );
buf ( n51656 , n51655 );
not ( n51657 , n51656 );
not ( n51658 , n44518 );
and ( n51659 , n51657 , n51658 );
and ( n51660 , n50880 , n44496 );
nor ( n51661 , n51659 , n51660 );
buf ( n51662 , n51661 );
not ( n51663 , n51662 );
or ( n51664 , n51641 , n51663 );
buf ( n51665 , n46246 );
not ( n51666 , n51665 );
buf ( n51667 , n50901 );
not ( n51668 , n51667 );
or ( n51669 , n51666 , n51668 );
buf ( n51670 , n45753 );
not ( n51671 , n51670 );
buf ( n51672 , n38098 );
not ( n51673 , n51672 );
or ( n51674 , n51671 , n51673 );
buf ( n51675 , n39340 );
buf ( n51676 , n45750 );
nand ( n51677 , n51675 , n51676 );
buf ( n51678 , n51677 );
buf ( n51679 , n51678 );
nand ( n51680 , n51674 , n51679 );
buf ( n51681 , n51680 );
buf ( n51682 , n51681 );
buf ( n51683 , n46225 );
nand ( n51684 , n51682 , n51683 );
buf ( n51685 , n51684 );
buf ( n51686 , n51685 );
nand ( n51687 , n51669 , n51686 );
buf ( n51688 , n51687 );
buf ( n51689 , n51688 );
nand ( n51690 , n51664 , n51689 );
buf ( n51691 , n51690 );
buf ( n51692 , n51691 );
not ( n51693 , n51661 );
buf ( n51694 , n51639 );
not ( n51695 , n51694 );
buf ( n51696 , n51695 );
nand ( n51697 , n51693 , n51696 );
buf ( n51698 , n51697 );
nand ( n51699 , n51692 , n51698 );
buf ( n51700 , n51699 );
buf ( n51701 , n51700 );
or ( n51702 , n51611 , n51701 );
buf ( n51703 , n51702 );
buf ( n51704 , n51703 );
xor ( n51705 , n50361 , n50385 );
xor ( n51706 , n51705 , n50411 );
buf ( n51707 , n51706 );
buf ( n51708 , n51707 );
xor ( n51709 , n50750 , n50772 );
xor ( n51710 , n51709 , n50801 );
buf ( n51711 , n51710 );
buf ( n51712 , n51711 );
buf ( n51713 , n46294 );
not ( n51714 , n51713 );
buf ( n51715 , n50790 );
not ( n51716 , n51715 );
or ( n51717 , n51714 , n51716 );
buf ( n51718 , n48357 );
not ( n51719 , n51718 );
buf ( n51720 , n28722 );
not ( n51721 , n51720 );
or ( n51722 , n51719 , n51721 );
buf ( n51723 , n41762 );
buf ( n51724 , n50045 );
nand ( n51725 , n51723 , n51724 );
buf ( n51726 , n51725 );
buf ( n51727 , n51726 );
nand ( n51728 , n51722 , n51727 );
buf ( n51729 , n51728 );
buf ( n51730 , n51729 );
buf ( n51731 , n43938 );
nand ( n51732 , n51730 , n51731 );
buf ( n51733 , n51732 );
buf ( n51734 , n51733 );
nand ( n51735 , n51717 , n51734 );
buf ( n51736 , n51735 );
buf ( n51737 , n51736 );
buf ( n51738 , n37863 );
buf ( n51739 , n51738 );
buf ( n51740 , n43063 );
not ( n51741 , n51740 );
buf ( n51742 , n37880 );
not ( n51743 , n51742 );
or ( n51744 , n51741 , n51743 );
buf ( n51745 , n41889 );
buf ( n51746 , n43064 );
nand ( n51747 , n51745 , n51746 );
buf ( n51748 , n51747 );
buf ( n51749 , n51748 );
nand ( n51750 , n51744 , n51749 );
buf ( n51751 , n51750 );
buf ( n51752 , n51751 );
nand ( n51753 , n51739 , n51752 );
buf ( n51754 , n51753 );
or ( n51755 , n51754 , n41905 );
nand ( n51756 , n50556 , n41905 );
nand ( n51757 , n51755 , n51756 );
buf ( n51758 , n51757 );
xor ( n51759 , n51737 , n51758 );
buf ( n51760 , n50610 );
not ( n51761 , n51760 );
buf ( n51762 , n51761 );
buf ( n51763 , n51762 );
buf ( n51764 , n48172 );
not ( n51765 , n51764 );
buf ( n51766 , n47031 );
not ( n51767 , n51766 );
or ( n51768 , n51765 , n51767 );
buf ( n51769 , n38979 );
buf ( n51770 , n42072 );
nand ( n51771 , n51769 , n51770 );
buf ( n51772 , n51771 );
buf ( n51773 , n51772 );
nand ( n51774 , n51768 , n51773 );
buf ( n51775 , n51774 );
buf ( n51776 , n51775 );
not ( n51777 , n51776 );
buf ( n51778 , n47014 );
not ( n51779 , n51778 );
or ( n51780 , n51777 , n51779 );
buf ( n51781 , n50636 );
buf ( n51782 , n50104 );
nand ( n51783 , n51781 , n51782 );
buf ( n51784 , n51783 );
buf ( n51785 , n51784 );
nand ( n51786 , n51780 , n51785 );
buf ( n51787 , n51786 );
buf ( n51788 , n51787 );
xor ( n51789 , n51763 , n51788 );
buf ( n51790 , n51260 );
not ( n51791 , n51790 );
buf ( n51792 , n47872 );
not ( n51793 , n51792 );
or ( n51794 , n51791 , n51793 );
not ( n51795 , n25159 );
buf ( n51796 , n29358 );
not ( n51797 , n51796 );
buf ( n51798 , n51797 );
not ( n51799 , n51798 );
or ( n51800 , n51795 , n51799 );
buf ( n51801 , n29360 );
buf ( n51802 , n25159 );
not ( n51803 , n51802 );
buf ( n51804 , n51803 );
buf ( n51805 , n51804 );
nand ( n51806 , n51801 , n51805 );
buf ( n51807 , n51806 );
nand ( n51808 , n51800 , n51807 );
buf ( n51809 , n51808 );
buf ( n51810 , n42631 );
nand ( n51811 , n51809 , n51810 );
buf ( n51812 , n51811 );
buf ( n51813 , n51812 );
nand ( n51814 , n51794 , n51813 );
buf ( n51815 , n51814 );
buf ( n51816 , n51815 );
and ( n51817 , n51789 , n51816 );
and ( n51818 , n51763 , n51788 );
or ( n51819 , n51817 , n51818 );
buf ( n51820 , n51819 );
buf ( n51821 , n51820 );
and ( n51822 , n51759 , n51821 );
and ( n51823 , n51737 , n51758 );
or ( n51824 , n51822 , n51823 );
buf ( n51825 , n51824 );
buf ( n51826 , n51825 );
xor ( n51827 , n51712 , n51826 );
buf ( n51828 , n42712 );
not ( n51829 , n51828 );
buf ( n51830 , n42672 );
buf ( n51831 , n42973 );
not ( n51832 , n51831 );
buf ( n51833 , n51832 );
buf ( n51834 , n51833 );
and ( n51835 , n51830 , n51834 );
not ( n51836 , n51830 );
buf ( n51837 , n42795 );
and ( n51838 , n51836 , n51837 );
nor ( n51839 , n51835 , n51838 );
buf ( n51840 , n51839 );
buf ( n51841 , n51840 );
not ( n51842 , n51841 );
or ( n51843 , n51829 , n51842 );
buf ( n51844 , n50935 );
buf ( n51845 , n42668 );
nand ( n51846 , n51844 , n51845 );
buf ( n51847 , n51846 );
buf ( n51848 , n51847 );
nand ( n51849 , n51843 , n51848 );
buf ( n51850 , n51849 );
buf ( n51851 , n51850 );
and ( n51852 , n51827 , n51851 );
and ( n51853 , n51712 , n51826 );
or ( n51854 , n51852 , n51853 );
buf ( n51855 , n51854 );
buf ( n51856 , n51855 );
or ( n51857 , n51708 , n51856 );
not ( n51858 , n50654 );
xor ( n51859 , n50681 , n51858 );
not ( n51860 , n50569 );
xor ( n51861 , n51859 , n51860 );
buf ( n51862 , n51861 );
not ( n51863 , n51862 );
not ( n51864 , n42252 );
buf ( n51865 , n42266 );
not ( n51866 , n51865 );
buf ( n51867 , n39240 );
not ( n51868 , n51867 );
or ( n51869 , n51866 , n51868 );
buf ( n51870 , n37686 );
buf ( n51871 , n51870 );
buf ( n51872 , n51871 );
buf ( n51873 , n51872 );
buf ( n51874 , n42263 );
nand ( n51875 , n51873 , n51874 );
buf ( n51876 , n51875 );
buf ( n51877 , n51876 );
nand ( n51878 , n51869 , n51877 );
buf ( n51879 , n51878 );
not ( n51880 , n51879 );
or ( n51881 , n51864 , n51880 );
buf ( n51882 , n51449 );
buf ( n51883 , n42315 );
nand ( n51884 , n51882 , n51883 );
buf ( n51885 , n51884 );
nand ( n51886 , n51881 , n51885 );
buf ( n51887 , n51886 );
not ( n51888 , n51887 );
or ( n51889 , n51863 , n51888 );
buf ( n51890 , n51886 );
buf ( n51891 , n51861 );
or ( n51892 , n51890 , n51891 );
xor ( n51893 , n50611 , n50621 );
xor ( n51894 , n51893 , n50650 );
buf ( n51895 , n51894 );
buf ( n51896 , n42008 );
not ( n51897 , n51896 );
buf ( n51898 , n37472 );
not ( n51899 , n51898 );
or ( n51900 , n51897 , n51899 );
not ( n51901 , n37472 );
buf ( n51902 , n51901 );
buf ( n51903 , n42017 );
nand ( n51904 , n51902 , n51903 );
buf ( n51905 , n51904 );
buf ( n51906 , n51905 );
nand ( n51907 , n51900 , n51906 );
buf ( n51908 , n51907 );
not ( n51909 , n51908 );
buf ( n51910 , n37514 );
not ( n51911 , n51910 );
buf ( n51912 , n51911 );
not ( n51913 , n51912 );
or ( n51914 , n51909 , n51913 );
buf ( n51915 , n50666 );
buf ( n51916 , n37446 );
nand ( n51917 , n51915 , n51916 );
buf ( n51918 , n51917 );
nand ( n51919 , n51914 , n51918 );
xor ( n51920 , n51895 , n51919 );
buf ( n51921 , n47716 );
not ( n51922 , n51921 );
buf ( n51923 , n39493 );
not ( n51924 , n51923 );
or ( n51925 , n51922 , n51924 );
buf ( n51926 , n43503 );
buf ( n51927 , n47725 );
nand ( n51928 , n51926 , n51927 );
buf ( n51929 , n51928 );
buf ( n51930 , n51929 );
nand ( n51931 , n51925 , n51930 );
buf ( n51932 , n51931 );
buf ( n51933 , n51932 );
not ( n51934 , n51933 );
buf ( n51935 , n36098 );
not ( n51936 , n51935 );
buf ( n51937 , n51936 );
buf ( n51938 , n51937 );
not ( n51939 , n51938 );
or ( n51940 , n51934 , n51939 );
buf ( n51941 , n32969 );
buf ( n51942 , n51032 );
nand ( n51943 , n51941 , n51942 );
buf ( n51944 , n51943 );
buf ( n51945 , n51944 );
nand ( n51946 , n51940 , n51945 );
buf ( n51947 , n51946 );
and ( n51948 , n51920 , n51947 );
and ( n51949 , n51895 , n51919 );
or ( n51950 , n51948 , n51949 );
buf ( n51951 , n51950 );
nand ( n51952 , n51892 , n51951 );
buf ( n51953 , n51952 );
buf ( n51954 , n51953 );
nand ( n51955 , n51889 , n51954 );
buf ( n51956 , n51955 );
buf ( n51957 , n51956 );
nand ( n51958 , n51857 , n51957 );
buf ( n51959 , n51958 );
buf ( n51960 , n51959 );
buf ( n51961 , n51707 );
buf ( n51962 , n51855 );
nand ( n51963 , n51961 , n51962 );
buf ( n51964 , n51963 );
buf ( n51965 , n51964 );
nand ( n51966 , n51960 , n51965 );
buf ( n51967 , n51966 );
buf ( n51968 , n51967 );
and ( n51969 , n51704 , n51968 );
buf ( n51970 , n51700 );
buf ( n51971 , n51610 );
and ( n51972 , n51970 , n51971 );
buf ( n51973 , n51972 );
buf ( n51974 , n51973 );
nor ( n51975 , n51969 , n51974 );
buf ( n51976 , n51975 );
buf ( n51977 , n51976 );
buf ( n51978 , n51057 );
buf ( n51979 , n51062 );
nand ( n51980 , n51978 , n51979 );
buf ( n51981 , n51980 );
and ( n51982 , n51069 , n50864 );
not ( n51983 , n51069 );
and ( n51984 , n51983 , n50863 );
nor ( n51985 , n51982 , n51984 );
xor ( n51986 , n51981 , n51985 );
buf ( n51987 , n51986 );
xor ( n51988 , n51977 , n51987 );
xor ( n51989 , n50355 , n50415 );
buf ( n51990 , n51989 );
buf ( n51991 , n50423 );
not ( n51992 , n51991 );
buf ( n51993 , n51992 );
buf ( n51994 , n51993 );
and ( n51995 , n51990 , n51994 );
not ( n51996 , n51990 );
buf ( n51997 , n50423 );
and ( n51998 , n51996 , n51997 );
nor ( n51999 , n51995 , n51998 );
buf ( n52000 , n51999 );
buf ( n52001 , n50890 );
not ( n52002 , n52001 );
buf ( n52003 , n51051 );
not ( n52004 , n52003 );
buf ( n52005 , n52004 );
buf ( n52006 , n52005 );
not ( n52007 , n52006 );
or ( n52008 , n52002 , n52007 );
buf ( n52009 , n50893 );
buf ( n52010 , n51051 );
nand ( n52011 , n52009 , n52010 );
buf ( n52012 , n52011 );
buf ( n52013 , n52012 );
nand ( n52014 , n52008 , n52013 );
buf ( n52015 , n52014 );
buf ( n52016 , n52015 );
buf ( n52017 , n50912 );
and ( n52018 , n52016 , n52017 );
not ( n52019 , n52016 );
buf ( n52020 , n50911 );
and ( n52021 , n52019 , n52020 );
nor ( n52022 , n52018 , n52021 );
buf ( n52023 , n52022 );
xor ( n52024 , n52000 , n52023 );
xor ( n52025 , n51216 , n51210 );
xnor ( n52026 , n52025 , n51378 );
and ( n52027 , n52024 , n52026 );
and ( n52028 , n52000 , n52023 );
or ( n52029 , n52027 , n52028 );
buf ( n52030 , n52029 );
and ( n52031 , n51988 , n52030 );
and ( n52032 , n51977 , n51987 );
or ( n52033 , n52031 , n52032 );
buf ( n52034 , n52033 );
not ( n52035 , n52034 );
and ( n52036 , n51608 , n52035 );
buf ( n52037 , n50949 );
buf ( n52038 , n52037 );
buf ( n52039 , n52038 );
buf ( n52040 , n52039 );
buf ( n52041 , n51049 );
not ( n52042 , n52041 );
buf ( n52043 , n50957 );
not ( n52044 , n52043 );
or ( n52045 , n52042 , n52044 );
buf ( n52046 , n51049 );
not ( n52047 , n52046 );
buf ( n52048 , n52047 );
buf ( n52049 , n52048 );
buf ( n52050 , n50942 );
nand ( n52051 , n52049 , n52050 );
buf ( n52052 , n52051 );
buf ( n52053 , n52052 );
nand ( n52054 , n52045 , n52053 );
buf ( n52055 , n52054 );
buf ( n52056 , n52055 );
xor ( n52057 , n52040 , n52056 );
buf ( n52058 , n52057 );
buf ( n52059 , n52058 );
not ( n52060 , n52059 );
buf ( n52061 , n52060 );
buf ( n52062 , n52061 );
not ( n52063 , n52062 );
xor ( n52064 , n50989 , n51024 );
xor ( n52065 , n52064 , n51045 );
buf ( n52066 , n52065 );
not ( n52067 , n44708 );
not ( n52068 , n44533 );
not ( n52069 , n39407 );
or ( n52070 , n52068 , n52069 );
not ( n52071 , n44533 );
not ( n52072 , n38218 );
nand ( n52073 , n52071 , n52072 );
nand ( n52074 , n52070 , n52073 );
not ( n52075 , n52074 );
or ( n52076 , n52067 , n52075 );
buf ( n52077 , n51653 );
buf ( n52078 , n44496 );
nand ( n52079 , n52077 , n52078 );
buf ( n52080 , n52079 );
nand ( n52081 , n52076 , n52080 );
or ( n52082 , n52066 , n52081 );
not ( n52083 , n12548 );
nand ( n52084 , n52083 , n12528 );
not ( n52085 , n12542 );
nor ( n52086 , n52085 , n12545 );
nand ( n52087 , n52086 , n12529 );
nand ( n52088 , n12528 , n12546 );
not ( n52089 , n12545 );
nor ( n52090 , n52089 , n12542 );
nand ( n52091 , n12529 , n52090 );
nand ( n52092 , n52084 , n52087 , n52088 , n52091 );
not ( n52093 , n52092 );
buf ( n52094 , n52093 );
buf ( n52095 , n52094 );
buf ( n52096 , n38834 );
and ( n52097 , n52095 , n52096 );
not ( n52098 , n52095 );
buf ( n52099 , n37649 );
and ( n52100 , n52098 , n52099 );
nor ( n52101 , n52097 , n52100 );
buf ( n52102 , n52101 );
buf ( n52103 , n36444 );
buf ( n52104 , n51016 );
nand ( n52105 , n52103 , n52104 );
buf ( n52106 , n52105 );
buf ( n52107 , n52106 );
nand ( n52108 , C1 , n52107 );
buf ( n52109 , n52108 );
buf ( n52110 , n52109 );
buf ( n52111 , n41647 );
not ( n52112 , n52111 );
buf ( n52113 , n50977 );
not ( n52114 , n52113 );
or ( n52115 , n52112 , n52114 );
not ( n52116 , n41660 );
not ( n52117 , n43446 );
or ( n52118 , n52116 , n52117 );
nand ( n52119 , n50040 , n48390 );
nand ( n52120 , n52118 , n52119 );
buf ( n52121 , n52120 );
buf ( n52122 , n50982 );
nand ( n52123 , n52121 , n52122 );
buf ( n52124 , n52123 );
buf ( n52125 , n52124 );
nand ( n52126 , n52115 , n52125 );
buf ( n52127 , n52126 );
buf ( n52128 , n52127 );
xor ( n52129 , n52110 , n52128 );
buf ( n52130 , n43938 );
not ( n52131 , n52130 );
buf ( n52132 , n50045 );
buf ( n52133 , n42119 );
and ( n52134 , n52132 , n52133 );
not ( n52135 , n52132 );
buf ( n52136 , n28305 );
and ( n52137 , n52135 , n52136 );
nor ( n52138 , n52134 , n52137 );
buf ( n52139 , n52138 );
buf ( n52140 , n52139 );
not ( n52141 , n52140 );
or ( n52142 , n52131 , n52141 );
buf ( n52143 , n51729 );
buf ( n52144 , n46294 );
nand ( n52145 , n52143 , n52144 );
buf ( n52146 , n52145 );
buf ( n52147 , n52146 );
nand ( n52148 , n52142 , n52147 );
buf ( n52149 , n52148 );
buf ( n52150 , n52149 );
buf ( n52151 , n38404 );
not ( n52152 , n52151 );
buf ( n52153 , n43108 );
not ( n52154 , n52153 );
buf ( n52155 , n38411 );
not ( n52156 , n52155 );
or ( n52157 , n52154 , n52156 );
buf ( n52158 , n47068 );
buf ( n52159 , n43099 );
nand ( n52160 , n52158 , n52159 );
buf ( n52161 , n52160 );
buf ( n52162 , n52161 );
nand ( n52163 , n52157 , n52162 );
buf ( n52164 , n52163 );
buf ( n52165 , n52164 );
not ( n52166 , n52165 );
or ( n52167 , n52152 , n52166 );
buf ( n52168 , n51280 );
buf ( n52169 , n46606 );
not ( n52170 , n52169 );
buf ( n52171 , n52170 );
buf ( n52172 , n52171 );
not ( n52173 , n52172 );
buf ( n52174 , n52173 );
buf ( n52175 , n52174 );
nand ( n52176 , n52168 , n52175 );
buf ( n52177 , n52176 );
buf ( n52178 , n52177 );
nand ( n52179 , n52167 , n52178 );
buf ( n52180 , n52179 );
buf ( n52181 , n52180 );
xor ( n52182 , n52150 , n52181 );
buf ( n52183 , n50982 );
not ( n52184 , n52183 );
buf ( n52185 , n48390 );
not ( n52186 , n52185 );
buf ( n52187 , n46641 );
not ( n52188 , n52187 );
or ( n52189 , n52186 , n52188 );
buf ( n52190 , n42398 );
buf ( n52191 , n41660 );
nand ( n52192 , n52190 , n52191 );
buf ( n52193 , n52192 );
buf ( n52194 , n52193 );
nand ( n52195 , n52189 , n52194 );
buf ( n52196 , n52195 );
buf ( n52197 , n52196 );
not ( n52198 , n52197 );
or ( n52199 , n52184 , n52198 );
nand ( n52200 , n52120 , n48671 );
buf ( n52201 , n52200 );
nand ( n52202 , n52199 , n52201 );
buf ( n52203 , n52202 );
buf ( n52204 , n52203 );
and ( n52205 , n52182 , n52204 );
and ( n52206 , n52150 , n52181 );
or ( n52207 , n52205 , n52206 );
buf ( n52208 , n52207 );
buf ( n52209 , n52208 );
and ( n52210 , n52129 , n52209 );
and ( n52211 , n52110 , n52128 );
or ( n52212 , n52210 , n52211 );
buf ( n52213 , n52212 );
nand ( n52214 , n52082 , n52213 );
buf ( n52215 , n52214 );
nand ( n52216 , n52081 , n52066 );
buf ( n52217 , n52216 );
nand ( n52218 , n52215 , n52217 );
buf ( n52219 , n52218 );
buf ( n52220 , n52219 );
not ( n52221 , n52220 );
or ( n52222 , n52063 , n52221 );
buf ( n52223 , n52061 );
buf ( n52224 , n52219 );
or ( n52225 , n52223 , n52224 );
not ( n52226 , n41608 );
buf ( n52227 , n50463 );
not ( n52228 , n52227 );
buf ( n52229 , n52228 );
not ( n52230 , n52229 );
or ( n52231 , n52226 , n52230 );
buf ( n52232 , n50463 );
buf ( n52233 , n41611 );
nand ( n52234 , n52232 , n52233 );
buf ( n52235 , n52234 );
nand ( n52236 , n52231 , n52235 );
and ( n52237 , n52236 , n44267 );
and ( n52238 , n51135 , n43868 );
nor ( n52239 , n52237 , n52238 );
not ( n52240 , n52239 );
not ( n52241 , n52240 );
buf ( n52242 , n50060 );
not ( n52243 , n52242 );
buf ( n52244 , n36527 );
not ( n52245 , n52244 );
buf ( n52246 , n52245 );
buf ( n52247 , n52246 );
not ( n52248 , n52247 );
or ( n52249 , n52243 , n52248 );
nand ( n52250 , n50067 , n41715 );
buf ( n52251 , n52250 );
nand ( n52252 , n52249 , n52251 );
buf ( n52253 , n52252 );
buf ( n52254 , n52253 );
not ( n52255 , n52254 );
buf ( n52256 , n50374 );
not ( n52257 , n52256 );
or ( n52258 , n52255 , n52257 );
buf ( n52259 , n36643 );
buf ( n52260 , n51345 );
nand ( n52261 , n52259 , n52260 );
buf ( n52262 , n52261 );
buf ( n52263 , n52262 );
nand ( n52264 , n52258 , n52263 );
buf ( n52265 , n52264 );
buf ( n52266 , n52265 );
or ( n52267 , n51181 , n44682 );
buf ( n52268 , n46117 );
buf ( n52269 , n42082 );
and ( n52270 , n52268 , n52269 );
not ( n52271 , n52268 );
buf ( n52272 , n42062 );
and ( n52273 , n52271 , n52272 );
nor ( n52274 , n52270 , n52273 );
buf ( n52275 , n52274 );
or ( n52276 , n52275 , n44670 );
nand ( n52277 , n52267 , n52276 );
buf ( n52278 , n52277 );
or ( n52279 , n52266 , n52278 );
buf ( n52280 , n52279 );
buf ( n52281 , n52280 );
and ( n52282 , n41769 , n41721 );
not ( n52283 , n41769 );
and ( n52284 , n52283 , n42504 );
or ( n52285 , n52282 , n52284 );
not ( n52286 , n52285 );
not ( n52287 , n37397 );
or ( n52288 , n52286 , n52287 );
buf ( n52289 , n42132 );
not ( n52290 , n52289 );
buf ( n52291 , n51303 );
nand ( n52292 , n52290 , n52291 );
buf ( n52293 , n52292 );
nand ( n52294 , n52288 , n52293 );
buf ( n52295 , n52294 );
not ( n52296 , n52295 );
buf ( n52297 , n41843 );
buf ( n52298 , n43966 );
nand ( n52299 , n52297 , n52298 );
buf ( n52300 , n52299 );
nand ( n52301 , n41993 , n37472 );
nand ( n52302 , n52300 , n52301 );
not ( n52303 , n52302 );
not ( n52304 , n50671 );
or ( n52305 , n52303 , n52304 );
nand ( n52306 , n37440 , n51908 );
nand ( n52307 , n52305 , n52306 );
buf ( n52308 , n52307 );
not ( n52309 , n52308 );
or ( n52310 , n52296 , n52309 );
buf ( n52311 , n52294 );
not ( n52312 , n52311 );
buf ( n52313 , n52312 );
buf ( n52314 , n52313 );
not ( n52315 , n52314 );
buf ( n52316 , n52307 );
not ( n52317 , n52316 );
buf ( n52318 , n52317 );
buf ( n52319 , n52318 );
not ( n52320 , n52319 );
or ( n52321 , n52315 , n52320 );
not ( n52322 , n41862 );
buf ( n52323 , n52322 );
not ( n52324 , n52323 );
buf ( n52325 , n42862 );
buf ( n52326 , n41947 );
and ( n52327 , n52325 , n52326 );
not ( n52328 , n52325 );
buf ( n52329 , n41894 );
and ( n52330 , n52328 , n52329 );
nor ( n52331 , n52327 , n52330 );
buf ( n52332 , n52331 );
buf ( n52333 , n52332 );
not ( n52334 , n52333 );
and ( n52335 , n52324 , n52334 );
buf ( n52336 , n51751 );
not ( n52337 , n52336 );
buf ( n52338 , n37916 );
nor ( n52339 , n52337 , n52338 );
buf ( n52340 , n52339 );
buf ( n52341 , n52340 );
nor ( n52342 , n52335 , n52341 );
buf ( n52343 , n52342 );
not ( n52344 , n52343 );
buf ( n52345 , n52344 );
nand ( n52346 , n52321 , n52345 );
buf ( n52347 , n52346 );
buf ( n52348 , n52347 );
nand ( n52349 , n52310 , n52348 );
buf ( n52350 , n52349 );
buf ( n52351 , n52350 );
and ( n52352 , n52281 , n52351 );
buf ( n52353 , n52265 );
buf ( n52354 , n52277 );
and ( n52355 , n52353 , n52354 );
buf ( n52356 , n52355 );
buf ( n52357 , n52356 );
nor ( n52358 , n52352 , n52357 );
buf ( n52359 , n52358 );
buf ( n52360 , n52359 );
not ( n52361 , n52360 );
buf ( n52362 , n52361 );
not ( n52363 , n52362 );
or ( n52364 , n52241 , n52363 );
buf ( n52365 , n52239 );
not ( n52366 , n52365 );
buf ( n52367 , n52359 );
not ( n52368 , n52367 );
or ( n52369 , n52366 , n52368 );
xor ( n52370 , n51168 , n51175 );
xor ( n52371 , n52370 , n51192 );
buf ( n52372 , n52371 );
buf ( n52373 , n52372 );
nand ( n52374 , n52369 , n52373 );
buf ( n52375 , n52374 );
nand ( n52376 , n52364 , n52375 );
buf ( n52377 , n52376 );
nand ( n52378 , n52225 , n52377 );
buf ( n52379 , n52378 );
buf ( n52380 , n52379 );
nand ( n52381 , n52222 , n52380 );
buf ( n52382 , n52381 );
buf ( n52383 , n42847 );
not ( n52384 , n52383 );
buf ( n52385 , n43371 );
not ( n52386 , n52385 );
or ( n52387 , n52384 , n52386 );
buf ( n52388 , n44004 );
buf ( n52389 , n46691 );
nand ( n52390 , n52388 , n52389 );
buf ( n52391 , n52390 );
buf ( n52392 , n52391 );
nand ( n52393 , n52387 , n52392 );
buf ( n52394 , n52393 );
buf ( n52395 , n52394 );
not ( n52396 , n52395 );
buf ( n52397 , n46165 );
not ( n52398 , n52397 );
or ( n52399 , n52396 , n52398 );
not ( n52400 , n51154 );
nand ( n52401 , n52400 , n38060 );
buf ( n52402 , n52401 );
nand ( n52403 , n52399 , n52402 );
buf ( n52404 , n52403 );
not ( n52405 , n42339 );
not ( n52406 , n51327 );
or ( n52407 , n52405 , n52406 );
buf ( n52408 , n42378 );
not ( n52409 , n42350 );
not ( n52410 , n38821 );
or ( n52411 , n52409 , n52410 );
nand ( n52412 , n42343 , n47932 );
nand ( n52413 , n52411 , n52412 );
buf ( n52414 , n52413 );
nand ( n52415 , n52408 , n52414 );
buf ( n52416 , n52415 );
nand ( n52417 , n52407 , n52416 );
or ( n52418 , n52404 , n52417 );
and ( n52419 , n51265 , n51287 );
not ( n52420 , n51265 );
and ( n52421 , n52420 , n51284 );
or ( n52422 , n52419 , n52421 );
and ( n52423 , n52422 , n51310 );
not ( n52424 , n52422 );
not ( n52425 , n51310 );
and ( n52426 , n52424 , n52425 );
nor ( n52427 , n52423 , n52426 );
and ( n52428 , n52418 , n52427 );
buf ( n52429 , n52417 );
buf ( n52430 , n52404 );
and ( n52431 , n52429 , n52430 );
buf ( n52432 , n52431 );
nor ( n52433 , n52428 , n52432 );
buf ( n52434 , n52433 );
buf ( n52435 , n51488 );
not ( n52436 , n52435 );
buf ( n52437 , n48836 );
not ( n52438 , n52437 );
buf ( n52439 , n36035 );
not ( n52440 , n52439 );
or ( n52441 , n52438 , n52440 );
buf ( n52442 , n43857 );
not ( n52443 , n52442 );
buf ( n52444 , n52443 );
buf ( n52445 , n52444 );
buf ( n52446 , n51493 );
nand ( n52447 , n52445 , n52446 );
buf ( n52448 , n52447 );
buf ( n52449 , n52448 );
nand ( n52450 , n52441 , n52449 );
buf ( n52451 , n52450 );
buf ( n52452 , n52451 );
not ( n52453 , n52452 );
or ( n52454 , n52436 , n52453 );
buf ( n52455 , n51508 );
not ( n52456 , n51473 );
buf ( n52457 , n52456 );
nand ( n52458 , n52455 , n52457 );
buf ( n52459 , n52458 );
buf ( n52460 , n52459 );
nand ( n52461 , n52454 , n52460 );
buf ( n52462 , n52461 );
buf ( n52463 , n52462 );
not ( n52464 , n52463 );
buf ( n52465 , n52464 );
buf ( n52466 , n52465 );
xor ( n52467 , n52434 , n52466 );
xor ( n52468 , n51316 , n51332 );
xor ( n52469 , n52468 , n51358 );
buf ( n52470 , n52469 );
and ( n52471 , n52467 , n52470 );
and ( n52472 , n52434 , n52466 );
or ( n52473 , n52471 , n52472 );
buf ( n52474 , n52473 );
buf ( n52475 , n52474 );
not ( n52476 , n52475 );
buf ( n52477 , n52476 );
buf ( n52478 , n52477 );
not ( n52479 , n52478 );
buf ( n52480 , n51123 );
buf ( n52481 , n51203 );
xor ( n52482 , n52480 , n52481 );
buf ( n52483 , n51196 );
xor ( n52484 , n52482 , n52483 );
buf ( n52485 , n52484 );
buf ( n52486 , n52485 );
not ( n52487 , n52486 );
or ( n52488 , n52479 , n52487 );
buf ( n52489 , n52474 );
not ( n52490 , n52489 );
buf ( n52491 , n52485 );
not ( n52492 , n52491 );
buf ( n52493 , n52492 );
buf ( n52494 , n52493 );
not ( n52495 , n52494 );
or ( n52496 , n52490 , n52495 );
xor ( n52497 , n51712 , n51826 );
xor ( n52498 , n52497 , n51851 );
buf ( n52499 , n52498 );
not ( n52500 , n46246 );
not ( n52501 , n51681 );
or ( n52502 , n52500 , n52501 );
buf ( n52503 , n45753 );
not ( n52504 , n52503 );
buf ( n52505 , n50871 );
not ( n52506 , n52505 );
or ( n52507 , n52504 , n52506 );
buf ( n52508 , n50876 );
buf ( n52509 , n45750 );
nand ( n52510 , n52508 , n52509 );
buf ( n52511 , n52510 );
buf ( n52512 , n52511 );
nand ( n52513 , n52507 , n52512 );
buf ( n52514 , n52513 );
buf ( n52515 , n52514 );
buf ( n52516 , n46225 );
nand ( n52517 , n52515 , n52516 );
buf ( n52518 , n52517 );
nand ( n52519 , n52502 , n52518 );
xor ( n52520 , n52499 , n52519 );
buf ( n52521 , n50624 );
not ( n52522 , n52521 );
buf ( n52523 , n50599 );
not ( n52524 , n52523 );
or ( n52525 , n52522 , n52524 );
buf ( n52526 , n50591 );
buf ( n52527 , n47436 );
nand ( n52528 , n52526 , n52527 );
buf ( n52529 , n52528 );
buf ( n52530 , n52529 );
nand ( n52531 , n52525 , n52530 );
buf ( n52532 , n52531 );
buf ( n52533 , n52532 );
not ( n52534 , n52533 );
buf ( n52535 , n39998 );
not ( n52536 , n52535 );
buf ( n52537 , n52536 );
buf ( n52538 , n52537 );
not ( n52539 , n52538 );
or ( n52540 , n52534 , n52539 );
buf ( n52541 , n50605 );
buf ( n52542 , n48705 );
nand ( n52543 , n52541 , n52542 );
buf ( n52544 , n52543 );
buf ( n52545 , n52544 );
nand ( n52546 , n52540 , n52545 );
buf ( n52547 , n52546 );
not ( n52548 , n52547 );
buf ( n52549 , n48172 );
not ( n52550 , n52549 );
not ( n52551 , n24092 );
buf ( n52552 , n52551 );
not ( n52553 , n52552 );
or ( n52554 , n52550 , n52553 );
nand ( n52555 , n50598 , n42072 );
buf ( n52556 , n52555 );
nand ( n52557 , n52554 , n52556 );
buf ( n52558 , n52557 );
buf ( n52559 , n52558 );
not ( n52560 , n52559 );
buf ( n52561 , n52537 );
not ( n52562 , n52561 );
or ( n52563 , n52560 , n52562 );
buf ( n52564 , n52532 );
buf ( n52565 , n48705 );
nand ( n52566 , n52564 , n52565 );
buf ( n52567 , n52566 );
buf ( n52568 , n52567 );
nand ( n52569 , n52563 , n52568 );
buf ( n52570 , n52569 );
buf ( n52571 , n52570 );
not ( n52572 , n52571 );
buf ( n52573 , n52572 );
nand ( n52574 , n52548 , n52573 );
not ( n52575 , n52574 );
buf ( n52576 , n42049 );
not ( n52577 , n52576 );
buf ( n52578 , n47031 );
not ( n52579 , n52578 );
or ( n52580 , n52577 , n52579 );
buf ( n52581 , n42468 );
buf ( n52582 , n42052 );
nand ( n52583 , n52581 , n52582 );
buf ( n52584 , n52583 );
buf ( n52585 , n52584 );
nand ( n52586 , n52580 , n52585 );
buf ( n52587 , n52586 );
buf ( n52588 , n52587 );
not ( n52589 , n52588 );
buf ( n52590 , n47050 );
not ( n52591 , n52590 );
or ( n52592 , n52589 , n52591 );
buf ( n52593 , n51775 );
not ( n52594 , n47018 );
not ( n52595 , n52594 );
buf ( n52596 , n52595 );
nand ( n52597 , n52593 , n52596 );
buf ( n52598 , n52597 );
buf ( n52599 , n52598 );
nand ( n52600 , n52592 , n52599 );
buf ( n52601 , n52600 );
not ( n52602 , n52601 );
or ( n52603 , n52575 , n52602 );
buf ( n52604 , n52547 );
buf ( n52605 , n52570 );
nand ( n52606 , n52604 , n52605 );
buf ( n52607 , n52606 );
nand ( n52608 , n52603 , n52607 );
buf ( n52609 , n42378 );
not ( n52610 , n52609 );
buf ( n52611 , n42343 );
buf ( n52612 , n30187 );
and ( n52613 , n52611 , n52612 );
not ( n52614 , n52611 );
buf ( n52615 , n43308 );
and ( n52616 , n52614 , n52615 );
nor ( n52617 , n52613 , n52616 );
buf ( n52618 , n52617 );
buf ( n52619 , n52618 );
not ( n52620 , n52619 );
or ( n52621 , n52610 , n52620 );
buf ( n52622 , n52413 );
buf ( n52623 , n42339 );
nand ( n52624 , n52622 , n52623 );
buf ( n52625 , n52624 );
buf ( n52626 , n52625 );
nand ( n52627 , n52621 , n52626 );
buf ( n52628 , n52627 );
xor ( n52629 , n52608 , n52628 );
xor ( n52630 , n51763 , n51788 );
xor ( n52631 , n52630 , n51816 );
buf ( n52632 , n52631 );
and ( n52633 , n52629 , n52632 );
and ( n52634 , n52608 , n52628 );
or ( n52635 , n52633 , n52634 );
buf ( n52636 , n52635 );
buf ( n52637 , n42315 );
not ( n52638 , n52637 );
buf ( n52639 , n51879 );
not ( n52640 , n52639 );
or ( n52641 , n52638 , n52640 );
buf ( n52642 , n42266 );
not ( n52643 , n52642 );
buf ( n52644 , n39518 );
not ( n52645 , n52644 );
or ( n52646 , n52643 , n52645 );
buf ( n52647 , n39522 );
buf ( n52648 , n42263 );
nand ( n52649 , n52647 , n52648 );
buf ( n52650 , n52649 );
buf ( n52651 , n52650 );
nand ( n52652 , n52646 , n52651 );
buf ( n52653 , n52652 );
buf ( n52654 , n52653 );
buf ( n52655 , n42252 );
nand ( n52656 , n52654 , n52655 );
buf ( n52657 , n52656 );
buf ( n52658 , n52657 );
nand ( n52659 , n52641 , n52658 );
buf ( n52660 , n52659 );
buf ( n52661 , n52660 );
xor ( n52662 , n52636 , n52661 );
buf ( n52663 , n47872 );
not ( n52664 , n52663 );
buf ( n52665 , n51808 );
not ( n52666 , n52665 );
or ( n52667 , n52664 , n52666 );
buf ( n52668 , n39973 );
not ( n52669 , n52668 );
buf ( n52670 , n52669 );
buf ( n52671 , n52670 );
not ( n52672 , n52671 );
buf ( n52673 , n52672 );
not ( n52674 , n52673 );
not ( n52675 , n47072 );
or ( n52676 , n52674 , n52675 );
nand ( n52677 , n50575 , n51804 );
nand ( n52678 , n52676 , n52677 );
buf ( n52679 , n52678 );
buf ( n52680 , n50128 );
nand ( n52681 , n52679 , n52680 );
buf ( n52682 , n52681 );
buf ( n52683 , n52682 );
nand ( n52684 , n52667 , n52683 );
buf ( n52685 , n52684 );
buf ( n52686 , n52685 );
buf ( n52687 , n41736 );
not ( n52688 , n52687 );
buf ( n52689 , n45069 );
not ( n52690 , n52689 );
or ( n52691 , n52688 , n52690 );
buf ( n52692 , n47068 );
buf ( n52693 , n41748 );
nand ( n52694 , n52692 , n52693 );
buf ( n52695 , n52694 );
buf ( n52696 , n52695 );
nand ( n52697 , n52691 , n52696 );
buf ( n52698 , n52697 );
buf ( n52699 , n52698 );
not ( n52700 , n52699 );
buf ( n52701 , n38404 );
not ( n52702 , n52701 );
or ( n52703 , n52700 , n52702 );
buf ( n52704 , n52164 );
buf ( n52705 , n46606 );
nand ( n52706 , n52704 , n52705 );
buf ( n52707 , n52706 );
buf ( n52708 , n52707 );
nand ( n52709 , n52703 , n52708 );
buf ( n52710 , n52709 );
buf ( n52711 , n52710 );
or ( n52712 , n52686 , n52711 );
buf ( n52713 , n46294 );
not ( n52714 , n52713 );
buf ( n52715 , n52139 );
not ( n52716 , n52715 );
or ( n52717 , n52714 , n52716 );
buf ( n52718 , n48357 );
not ( n52719 , n52718 );
buf ( n52720 , n29325 );
not ( n52721 , n52720 );
or ( n52722 , n52719 , n52721 );
buf ( n52723 , n29328 );
not ( n52724 , n42559 );
not ( n52725 , n52724 );
buf ( n52726 , n52725 );
nand ( n52727 , n52723 , n52726 );
buf ( n52728 , n52727 );
buf ( n52729 , n52728 );
nand ( n52730 , n52722 , n52729 );
buf ( n52731 , n52730 );
buf ( n52732 , n52731 );
buf ( n52733 , n43938 );
nand ( n52734 , n52732 , n52733 );
buf ( n52735 , n52734 );
buf ( n52736 , n52735 );
nand ( n52737 , n52717 , n52736 );
buf ( n52738 , n52737 );
buf ( n52739 , n52738 );
nand ( n52740 , n52712 , n52739 );
buf ( n52741 , n52740 );
buf ( n52742 , n52741 );
buf ( n52743 , n52710 );
buf ( n52744 , n52685 );
nand ( n52745 , n52743 , n52744 );
buf ( n52746 , n52745 );
buf ( n52747 , n52746 );
nand ( n52748 , n52742 , n52747 );
buf ( n52749 , n52748 );
buf ( n52750 , n48323 );
not ( n52751 , n52750 );
buf ( n52752 , n39493 );
not ( n52753 , n52752 );
or ( n52754 , n52751 , n52753 );
buf ( n52755 , n43265 );
buf ( n52756 , n48320 );
nand ( n52757 , n52755 , n52756 );
buf ( n52758 , n52757 );
buf ( n52759 , n52758 );
nand ( n52760 , n52754 , n52759 );
buf ( n52761 , n52760 );
buf ( n52762 , n52761 );
not ( n52763 , n52762 );
buf ( n52764 , n36101 );
not ( n52765 , n52764 );
or ( n52766 , n52763 , n52765 );
buf ( n52767 , n42530 );
buf ( n52768 , n51932 );
nand ( n52769 , n52767 , n52768 );
buf ( n52770 , n52769 );
buf ( n52771 , n52770 );
nand ( n52772 , n52766 , n52771 );
buf ( n52773 , n52772 );
xor ( n52774 , n52749 , n52773 );
xor ( n52775 , n12439 , n12506 );
xor ( n52776 , n52775 , n12524 );
buf ( n52777 , n52776 );
buf ( n52778 , n52777 );
buf ( n52779 , n52778 );
buf ( n52780 , n52779 );
buf ( n52781 , n52780 );
not ( n52782 , n52781 );
buf ( n52783 , n38837 );
not ( n52784 , n52783 );
or ( n52785 , n52782 , n52784 );
buf ( n52786 , n38798 );
buf ( n52787 , n52780 );
not ( n52788 , n52787 );
buf ( n52789 , n52788 );
buf ( n52790 , n52789 );
nand ( n52791 , n52786 , n52790 );
buf ( n52792 , n52791 );
buf ( n52793 , n52792 );
nand ( n52794 , n52785 , n52793 );
buf ( n52795 , n52794 );
buf ( n52796 , n42004 );
buf ( n52797 , n52102 );
or ( n52798 , n52796 , n52797 );
nand ( n52799 , C1 , n52798 );
buf ( n52800 , n52799 );
and ( n52801 , n52774 , n52800 );
and ( n52802 , n52749 , n52773 );
or ( n52803 , n52801 , n52802 );
buf ( n52804 , n52803 );
and ( n52805 , n52662 , n52804 );
and ( n52806 , n52636 , n52661 );
or ( n52807 , n52805 , n52806 );
buf ( n52808 , n52807 );
and ( n52809 , n52520 , n52808 );
and ( n52810 , n52499 , n52519 );
or ( n52811 , n52809 , n52810 );
buf ( n52812 , n52811 );
nand ( n52813 , n52496 , n52812 );
buf ( n52814 , n52813 );
buf ( n52815 , n52814 );
nand ( n52816 , n52488 , n52815 );
buf ( n52817 , n52816 );
xor ( n52818 , n52382 , n52817 );
buf ( n52819 , n51519 );
buf ( n52820 , n51544 );
xor ( n52821 , n52819 , n52820 );
buf ( n52822 , n51530 );
xor ( n52823 , n52821 , n52822 );
buf ( n52824 , n52823 );
and ( n52825 , n52818 , n52824 );
and ( n52826 , n52382 , n52817 );
or ( n52827 , n52825 , n52826 );
not ( n52828 , n52827 );
xor ( n52829 , n51550 , n51403 );
xor ( n52830 , n52829 , n51557 );
buf ( n52831 , n51106 );
buf ( n52832 , n51113 );
xor ( n52833 , n52831 , n52832 );
buf ( n52834 , n51387 );
xor ( n52835 , n52833 , n52834 );
buf ( n52836 , n52835 );
nand ( n52837 , n52830 , n52836 );
not ( n52838 , n52837 );
or ( n52839 , n52828 , n52838 );
buf ( n52840 , n52836 );
not ( n52841 , n52840 );
not ( n52842 , n52830 );
buf ( n52843 , n52842 );
nand ( n52844 , n52841 , n52843 );
buf ( n52845 , n52844 );
nand ( n52846 , n52839 , n52845 );
buf ( n52847 , n51607 );
buf ( n52848 , n52034 );
nand ( n52849 , n52847 , n52848 );
buf ( n52850 , n52849 );
and ( n52851 , n52846 , n52850 );
nor ( n52852 , n52036 , n52851 );
buf ( n52853 , n52852 );
not ( n52854 , n52853 );
buf ( n52855 , n52854 );
nand ( n52856 , n51601 , n52855 );
nand ( n52857 , n51597 , n52856 );
not ( n52858 , n52857 );
nand ( n52859 , n51584 , n52858 );
xor ( n52860 , n51572 , n51573 );
buf ( n52861 , n52860 );
buf ( n52862 , n52861 );
buf ( n52863 , n51569 );
xor ( n52864 , n52862 , n52863 );
buf ( n52865 , n52864 );
buf ( n52866 , n52865 );
xor ( n52867 , n51977 , n51987 );
xor ( n52868 , n52867 , n52030 );
buf ( n52869 , n52868 );
not ( n52870 , n52869 );
xor ( n52871 , n51970 , n51971 );
buf ( n52872 , n52871 );
xnor ( n52873 , n52872 , n51967 );
buf ( n52874 , n52873 );
not ( n52875 , n52874 );
buf ( n52876 , n52875 );
buf ( n52877 , n52876 );
not ( n52878 , n52877 );
xor ( n52879 , n52000 , n52023 );
xor ( n52880 , n52879 , n52026 );
not ( n52881 , n52880 );
buf ( n52882 , n52881 );
not ( n52883 , n52882 );
or ( n52884 , n52878 , n52883 );
buf ( n52885 , n52873 );
not ( n52886 , n52885 );
buf ( n52887 , n52880 );
not ( n52888 , n52887 );
or ( n52889 , n52886 , n52888 );
xor ( n52890 , n51433 , n51511 );
not ( n52891 , n51457 );
xor ( n52892 , n52890 , n52891 );
buf ( n52893 , n52892 );
xor ( n52894 , n51376 , n51243 );
xor ( n52895 , n52894 , n51361 );
buf ( n52896 , n52895 );
xor ( n52897 , n52893 , n52896 );
xor ( n52898 , n51737 , n51758 );
xor ( n52899 , n52898 , n51821 );
buf ( n52900 , n52899 );
buf ( n52901 , n52900 );
buf ( n52902 , n42668 );
not ( n52903 , n52902 );
buf ( n52904 , n51840 );
not ( n52905 , n52904 );
or ( n52906 , n52903 , n52905 );
buf ( n52907 , n42672 );
not ( n52908 , n52907 );
buf ( n52909 , n37595 );
not ( n52910 , n52909 );
or ( n52911 , n52908 , n52910 );
buf ( n52912 , n37586 );
buf ( n52913 , n42679 );
nand ( n52914 , n52912 , n52913 );
buf ( n52915 , n52914 );
buf ( n52916 , n52915 );
nand ( n52917 , n52911 , n52916 );
buf ( n52918 , n52917 );
buf ( n52919 , n52918 );
buf ( n52920 , n42712 );
nand ( n52921 , n52919 , n52920 );
buf ( n52922 , n52921 );
buf ( n52923 , n52922 );
nand ( n52924 , n52906 , n52923 );
buf ( n52925 , n52924 );
buf ( n52926 , n52925 );
xor ( n52927 , n52901 , n52926 );
xor ( n52928 , n52110 , n52128 );
xor ( n52929 , n52928 , n52209 );
buf ( n52930 , n52929 );
buf ( n52931 , n52930 );
and ( n52932 , n52927 , n52931 );
and ( n52933 , n52901 , n52926 );
or ( n52934 , n52932 , n52933 );
buf ( n52935 , n52934 );
buf ( n52936 , n52935 );
buf ( n52937 , n48855 );
not ( n52938 , n52937 );
buf ( n52939 , n48808 );
not ( n52940 , n52939 );
buf ( n52941 , n39930 );
not ( n52942 , n52941 );
or ( n52943 , n52940 , n52942 );
buf ( n52944 , n39924 );
buf ( n52945 , n48818 );
nand ( n52946 , n52944 , n52945 );
buf ( n52947 , n52946 );
buf ( n52948 , n52947 );
nand ( n52949 , n52943 , n52948 );
buf ( n52950 , n52949 );
buf ( n52951 , n52950 );
not ( n52952 , n52951 );
or ( n52953 , n52938 , n52952 );
buf ( n52954 , n51426 );
buf ( n52955 , n48868 );
nand ( n52956 , n52954 , n52955 );
buf ( n52957 , n52956 );
buf ( n52958 , n52957 );
nand ( n52959 , n52953 , n52958 );
buf ( n52960 , n52959 );
buf ( n52961 , n52960 );
xor ( n52962 , n52936 , n52961 );
buf ( n52963 , n44952 );
buf ( n52964 , n43371 );
and ( n52965 , n52963 , n52964 );
not ( n52966 , n52963 );
buf ( n52967 , n45376 );
and ( n52968 , n52966 , n52967 );
nor ( n52969 , n52965 , n52968 );
buf ( n52970 , n52969 );
buf ( n52971 , n52970 );
not ( n52972 , n52971 );
buf ( n52973 , n52972 );
buf ( n52974 , n52973 );
not ( n52975 , n52974 );
buf ( n52976 , n43386 );
not ( n52977 , n52976 );
or ( n52978 , n52975 , n52977 );
buf ( n52979 , n52394 );
buf ( n52980 , n45144 );
nand ( n52981 , n52979 , n52980 );
buf ( n52982 , n52981 );
buf ( n52983 , n52982 );
nand ( n52984 , n52978 , n52983 );
buf ( n52985 , n52984 );
buf ( n52986 , n52985 );
not ( n52987 , n52986 );
buf ( n52988 , n52987 );
buf ( n52989 , n52988 );
not ( n52990 , n52989 );
not ( n52991 , n42712 );
buf ( n52992 , n42672 );
not ( n52993 , n52992 );
buf ( n52994 , n39701 );
not ( n52995 , n52994 );
or ( n52996 , n52993 , n52995 );
buf ( n52997 , n37641 );
buf ( n52998 , n42679 );
nand ( n52999 , n52997 , n52998 );
buf ( n53000 , n52999 );
buf ( n53001 , n53000 );
nand ( n53002 , n52996 , n53001 );
buf ( n53003 , n53002 );
not ( n53004 , n53003 );
or ( n53005 , n52991 , n53004 );
buf ( n53006 , n52918 );
buf ( n53007 , n42668 );
nand ( n53008 , n53006 , n53007 );
buf ( n53009 , n53008 );
nand ( n53010 , n53005 , n53009 );
not ( n53011 , n53010 );
buf ( n53012 , n53011 );
not ( n53013 , n53012 );
or ( n53014 , n52990 , n53013 );
xor ( n53015 , n52150 , n52181 );
xor ( n53016 , n53015 , n52204 );
buf ( n53017 , n53016 );
buf ( n53018 , n53017 );
nand ( n53019 , n53014 , n53018 );
buf ( n53020 , n53019 );
buf ( n53021 , n53020 );
buf ( n53022 , n53010 );
buf ( n53023 , n52985 );
nand ( n53024 , n53022 , n53023 );
buf ( n53025 , n53024 );
buf ( n53026 , n53025 );
nand ( n53027 , n53021 , n53026 );
buf ( n53028 , n53027 );
buf ( n53029 , n53028 );
xor ( n53030 , n51895 , n51919 );
xor ( n53031 , n53030 , n51947 );
buf ( n53032 , n53031 );
xor ( n53033 , n53029 , n53032 );
not ( n53034 , n44496 );
not ( n53035 , n52074 );
or ( n53036 , n53034 , n53035 );
not ( n53037 , n44518 );
buf ( n53038 , n44533 );
buf ( n53039 , n38247 );
and ( n53040 , n53038 , n53039 );
not ( n53041 , n53038 );
buf ( n53042 , n38247 );
not ( n53043 , n53042 );
buf ( n53044 , n53043 );
buf ( n53045 , n53044 );
and ( n53046 , n53041 , n53045 );
nor ( n53047 , n53040 , n53046 );
buf ( n53048 , n53047 );
nand ( n53049 , n53037 , n53048 );
nand ( n53050 , n53036 , n53049 );
buf ( n53051 , n53050 );
and ( n53052 , n53033 , n53051 );
and ( n53053 , n53029 , n53032 );
or ( n53054 , n53052 , n53053 );
buf ( n53055 , n53054 );
buf ( n53056 , n53055 );
and ( n53057 , n52962 , n53056 );
and ( n53058 , n52936 , n52961 );
or ( n53059 , n53057 , n53058 );
buf ( n53060 , n53059 );
buf ( n53061 , n53060 );
and ( n53062 , n52897 , n53061 );
and ( n53063 , n52893 , n52896 );
or ( n53064 , n53062 , n53063 );
buf ( n53065 , n53064 );
buf ( n53066 , n53065 );
nand ( n53067 , n52889 , n53066 );
buf ( n53068 , n53067 );
buf ( n53069 , n53068 );
nand ( n53070 , n52884 , n53069 );
buf ( n53071 , n53070 );
buf ( n53072 , n53071 );
not ( n53073 , n53072 );
buf ( n53074 , n53073 );
not ( n53075 , n53074 );
or ( n53076 , n52870 , n53075 );
buf ( n53077 , n51855 );
buf ( n53078 , n51707 );
xor ( n53079 , n53077 , n53078 );
buf ( n53080 , n51956 );
xnor ( n53081 , n53079 , n53080 );
buf ( n53082 , n53081 );
buf ( n53083 , n53082 );
xor ( n53084 , n52213 , n52066 );
xnor ( n53085 , n53084 , n52081 );
not ( n53086 , n53085 );
not ( n53087 , n47331 );
buf ( n53088 , n36396 );
buf ( n53089 , n46890 );
nand ( n53090 , n53088 , n53089 );
buf ( n53091 , n53090 );
nand ( n53092 , n51622 , n39891 );
nand ( n53093 , n53091 , n53092 );
not ( n53094 , n53093 );
or ( n53095 , n53087 , n53094 );
buf ( n53096 , n51634 );
buf ( n53097 , n46912 );
nand ( n53098 , n53096 , n53097 );
buf ( n53099 , n53098 );
nand ( n53100 , n53095 , n53099 );
not ( n53101 , n53100 );
not ( n53102 , n53101 );
and ( n53103 , n53086 , n53102 );
buf ( n53104 , n53085 );
buf ( n53105 , n53101 );
nand ( n53106 , n53104 , n53105 );
buf ( n53107 , n53106 );
and ( n53108 , n51886 , n51861 );
not ( n53109 , n51886 );
not ( n53110 , n51861 );
and ( n53111 , n53109 , n53110 );
nor ( n53112 , n53108 , n53111 );
and ( n53113 , n53112 , n51950 );
not ( n53114 , n53112 );
not ( n53115 , n51950 );
and ( n53116 , n53114 , n53115 );
nor ( n53117 , n53113 , n53116 );
not ( n53118 , n53117 );
not ( n53119 , n53118 );
and ( n53120 , n53107 , n53119 );
nor ( n53121 , n53103 , n53120 );
buf ( n53122 , n53121 );
xor ( n53123 , n53083 , n53122 );
xor ( n53124 , n52219 , n52058 );
xor ( n53125 , n53124 , n52376 );
buf ( n53126 , n53125 );
and ( n53127 , n53123 , n53126 );
and ( n53128 , n53083 , n53122 );
or ( n53129 , n53127 , n53128 );
buf ( n53130 , n53129 );
not ( n53131 , n53130 );
xor ( n53132 , n51661 , n51696 );
xor ( n53133 , n53132 , n51688 );
buf ( n53134 , n53133 );
xor ( n53135 , n52434 , n52466 );
xor ( n53136 , n53135 , n52470 );
buf ( n53137 , n53136 );
not ( n53138 , n53137 );
buf ( n53139 , n52456 );
not ( n53140 , n53139 );
buf ( n53141 , n52451 );
not ( n53142 , n53141 );
or ( n53143 , n53140 , n53142 );
not ( n53144 , n51496 );
not ( n53145 , n39582 );
or ( n53146 , n53144 , n53145 );
buf ( n53147 , n36611 );
buf ( n53148 , n51493 );
nand ( n53149 , n53147 , n53148 );
buf ( n53150 , n53149 );
nand ( n53151 , n53146 , n53150 );
nand ( n53152 , n53151 , n51488 );
buf ( n53153 , n53152 );
nand ( n53154 , n53143 , n53153 );
buf ( n53155 , n53154 );
not ( n53156 , n53155 );
buf ( n53157 , n44538 );
not ( n53158 , n53157 );
buf ( n53159 , n53158 );
buf ( n53160 , C1 );
or ( n53161 , n53156 , C0 );
xor ( n53162 , n52353 , n52354 );
buf ( n53163 , n53162 );
xor ( n53164 , n52350 , n53163 );
nand ( n53165 , C1 , n53164 );
nand ( n53166 , n53161 , n53165 );
not ( n53167 , n53166 );
not ( n53168 , n53167 );
or ( n53169 , n53138 , n53168 );
nor ( n53170 , n53167 , n53137 );
not ( n53171 , n43868 );
not ( n53172 , n52236 );
or ( n53173 , n53171 , n53172 );
buf ( n53174 , n41608 );
not ( n53175 , n53174 );
buf ( n53176 , n38286 );
not ( n53177 , n53176 );
or ( n53178 , n53175 , n53177 );
buf ( n53179 , n37293 );
buf ( n53180 , n41611 );
nand ( n53181 , n53179 , n53180 );
buf ( n53182 , n53181 );
buf ( n53183 , n53182 );
nand ( n53184 , n53178 , n53183 );
buf ( n53185 , n53184 );
buf ( n53186 , n53185 );
buf ( n53187 , n44267 );
nand ( n53188 , n53186 , n53187 );
buf ( n53189 , n53188 );
nand ( n53190 , n53173 , n53189 );
buf ( n53191 , n53190 );
xor ( n53192 , n52429 , n52430 );
buf ( n53193 , n53192 );
and ( n53194 , n53193 , n52427 );
not ( n53195 , n53193 );
not ( n53196 , n52427 );
and ( n53197 , n53195 , n53196 );
nor ( n53198 , n53194 , n53197 );
buf ( n53199 , n53198 );
xor ( n53200 , n53191 , n53199 );
not ( n53201 , n44141 );
not ( n53202 , n52253 );
or ( n53203 , n53201 , n53202 );
and ( n53204 , n51004 , n43959 );
not ( n53205 , n51004 );
and ( n53206 , n53205 , n36527 );
or ( n53207 , n53204 , n53206 );
nand ( n53208 , n39803 , n53207 );
nand ( n53209 , n53203 , n53208 );
buf ( n53210 , n53209 );
buf ( n53211 , n46390 );
buf ( n53212 , n42062 );
not ( n53213 , n53212 );
xor ( n53214 , n53211 , n53213 );
buf ( n53215 , n53214 );
buf ( n53216 , n53215 );
not ( n53217 , n53216 );
buf ( n53218 , n53217 );
buf ( n53219 , n53218 );
not ( n53220 , n53219 );
buf ( n53221 , n45158 );
not ( n53222 , n53221 );
or ( n53223 , n53220 , n53222 );
buf ( n53224 , n52275 );
not ( n53225 , n53224 );
buf ( n53226 , n44679 );
nand ( n53227 , n53225 , n53226 );
buf ( n53228 , n53227 );
buf ( n53229 , n53228 );
nand ( n53230 , n53223 , n53229 );
buf ( n53231 , n53230 );
buf ( n53232 , n53231 );
xor ( n53233 , n53210 , n53232 );
buf ( n53234 , n42008 );
not ( n53235 , n53234 );
buf ( n53236 , n43442 );
not ( n53237 , n53236 );
or ( n53238 , n53235 , n53237 );
buf ( n53239 , n41779 );
buf ( n53240 , n42017 );
nand ( n53241 , n53239 , n53240 );
buf ( n53242 , n53241 );
buf ( n53243 , n53242 );
nand ( n53244 , n53238 , n53243 );
buf ( n53245 , n53244 );
buf ( n53246 , n53245 );
not ( n53247 , n53246 );
buf ( n53248 , n37397 );
not ( n53249 , n53248 );
or ( n53250 , n53247 , n53249 );
nand ( n53251 , n45108 , n52285 );
buf ( n53252 , n53251 );
nand ( n53253 , n53250 , n53252 );
buf ( n53254 , n53253 );
buf ( n53255 , n53254 );
buf ( n53256 , n48671 );
not ( n53257 , n53256 );
buf ( n53258 , n52196 );
not ( n53259 , n53258 );
or ( n53260 , n53257 , n53259 );
buf ( n53261 , n41762 );
not ( n53262 , n53261 );
buf ( n53263 , n41660 );
not ( n53264 , n53263 );
and ( n53265 , n53262 , n53264 );
buf ( n53266 , n41782 );
buf ( n53267 , n41660 );
and ( n53268 , n53266 , n53267 );
nor ( n53269 , n53265 , n53268 );
buf ( n53270 , n53269 );
buf ( n53271 , n53270 );
not ( n53272 , n53271 );
buf ( n53273 , n50982 );
nand ( n53274 , n53272 , n53273 );
buf ( n53275 , n53274 );
buf ( n53276 , n53275 );
nand ( n53277 , n53260 , n53276 );
buf ( n53278 , n53277 );
buf ( n53279 , n53278 );
xor ( n53280 , n53255 , n53279 );
buf ( n53281 , n43063 );
not ( n53282 , n53281 );
buf ( n53283 , n48207 );
not ( n53284 , n53283 );
or ( n53285 , n53282 , n53284 );
buf ( n53286 , n37473 );
buf ( n53287 , n43064 );
nand ( n53288 , n53286 , n53287 );
buf ( n53289 , n53288 );
buf ( n53290 , n53289 );
nand ( n53291 , n53285 , n53290 );
buf ( n53292 , n53291 );
buf ( n53293 , n53292 );
not ( n53294 , n53293 );
buf ( n53295 , n44338 );
not ( n53296 , n53295 );
or ( n53297 , n53294 , n53296 );
nand ( n53298 , n52302 , n41852 );
buf ( n53299 , n53298 );
nand ( n53300 , n53297 , n53299 );
buf ( n53301 , n53300 );
buf ( n53302 , n53301 );
and ( n53303 , n53280 , n53302 );
and ( n53304 , n53255 , n53279 );
or ( n53305 , n53303 , n53304 );
buf ( n53306 , n53305 );
buf ( n53307 , n53306 );
and ( n53308 , n53233 , n53307 );
and ( n53309 , n53210 , n53232 );
or ( n53310 , n53308 , n53309 );
buf ( n53311 , n53310 );
buf ( n53312 , n53311 );
and ( n53313 , n53200 , n53312 );
and ( n53314 , n53191 , n53199 );
or ( n53315 , n53313 , n53314 );
buf ( n53316 , n53315 );
or ( n53317 , n53170 , n53316 );
nand ( n53318 , n53169 , n53317 );
buf ( n53319 , n53318 );
xor ( n53320 , n53134 , n53319 );
buf ( n53321 , n52485 );
buf ( n53322 , n52477 );
and ( n53323 , n53321 , n53322 );
not ( n53324 , n53321 );
buf ( n53325 , n52474 );
and ( n53326 , n53324 , n53325 );
nor ( n53327 , n53323 , n53326 );
buf ( n53328 , n53327 );
xnor ( n53329 , n53328 , n52811 );
buf ( n53330 , n53329 );
and ( n53331 , n53320 , n53330 );
and ( n53332 , n53134 , n53319 );
or ( n53333 , n53331 , n53332 );
buf ( n53334 , n53333 );
not ( n53335 , n53334 );
or ( n53336 , n53131 , n53335 );
xor ( n53337 , n52382 , n52817 );
xor ( n53338 , n53337 , n52824 );
nand ( n53339 , n53336 , n53338 );
not ( n53340 , n53130 );
buf ( n53341 , n53334 );
not ( n53342 , n53341 );
buf ( n53343 , n53342 );
nand ( n53344 , n53340 , n53343 );
nand ( n53345 , n53339 , n53344 );
nand ( n53346 , n53076 , n53345 );
buf ( n53347 , n53346 );
buf ( n53348 , n52869 );
not ( n53349 , n53348 );
buf ( n53350 , n53071 );
nand ( n53351 , n53349 , n53350 );
buf ( n53352 , n53351 );
buf ( n53353 , n53352 );
nand ( n53354 , n53347 , n53353 );
buf ( n53355 , n53354 );
buf ( n53356 , n53355 );
xor ( n53357 , n52866 , n53356 );
buf ( n53358 , n52846 );
not ( n53359 , n53358 );
xnor ( n53360 , n51607 , n52034 );
buf ( n53361 , n53360 );
not ( n53362 , n53361 );
or ( n53363 , n53359 , n53362 );
buf ( n53364 , n52846 );
buf ( n53365 , n53360 );
or ( n53366 , n53364 , n53365 );
nand ( n53367 , n53363 , n53366 );
buf ( n53368 , n53367 );
buf ( n53369 , n53368 );
and ( n53370 , n53357 , n53369 );
and ( n53371 , n52866 , n53356 );
or ( n53372 , n53370 , n53371 );
buf ( n53373 , n53372 );
buf ( n53374 , n53373 );
not ( n53375 , n53374 );
buf ( n53376 , n53375 );
not ( n53377 , n51590 );
not ( n53378 , n52852 );
not ( n53379 , n53378 );
or ( n53380 , n53377 , n53379 );
nand ( n53381 , n51598 , n52852 );
nand ( n53382 , n53380 , n53381 );
not ( n53383 , n51594 );
and ( n53384 , n53382 , n53383 );
not ( n53385 , n53382 );
not ( n53386 , n51595 );
and ( n53387 , n53385 , n53386 );
nor ( n53388 , n53384 , n53387 );
nand ( n53389 , n53376 , n53388 );
nand ( n53390 , n52859 , n53389 );
not ( n53391 , n53390 );
buf ( n53392 , n53391 );
buf ( n53393 , n47238 );
buf ( n53394 , n47370 );
xor ( n53395 , n53393 , n53394 );
buf ( n53396 , n47243 );
xnor ( n53397 , n53395 , n53396 );
buf ( n53398 , n53397 );
buf ( n53399 , n53398 );
buf ( n53400 , n50219 );
not ( n53401 , n53400 );
buf ( n53402 , n49715 );
not ( n53403 , n53402 );
or ( n53404 , n53401 , n53403 );
buf ( n53405 , n50845 );
buf ( n53406 , n49715 );
not ( n53407 , n53406 );
buf ( n53408 , n50224 );
nand ( n53409 , n53407 , n53408 );
buf ( n53410 , n53409 );
buf ( n53411 , n53410 );
nand ( n53412 , n53405 , n53411 );
buf ( n53413 , n53412 );
buf ( n53414 , n53413 );
nand ( n53415 , n53404 , n53414 );
buf ( n53416 , n53415 );
buf ( n53417 , n53416 );
not ( n53418 , n53417 );
buf ( n53419 , n53418 );
buf ( n53420 , n53419 );
xor ( n53421 , n53399 , n53420 );
xor ( n53422 , n48143 , n48566 );
xor ( n53423 , n53422 , n49119 );
buf ( n53424 , n53423 );
buf ( n53425 , n53424 );
xor ( n53426 , n53421 , n53425 );
buf ( n53427 , n53426 );
xor ( n53428 , n49696 , n50850 );
and ( n53429 , n53428 , n51583 );
and ( n53430 , n49696 , n50850 );
or ( n53431 , n53429 , n53430 );
nand ( n53432 , n53427 , n53431 );
xor ( n53433 , n48125 , n48135 );
xor ( n53434 , n53433 , n49124 );
buf ( n53435 , n53434 );
xor ( n53436 , n53399 , n53420 );
and ( n53437 , n53436 , n53425 );
and ( n53438 , n53399 , n53420 );
or ( n53439 , n53437 , n53438 );
buf ( n53440 , n53439 );
nand ( n53441 , n53435 , n53440 );
and ( n53442 , n53432 , n53441 );
buf ( n53443 , n53442 );
and ( n53444 , n53392 , n53443 );
buf ( n53445 , n53444 );
nand ( n53446 , n49693 , n53445 );
not ( n53447 , n53446 );
not ( n53448 , n52836 );
and ( n53449 , n52827 , n53448 );
not ( n53450 , n52827 );
and ( n53451 , n53450 , n52836 );
nor ( n53452 , n53449 , n53451 );
buf ( n53453 , n53452 );
not ( n53454 , n52842 );
buf ( n53455 , n53454 );
and ( n53456 , n53453 , n53455 );
not ( n53457 , n53453 );
buf ( n53458 , n52842 );
and ( n53459 , n53457 , n53458 );
nor ( n53460 , n53456 , n53459 );
buf ( n53461 , n53460 );
not ( n53462 , n52869 );
not ( n53463 , n53462 );
not ( n53464 , n53074 );
or ( n53465 , n53463 , n53464 );
nand ( n53466 , n52869 , n53071 );
nand ( n53467 , n53465 , n53466 );
not ( n53468 , n53345 );
and ( n53469 , n53467 , n53468 );
not ( n53470 , n53467 );
and ( n53471 , n53470 , n53345 );
nor ( n53472 , n53469 , n53471 );
xor ( n53473 , n53461 , n53472 );
xor ( n53474 , n52893 , n52896 );
xor ( n53475 , n53474 , n53061 );
buf ( n53476 , n53475 );
buf ( n53477 , n53476 );
xor ( n53478 , n52239 , n52372 );
xnor ( n53479 , n53478 , n52362 );
buf ( n53480 , n53479 );
xor ( n53481 , n52499 , n52519 );
xor ( n53482 , n53481 , n52808 );
buf ( n53483 , n53482 );
xor ( n53484 , n53480 , n53483 );
buf ( n53485 , n46246 );
not ( n53486 , n53485 );
buf ( n53487 , n52514 );
not ( n53488 , n53487 );
or ( n53489 , n53486 , n53488 );
buf ( n53490 , n45747 );
not ( n53491 , n53490 );
buf ( n53492 , n53491 );
buf ( n53493 , n53492 );
not ( n53494 , n53493 );
buf ( n53495 , n42926 );
not ( n53496 , n53495 );
or ( n53497 , n53494 , n53496 );
buf ( n53498 , n49804 );
buf ( n53499 , n45747 );
nand ( n53500 , n53498 , n53499 );
buf ( n53501 , n53500 );
buf ( n53502 , n53501 );
nand ( n53503 , n53497 , n53502 );
buf ( n53504 , n53503 );
buf ( n53505 , n53504 );
buf ( n53506 , n46225 );
nand ( n53507 , n53505 , n53506 );
buf ( n53508 , n53507 );
buf ( n53509 , n53508 );
nand ( n53510 , n53489 , n53509 );
buf ( n53511 , n53510 );
buf ( n53512 , n53511 );
not ( n53513 , n42339 );
not ( n53514 , n52618 );
or ( n53515 , n53513 , n53514 );
buf ( n53516 , n42343 );
not ( n53517 , n53516 );
buf ( n53518 , n42437 );
not ( n53519 , n53518 );
or ( n53520 , n53517 , n53519 );
buf ( n53521 , n43446 );
buf ( n53522 , n46855 );
nand ( n53523 , n53521 , n53522 );
buf ( n53524 , n53523 );
buf ( n53525 , n53524 );
nand ( n53526 , n53520 , n53525 );
buf ( n53527 , n53526 );
buf ( n53528 , n53527 );
buf ( n53529 , n42378 );
nand ( n53530 , n53528 , n53529 );
buf ( n53531 , n53530 );
nand ( n53532 , n53515 , n53531 );
not ( n53533 , n53532 );
xor ( n53534 , n12447 , n12489 );
xor ( n53535 , n53534 , n12502 );
buf ( n53536 , n53535 );
buf ( n53537 , n53536 );
buf ( n53538 , n53537 );
buf ( n53539 , n53538 );
buf ( n53540 , n53539 );
not ( n53541 , n53540 );
buf ( n53542 , n38837 );
not ( n53543 , n53542 );
or ( n53544 , n53541 , n53543 );
buf ( n53545 , n36360 );
buf ( n53546 , n53539 );
not ( n53547 , n53546 );
buf ( n53548 , n53547 );
buf ( n53549 , n53548 );
nand ( n53550 , n53545 , n53549 );
buf ( n53551 , n53550 );
buf ( n53552 , n53551 );
nand ( n53553 , n53544 , n53552 );
buf ( n53554 , n53553 );
buf ( n53555 , n36444 );
buf ( n53556 , n52795 );
nand ( n53557 , n53555 , n53556 );
buf ( n53558 , n53557 );
nand ( n53559 , C1 , n53558 );
not ( n53560 , n53559 );
or ( n53561 , n53533 , n53560 );
or ( n53562 , n53532 , n53559 );
and ( n53563 , n52547 , n52570 );
not ( n53564 , n52547 );
and ( n53565 , n53564 , n52573 );
or ( n53566 , n53563 , n53565 );
not ( n53567 , n52601 );
and ( n53568 , n53566 , n53567 );
not ( n53569 , n53566 );
and ( n53570 , n53569 , n52601 );
nor ( n53571 , n53568 , n53570 );
nand ( n53572 , n53562 , n53571 );
nand ( n53573 , n53561 , n53572 );
buf ( n53574 , n53573 );
buf ( n53575 , n50128 );
not ( n53576 , n53575 );
buf ( n53577 , n25159 );
not ( n53578 , n53577 );
not ( n53579 , n42146 );
buf ( n53580 , n53579 );
not ( n53581 , n53580 );
or ( n53582 , n53578 , n53581 );
buf ( n53583 , n42146 );
buf ( n53584 , n52670 );
nand ( n53585 , n53583 , n53584 );
buf ( n53586 , n53585 );
buf ( n53587 , n53586 );
nand ( n53588 , n53582 , n53587 );
buf ( n53589 , n53588 );
buf ( n53590 , n53589 );
not ( n53591 , n53590 );
or ( n53592 , n53576 , n53591 );
buf ( n53593 , n52678 );
buf ( n53594 , n42564 );
nand ( n53595 , n53593 , n53594 );
buf ( n53596 , n53595 );
buf ( n53597 , n53596 );
nand ( n53598 , n53592 , n53597 );
buf ( n53599 , n53598 );
buf ( n53600 , n53599 );
buf ( n53601 , n13653 );
not ( n53602 , n53601 );
buf ( n53603 , n47031 );
not ( n53604 , n53603 );
or ( n53605 , n53602 , n53604 );
buf ( n53606 , n42468 );
buf ( n53607 , n43099 );
nand ( n53608 , n53606 , n53607 );
buf ( n53609 , n53608 );
buf ( n53610 , n53609 );
nand ( n53611 , n53605 , n53610 );
buf ( n53612 , n53611 );
buf ( n53613 , n53612 );
not ( n53614 , n53613 );
buf ( n53615 , n47014 );
not ( n53616 , n53615 );
or ( n53617 , n53614 , n53616 );
buf ( n53618 , n47019 );
not ( n53619 , n53618 );
buf ( n53620 , n52587 );
nand ( n53621 , n53619 , n53620 );
buf ( n53622 , n53621 );
buf ( n53623 , n53622 );
nand ( n53624 , n53617 , n53623 );
buf ( n53625 , n53624 );
buf ( n53626 , n53625 );
or ( n53627 , n53600 , n53626 );
not ( n53628 , n43931 );
buf ( n53629 , n53628 );
not ( n53630 , n53629 );
buf ( n53631 , n52724 );
not ( n53632 , n53631 );
buf ( n53633 , n47001 );
not ( n53634 , n53633 );
or ( n53635 , n53632 , n53634 );
buf ( n53636 , n29358 );
buf ( n53637 , n52725 );
nand ( n53638 , n53636 , n53637 );
buf ( n53639 , n53638 );
buf ( n53640 , n53639 );
nand ( n53641 , n53635 , n53640 );
buf ( n53642 , n53641 );
buf ( n53643 , n53642 );
not ( n53644 , n53643 );
or ( n53645 , n53630 , n53644 );
buf ( n53646 , n52731 );
buf ( n53647 , n43904 );
not ( n53648 , n53647 );
buf ( n53649 , n53648 );
buf ( n53650 , n53649 );
nand ( n53651 , n53646 , n53650 );
buf ( n53652 , n53651 );
buf ( n53653 , n53652 );
nand ( n53654 , n53645 , n53653 );
buf ( n53655 , n53654 );
buf ( n53656 , n53655 );
nand ( n53657 , n53627 , n53656 );
buf ( n53658 , n53657 );
buf ( n53659 , n53658 );
buf ( n53660 , n53625 );
buf ( n53661 , n53599 );
nand ( n53662 , n53660 , n53661 );
buf ( n53663 , n53662 );
buf ( n53664 , n53663 );
nand ( n53665 , n53659 , n53664 );
buf ( n53666 , n53665 );
buf ( n53667 , n53666 );
buf ( n53668 , n42847 );
not ( n53669 , n53668 );
buf ( n53670 , n41925 );
not ( n53671 , n53670 );
or ( n53672 , n53669 , n53671 );
nand ( n53673 , n41895 , n46691 );
buf ( n53674 , n53673 );
nand ( n53675 , n53672 , n53674 );
buf ( n53676 , n53675 );
buf ( n53677 , n53676 );
not ( n53678 , n53677 );
buf ( n53679 , n37872 );
not ( n53680 , n53679 );
or ( n53681 , n53678 , n53680 );
buf ( n53682 , n52332 );
not ( n53683 , n53682 );
buf ( n53684 , n45617 );
nand ( n53685 , n53683 , n53684 );
buf ( n53686 , n53685 );
buf ( n53687 , n53686 );
nand ( n53688 , n53681 , n53687 );
buf ( n53689 , n53688 );
buf ( n53690 , n53689 );
xor ( n53691 , n53667 , n53690 );
buf ( n53692 , n50060 );
not ( n53693 , n53692 );
buf ( n53694 , n39478 );
not ( n53695 , n53694 );
or ( n53696 , n53693 , n53695 );
buf ( n53697 , n33076 );
buf ( n53698 , n50067 );
nand ( n53699 , n53697 , n53698 );
buf ( n53700 , n53699 );
buf ( n53701 , n53700 );
nand ( n53702 , n53696 , n53701 );
buf ( n53703 , n53702 );
buf ( n53704 , n53703 );
not ( n53705 , n53704 );
buf ( n53706 , n42521 );
not ( n53707 , n53706 );
or ( n53708 , n53705 , n53707 );
buf ( n53709 , n52761 );
buf ( n53710 , n42530 );
nand ( n53711 , n53709 , n53710 );
buf ( n53712 , n53711 );
buf ( n53713 , n53712 );
nand ( n53714 , n53708 , n53713 );
buf ( n53715 , n53714 );
buf ( n53716 , n53715 );
and ( n53717 , n53691 , n53716 );
and ( n53718 , n53667 , n53690 );
or ( n53719 , n53717 , n53718 );
buf ( n53720 , n53719 );
buf ( n53721 , n53720 );
xor ( n53722 , n53574 , n53721 );
buf ( n53723 , n42252 );
not ( n53724 , n53723 );
buf ( n53725 , n42266 );
not ( n53726 , n53725 );
buf ( n53727 , n47626 );
not ( n53728 , n53727 );
or ( n53729 , n53726 , n53728 );
buf ( n53730 , n37783 );
buf ( n53731 , n42263 );
nand ( n53732 , n53730 , n53731 );
buf ( n53733 , n53732 );
buf ( n53734 , n53733 );
nand ( n53735 , n53729 , n53734 );
buf ( n53736 , n53735 );
buf ( n53737 , n53736 );
not ( n53738 , n53737 );
or ( n53739 , n53724 , n53738 );
buf ( n53740 , n52653 );
buf ( n53741 , n42315 );
nand ( n53742 , n53740 , n53741 );
buf ( n53743 , n53742 );
buf ( n53744 , n53743 );
nand ( n53745 , n53739 , n53744 );
buf ( n53746 , n53745 );
buf ( n53747 , n53746 );
and ( n53748 , n53722 , n53747 );
and ( n53749 , n53574 , n53721 );
or ( n53750 , n53748 , n53749 );
buf ( n53751 , n53750 );
buf ( n53752 , n53751 );
xor ( n53753 , n53512 , n53752 );
buf ( n53754 , n46912 );
not ( n53755 , n53754 );
buf ( n53756 , n53093 );
not ( n53757 , n53756 );
or ( n53758 , n53755 , n53757 );
buf ( n53759 , n51622 );
not ( n53760 , n53759 );
buf ( n53761 , n38098 );
not ( n53762 , n53761 );
or ( n53763 , n53760 , n53762 );
buf ( n53764 , n38098 );
not ( n53765 , n53764 );
buf ( n53766 , n46890 );
nand ( n53767 , n53765 , n53766 );
buf ( n53768 , n53767 );
buf ( n53769 , n53768 );
nand ( n53770 , n53763 , n53769 );
buf ( n53771 , n53770 );
buf ( n53772 , n53771 );
buf ( n53773 , n47331 );
nand ( n53774 , n53772 , n53773 );
buf ( n53775 , n53774 );
buf ( n53776 , n53775 );
nand ( n53777 , n53758 , n53776 );
buf ( n53778 , n53777 );
buf ( n53779 , n53778 );
and ( n53780 , n53753 , n53779 );
and ( n53781 , n53512 , n53752 );
or ( n53782 , n53780 , n53781 );
buf ( n53783 , n53782 );
buf ( n53784 , n53783 );
and ( n53785 , n53484 , n53784 );
and ( n53786 , n53480 , n53483 );
or ( n53787 , n53785 , n53786 );
buf ( n53788 , n53787 );
buf ( n53789 , n53788 );
xor ( n53790 , n53477 , n53789 );
xor ( n53791 , n52901 , n52926 );
xor ( n53792 , n53791 , n52931 );
buf ( n53793 , n53792 );
buf ( n53794 , n53793 );
xor ( n53795 , n52608 , n52628 );
xor ( n53796 , n53795 , n52632 );
not ( n53797 , n52970 );
not ( n53798 , n38057 );
and ( n53799 , n53797 , n53798 );
buf ( n53800 , n46117 );
not ( n53801 , n53800 );
buf ( n53802 , n38068 );
not ( n53803 , n53802 );
or ( n53804 , n53801 , n53803 );
buf ( n53805 , n43400 );
buf ( n53806 , n46126 );
nand ( n53807 , n53805 , n53806 );
buf ( n53808 , n53807 );
buf ( n53809 , n53808 );
nand ( n53810 , n53804 , n53809 );
buf ( n53811 , n53810 );
not ( n53812 , n53811 );
buf ( n53813 , n38121 );
buf ( n53814 , n38115 );
buf ( n53815 , n38051 );
nand ( n53816 , n53813 , n53814 , n53815 );
buf ( n53817 , n53816 );
nor ( n53818 , n53812 , n53817 );
nor ( n53819 , n53799 , n53818 );
buf ( n53820 , n53819 );
not ( n53821 , n53820 );
buf ( n53822 , n53821 );
not ( n53823 , n53822 );
buf ( n53824 , n52685 );
buf ( n53825 , n52738 );
xor ( n53826 , n53824 , n53825 );
buf ( n53827 , n52710 );
xnor ( n53828 , n53826 , n53827 );
buf ( n53829 , n53828 );
buf ( n53830 , n53829 );
not ( n53831 , n53830 );
buf ( n53832 , n53831 );
not ( n53833 , n53832 );
or ( n53834 , n53823 , n53833 );
buf ( n53835 , n53829 );
not ( n53836 , n53835 );
buf ( n53837 , n53819 );
not ( n53838 , n53837 );
or ( n53839 , n53836 , n53838 );
not ( n53840 , n53270 );
not ( n53841 , n41644 );
and ( n53842 , n53840 , n53841 );
buf ( n53843 , n48390 );
not ( n53844 , n53843 );
buf ( n53845 , n44025 );
not ( n53846 , n53845 );
or ( n53847 , n53844 , n53846 );
buf ( n53848 , n28306 );
buf ( n53849 , n41660 );
nand ( n53850 , n53848 , n53849 );
buf ( n53851 , n53850 );
buf ( n53852 , n53851 );
nand ( n53853 , n53847 , n53852 );
buf ( n53854 , n53853 );
and ( n53855 , n53854 , n50982 );
nor ( n53856 , n53842 , n53855 );
not ( n53857 , n53856 );
not ( n53858 , n53857 );
buf ( n53859 , n37327 );
buf ( n53860 , n53859 );
buf ( n53861 , n53860 );
and ( n53862 , n53861 , n43966 );
not ( n53863 , n53861 );
and ( n53864 , n53863 , n41993 );
or ( n53865 , n53862 , n53864 );
not ( n53866 , n53865 );
not ( n53867 , n37397 );
or ( n53868 , n53866 , n53867 );
buf ( n53869 , n42132 );
not ( n53870 , n53869 );
buf ( n53871 , n53245 );
nand ( n53872 , n53870 , n53871 );
buf ( n53873 , n53872 );
nand ( n53874 , n53868 , n53873 );
not ( n53875 , n53874 );
or ( n53876 , n53858 , n53875 );
buf ( n53877 , n53856 );
not ( n53878 , n53877 );
buf ( n53879 , n53874 );
not ( n53880 , n53879 );
buf ( n53881 , n53880 );
buf ( n53882 , n53881 );
not ( n53883 , n53882 );
or ( n53884 , n53878 , n53883 );
not ( n53885 , n42378 );
buf ( n53886 , n42343 );
not ( n53887 , n53886 );
buf ( n53888 , n39656 );
not ( n53889 , n53888 );
or ( n53890 , n53887 , n53889 );
buf ( n53891 , n39653 );
buf ( n53892 , n46855 );
nand ( n53893 , n53891 , n53892 );
buf ( n53894 , n53893 );
buf ( n53895 , n53894 );
nand ( n53896 , n53890 , n53895 );
buf ( n53897 , n53896 );
not ( n53898 , n53897 );
or ( n53899 , n53885 , n53898 );
buf ( n53900 , n53527 );
buf ( n53901 , n42339 );
nand ( n53902 , n53900 , n53901 );
buf ( n53903 , n53902 );
nand ( n53904 , n53899 , n53903 );
buf ( n53905 , n53904 );
nand ( n53906 , n53884 , n53905 );
buf ( n53907 , n53906 );
nand ( n53908 , n53876 , n53907 );
buf ( n53909 , n53908 );
nand ( n53910 , n53839 , n53909 );
buf ( n53911 , n53910 );
nand ( n53912 , n53834 , n53911 );
xor ( n53913 , n53796 , n53912 );
not ( n53914 , n46225 );
buf ( n53915 , n53492 );
not ( n53916 , n53915 );
buf ( n53917 , n39406 );
not ( n53918 , n53917 );
or ( n53919 , n53916 , n53918 );
not ( n53920 , n38218 );
not ( n53921 , n45753 );
nand ( n53922 , n53920 , n53921 );
buf ( n53923 , n53922 );
nand ( n53924 , n53919 , n53923 );
buf ( n53925 , n53924 );
not ( n53926 , n53925 );
or ( n53927 , n53914 , n53926 );
buf ( n53928 , n53504 );
buf ( n53929 , n46246 );
nand ( n53930 , n53928 , n53929 );
buf ( n53931 , n53930 );
nand ( n53932 , n53927 , n53931 );
and ( n53933 , n53913 , n53932 );
and ( n53934 , n53796 , n53912 );
or ( n53935 , n53933 , n53934 );
buf ( n53936 , n53935 );
xor ( n53937 , n53794 , n53936 );
xor ( n53938 , n53255 , n53279 );
xor ( n53939 , n53938 , n53302 );
buf ( n53940 , n53939 );
buf ( n53941 , n53940 );
buf ( n53942 , n39803 );
not ( n53943 , n53942 );
buf ( n53944 , n52094 );
not ( n53945 , n53944 );
buf ( n53946 , n53945 );
not ( n53947 , n53946 );
xor ( n53948 , n39726 , n53947 );
buf ( n53949 , n53948 );
not ( n53950 , n53949 );
or ( n53951 , n53943 , n53950 );
nand ( n53952 , n53207 , n43982 );
buf ( n53953 , n53952 );
nand ( n53954 , n53951 , n53953 );
buf ( n53955 , n53954 );
buf ( n53956 , n53955 );
or ( n53957 , n53941 , n53956 );
buf ( n53958 , n53957 );
buf ( n53959 , n42865 );
not ( n53960 , n53959 );
buf ( n53961 , n41977 );
not ( n53962 , n53961 );
or ( n53963 , n53960 , n53962 );
buf ( n53964 , n51901 );
buf ( n53965 , n42862 );
nand ( n53966 , n53964 , n53965 );
buf ( n53967 , n53966 );
buf ( n53968 , n53967 );
nand ( n53969 , n53963 , n53968 );
buf ( n53970 , n53969 );
buf ( n53971 , n53970 );
not ( n53972 , n53971 );
buf ( n53973 , n41966 );
not ( n53974 , n53973 );
or ( n53975 , n53972 , n53974 );
buf ( n53976 , n53292 );
buf ( n53977 , n37446 );
nand ( n53978 , n53976 , n53977 );
buf ( n53979 , n53978 );
buf ( n53980 , n53979 );
nand ( n53981 , n53975 , n53980 );
buf ( n53982 , n53981 );
buf ( n53983 , n53982 );
not ( n53984 , n53983 );
and ( n53985 , n44949 , n41947 );
not ( n53986 , n44949 );
and ( n53987 , n53986 , n44381 );
or ( n53988 , n53985 , n53987 );
not ( n53989 , n53988 );
not ( n53990 , n37872 );
or ( n53991 , n53989 , n53990 );
buf ( n53992 , n45617 );
buf ( n53993 , n53676 );
nand ( n53994 , n53992 , n53993 );
buf ( n53995 , n53994 );
nand ( n53996 , n53991 , n53995 );
buf ( n53997 , n53996 );
not ( n53998 , n53997 );
or ( n53999 , n53984 , n53998 );
buf ( n54000 , n53982 );
buf ( n54001 , n53996 );
or ( n54002 , n54000 , n54001 );
buf ( n54003 , n42049 );
not ( n54004 , n54003 );
buf ( n54005 , n50599 );
not ( n54006 , n54005 );
or ( n54007 , n54004 , n54006 );
buf ( n54008 , n50591 );
buf ( n54009 , n42052 );
nand ( n54010 , n54008 , n54009 );
buf ( n54011 , n54010 );
buf ( n54012 , n54011 );
nand ( n54013 , n54007 , n54012 );
buf ( n54014 , n54013 );
buf ( n54015 , n54014 );
not ( n54016 , n54015 );
buf ( n54017 , n50608 );
not ( n54018 , n54017 );
or ( n54019 , n54016 , n54018 );
buf ( n54020 , n52558 );
buf ( n54021 , n46633 );
nand ( n54022 , n54020 , n54021 );
buf ( n54023 , n54022 );
buf ( n54024 , n54023 );
nand ( n54025 , n54019 , n54024 );
buf ( n54026 , n54025 );
buf ( n54027 , n54026 );
not ( n54028 , n54027 );
buf ( n54029 , n41736 );
not ( n54030 , n54029 );
buf ( n54031 , n42471 );
not ( n54032 , n54031 );
or ( n54033 , n54030 , n54032 );
buf ( n54034 , n42468 );
buf ( n54035 , n41733 );
nand ( n54036 , n54034 , n54035 );
buf ( n54037 , n54036 );
buf ( n54038 , n54037 );
nand ( n54039 , n54033 , n54038 );
buf ( n54040 , n54039 );
buf ( n54041 , n54040 );
not ( n54042 , n54041 );
buf ( n54043 , n47050 );
not ( n54044 , n54043 );
or ( n54045 , n54042 , n54044 );
buf ( n54046 , n53612 );
buf ( n54047 , n50104 );
nand ( n54048 , n54046 , n54047 );
buf ( n54049 , n54048 );
buf ( n54050 , n54049 );
nand ( n54051 , n54045 , n54050 );
buf ( n54052 , n54051 );
buf ( n54053 , n54052 );
not ( n54054 , n54053 );
or ( n54055 , n54028 , n54054 );
buf ( n54056 , n54052 );
buf ( n54057 , n54026 );
or ( n54058 , n54056 , n54057 );
buf ( n54059 , n53649 );
not ( n54060 , n54059 );
buf ( n54061 , n53642 );
not ( n54062 , n54061 );
or ( n54063 , n54060 , n54062 );
not ( n54064 , n52725 );
not ( n54065 , n47063 );
or ( n54066 , n54064 , n54065 );
buf ( n54067 , n42559 );
not ( n54068 , n54067 );
nand ( n54069 , n54068 , n47072 );
nand ( n54070 , n54066 , n54069 );
nand ( n54071 , n54070 , n43938 );
buf ( n54072 , n54071 );
nand ( n54073 , n54063 , n54072 );
buf ( n54074 , n54073 );
buf ( n54075 , n54074 );
nand ( n54076 , n54058 , n54075 );
buf ( n54077 , n54076 );
buf ( n54078 , n54077 );
nand ( n54079 , n54055 , n54078 );
buf ( n54080 , n54079 );
buf ( n54081 , n54080 );
nand ( n54082 , n54002 , n54081 );
buf ( n54083 , n54082 );
buf ( n54084 , n54083 );
nand ( n54085 , n53999 , n54084 );
buf ( n54086 , n54085 );
and ( n54087 , n53958 , n54086 );
buf ( n54088 , n53955 );
buf ( n54089 , n53940 );
and ( n54090 , n54088 , n54089 );
buf ( n54091 , n54090 );
nor ( n54092 , n54087 , n54091 );
buf ( n54093 , n54092 );
not ( n54094 , n54093 );
not ( n54095 , n52985 );
not ( n54096 , n53011 );
or ( n54097 , n54095 , n54096 );
buf ( n54098 , n52988 );
buf ( n54099 , n53010 );
nand ( n54100 , n54098 , n54099 );
buf ( n54101 , n54100 );
nand ( n54102 , n54097 , n54101 );
buf ( n54103 , n53017 );
not ( n54104 , n54103 );
buf ( n54105 , n54104 );
and ( n54106 , n54102 , n54105 );
not ( n54107 , n54102 );
and ( n54108 , n54107 , n53017 );
nor ( n54109 , n54106 , n54108 );
buf ( n54110 , n54109 );
not ( n54111 , n54110 );
buf ( n54112 , n54111 );
buf ( n54113 , n54112 );
nand ( n54114 , n54094 , n54113 );
buf ( n54115 , n54114 );
not ( n54116 , n54109 );
not ( n54117 , n54092 );
or ( n54118 , n54116 , n54117 );
buf ( n54119 , n52573 );
buf ( n54120 , n53589 );
not ( n54121 , n54120 );
buf ( n54122 , n42563 );
nor ( n54123 , n54121 , n54122 );
buf ( n54124 , n54123 );
not ( n54125 , n54124 );
buf ( n54126 , n25159 );
buf ( n54127 , n43362 );
and ( n54128 , n54126 , n54127 );
not ( n54129 , n54126 );
buf ( n54130 , n50624 );
and ( n54131 , n54129 , n54130 );
nor ( n54132 , n54128 , n54131 );
buf ( n54133 , n54132 );
nor ( n54134 , n42625 , n54133 );
nand ( n54135 , n611 , n613 );
nand ( n54136 , n610 , n614 );
and ( n54137 , n54135 , n54136 );
not ( n54138 , n54135 );
not ( n54139 , n54136 );
and ( n54140 , n54138 , n54139 );
nor ( n54141 , n54137 , n54140 );
nand ( n54142 , n608 , n616 );
and ( n54143 , n54141 , n54142 );
nor ( n54144 , n54141 , n54142 );
nor ( n54145 , n54143 , n54144 );
nand ( n54146 , n609 , n615 );
nand ( n54147 , n610 , n615 );
not ( n54148 , n54147 );
nand ( n54149 , n612 , n54148 );
nand ( n54150 , n612 , n613 );
and ( n54151 , n54149 , n54150 );
xor ( n54152 , n54146 , n54151 );
nand ( n54153 , n611 , n614 );
nand ( n54154 , n609 , n616 );
xor ( n54155 , n54153 , n54154 );
nand ( n54156 , n608 , n617 );
and ( n54157 , n54155 , n54156 );
and ( n54158 , n54153 , n54154 );
or ( n54159 , n54157 , n54158 );
xor ( n54160 , n54152 , n54159 );
xor ( n54161 , n54145 , n54160 );
nand ( n54162 , n612 , n614 );
nand ( n54163 , n611 , n615 );
xor ( n54164 , n54162 , n54163 );
nand ( n54165 , n609 , n617 );
and ( n54166 , n54164 , n54165 );
and ( n54167 , n54162 , n54163 );
or ( n54168 , n54166 , n54167 );
and ( n54169 , n54150 , n612 );
nor ( n54170 , C0 , n54169 );
and ( n54171 , n54170 , n54148 );
not ( n54172 , n54170 );
and ( n54173 , n54172 , n54147 );
nor ( n54174 , n54171 , n54173 );
xor ( n54175 , n54168 , n54174 );
xor ( n54176 , n54153 , n54154 );
xor ( n54177 , n54176 , n54156 );
and ( n54178 , n54175 , n54177 );
and ( n54179 , n54168 , n54174 );
or ( n54180 , n54178 , n54179 );
and ( n54181 , n54161 , n54180 );
and ( n54182 , n54145 , n54160 );
or ( n54183 , n54181 , n54182 );
nand ( n54184 , n610 , n613 );
nand ( n54185 , n608 , n615 );
xor ( n54186 , n54184 , n54185 );
not ( n54187 , n54139 );
not ( n54188 , n54135 );
not ( n54189 , n54188 );
or ( n54190 , n54187 , n54189 );
not ( n54191 , n54136 );
not ( n54192 , n54135 );
or ( n54193 , n54191 , n54192 );
not ( n54194 , n54142 );
nand ( n54195 , n54193 , n54194 );
nand ( n54196 , n54190 , n54195 );
not ( n54197 , n54196 );
xor ( n54198 , n54186 , n54197 );
nand ( n54199 , n609 , n614 );
nand ( n54200 , n611 , n612 );
xor ( n54201 , n54199 , n54200 );
not ( n54202 , n611 );
xor ( n54203 , n54201 , n54202 );
xor ( n54204 , n54146 , n54151 );
and ( n54205 , n54204 , n54159 );
and ( n54206 , n54146 , n54151 );
or ( n54207 , n54205 , n54206 );
xor ( n54208 , n54203 , n54207 );
xor ( n54209 , n54198 , n54208 );
nand ( n54210 , n54183 , n54209 );
xor ( n54211 , n54184 , n54185 );
xor ( n54212 , n54211 , n54197 );
and ( n54213 , n54203 , n54212 );
xor ( n54214 , n54184 , n54185 );
xor ( n54215 , n54214 , n54197 );
and ( n54216 , n54207 , n54215 );
and ( n54217 , n54203 , n54207 );
or ( n54218 , n54213 , n54216 , n54217 );
nand ( n54219 , n609 , n613 );
nand ( n54220 , n610 , n612 );
xor ( n54221 , n54219 , n54220 );
nand ( n54222 , n608 , n614 );
xor ( n54223 , n54221 , n54222 );
xor ( n54224 , n54199 , n54200 );
and ( n54225 , n54224 , n54202 );
and ( n54226 , n54199 , n54200 );
or ( n54227 , n54225 , n54226 );
xor ( n54228 , n54184 , n54185 );
and ( n54229 , n54228 , n54197 );
and ( n54230 , n54184 , n54185 );
or ( n54231 , n54229 , n54230 );
xor ( n54232 , n54227 , n54231 );
xor ( n54233 , n54223 , n54232 );
nand ( n54234 , n54218 , n54233 );
and ( n54235 , n54210 , n54234 );
xor ( n54236 , n54219 , n54220 );
and ( n54237 , n54236 , n54222 );
and ( n54238 , n54219 , n54220 );
or ( n54239 , n54237 , n54238 );
nand ( n54240 , n609 , n612 );
xor ( n54241 , n54239 , n54240 );
nand ( n54242 , n608 , n613 );
nand ( n54243 , n610 , n611 );
xor ( n54244 , n54242 , n54243 );
not ( n54245 , n610 );
xor ( n54246 , n54244 , n54245 );
and ( n54247 , n54241 , n54246 );
and ( n54248 , n54239 , n54240 );
or ( n54249 , n54247 , n54248 );
nand ( n54250 , n609 , n611 );
nand ( n54251 , n608 , n612 );
xor ( n54252 , n54250 , n54251 );
xor ( n54253 , n54242 , n54243 );
and ( n54254 , n54253 , n54245 );
and ( n54255 , n54242 , n54243 );
or ( n54256 , n54254 , n54255 );
xor ( n54257 , n54252 , n54256 );
nand ( n54258 , n54249 , n54257 );
not ( n54259 , n54258 );
xor ( n54260 , n54250 , n54251 );
and ( n54261 , n54260 , n54256 );
and ( n54262 , n54250 , n54251 );
or ( n54263 , n54261 , n54262 );
nand ( n54264 , n608 , n611 );
nand ( n54265 , n609 , n610 );
xor ( n54266 , n54264 , n54265 );
not ( n54267 , n609 );
xor ( n54268 , n54266 , n54267 );
nand ( n54269 , n54263 , n54268 );
xor ( n54270 , n54264 , n54265 );
and ( n54271 , n54270 , n54267 );
and ( n54272 , n54264 , n54265 );
or ( n54273 , n54271 , n54272 );
nand ( n54274 , n608 , n610 );
nand ( n54275 , n54273 , n54274 );
nand ( n54276 , n54269 , n54275 );
nor ( n54277 , n54259 , n54276 );
xor ( n54278 , n54219 , n54220 );
xor ( n54279 , n54278 , n54222 );
and ( n54280 , n54227 , n54279 );
xor ( n54281 , n54219 , n54220 );
xor ( n54282 , n54281 , n54222 );
and ( n54283 , n54231 , n54282 );
and ( n54284 , n54227 , n54231 );
or ( n54285 , n54280 , n54283 , n54284 );
xor ( n54286 , n54239 , n54240 );
xor ( n54287 , n54286 , n54246 );
nand ( n54288 , n54285 , n54287 );
and ( n54289 , n54235 , n54277 , n54288 );
not ( n54290 , n54289 );
nand ( n54291 , n610 , n616 );
nand ( n54292 , n608 , n618 );
xor ( n54293 , n54291 , n54292 );
nand ( n54294 , n612 , n615 );
nand ( n54295 , n610 , n617 );
xor ( n54296 , n54294 , n54295 );
nand ( n54297 , n609 , n618 );
and ( n54298 , n54296 , n54297 );
and ( n54299 , n54294 , n54295 );
or ( n54300 , n54298 , n54299 );
xor ( n54301 , n54293 , n54300 );
and ( n54302 , n608 , n619 );
not ( n54303 , n54302 );
nand ( n54304 , n609 , n619 );
not ( n54305 , n54304 );
nand ( n54306 , n611 , n617 );
not ( n54307 , n54306 );
or ( n54308 , n54305 , n54307 );
nand ( n54309 , n608 , n620 );
not ( n54310 , n54309 );
nand ( n54311 , n54308 , n54310 );
not ( n54312 , n54304 );
not ( n54313 , n54306 );
nand ( n54314 , n54312 , n54313 );
nand ( n54315 , n54311 , n54314 );
not ( n54316 , n54315 );
or ( n54317 , n54303 , n54316 );
or ( n54318 , n54315 , n54302 );
nand ( n54319 , n612 , n616 );
nand ( n54320 , n613 , n615 );
xor ( n54321 , n54319 , n54320 );
nand ( n54322 , n610 , n618 );
and ( n54323 , n54321 , n54322 );
and ( n54324 , n54319 , n54320 );
nor ( n54325 , n54323 , n54324 );
nand ( n54326 , n54318 , n54325 );
nand ( n54327 , n54317 , n54326 );
nand ( n54328 , n613 , n614 );
and ( n54329 , n611 , n616 );
nand ( n54330 , n613 , n54329 );
nand ( n54331 , n54328 , n54330 );
not ( n54332 , n54331 );
xor ( n54333 , n54162 , n54163 );
xor ( n54334 , n54333 , n54165 );
not ( n54335 , n54334 );
or ( n54336 , n54332 , n54335 );
or ( n54337 , n54334 , n54331 );
nand ( n54338 , n54336 , n54337 );
xnor ( n54339 , n54327 , n54338 );
and ( n54340 , n54328 , n613 );
nor ( n54341 , C0 , n54340 );
xor ( n54342 , n54341 , n54329 );
xor ( n54343 , n54294 , n54295 );
xor ( n54344 , n54343 , n54297 );
xor ( n54345 , n54342 , n54344 );
xor ( n54346 , n54302 , n54325 );
xnor ( n54347 , n54346 , n54315 );
and ( n54348 , n54345 , n54347 );
and ( n54349 , n54342 , n54344 );
or ( n54350 , n54348 , n54349 );
xor ( n54351 , n54339 , n54350 );
xor ( n54352 , n54301 , n54351 );
nand ( n54353 , n611 , n618 );
nand ( n54354 , n608 , n621 );
xor ( n54355 , n54353 , n54354 );
nand ( n54356 , n613 , n616 );
and ( n54357 , n54355 , n54356 );
and ( n54358 , n54353 , n54354 );
or ( n54359 , n54357 , n54358 );
nand ( n54360 , n614 , n615 );
nand ( n54361 , n612 , n617 );
xor ( n54362 , n54360 , n54361 );
not ( n54363 , n614 );
and ( n54364 , n54362 , n54363 );
and ( n54365 , n54360 , n54361 );
or ( n54366 , n54364 , n54365 );
xor ( n54367 , n54359 , n54366 );
xor ( n54368 , n54319 , n54320 );
xor ( n54369 , n54368 , n54322 );
and ( n54370 , n54367 , n54369 );
and ( n54371 , n54359 , n54366 );
or ( n54372 , n54370 , n54371 );
xor ( n54373 , n54342 , n54344 );
xor ( n54374 , n54373 , n54347 );
xor ( n54375 , n54372 , n54374 );
xor ( n54376 , n54360 , n54361 );
xor ( n54377 , n54376 , n54363 );
not ( n54378 , n54377 );
nand ( n54379 , n612 , n618 );
nand ( n54380 , n610 , n620 );
xor ( n54381 , n54379 , n54380 );
nand ( n54382 , n609 , n621 );
and ( n54383 , n54381 , n54382 );
and ( n54384 , n54379 , n54380 );
or ( n54385 , n54383 , n54384 );
not ( n54386 , n54385 );
or ( n54387 , n54378 , n54386 );
not ( n54388 , n54385 );
not ( n54389 , n54388 );
not ( n54390 , n54377 );
not ( n54391 , n54390 );
or ( n54392 , n54389 , n54391 );
xor ( n54393 , n54353 , n54354 );
xor ( n54394 , n54393 , n54356 );
nand ( n54395 , n54392 , n54394 );
nand ( n54396 , n54387 , n54395 );
not ( n54397 , n54396 );
nand ( n54398 , n610 , n619 );
nand ( n54399 , n609 , n620 );
xor ( n54400 , n54398 , n54399 );
nand ( n54401 , n614 , n616 );
nand ( n54402 , n611 , n619 );
xor ( n54403 , n54401 , n54402 );
nand ( n54404 , n613 , n617 );
and ( n54405 , n54403 , n54404 );
and ( n54406 , n54401 , n54402 );
or ( n54407 , n54405 , n54406 );
and ( n54408 , n54400 , n54407 );
and ( n54409 , n54398 , n54399 );
or ( n54410 , n54408 , n54409 );
not ( n54411 , n54410 );
not ( n54412 , n54304 );
not ( n54413 , n54313 );
or ( n54414 , n54412 , n54413 );
or ( n54415 , n54304 , n54313 );
nand ( n54416 , n54414 , n54415 );
not ( n54417 , n54416 );
not ( n54418 , n54309 );
and ( n54419 , n54417 , n54418 );
and ( n54420 , n54416 , n54309 );
nor ( n54421 , n54419 , n54420 );
not ( n54422 , n54421 );
nand ( n54423 , n54411 , n54422 );
not ( n54424 , n54423 );
or ( n54425 , n54397 , n54424 );
nand ( n54426 , n54410 , n54421 );
nand ( n54427 , n54425 , n54426 );
and ( n54428 , n54375 , n54427 );
and ( n54429 , n54372 , n54374 );
or ( n54430 , n54428 , n54429 );
nand ( n54431 , n54352 , n54430 );
xor ( n54432 , n54291 , n54292 );
xor ( n54433 , n54432 , n54300 );
and ( n54434 , n54339 , n54433 );
xor ( n54435 , n54291 , n54292 );
xor ( n54436 , n54435 , n54300 );
and ( n54437 , n54350 , n54436 );
and ( n54438 , n54339 , n54350 );
or ( n54439 , n54434 , n54437 , n54438 );
xor ( n54440 , n54168 , n54174 );
xor ( n54441 , n54440 , n54177 );
xor ( n54442 , n54291 , n54292 );
and ( n54443 , n54442 , n54300 );
and ( n54444 , n54291 , n54292 );
or ( n54445 , n54443 , n54444 );
not ( n54446 , n54331 );
nand ( n54447 , n54446 , n54334 );
not ( n54448 , n54447 );
not ( n54449 , n54327 );
or ( n54450 , n54448 , n54449 );
not ( n54451 , n54334 );
nand ( n54452 , n54451 , n54331 );
nand ( n54453 , n54450 , n54452 );
not ( n54454 , n54453 );
xor ( n54455 , n54445 , n54454 );
xor ( n54456 , n54441 , n54455 );
nand ( n54457 , n54439 , n54456 );
and ( n54458 , n54431 , n54457 );
xor ( n54459 , n54168 , n54174 );
xor ( n54460 , n54459 , n54177 );
and ( n54461 , n54445 , n54460 );
xor ( n54462 , n54168 , n54174 );
xor ( n54463 , n54462 , n54177 );
and ( n54464 , n54454 , n54463 );
and ( n54465 , n54445 , n54454 );
or ( n54466 , n54461 , n54464 , n54465 );
xor ( n54467 , n54145 , n54160 );
xor ( n54468 , n54467 , n54180 );
nand ( n54469 , n54466 , n54468 );
and ( n54470 , n54458 , n54469 );
not ( n54471 , n54470 );
not ( n54472 , n54396 );
not ( n54473 , n54410 );
not ( n54474 , n54422 );
or ( n54475 , n54473 , n54474 );
nand ( n54476 , n54411 , n54421 );
nand ( n54477 , n54475 , n54476 );
nand ( n54478 , n54472 , n54477 );
nand ( n54479 , n54410 , n54396 , n54421 );
nand ( n54480 , n54411 , n54396 , n54422 );
nand ( n54481 , n54478 , n54479 , n54480 );
xor ( n54482 , n54359 , n54366 );
xor ( n54483 , n54482 , n54369 );
and ( n54484 , n54481 , n54483 );
xor ( n54485 , n54398 , n54399 );
xor ( n54486 , n54485 , n54407 );
nand ( n54487 , n608 , n622 );
nand ( n54488 , n615 , n616 );
xor ( n54489 , n54487 , n54488 );
nand ( n54490 , n609 , n622 );
nand ( n54491 , n608 , n623 );
xor ( n54492 , n54490 , n54491 );
nand ( n54493 , n613 , n618 );
and ( n54494 , n54492 , n54493 );
and ( n54495 , n54490 , n54491 );
or ( n54496 , n54494 , n54495 );
and ( n54497 , n54489 , n54496 );
and ( n54498 , n54487 , n54488 );
or ( n54499 , n54497 , n54498 );
xor ( n54500 , n54486 , n54499 );
nand ( n54501 , n614 , n617 );
nand ( n54502 , n611 , n620 );
xor ( n54503 , n54501 , n54502 );
nand ( n54504 , n612 , n619 );
and ( n54505 , n54503 , n54504 );
and ( n54506 , n54501 , n54502 );
or ( n54507 , n54505 , n54506 );
xor ( n54508 , n54379 , n54380 );
xor ( n54509 , n54508 , n54382 );
xor ( n54510 , n54507 , n54509 );
xor ( n54511 , n54401 , n54402 );
xor ( n54512 , n54511 , n54404 );
and ( n54513 , n54510 , n54512 );
and ( n54514 , n54507 , n54509 );
or ( n54515 , n54513 , n54514 );
and ( n54516 , n54500 , n54515 );
and ( n54517 , n54486 , n54499 );
or ( n54518 , n54516 , n54517 );
xor ( n54519 , n54359 , n54366 );
xor ( n54520 , n54519 , n54369 );
and ( n54521 , n54518 , n54520 );
and ( n54522 , n54481 , n54518 );
or ( n54523 , n54484 , n54521 , n54522 );
xor ( n54524 , n54372 , n54374 );
xor ( n54525 , n54524 , n54427 );
nand ( n54526 , n54523 , n54525 );
xor ( n54527 , n54359 , n54366 );
xor ( n54528 , n54527 , n54369 );
xor ( n54529 , n54481 , n54518 );
xor ( n54530 , n54528 , n54529 );
and ( n54531 , n54390 , n54394 , n54388 );
and ( n54532 , n54377 , n54385 , n54394 );
nor ( n54533 , n54531 , n54532 );
nor ( n54534 , n54394 , n54385 );
and ( n54535 , n54534 , n54377 );
nor ( n54536 , n54377 , n54388 , n54394 );
nor ( n54537 , n54535 , n54536 );
nand ( n54538 , n54533 , n54537 );
nand ( n54539 , n610 , n621 );
nand ( n54540 , n615 , n617 , n614 , n618 );
xor ( n54541 , n54539 , n54540 );
not ( n54542 , n616 );
nand ( n54543 , n54542 , n615 );
and ( n54544 , n54541 , n54543 );
and ( n54545 , n54539 , n54540 );
or ( n54546 , n54544 , n54545 );
xor ( n54547 , n54487 , n54488 );
xor ( n54548 , n54547 , n54496 );
xor ( n54549 , n54546 , n54548 );
nand ( n54550 , n613 , n619 );
nand ( n54551 , n611 , n621 );
xor ( n54552 , n54550 , n54551 );
nand ( n54553 , n612 , n620 );
and ( n54554 , n54552 , n54553 );
and ( n54555 , n54550 , n54551 );
or ( n54556 , n54554 , n54555 );
xor ( n54557 , n54501 , n54502 );
xor ( n54558 , n54557 , n54504 );
xor ( n54559 , n54556 , n54558 );
xor ( n54560 , n54490 , n54491 );
xor ( n54561 , n54560 , n54493 );
and ( n54562 , n54559 , n54561 );
and ( n54563 , n54556 , n54558 );
or ( n54564 , n54562 , n54563 );
and ( n54565 , n54549 , n54564 );
and ( n54566 , n54546 , n54548 );
or ( n54567 , n54565 , n54566 );
xor ( n54568 , n54538 , n54567 );
xor ( n54569 , n54486 , n54499 );
xor ( n54570 , n54569 , n54515 );
and ( n54571 , n54568 , n54570 );
and ( n54572 , n54538 , n54567 );
or ( n54573 , n54571 , n54572 );
nand ( n54574 , n54530 , n54573 );
and ( n54575 , n54526 , n54574 );
not ( n54576 , n54575 );
nand ( n54577 , n610 , n622 );
nand ( n54578 , n609 , n623 );
xor ( n54579 , n54577 , n54578 );
and ( n54580 , n614 , n618 );
not ( n54581 , n54580 );
nand ( n54582 , n615 , n617 );
not ( n54583 , n54582 );
and ( n54584 , n54581 , n54583 );
and ( n54585 , n54582 , n54580 );
nor ( n54586 , n54584 , n54585 );
xor ( n54587 , n54579 , n54586 );
xor ( n54588 , n54550 , n54551 );
xor ( n54589 , n54588 , n54553 );
and ( n54590 , n54587 , n54589 );
nand ( n54591 , n615 , n619 );
not ( n54592 , n54591 );
and ( n54593 , n616 , n618 );
nand ( n54594 , n54592 , n54593 );
nand ( n54595 , n616 , n617 );
and ( n54596 , n54595 , n616 );
nor ( n54597 , C0 , n54596 );
xor ( n54598 , n54594 , n54597 );
nand ( n54599 , n612 , n622 );
not ( n54600 , n54599 );
nand ( n54601 , n614 , n620 );
not ( n54602 , n54601 );
or ( n54603 , n54600 , n54602 );
and ( n54604 , n613 , n621 );
nand ( n54605 , n54603 , n54604 );
not ( n54606 , n54599 );
not ( n54607 , n54601 );
nand ( n54608 , n54606 , n54607 );
and ( n54609 , n54605 , n54608 );
and ( n54610 , n54598 , n54609 );
and ( n54611 , n54594 , n54597 );
or ( n54612 , n54610 , n54611 );
xor ( n54613 , n54550 , n54551 );
xor ( n54614 , n54613 , n54553 );
and ( n54615 , n54612 , n54614 );
and ( n54616 , n54587 , n54612 );
or ( n54617 , n54590 , n54615 , n54616 );
xor ( n54618 , n54556 , n54558 );
xor ( n54619 , n54618 , n54561 );
xor ( n54620 , n54617 , n54619 );
xor ( n54621 , n54577 , n54578 );
and ( n54622 , n54621 , n54586 );
and ( n54623 , n54577 , n54578 );
or ( n54624 , n54622 , n54623 );
xor ( n54625 , n54539 , n54540 );
xor ( n54626 , n54625 , n54543 );
xor ( n54627 , n54624 , n54626 );
nand ( n54628 , n611 , n622 );
not ( n54629 , n54628 );
not ( n54630 , n54629 );
nand ( n54631 , n612 , n621 );
not ( n54632 , n54631 );
not ( n54633 , n54632 );
or ( n54634 , n54630 , n54633 );
not ( n54635 , n54628 );
not ( n54636 , n54631 );
or ( n54637 , n54635 , n54636 );
and ( n54638 , n615 , n618 );
nand ( n54639 , n54637 , n54638 );
nand ( n54640 , n54634 , n54639 );
not ( n54641 , n54640 );
xor ( n54642 , n54595 , n54641 );
nand ( n54643 , n610 , n623 );
not ( n54644 , n54643 );
not ( n54645 , n54644 );
nand ( n54646 , n613 , n620 );
not ( n54647 , n54646 );
not ( n54648 , n54647 );
or ( n54649 , n54645 , n54648 );
not ( n54650 , n54643 );
not ( n54651 , n54646 );
or ( n54652 , n54650 , n54651 );
and ( n54653 , n614 , n619 );
nand ( n54654 , n54652 , n54653 );
nand ( n54655 , n54649 , n54654 );
not ( n54656 , n54655 );
and ( n54657 , n54642 , n54656 );
and ( n54658 , n54595 , n54641 );
or ( n54659 , n54657 , n54658 );
xor ( n54660 , n54627 , n54659 );
xor ( n54661 , n54620 , n54660 );
xor ( n54662 , n54595 , n54641 );
xor ( n54663 , n54662 , n54656 );
not ( n54664 , n54643 );
not ( n54665 , n54653 );
or ( n54666 , n54664 , n54665 );
or ( n54667 , n54643 , n54653 );
nand ( n54668 , n54666 , n54667 );
and ( n54669 , n54668 , n54647 );
not ( n54670 , n54668 );
and ( n54671 , n54670 , n54646 );
nor ( n54672 , n54669 , n54671 );
not ( n54673 , n54672 );
not ( n54674 , n54673 );
not ( n54675 , n54631 );
not ( n54676 , n54638 );
or ( n54677 , n54675 , n54676 );
or ( n54678 , n54631 , n54638 );
nand ( n54679 , n54677 , n54678 );
and ( n54680 , n54679 , n54628 );
not ( n54681 , n54679 );
and ( n54682 , n54681 , n54629 );
nor ( n54683 , n54680 , n54682 );
not ( n54684 , n54683 );
or ( n54685 , n54674 , n54684 );
nand ( n54686 , n611 , n623 );
nand ( n54687 , n617 , n618 );
xor ( n54688 , n54686 , n54687 );
not ( n54689 , n54591 );
not ( n54690 , n54593 );
or ( n54691 , n54689 , n54690 );
or ( n54692 , n54591 , n54593 );
nand ( n54693 , n54691 , n54692 );
not ( n54694 , n54693 );
and ( n54695 , n54688 , n54694 );
and ( n54696 , n54686 , n54687 );
or ( n54697 , n54695 , n54696 );
not ( n54698 , n54697 );
nand ( n54699 , n54685 , n54698 );
not ( n54700 , n54683 );
nand ( n54701 , n54700 , n54672 );
and ( n54702 , n54699 , n54701 );
xor ( n54703 , n54663 , n54702 );
xor ( n54704 , n54550 , n54551 );
xor ( n54705 , n54704 , n54553 );
xor ( n54706 , n54587 , n54612 );
xor ( n54707 , n54705 , n54706 );
and ( n54708 , n54703 , n54707 );
and ( n54709 , n54663 , n54702 );
or ( n54710 , n54708 , n54709 );
nand ( n54711 , n54661 , n54710 );
xor ( n54712 , n54617 , n54619 );
and ( n54713 , n54712 , n54660 );
and ( n54714 , n54617 , n54619 );
or ( n54715 , n54713 , n54714 );
xor ( n54716 , n54507 , n54509 );
xor ( n54717 , n54716 , n54512 );
xor ( n54718 , n54546 , n54548 );
xor ( n54719 , n54718 , n54564 );
xor ( n54720 , n54717 , n54719 );
xor ( n54721 , n54624 , n54626 );
and ( n54722 , n54721 , n54659 );
and ( n54723 , n54624 , n54626 );
or ( n54724 , n54722 , n54723 );
xor ( n54725 , n54720 , n54724 );
nand ( n54726 , n54715 , n54725 );
xor ( n54727 , n54538 , n54567 );
xor ( n54728 , n54727 , n54570 );
xor ( n54729 , n54717 , n54719 );
and ( n54730 , n54729 , n54724 );
and ( n54731 , n54717 , n54719 );
or ( n54732 , n54730 , n54731 );
nand ( n54733 , n54728 , n54732 );
and ( n54734 , n54711 , n54726 , n54733 );
not ( n54735 , n54734 );
xor ( n54736 , n54663 , n54702 );
xor ( n54737 , n54736 , n54707 );
xor ( n54738 , n54594 , n54597 );
xor ( n54739 , n54738 , n54609 );
nand ( n54740 , n616 , n619 );
nand ( n54741 , n614 , n621 );
xor ( n54742 , n54740 , n54741 );
nand ( n54743 , n615 , n620 );
and ( n54744 , n54742 , n54743 );
and ( n54745 , n54740 , n54741 );
or ( n54746 , n54744 , n54745 );
not ( n54747 , n54599 );
not ( n54748 , n54604 );
or ( n54749 , n54747 , n54748 );
or ( n54750 , n54599 , n54604 );
nand ( n54751 , n54749 , n54750 );
and ( n54752 , n54751 , n54601 );
not ( n54753 , n54751 );
and ( n54754 , n54753 , n54607 );
nor ( n54755 , n54752 , n54754 );
xor ( n54756 , n54746 , n54755 );
nand ( n54757 , n613 , n622 );
nand ( n54758 , n612 , n623 );
nand ( n54759 , n54757 , n54758 );
not ( n54760 , n54759 );
nand ( n54761 , n616 , n620 );
nand ( n54762 , n617 , n619 );
nor ( n54763 , n54761 , n54762 );
not ( n54764 , n54763 );
or ( n54765 , n54760 , n54764 );
not ( n54766 , n54758 );
not ( n54767 , n54757 );
nand ( n54768 , n54766 , n54767 );
nand ( n54769 , n54765 , n54768 );
not ( n54770 , n54769 );
and ( n54771 , n54756 , n54770 );
and ( n54772 , n54746 , n54755 );
or ( n54773 , n54771 , n54772 );
xor ( n54774 , n54739 , n54773 );
not ( n54775 , n54683 );
not ( n54776 , n54672 );
or ( n54777 , n54775 , n54776 );
or ( n54778 , n54683 , n54672 );
nand ( n54779 , n54777 , n54778 );
xnor ( n54780 , n54779 , n54698 );
and ( n54781 , n54774 , n54780 );
and ( n54782 , n54739 , n54773 );
or ( n54783 , n54781 , n54782 );
nand ( n54784 , n54737 , n54783 );
not ( n54785 , n54784 );
xor ( n54786 , n54739 , n54773 );
xor ( n54787 , n54786 , n54780 );
xor ( n54788 , n54686 , n54687 );
not ( n54789 , n54693 );
xor ( n54790 , n54788 , n54789 );
and ( n54791 , n54687 , n617 );
nor ( n54792 , C0 , n54791 );
nand ( n54793 , n613 , n623 );
not ( n54794 , n54793 );
nand ( n54795 , n615 , n621 );
not ( n54796 , n54795 );
or ( n54797 , n54794 , n54796 );
and ( n54798 , n614 , n622 );
nand ( n54799 , n54797 , n54798 );
not ( n54800 , n54793 );
not ( n54801 , n54795 );
nand ( n54802 , n54800 , n54801 );
and ( n54803 , n54799 , n54802 );
xor ( n54804 , n54792 , n54803 );
xor ( n54805 , n54740 , n54741 );
xor ( n54806 , n54805 , n54743 );
and ( n54807 , n54804 , n54806 );
and ( n54808 , n54792 , n54803 );
or ( n54809 , n54807 , n54808 );
xor ( n54810 , n54790 , n54809 );
xor ( n54811 , n54746 , n54755 );
xor ( n54812 , n54811 , n54770 );
and ( n54813 , n54810 , n54812 );
and ( n54814 , n54790 , n54809 );
or ( n54815 , n54813 , n54814 );
and ( n54816 , n54787 , n54815 );
nor ( n54817 , n54785 , n54816 );
not ( n54818 , n54817 );
xor ( n54819 , n54790 , n54809 );
xor ( n54820 , n54819 , n54812 );
not ( n54821 , n54767 );
not ( n54822 , n54758 );
and ( n54823 , n54821 , n54822 );
and ( n54824 , n54758 , n54767 );
nor ( n54825 , n54823 , n54824 );
not ( n54826 , n54825 );
not ( n54827 , n54763 );
and ( n54828 , n54826 , n54827 );
and ( n54829 , n54763 , n54825 );
nor ( n54830 , n54828 , n54829 );
nand ( n54831 , n618 , n619 );
xnor ( n54832 , n54762 , n54761 );
xor ( n54833 , n54831 , n54832 );
nand ( n54834 , n616 , n621 );
nand ( n54835 , n615 , n622 );
xor ( n54836 , n54834 , n54835 );
nand ( n54837 , n617 , n620 );
and ( n54838 , n54836 , n54837 );
and ( n54839 , n54834 , n54835 );
or ( n54840 , n54838 , n54839 );
and ( n54841 , n54833 , n54840 );
and ( n54842 , n54831 , n54832 );
or ( n54843 , n54841 , n54842 );
xor ( n54844 , n54830 , n54843 );
xor ( n54845 , n54792 , n54803 );
xor ( n54846 , n54845 , n54806 );
and ( n54847 , n54844 , n54846 );
and ( n54848 , n54830 , n54843 );
or ( n54849 , n54847 , n54848 );
nand ( n54850 , n54820 , n54849 );
not ( n54851 , n54850 );
xor ( n54852 , n54830 , n54843 );
xor ( n54853 , n54852 , n54846 );
not ( n54854 , n54793 );
not ( n54855 , n54798 );
or ( n54856 , n54854 , n54855 );
or ( n54857 , n54793 , n54798 );
nand ( n54858 , n54856 , n54857 );
and ( n54859 , n54858 , n54795 );
not ( n54860 , n54858 );
and ( n54861 , n54860 , n54801 );
nor ( n54862 , n54859 , n54861 );
nand ( n54863 , n614 , n623 );
not ( n54864 , n54863 );
nand ( n54865 , n618 , n620 );
nand ( n54866 , n617 , n621 );
nor ( n54867 , n54865 , n54866 );
not ( n54868 , n54867 );
not ( n54869 , n54868 );
or ( n54870 , n54864 , n54869 );
and ( n54871 , n54831 , n618 );
nor ( n54872 , C0 , n54871 );
not ( n54873 , n54872 );
nand ( n54874 , n54870 , n54873 );
not ( n54875 , n54863 );
nand ( n54876 , n54875 , n54867 );
and ( n54877 , n54874 , n54876 );
xor ( n54878 , n54862 , n54877 );
xor ( n54879 , n54831 , n54832 );
xor ( n54880 , n54879 , n54840 );
and ( n54881 , n54878 , n54880 );
and ( n54882 , n54862 , n54877 );
or ( n54883 , n54881 , n54882 );
and ( n54884 , n54853 , n54883 );
nor ( n54885 , n54851 , n54884 );
not ( n54886 , n54885 );
xor ( n54887 , n54862 , n54877 );
xor ( n54888 , n54887 , n54880 );
nand ( n54889 , n616 , n622 );
nand ( n54890 , n615 , n623 );
xor ( n54891 , n54889 , n54890 );
nand ( n54892 , n619 , n620 );
and ( n54893 , n54891 , n54892 );
and ( n54894 , n54889 , n54890 );
or ( n54895 , n54893 , n54894 );
xor ( n54896 , n54834 , n54835 );
xor ( n54897 , n54896 , n54837 );
xor ( n54898 , n54895 , n54897 );
xor ( n54899 , n54863 , n54867 );
xnor ( n54900 , n54899 , n54872 );
and ( n54901 , n54898 , n54900 );
and ( n54902 , n54895 , n54897 );
or ( n54903 , n54901 , n54902 );
nand ( n54904 , n54888 , n54903 );
xor ( n54905 , n54895 , n54897 );
xor ( n54906 , n54905 , n54900 );
xnor ( n54907 , n54865 , n54866 );
nand ( n54908 , n616 , n623 );
not ( n54909 , n54908 );
nand ( n54910 , n617 , n622 );
not ( n54911 , n54910 );
or ( n54912 , n54909 , n54911 );
nand ( n54913 , n618 , n621 );
not ( n54914 , n54913 );
nand ( n54915 , n54912 , n54914 );
not ( n54916 , n54908 );
not ( n54917 , n54910 );
nand ( n54918 , n54916 , n54917 );
and ( n54919 , n54915 , n54918 );
xor ( n54920 , n54907 , n54919 );
xor ( n54921 , n54889 , n54890 );
xor ( n54922 , n54921 , n54892 );
and ( n54923 , n54920 , n54922 );
and ( n54924 , n54907 , n54919 );
or ( n54925 , n54923 , n54924 );
nand ( n54926 , n54906 , n54925 );
and ( n54927 , n54904 , n54926 );
not ( n54928 , n54927 );
and ( n54929 , n618 , n622 );
and ( n54930 , n619 , n621 );
and ( n54931 , n54929 , n54930 );
not ( n54932 , n619 );
not ( n54933 , n54892 );
or ( n54934 , n54932 , n54933 );
nand ( n54935 , n54934 , C1 );
xor ( n54936 , n54931 , n54935 );
not ( n54937 , n54908 );
not ( n54938 , n54917 );
or ( n54939 , n54937 , n54938 );
or ( n54940 , n54908 , n54917 );
nand ( n54941 , n54939 , n54940 );
and ( n54942 , n54941 , n54914 );
not ( n54943 , n54941 );
and ( n54944 , n54943 , n54913 );
nor ( n54945 , n54942 , n54944 );
and ( n54946 , n54936 , n54945 );
and ( n54947 , n54931 , n54935 );
or ( n54948 , n54946 , n54947 );
not ( n54949 , n54948 );
xor ( n54950 , n54907 , n54919 );
xor ( n54951 , n54950 , n54922 );
nand ( n54952 , n54949 , n54951 );
not ( n54953 , n54952 );
nand ( n54954 , n617 , n623 );
not ( n54955 , n54954 );
not ( n54956 , n54955 );
nand ( n54957 , n620 , n621 );
not ( n54958 , n54957 );
not ( n54959 , n54958 );
or ( n54960 , n54956 , n54959 );
not ( n54961 , n54954 );
not ( n54962 , n54957 );
or ( n54963 , n54961 , n54962 );
xor ( n54964 , n54929 , n54930 );
nand ( n54965 , n54963 , n54964 );
nand ( n54966 , n54960 , n54965 );
xor ( n54967 , n54931 , n54935 );
xor ( n54968 , n54967 , n54945 );
xor ( n54969 , n54966 , n54968 );
and ( n54970 , n54964 , n54954 );
not ( n54971 , n54964 );
and ( n54972 , n54971 , n54955 );
or ( n54973 , n54970 , n54972 );
xnor ( n54974 , n54958 , n54973 );
and ( n54975 , n619 , n622 );
and ( n54976 , n618 , n623 );
xor ( n54977 , n54975 , n54976 );
not ( n54978 , n620 );
not ( n54979 , n54957 );
or ( n54980 , n54978 , n54979 );
nand ( n54981 , n54980 , C1 );
and ( n54982 , n54977 , n54981 );
and ( n54983 , n54975 , n54976 );
or ( n54984 , n54982 , n54983 );
not ( n54985 , n54984 );
nand ( n54986 , n54974 , n54985 );
not ( n54987 , n54986 );
nand ( n54988 , n621 , n623 );
nand ( n54989 , n622 , n623 );
nor ( n54990 , n54988 , n54989 );
not ( n54991 , n54990 );
not ( n54992 , n54991 );
not ( n54993 , n54957 );
nand ( n54994 , n54993 , n623 );
not ( n54995 , n54994 );
and ( n54996 , n620 , n622 );
not ( n54997 , n54996 );
nand ( n54998 , n619 , n623 );
not ( n54999 , n54998 );
and ( n55000 , n54997 , n54999 );
and ( n55001 , n54996 , n54998 );
nor ( n55002 , n55000 , n55001 );
not ( n55003 , n55002 );
nor ( n55004 , n54995 , n55003 );
not ( n55005 , n55004 );
and ( n55006 , n54992 , n55005 );
not ( n55007 , n55002 );
nand ( n55008 , n620 , n623 );
nand ( n55009 , n55008 , n621 );
nand ( n55010 , n621 , n622 );
nor ( n55011 , n55009 , n55010 );
nand ( n55012 , n55007 , n55011 );
nand ( n55013 , n55003 , n54995 );
nand ( n55014 , n55012 , n55013 );
nor ( n55015 , n55006 , n55014 );
xor ( n55016 , n54975 , n54976 );
xor ( n55017 , n55016 , n54981 );
nor ( n55018 , n54892 , n54989 );
nor ( n55019 , n55017 , n55018 );
or ( n55020 , n55015 , n55019 );
nand ( n55021 , n55017 , n55018 );
nand ( n55022 , n55020 , n55021 );
not ( n55023 , n55022 );
or ( n55024 , n54987 , n55023 );
nor ( n55025 , n54974 , n54985 );
not ( n55026 , n55025 );
nand ( n55027 , n55024 , n55026 );
and ( n55028 , n54969 , n55027 );
and ( n55029 , n54966 , n54968 );
or ( n55030 , n55028 , n55029 );
not ( n55031 , n55030 );
or ( n55032 , n54953 , n55031 );
not ( n55033 , n54951 );
nand ( n55034 , n55033 , n54948 );
nand ( n55035 , n55032 , n55034 );
not ( n55036 , n55035 );
or ( n55037 , n54928 , n55036 );
nor ( n55038 , n54906 , n54925 );
nand ( n55039 , n54904 , n55038 );
or ( n55040 , n54888 , n54903 );
and ( n55041 , n55039 , n55040 );
nand ( n55042 , n55037 , n55041 );
not ( n55043 , n55042 );
or ( n55044 , n54886 , n55043 );
nor ( n55045 , n54883 , n54853 );
nand ( n55046 , n54850 , n55045 );
or ( n55047 , n54820 , n54849 );
and ( n55048 , n55046 , n55047 );
nand ( n55049 , n55044 , n55048 );
not ( n55050 , n55049 );
or ( n55051 , n54818 , n55050 );
nor ( n55052 , n54787 , n54815 );
nand ( n55053 , n55052 , n54784 );
or ( n55054 , n54783 , n54737 );
and ( n55055 , n55053 , n55054 );
nand ( n55056 , n55051 , n55055 );
not ( n55057 , n55056 );
or ( n55058 , n54735 , n55057 );
not ( n55059 , n54726 );
nor ( n55060 , n54661 , n54710 );
not ( n55061 , n55060 );
or ( n55062 , n55059 , n55061 );
or ( n55063 , n54715 , n54725 );
nand ( n55064 , n55062 , n55063 );
and ( n55065 , n54733 , n55064 );
nor ( n55066 , n54728 , n54732 );
nor ( n55067 , n55065 , n55066 );
nand ( n55068 , n55058 , n55067 );
not ( n55069 , n55068 );
or ( n55070 , n54576 , n55069 );
nor ( n55071 , n54530 , n54573 );
and ( n55072 , n54526 , n55071 );
nor ( n55073 , n54523 , n54525 );
nor ( n55074 , n55072 , n55073 );
nand ( n55075 , n55070 , n55074 );
not ( n55076 , n55075 );
or ( n55077 , n54471 , n55076 );
nor ( n55078 , n54352 , n54430 );
and ( n55079 , n55078 , n54457 );
nor ( n55080 , n54439 , n54456 );
nor ( n55081 , n55079 , n55080 );
not ( n55082 , n55081 );
and ( n55083 , n55082 , n54469 );
nor ( n55084 , n54466 , n54468 );
nor ( n55085 , n55083 , n55084 );
nand ( n55086 , n55077 , n55085 );
not ( n55087 , n55086 );
or ( n55088 , n54290 , n55087 );
nor ( n55089 , n54183 , n54209 );
and ( n55090 , n55089 , n54234 );
nor ( n55091 , n54218 , n54233 );
nor ( n55092 , n55090 , n55091 );
not ( n55093 , n54288 );
or ( n55094 , n55092 , n55093 );
nor ( n55095 , n54285 , n54287 );
not ( n55096 , n55095 );
nand ( n55097 , n55094 , n55096 );
and ( n55098 , n55097 , n54277 );
nor ( n55099 , n54249 , n54257 );
and ( n55100 , n55099 , n54269 );
nor ( n55101 , n54263 , n54268 );
nor ( n55102 , n55100 , n55101 );
not ( n55103 , n54275 );
or ( n55104 , n55102 , n55103 );
or ( n55105 , n54273 , n54274 );
nand ( n55106 , n55104 , n55105 );
nor ( n55107 , n55098 , n55106 );
nand ( n55108 , n55088 , n55107 );
nand ( n55109 , n54267 , n608 );
nor ( n55110 , n55108 , n55109 );
not ( n55111 , n55110 );
nand ( n55112 , n55108 , n55109 );
nand ( n55113 , n55111 , n55112 );
buf ( n55114 , n55113 );
buf ( n55115 , n15731 );
buf ( n55116 , n15269 );
not ( n55117 , n55116 );
buf ( n55118 , n55117 );
buf ( n55119 , n55118 );
and ( n55120 , n55115 , n55119 );
not ( n55121 , n55115 );
buf ( n55122 , n15269 );
and ( n55123 , n55121 , n55122 );
nor ( n55124 , n55120 , n55123 );
buf ( n55125 , n55124 );
buf ( n55126 , n55125 );
buf ( n55127 , n15731 );
nand ( n55128 , n55126 , n55127 );
buf ( n55129 , n55128 );
buf ( n55130 , n55129 );
not ( n55131 , n55130 );
buf ( n55132 , n55131 );
buf ( n55133 , n55132 );
and ( n55134 , n55114 , n55133 );
not ( n55135 , n608 );
nor ( n55136 , n55135 , n54276 );
not ( n55137 , n55136 );
and ( n55138 , n54235 , n54288 , n54258 );
not ( n55139 , n55138 );
not ( n55140 , n55086 );
or ( n55141 , n55139 , n55140 );
and ( n55142 , n55097 , n54258 );
nor ( n55143 , n55142 , n55099 );
nand ( n55144 , n55141 , n55143 );
not ( n55145 , n55144 );
or ( n55146 , n55137 , n55145 );
and ( n55147 , n55101 , n54275 );
not ( n55148 , n55105 );
nor ( n55149 , n55147 , n55148 , n609 );
not ( n55150 , n55149 );
nand ( n55151 , n55150 , n608 );
nand ( n55152 , n55146 , n55151 );
buf ( n55153 , n55152 );
buf ( n55154 , n55125 );
not ( n55155 , n55154 );
buf ( n55156 , n55155 );
buf ( n55157 , n55156 );
and ( n55158 , n55153 , n55157 );
nor ( n55159 , n55134 , n55158 );
buf ( n55160 , n55159 );
buf ( n55161 , n55160 );
buf ( n55162 , n7276 );
buf ( n55163 , n55162 );
buf ( n55164 , n16472 );
xnor ( n55165 , n55163 , n55164 );
buf ( n55166 , n55165 );
buf ( n55167 , n55166 );
buf ( n55168 , n55118 );
nor ( n55169 , n55167 , n55168 );
buf ( n55170 , n55169 );
buf ( n55171 , n55170 );
not ( n55172 , n55171 );
buf ( n55173 , n55166 );
buf ( n55174 , n55162 );
buf ( n55175 , n15269 );
xor ( n55176 , n55174 , n55175 );
buf ( n55177 , n55176 );
buf ( n55178 , n55177 );
and ( n55179 , n55173 , n55178 );
buf ( n55180 , n55179 );
buf ( n55181 , n55180 );
buf ( n55182 , n15269 );
buf ( n55183 , n55182 );
buf ( n55184 , n55183 );
buf ( n55185 , n55184 );
nand ( n55186 , n55181 , n55185 );
buf ( n55187 , n55186 );
buf ( n55188 , n55187 );
nand ( n55189 , n55172 , n55188 );
buf ( n55190 , n55189 );
buf ( n55191 , n55190 );
xor ( n55192 , n55161 , n55191 );
buf ( n55193 , n55118 );
buf ( n55194 , n55193 );
buf ( n55195 , n55194 );
buf ( n55196 , n55195 );
not ( n55197 , n55196 );
buf ( n55198 , n55197 );
buf ( n55199 , n55198 );
buf ( n55200 , n55199 );
buf ( n55201 , n55200 );
buf ( n55202 , n55201 );
buf ( n55203 , n55152 );
not ( n55204 , n55203 );
buf ( n55205 , n55204 );
buf ( n55206 , n55205 );
and ( n55207 , n55202 , n55206 );
not ( n55208 , n55202 );
buf ( n55209 , n55152 );
and ( n55210 , n55208 , n55209 );
nor ( n55211 , n55207 , n55210 );
buf ( n55212 , n55211 );
buf ( n55213 , n55212 );
not ( n55214 , n55213 );
buf ( n55215 , n55214 );
buf ( n55216 , n55215 );
buf ( n55217 , n55180 );
and ( n55218 , n55216 , n55217 );
buf ( n55219 , n55170 );
nor ( n55220 , n55218 , n55219 );
buf ( n55221 , n55220 );
buf ( n55222 , n55221 );
not ( n55223 , n54269 );
nor ( n55224 , n54259 , n55093 , n55223 );
and ( n55225 , n54469 , n54235 , n55224 );
not ( n55226 , n55225 );
not ( n55227 , n54458 );
not ( n55228 , n55075 );
or ( n55229 , n55227 , n55228 );
nand ( n55230 , n55229 , n55081 );
not ( n55231 , n55230 );
or ( n55232 , n55226 , n55231 );
not ( n55233 , n54235 );
not ( n55234 , n55084 );
or ( n55235 , n55233 , n55234 );
nand ( n55236 , n55235 , n55092 );
and ( n55237 , n55236 , n55224 );
and ( n55238 , n55095 , n54258 );
nor ( n55239 , n55238 , n55099 );
or ( n55240 , n55239 , n55223 );
not ( n55241 , n55101 );
nand ( n55242 , n55240 , n55241 );
nor ( n55243 , n55237 , n55242 );
nand ( n55244 , n55232 , n55243 );
nand ( n55245 , n54275 , n55105 );
nor ( n55246 , n55244 , n55245 );
not ( n55247 , n55246 );
nand ( n55248 , n55244 , n55245 );
nand ( n55249 , n55247 , n55248 );
buf ( n55250 , n55249 );
buf ( n55251 , n55132 );
and ( n55252 , n55250 , n55251 );
buf ( n55253 , n55113 );
buf ( n55254 , n55156 );
and ( n55255 , n55253 , n55254 );
nor ( n55256 , n55252 , n55255 );
buf ( n55257 , n55256 );
buf ( n55258 , n55257 );
nand ( n55259 , n55222 , n55258 );
buf ( n55260 , n55259 );
buf ( n55261 , n55260 );
not ( n55262 , n55261 );
buf ( n55263 , n55262 );
buf ( n55264 , n55263 );
and ( n55265 , n55192 , n55264 );
and ( n55266 , n55161 , n55191 );
or ( n55267 , n55265 , n55266 );
buf ( n55268 , n55267 );
buf ( n55269 , n55268 );
buf ( n55270 , n55152 );
buf ( n55271 , n55132 );
nand ( n55272 , n55270 , n55271 );
buf ( n55273 , n55272 );
buf ( n55274 , n55273 );
nand ( n55275 , n55269 , n55274 );
buf ( n55276 , n55275 );
nor ( n55277 , n54134 , n55276 );
nand ( n55278 , n54125 , n55277 );
buf ( n55279 , n55278 );
xor ( n55280 , n54119 , n55279 );
buf ( n55281 , n44039 );
buf ( n55282 , n42504 );
buf ( n55283 , n38412 );
and ( n55284 , n55282 , n55283 );
not ( n55285 , n55282 );
buf ( n55286 , n46623 );
and ( n55287 , n55285 , n55286 );
nor ( n55288 , n55284 , n55287 );
buf ( n55289 , n55288 );
buf ( n55290 , n55289 );
or ( n55291 , n55281 , n55290 );
buf ( n55292 , n52698 );
not ( n55293 , n55292 );
buf ( n55294 , n55293 );
buf ( n55295 , n55294 );
buf ( n55296 , n52171 );
or ( n55297 , n55295 , n55296 );
nand ( n55298 , n55291 , n55297 );
buf ( n55299 , n55298 );
buf ( n55300 , n55299 );
and ( n55301 , n55280 , n55300 );
and ( n55302 , n54119 , n55279 );
or ( n55303 , n55301 , n55302 );
buf ( n55304 , n55303 );
buf ( n55305 , n55304 );
buf ( n55306 , n42668 );
not ( n55307 , n55306 );
buf ( n55308 , n53003 );
not ( n55309 , n55308 );
or ( n55310 , n55307 , n55309 );
buf ( n55311 , n42672 );
not ( n55312 , n55311 );
buf ( n55313 , n47932 );
not ( n55314 , n55313 );
or ( n55315 , n55312 , n55314 );
buf ( n55316 , n38821 );
buf ( n55317 , n42671 );
nand ( n55318 , n55316 , n55317 );
buf ( n55319 , n55318 );
buf ( n55320 , n55319 );
nand ( n55321 , n55315 , n55320 );
buf ( n55322 , n55321 );
buf ( n55323 , n55322 );
buf ( n55324 , n42712 );
nand ( n55325 , n55323 , n55324 );
buf ( n55326 , n55325 );
buf ( n55327 , n55326 );
nand ( n55328 , n55310 , n55327 );
buf ( n55329 , n55328 );
buf ( n55330 , n55329 );
xor ( n55331 , n55305 , n55330 );
buf ( n55332 , n47716 );
buf ( n55333 , n42062 );
and ( n55334 , n55332 , n55333 );
not ( n55335 , n55332 );
buf ( n55336 , n49425 );
and ( n55337 , n55335 , n55336 );
nor ( n55338 , n55334 , n55337 );
buf ( n55339 , n55338 );
buf ( n55340 , n55339 );
not ( n55341 , n55340 );
buf ( n55342 , n44776 );
not ( n55343 , n55342 );
or ( n55344 , n55341 , n55343 );
buf ( n55345 , n53215 );
not ( n55346 , n55345 );
buf ( n55347 , n36912 );
nand ( n55348 , n55346 , n55347 );
buf ( n55349 , n55348 );
buf ( n55350 , n55349 );
nand ( n55351 , n55344 , n55350 );
buf ( n55352 , n55351 );
buf ( n55353 , n55352 );
and ( n55354 , n55331 , n55353 );
and ( n55355 , n55305 , n55330 );
or ( n55356 , n55354 , n55355 );
buf ( n55357 , n55356 );
nand ( n55358 , n54118 , n55357 );
nand ( n55359 , n54115 , n55358 );
buf ( n55360 , n55359 );
and ( n55361 , n53937 , n55360 );
and ( n55362 , n53794 , n53936 );
or ( n55363 , n55361 , n55362 );
buf ( n55364 , n55363 );
buf ( n55365 , n55364 );
buf ( n55366 , n48855 );
not ( n55367 , n55366 );
buf ( n55368 , n48808 );
not ( n55369 , n55368 );
buf ( n55370 , n36430 );
not ( n55371 , n55370 );
or ( n55372 , n55369 , n55371 );
buf ( n55373 , n40067 );
not ( n55374 , n55373 );
buf ( n55375 , n48818 );
nand ( n55376 , n55374 , n55375 );
buf ( n55377 , n55376 );
buf ( n55378 , n55377 );
nand ( n55379 , n55372 , n55378 );
buf ( n55380 , n55379 );
buf ( n55381 , n55380 );
not ( n55382 , n55381 );
or ( n55383 , n55367 , n55382 );
buf ( n55384 , n52950 );
buf ( n55385 , n48868 );
nand ( n55386 , n55384 , n55385 );
buf ( n55387 , n55386 );
buf ( n55388 , n55387 );
nand ( n55389 , n55383 , n55388 );
buf ( n55390 , n55389 );
buf ( n55391 , n55390 );
xor ( n55392 , n52636 , n52661 );
xor ( n55393 , n55392 , n52804 );
buf ( n55394 , n55393 );
buf ( n55395 , n55394 );
xor ( n55396 , n55391 , n55395 );
not ( n55397 , n52343 );
buf ( n55398 , n52294 );
buf ( n55399 , n52307 );
and ( n55400 , n55398 , n55399 );
not ( n55401 , n55398 );
buf ( n55402 , n52318 );
and ( n55403 , n55401 , n55402 );
nor ( n55404 , n55400 , n55403 );
buf ( n55405 , n55404 );
not ( n55406 , n55405 );
not ( n55407 , n55406 );
or ( n55408 , n55397 , n55407 );
nand ( n55409 , n55405 , n52344 );
nand ( n55410 , n55408 , n55409 );
buf ( n55411 , n55410 );
not ( n55412 , n55411 );
buf ( n55413 , n55412 );
buf ( n55414 , n55413 );
not ( n55415 , n55414 );
not ( n55416 , n44267 );
not ( n55417 , n37686 );
not ( n55418 , n41611 );
or ( n55419 , n55417 , n55418 );
nand ( n55420 , n41608 , n37708 );
nand ( n55421 , n55419 , n55420 );
not ( n55422 , n55421 );
or ( n55423 , n55416 , n55422 );
buf ( n55424 , n53185 );
buf ( n55425 , n43868 );
nand ( n55426 , n55424 , n55425 );
buf ( n55427 , n55426 );
nand ( n55428 , n55423 , n55427 );
buf ( n55429 , n55428 );
not ( n55430 , n55429 );
or ( n55431 , n55415 , n55430 );
xor ( n55432 , n52749 , n52773 );
xor ( n55433 , n55432 , n52800 );
buf ( n55434 , n55433 );
buf ( n55435 , n55428 );
not ( n55436 , n55435 );
buf ( n55437 , n55410 );
nand ( n55438 , n55436 , n55437 );
buf ( n55439 , n55438 );
buf ( n55440 , n55439 );
nand ( n55441 , n55434 , n55440 );
buf ( n55442 , n55441 );
buf ( n55443 , n55442 );
nand ( n55444 , n55431 , n55443 );
buf ( n55445 , n55444 );
buf ( n55446 , n55445 );
and ( n55447 , n55396 , n55446 );
and ( n55448 , n55391 , n55395 );
or ( n55449 , n55447 , n55448 );
buf ( n55450 , n55449 );
buf ( n55451 , n55450 );
xor ( n55452 , n55365 , n55451 );
not ( n55453 , n53118 );
not ( n55454 , n53100 );
and ( n55455 , n55453 , n55454 );
and ( n55456 , n53118 , n53100 );
nor ( n55457 , n55455 , n55456 );
and ( n55458 , n55457 , n53085 );
not ( n55459 , n55457 );
not ( n55460 , n53085 );
and ( n55461 , n55459 , n55460 );
nor ( n55462 , n55458 , n55461 );
buf ( n55463 , n55462 );
and ( n55464 , n55452 , n55463 );
and ( n55465 , n55365 , n55451 );
or ( n55466 , n55464 , n55465 );
buf ( n55467 , n55466 );
buf ( n55468 , n55467 );
and ( n55469 , n53790 , n55468 );
and ( n55470 , n53477 , n53789 );
or ( n55471 , n55469 , n55470 );
buf ( n55472 , n55471 );
buf ( n55473 , n55472 );
not ( n55474 , n55473 );
buf ( n55475 , n55474 );
buf ( n55476 , n55475 );
buf ( n55477 , n53065 );
buf ( n55478 , n52873 );
and ( n55479 , n55477 , n55478 );
not ( n55480 , n55477 );
buf ( n55481 , n52876 );
and ( n55482 , n55480 , n55481 );
nor ( n55483 , n55479 , n55482 );
buf ( n55484 , n55483 );
buf ( n55485 , n52881 );
and ( n55486 , n55484 , n55485 );
not ( n55487 , n55484 );
not ( n55488 , n55485 );
and ( n55489 , n55487 , n55488 );
nor ( n55490 , n55486 , n55489 );
buf ( n55491 , n55490 );
xor ( n55492 , n55476 , n55491 );
xor ( n55493 , n53130 , n53338 );
xor ( n55494 , n55493 , n53343 );
buf ( n55495 , n55494 );
and ( n55496 , n55492 , n55495 );
and ( n55497 , n55476 , n55491 );
or ( n55498 , n55496 , n55497 );
buf ( n55499 , n55498 );
xor ( n55500 , n53473 , n55499 );
xor ( n55501 , n53083 , n53122 );
xor ( n55502 , n55501 , n53126 );
buf ( n55503 , n55502 );
buf ( n55504 , n55503 );
xor ( n55505 , n53134 , n53319 );
xor ( n55506 , n55505 , n53330 );
buf ( n55507 , n55506 );
buf ( n55508 , n55507 );
xor ( n55509 , n55504 , n55508 );
buf ( n55510 , n53166 );
buf ( n55511 , n53316 );
xor ( n55512 , n55510 , n55511 );
buf ( n55513 , n53137 );
xnor ( n55514 , n55512 , n55513 );
buf ( n55515 , n55514 );
xor ( n55516 , n52936 , n52961 );
xor ( n55517 , n55516 , n53056 );
buf ( n55518 , n55517 );
or ( n55519 , n55515 , n55518 );
xor ( n55520 , n53029 , n53032 );
xor ( n55521 , n55520 , n53051 );
buf ( n55522 , n55521 );
buf ( n55523 , n55522 );
buf ( n55524 , n44708 );
not ( n55525 , n55524 );
buf ( n55526 , n44533 );
not ( n55527 , n55526 );
buf ( n55528 , n37268 );
not ( n55529 , n55528 );
or ( n55530 , n55527 , n55529 );
buf ( n55531 , n50463 );
buf ( n55532 , n44530 );
nand ( n55533 , n55531 , n55532 );
buf ( n55534 , n55533 );
buf ( n55535 , n55534 );
nand ( n55536 , n55530 , n55535 );
buf ( n55537 , n55536 );
buf ( n55538 , n55537 );
not ( n55539 , n55538 );
or ( n55540 , n55525 , n55539 );
buf ( n55541 , n53048 );
buf ( n55542 , n44496 );
nand ( n55543 , n55541 , n55542 );
buf ( n55544 , n55543 );
buf ( n55545 , n55544 );
nand ( n55546 , n55540 , n55545 );
buf ( n55547 , n55546 );
buf ( n55548 , n55547 );
buf ( n55549 , C0 );
buf ( n55550 , n55549 );
xor ( n55551 , n55548 , n55550 );
buf ( n55552 , n46912 );
not ( n55553 , n55552 );
buf ( n55554 , n53771 );
not ( n55555 , n55554 );
or ( n55556 , n55553 , n55555 );
buf ( n55557 , n51622 );
not ( n55558 , n55557 );
buf ( n55559 , n50871 );
not ( n55560 , n55559 );
or ( n55561 , n55558 , n55560 );
buf ( n55562 , n50876 );
buf ( n55563 , n46890 );
nand ( n55564 , n55562 , n55563 );
buf ( n55565 , n55564 );
buf ( n55566 , n55565 );
nand ( n55567 , n55561 , n55566 );
buf ( n55568 , n55567 );
buf ( n55569 , n55568 );
buf ( n55570 , n47331 );
nand ( n55571 , n55569 , n55570 );
buf ( n55572 , n55571 );
buf ( n55573 , n55572 );
nand ( n55574 , n55556 , n55573 );
buf ( n55575 , n55574 );
buf ( n55576 , n55575 );
and ( n55577 , n55551 , n55576 );
or ( n55578 , n55577 , C0 );
buf ( n55579 , n55578 );
buf ( n55580 , n55579 );
xor ( n55581 , n55523 , n55580 );
xor ( n55582 , n53160 , n53156 );
xnor ( n55583 , n55582 , n53164 );
buf ( n55584 , n55583 );
and ( n55585 , n55581 , n55584 );
and ( n55586 , n55523 , n55580 );
or ( n55587 , n55585 , n55586 );
buf ( n55588 , n55587 );
nand ( n55589 , n55519 , n55588 );
buf ( n55590 , n55515 );
buf ( n55591 , n55518 );
nand ( n55592 , n55590 , n55591 );
buf ( n55593 , n55592 );
and ( n55594 , n55589 , n55593 );
buf ( n55595 , n55594 );
and ( n55596 , n55509 , n55595 );
and ( n55597 , n55504 , n55508 );
or ( n55598 , n55596 , n55597 );
buf ( n55599 , n55598 );
buf ( n55600 , n55599 );
xor ( n55601 , n53477 , n53789 );
xor ( n55602 , n55601 , n55468 );
buf ( n55603 , n55602 );
buf ( n55604 , n55603 );
not ( n55605 , n55604 );
xor ( n55606 , n53191 , n53199 );
xor ( n55607 , n55606 , n53312 );
buf ( n55608 , n55607 );
buf ( n55609 , n55608 );
not ( n55610 , n53151 );
not ( n55611 , n55610 );
not ( n55612 , n51473 );
and ( n55613 , n55611 , n55612 );
and ( n55614 , n51493 , n42280 );
not ( n55615 , n51493 );
and ( n55616 , n55615 , n39927 );
or ( n55617 , n55614 , n55616 );
and ( n55618 , n55617 , n51488 );
nor ( n55619 , n55613 , n55618 );
not ( n55620 , n55619 );
not ( n55621 , n55620 );
xor ( n55622 , n53210 , n53232 );
xor ( n55623 , n55622 , n53307 );
buf ( n55624 , n55623 );
not ( n55625 , n55624 );
or ( n55626 , n55621 , n55625 );
not ( n55627 , n55624 );
buf ( n55628 , n55627 );
not ( n55629 , n55628 );
buf ( n55630 , n55619 );
not ( n55631 , n55630 );
or ( n55632 , n55629 , n55631 );
not ( n55633 , n43868 );
not ( n55634 , n55421 );
or ( n55635 , n55633 , n55634 );
buf ( n55636 , n41608 );
not ( n55637 , n55636 );
buf ( n55638 , n37745 );
not ( n55639 , n55638 );
or ( n55640 , n55637 , n55639 );
buf ( n55641 , n42596 );
buf ( n55642 , n41611 );
nand ( n55643 , n55641 , n55642 );
buf ( n55644 , n55643 );
buf ( n55645 , n55644 );
nand ( n55646 , n55640 , n55645 );
buf ( n55647 , n55646 );
buf ( n55648 , n55647 );
buf ( n55649 , n44267 );
nand ( n55650 , n55648 , n55649 );
buf ( n55651 , n55650 );
nand ( n55652 , n55635 , n55651 );
buf ( n55653 , n55652 );
buf ( n55654 , n42315 );
not ( n55655 , n55654 );
buf ( n55656 , n53736 );
not ( n55657 , n55656 );
or ( n55658 , n55655 , n55657 );
xor ( n55659 , n37586 , n42263 );
buf ( n55660 , n55659 );
not ( n55661 , n55660 );
buf ( n55662 , n42252 );
nand ( n55663 , n55661 , n55662 );
buf ( n55664 , n55663 );
buf ( n55665 , n55664 );
nand ( n55666 , n55658 , n55665 );
buf ( n55667 , n55666 );
buf ( n55668 , n55667 );
xor ( n55669 , n55653 , n55668 );
buf ( n55670 , n53599 );
buf ( n55671 , n53655 );
xor ( n55672 , n55670 , n55671 );
buf ( n55673 , n53625 );
xnor ( n55674 , n55672 , n55673 );
buf ( n55675 , n55674 );
not ( n55676 , n55675 );
not ( n55677 , n55676 );
not ( n55678 , n42668 );
not ( n55679 , n55322 );
or ( n55680 , n55678 , n55679 );
buf ( n55681 , n42672 );
not ( n55682 , n55681 );
buf ( n55683 , n42485 );
not ( n55684 , n55683 );
or ( n55685 , n55682 , n55684 );
buf ( n55686 , n30187 );
buf ( n55687 , n42671 );
nand ( n55688 , n55686 , n55687 );
buf ( n55689 , n55688 );
buf ( n55690 , n55689 );
nand ( n55691 , n55685 , n55690 );
buf ( n55692 , n55691 );
buf ( n55693 , n55692 );
buf ( n55694 , n42712 );
nand ( n55695 , n55693 , n55694 );
buf ( n55696 , n55695 );
nand ( n55697 , n55680 , n55696 );
not ( n55698 , n55697 );
or ( n55699 , n55677 , n55698 );
not ( n55700 , n55675 );
not ( n55701 , n55697 );
not ( n55702 , n55701 );
or ( n55703 , n55700 , n55702 );
or ( n55704 , n54134 , n54124 );
nand ( n55705 , n55704 , n55276 );
nand ( n55706 , n55705 , n55278 );
buf ( n55707 , n55706 );
not ( n55708 , n42008 );
and ( n55709 , n55708 , n47068 );
not ( n55710 , n55708 );
and ( n55711 , n55710 , n42403 );
or ( n55712 , n55709 , n55711 );
not ( n55713 , n55712 );
not ( n55714 , n46620 );
or ( n55715 , n55713 , n55714 );
not ( n55716 , n55289 );
nand ( n55717 , n55716 , n52174 );
nand ( n55718 , n55715 , n55717 );
buf ( n55719 , n55718 );
xor ( n55720 , n55707 , n55719 );
buf ( n55721 , n55268 );
buf ( n55722 , n55273 );
or ( n55723 , n55721 , n55722 );
buf ( n55724 , n55276 );
nand ( n55725 , n55723 , n55724 );
buf ( n55726 , n55725 );
not ( n55727 , n53649 );
not ( n55728 , n54070 );
or ( n55729 , n55727 , n55728 );
not ( n55730 , n48357 );
not ( n55731 , n53579 );
or ( n55732 , n55730 , n55731 );
buf ( n55733 , n42149 );
buf ( n55734 , n54067 );
nand ( n55735 , n55733 , n55734 );
buf ( n55736 , n55735 );
nand ( n55737 , n55732 , n55736 );
nand ( n55738 , n55737 , n53628 );
nand ( n55739 , n55729 , n55738 );
xor ( n55740 , n55726 , n55739 );
buf ( n55741 , n13653 );
not ( n55742 , n55741 );
not ( n55743 , n50591 );
buf ( n55744 , n55743 );
not ( n55745 , n55744 );
or ( n55746 , n55742 , n55745 );
buf ( n55747 , n50591 );
buf ( n55748 , n43099 );
nand ( n55749 , n55747 , n55748 );
buf ( n55750 , n55749 );
buf ( n55751 , n55750 );
nand ( n55752 , n55746 , n55751 );
buf ( n55753 , n55752 );
buf ( n55754 , n55753 );
not ( n55755 , n55754 );
buf ( n55756 , n39999 );
not ( n55757 , n55756 );
or ( n55758 , n55755 , n55757 );
buf ( n55759 , n54014 );
buf ( n55760 , n48705 );
nand ( n55761 , n55759 , n55760 );
buf ( n55762 , n55761 );
buf ( n55763 , n55762 );
nand ( n55764 , n55758 , n55763 );
buf ( n55765 , n55764 );
and ( n55766 , n55740 , n55765 );
and ( n55767 , n55726 , n55739 );
or ( n55768 , n55766 , n55767 );
buf ( n55769 , n55768 );
and ( n55770 , n55720 , n55769 );
and ( n55771 , n55707 , n55719 );
or ( n55772 , n55770 , n55771 );
buf ( n55773 , n55772 );
nand ( n55774 , n55703 , n55773 );
nand ( n55775 , n55699 , n55774 );
buf ( n55776 , n55775 );
and ( n55777 , n55669 , n55776 );
and ( n55778 , n55653 , n55668 );
or ( n55779 , n55777 , n55778 );
buf ( n55780 , n55779 );
buf ( n55781 , n55780 );
nand ( n55782 , n55632 , n55781 );
buf ( n55783 , n55782 );
nand ( n55784 , n55626 , n55783 );
buf ( n55785 , n55784 );
xor ( n55786 , n55609 , n55785 );
xor ( n55787 , n53512 , n53752 );
xor ( n55788 , n55787 , n53779 );
buf ( n55789 , n55788 );
buf ( n55790 , n55789 );
and ( n55791 , n55786 , n55790 );
and ( n55792 , n55609 , n55785 );
or ( n55793 , n55791 , n55792 );
buf ( n55794 , n55793 );
buf ( n55795 , n55794 );
xor ( n55796 , n53574 , n53721 );
xor ( n55797 , n55796 , n53747 );
buf ( n55798 , n55797 );
buf ( n55799 , n55798 );
not ( n55800 , n55799 );
buf ( n55801 , n48868 );
not ( n55802 , n55801 );
buf ( n55803 , n55380 );
not ( n55804 , n55803 );
or ( n55805 , n55802 , n55804 );
buf ( n55806 , n48808 );
not ( n55807 , n55806 );
buf ( n55808 , n39891 );
not ( n55809 , n55808 );
or ( n55810 , n55807 , n55809 );
buf ( n55811 , n39891 );
not ( n55812 , n55811 );
buf ( n55813 , n55812 );
buf ( n55814 , n55813 );
buf ( n55815 , n48818 );
nand ( n55816 , n55814 , n55815 );
buf ( n55817 , n55816 );
buf ( n55818 , n55817 );
nand ( n55819 , n55810 , n55818 );
buf ( n55820 , n55819 );
buf ( n55821 , n55820 );
buf ( n55822 , n48855 );
nand ( n55823 , n55821 , n55822 );
buf ( n55824 , n55823 );
buf ( n55825 , n55824 );
nand ( n55826 , n55805 , n55825 );
buf ( n55827 , n55826 );
buf ( n55828 , n55827 );
not ( n55829 , n55828 );
or ( n55830 , n55800 , n55829 );
buf ( n55831 , n55798 );
buf ( n55832 , n55827 );
or ( n55833 , n55831 , n55832 );
not ( n55834 , n12488 );
buf ( n55835 , n12485 );
buf ( n55836 , n12470 );
nand ( n55837 , n55835 , n55836 );
buf ( n55838 , n55837 );
nand ( n55839 , n55834 , n55838 );
buf ( n55840 , n55839 );
not ( n55841 , n55840 );
buf ( n55842 , n55841 );
not ( n55843 , n55842 );
buf ( n55844 , n37602 );
not ( n55845 , n55844 );
or ( n55846 , n55843 , n55845 );
buf ( n55847 , n36360 );
buf ( n55848 , n55840 );
nand ( n55849 , n55847 , n55848 );
buf ( n55850 , n55849 );
buf ( n55851 , n55850 );
nand ( n55852 , n55846 , n55851 );
buf ( n55853 , n55852 );
buf ( n55854 , n43053 );
buf ( n55855 , n53554 );
nand ( n55856 , n55854 , n55855 );
buf ( n55857 , n55856 );
buf ( n55858 , n55857 );
nand ( n55859 , C1 , n55858 );
buf ( n55860 , n55859 );
buf ( n55861 , n55860 );
not ( n55862 , n55861 );
buf ( n55863 , n55862 );
not ( n55864 , n55863 );
buf ( n55865 , n46390 );
not ( n55866 , n55865 );
buf ( n55867 , n38068 );
not ( n55868 , n55867 );
or ( n55869 , n55866 , n55868 );
buf ( n55870 , n43400 );
buf ( n55871 , n46393 );
nand ( n55872 , n55870 , n55871 );
buf ( n55873 , n55872 );
buf ( n55874 , n55873 );
nand ( n55875 , n55869 , n55874 );
buf ( n55876 , n55875 );
buf ( n55877 , n55876 );
not ( n55878 , n55877 );
buf ( n55879 , n53817 );
not ( n55880 , n55879 );
buf ( n55881 , n55880 );
buf ( n55882 , n55881 );
not ( n55883 , n55882 );
or ( n55884 , n55878 , n55883 );
buf ( n55885 , n53811 );
buf ( n55886 , n38054 );
nand ( n55887 , n55885 , n55886 );
buf ( n55888 , n55887 );
buf ( n55889 , n55888 );
nand ( n55890 , n55884 , n55889 );
buf ( n55891 , n55890 );
buf ( n55892 , n55891 );
not ( n55893 , n55892 );
buf ( n55894 , n55893 );
not ( n55895 , n55894 );
and ( n55896 , n55864 , n55895 );
buf ( n55897 , n55863 );
buf ( n55898 , n55894 );
nand ( n55899 , n55897 , n55898 );
buf ( n55900 , n55899 );
buf ( n55901 , n51004 );
not ( n55902 , n55901 );
buf ( n55903 , n36500 );
not ( n55904 , n55903 );
or ( n55905 , n55902 , n55904 );
buf ( n55906 , n33076 );
buf ( n55907 , n51001 );
nand ( n55908 , n55906 , n55907 );
buf ( n55909 , n55908 );
buf ( n55910 , n55909 );
nand ( n55911 , n55905 , n55910 );
buf ( n55912 , n55911 );
not ( n55913 , n55912 );
not ( n55914 , n43250 );
or ( n55915 , n55913 , n55914 );
buf ( n55916 , n53703 );
buf ( n55917 , n42527 );
nand ( n55918 , n55916 , n55917 );
buf ( n55919 , n55918 );
nand ( n55920 , n55915 , n55919 );
buf ( n55921 , n55920 );
and ( n55922 , n55900 , n55921 );
nor ( n55923 , n55896 , n55922 );
buf ( n55924 , n55923 );
not ( n55925 , n55924 );
xor ( n55926 , n53667 , n53690 );
xor ( n55927 , n55926 , n53716 );
buf ( n55928 , n55927 );
buf ( n55929 , n55928 );
not ( n55930 , n55929 );
buf ( n55931 , n55930 );
buf ( n55932 , n55931 );
not ( n55933 , n55932 );
or ( n55934 , n55925 , n55933 );
not ( n55935 , n53532 );
not ( n55936 , n53571 );
and ( n55937 , n55935 , n55936 );
and ( n55938 , n53532 , n53571 );
nor ( n55939 , n55937 , n55938 );
not ( n55940 , n53559 );
and ( n55941 , n55939 , n55940 );
not ( n55942 , n55939 );
and ( n55943 , n55942 , n53559 );
nor ( n55944 , n55941 , n55943 );
buf ( n55945 , n55944 );
not ( n55946 , n55945 );
buf ( n55947 , n55946 );
buf ( n55948 , n55947 );
nand ( n55949 , n55934 , n55948 );
buf ( n55950 , n55949 );
buf ( n55951 , n55950 );
buf ( n55952 , n55923 );
not ( n55953 , n55952 );
buf ( n55954 , n55928 );
nand ( n55955 , n55953 , n55954 );
buf ( n55956 , n55955 );
buf ( n55957 , n55956 );
nand ( n55958 , n55951 , n55957 );
buf ( n55959 , n55958 );
buf ( n55960 , n55959 );
nand ( n55961 , n55833 , n55960 );
buf ( n55962 , n55961 );
buf ( n55963 , n55962 );
nand ( n55964 , n55830 , n55963 );
buf ( n55965 , n55964 );
buf ( n55966 , n55965 );
not ( n55967 , n55966 );
xor ( n55968 , n53794 , n53936 );
xor ( n55969 , n55968 , n55360 );
buf ( n55970 , n55969 );
buf ( n55971 , n55970 );
not ( n55972 , n55971 );
or ( n55973 , n55967 , n55972 );
buf ( n55974 , n55970 );
buf ( n55975 , n55965 );
or ( n55976 , n55974 , n55975 );
not ( n55977 , n55428 );
not ( n55978 , n55410 );
or ( n55979 , n55977 , n55978 );
or ( n55980 , n55428 , n55410 );
nand ( n55981 , n55979 , n55980 );
not ( n55982 , n55433 );
and ( n55983 , n55981 , n55982 );
not ( n55984 , n55981 );
and ( n55985 , n55984 , n55433 );
nor ( n55986 , n55983 , n55985 );
buf ( n55987 , n55986 );
not ( n55988 , n55987 );
buf ( n55989 , n55988 );
buf ( n55990 , n55989 );
not ( n55991 , n55990 );
xor ( n55992 , n53796 , n53912 );
xor ( n55993 , n55992 , n53932 );
not ( n55994 , n55993 );
not ( n55995 , n55994 );
buf ( n55996 , n55995 );
not ( n55997 , n55996 );
or ( n55998 , n55991 , n55997 );
buf ( n55999 , n55986 );
not ( n56000 , n55999 );
buf ( n56001 , n55994 );
not ( n56002 , n56001 );
or ( n56003 , n56000 , n56002 );
buf ( n56004 , C1 );
not ( n56005 , n53819 );
not ( n56006 , n53832 );
or ( n56007 , n56005 , n56006 );
buf ( n56008 , n53829 );
buf ( n56009 , n53822 );
nand ( n56010 , n56008 , n56009 );
buf ( n56011 , n56010 );
nand ( n56012 , n56007 , n56011 );
buf ( n56013 , n53908 );
not ( n56014 , n56013 );
buf ( n56015 , n56014 );
not ( n56016 , n56015 );
and ( n56017 , n56012 , n56016 );
not ( n56018 , n56012 );
and ( n56019 , n56018 , n56015 );
nor ( n56020 , n56017 , n56019 );
xor ( n56021 , n56004 , n56020 );
xor ( n56022 , n54119 , n55279 );
xor ( n56023 , n56022 , n55300 );
buf ( n56024 , n56023 );
buf ( n56025 , n52780 );
not ( n56026 , n56025 );
buf ( n56027 , n41718 );
not ( n56028 , n56027 );
or ( n56029 , n56026 , n56028 );
buf ( n56030 , n41715 );
buf ( n56031 , n52789 );
nand ( n56032 , n56030 , n56031 );
buf ( n56033 , n56032 );
buf ( n56034 , n56033 );
nand ( n56035 , n56029 , n56034 );
buf ( n56036 , n56035 );
buf ( n56037 , n56036 );
not ( n56038 , n56037 );
buf ( n56039 , n50374 );
not ( n56040 , n56039 );
or ( n56041 , n56038 , n56040 );
buf ( n56042 , n36643 );
buf ( n56043 , n53948 );
nand ( n56044 , n56042 , n56043 );
buf ( n56045 , n56044 );
buf ( n56046 , n56045 );
nand ( n56047 , n56041 , n56046 );
buf ( n56048 , n56047 );
xor ( n56049 , n56024 , n56048 );
xor ( n56050 , n53856 , n53874 );
xnor ( n56051 , n56050 , n53904 );
and ( n56052 , n56049 , n56051 );
and ( n56053 , n56024 , n56048 );
or ( n56054 , n56052 , n56053 );
and ( n56055 , n56021 , n56054 );
and ( n56056 , n56004 , n56020 );
or ( n56057 , n56055 , n56056 );
buf ( n56058 , n56057 );
nand ( n56059 , n56003 , n56058 );
buf ( n56060 , n56059 );
buf ( n56061 , n56060 );
nand ( n56062 , n55998 , n56061 );
buf ( n56063 , n56062 );
buf ( n56064 , n56063 );
nand ( n56065 , n55976 , n56064 );
buf ( n56066 , n56065 );
buf ( n56067 , n56066 );
nand ( n56068 , n55973 , n56067 );
buf ( n56069 , n56068 );
buf ( n56070 , n56069 );
xor ( n56071 , n55795 , n56070 );
xor ( n56072 , n53480 , n53483 );
xor ( n56073 , n56072 , n53784 );
buf ( n56074 , n56073 );
buf ( n56075 , n56074 );
and ( n56076 , n56071 , n56075 );
and ( n56077 , n55795 , n56070 );
or ( n56078 , n56076 , n56077 );
buf ( n56079 , n56078 );
buf ( n56080 , n56079 );
not ( n56081 , n56080 );
or ( n56082 , n55605 , n56081 );
buf ( n56083 , n56079 );
not ( n56084 , n56083 );
buf ( n56085 , n56084 );
buf ( n56086 , n56085 );
not ( n56087 , n56086 );
buf ( n56088 , n55603 );
not ( n56089 , n56088 );
buf ( n56090 , n56089 );
buf ( n56091 , n56090 );
not ( n56092 , n56091 );
or ( n56093 , n56087 , n56092 );
xor ( n56094 , n55365 , n55451 );
xor ( n56095 , n56094 , n55463 );
buf ( n56096 , n56095 );
xor ( n56097 , n55391 , n55395 );
xor ( n56098 , n56097 , n55446 );
buf ( n56099 , n56098 );
not ( n56100 , n56099 );
buf ( n56101 , n53925 );
buf ( n56102 , n46246 );
and ( n56103 , n56101 , n56102 );
and ( n56104 , n38244 , n45747 );
not ( n56105 , n38244 );
and ( n56106 , n56105 , n45753 );
or ( n56107 , n56104 , n56106 );
buf ( n56108 , n56107 );
buf ( n56109 , n46225 );
and ( n56110 , n56108 , n56109 );
buf ( n56111 , n56110 );
buf ( n56112 , n56111 );
nor ( n56113 , n56103 , n56112 );
buf ( n56114 , n56113 );
buf ( n56115 , n56114 );
buf ( n56116 , n48671 );
not ( n56117 , n56116 );
buf ( n56118 , n53854 );
not ( n56119 , n56118 );
or ( n56120 , n56117 , n56119 );
not ( n56121 , n41821 );
not ( n56122 , n41660 );
or ( n56123 , n56121 , n56122 );
nand ( n56124 , n29325 , n48390 );
nand ( n56125 , n56123 , n56124 );
buf ( n56126 , n56125 );
buf ( n56127 , n50982 );
nand ( n56128 , n56126 , n56127 );
buf ( n56129 , n56128 );
buf ( n56130 , n56129 );
nand ( n56131 , n56120 , n56130 );
buf ( n56132 , n56131 );
buf ( n56133 , n56132 );
not ( n56134 , n36335 );
not ( n56135 , n56134 );
nand ( n56136 , n56135 , n36495 );
buf ( n56137 , n56136 );
buf ( n56138 , n12481 );
and ( n56139 , n56137 , n56138 );
not ( n56140 , n56134 );
not ( n56141 , n36492 );
or ( n56142 , n56140 , n56141 );
nand ( n56143 , n56142 , n38834 );
buf ( n56144 , n56143 );
nor ( n56145 , n56139 , n56144 );
buf ( n56146 , n56145 );
buf ( n56147 , n56146 );
xor ( n56148 , n56133 , n56147 );
buf ( n56149 , n43063 );
not ( n56150 , n56149 );
buf ( n56151 , n41778 );
not ( n56152 , n56151 );
or ( n56153 , n56150 , n56152 );
buf ( n56154 , n41769 );
buf ( n56155 , n43064 );
nand ( n56156 , n56154 , n56155 );
buf ( n56157 , n56156 );
buf ( n56158 , n56157 );
nand ( n56159 , n56153 , n56158 );
buf ( n56160 , n56159 );
buf ( n56161 , n56160 );
not ( n56162 , n56161 );
buf ( n56163 , n37400 );
not ( n56164 , n56163 );
or ( n56165 , n56162 , n56164 );
buf ( n56166 , n53865 );
buf ( n56167 , n37413 );
nand ( n56168 , n56166 , n56167 );
buf ( n56169 , n56168 );
buf ( n56170 , n56169 );
nand ( n56171 , n56165 , n56170 );
buf ( n56172 , n56171 );
buf ( n56173 , n56172 );
and ( n56174 , n56148 , n56173 );
and ( n56175 , n56133 , n56147 );
or ( n56176 , n56174 , n56175 );
buf ( n56177 , n56176 );
not ( n56178 , n56177 );
buf ( n56179 , n55659 );
not ( n56180 , n56179 );
buf ( n56181 , n42312 );
not ( n56182 , n56181 );
and ( n56183 , n56180 , n56182 );
buf ( n56184 , n42263 );
not ( n56185 , n56184 );
buf ( n56186 , n39205 );
not ( n56187 , n56186 );
or ( n56188 , n56185 , n56187 );
buf ( n56189 , n37641 );
buf ( n56190 , n42263 );
or ( n56191 , n56189 , n56190 );
buf ( n56192 , n56191 );
buf ( n56193 , n56192 );
nand ( n56194 , n56188 , n56193 );
buf ( n56195 , n56194 );
buf ( n56196 , n56195 );
buf ( n56197 , n42252 );
and ( n56198 , n56196 , n56197 );
nor ( n56199 , n56183 , n56198 );
buf ( n56200 , n56199 );
buf ( n56201 , n48323 );
not ( n56202 , n56201 );
buf ( n56203 , n49425 );
not ( n56204 , n56203 );
or ( n56205 , n56202 , n56204 );
buf ( n56206 , n39136 );
buf ( n56207 , n48320 );
nand ( n56208 , n56206 , n56207 );
buf ( n56209 , n56208 );
buf ( n56210 , n56209 );
nand ( n56211 , n56205 , n56210 );
buf ( n56212 , n56211 );
buf ( n56213 , n56212 );
not ( n56214 , n56213 );
buf ( n56215 , n36976 );
not ( n56216 , n56215 );
or ( n56217 , n56214 , n56216 );
buf ( n56218 , n44676 );
buf ( n56219 , n55339 );
nand ( n56220 , n56218 , n56219 );
buf ( n56221 , n56220 );
buf ( n56222 , n56221 );
nand ( n56223 , n56217 , n56222 );
buf ( n56224 , n56223 );
not ( n56225 , n56224 );
nand ( n56226 , n56200 , n56225 );
not ( n56227 , n56226 );
or ( n56228 , n56178 , n56227 );
buf ( n56229 , n56224 );
buf ( n56230 , n56200 );
not ( n56231 , n56230 );
buf ( n56232 , n56231 );
buf ( n56233 , n56232 );
nand ( n56234 , n56229 , n56233 );
buf ( n56235 , n56234 );
nand ( n56236 , n56228 , n56235 );
not ( n56237 , n56236 );
buf ( n56238 , n56237 );
and ( n56239 , n56115 , n56238 );
buf ( n56240 , n56239 );
buf ( n56241 , n56240 );
xor ( n56242 , n55305 , n55330 );
xor ( n56243 , n56242 , n55353 );
buf ( n56244 , n56243 );
buf ( n56245 , n56244 );
not ( n56246 , n56245 );
buf ( n56247 , n56246 );
buf ( n56248 , n56247 );
or ( n56249 , n56241 , n56248 );
buf ( n56250 , n56237 );
buf ( n56251 , n56114 );
or ( n56252 , n56250 , n56251 );
buf ( n56253 , n56252 );
buf ( n56254 , n56253 );
nand ( n56255 , n56249 , n56254 );
buf ( n56256 , n56255 );
buf ( n56257 , n56256 );
xor ( n56258 , n55548 , n55550 );
xor ( n56259 , n56258 , n55576 );
buf ( n56260 , n56259 );
buf ( n56261 , n56260 );
xor ( n56262 , n56257 , n56261 );
xor ( n56263 , n54088 , n54089 );
buf ( n56264 , n56263 );
xor ( n56265 , n54086 , n56264 );
buf ( n56266 , n56265 );
buf ( n56267 , n45916 );
not ( n56268 , n56267 );
buf ( n56269 , n41611 );
not ( n56270 , n56269 );
and ( n56271 , n56268 , n56270 );
buf ( n56272 , n45916 );
buf ( n56273 , n41611 );
and ( n56274 , n56272 , n56273 );
nor ( n56275 , n56271 , n56274 );
buf ( n56276 , n56275 );
buf ( n56277 , n56276 );
not ( n56278 , n56277 );
buf ( n56279 , n41599 );
not ( n56280 , n56279 );
and ( n56281 , n56278 , n56280 );
buf ( n56282 , n55647 );
buf ( n56283 , n41574 );
and ( n56284 , n56282 , n56283 );
nor ( n56285 , n56281 , n56284 );
buf ( n56286 , n56285 );
buf ( n56287 , n56286 );
not ( n56288 , n56287 );
not ( n56289 , n52093 );
buf ( n56290 , n56289 );
not ( n56291 , n56290 );
buf ( n56292 , n36500 );
not ( n56293 , n56292 );
or ( n56294 , n56291 , n56293 );
buf ( n56295 , n43265 );
buf ( n56296 , n52094 );
nand ( n56297 , n56295 , n56296 );
buf ( n56298 , n56297 );
buf ( n56299 , n56298 );
nand ( n56300 , n56294 , n56299 );
buf ( n56301 , n56300 );
buf ( n56302 , n56301 );
not ( n56303 , n56302 );
buf ( n56304 , n46340 );
not ( n56305 , n56304 );
or ( n56306 , n56303 , n56305 );
buf ( n56307 , n55912 );
buf ( n56308 , n42527 );
nand ( n56309 , n56307 , n56308 );
buf ( n56310 , n56309 );
buf ( n56311 , n56310 );
nand ( n56312 , n56306 , n56311 );
buf ( n56313 , n56312 );
buf ( n56314 , n56313 );
not ( n56315 , n56314 );
buf ( n56316 , n56315 );
not ( n56317 , n56316 );
not ( n56318 , n42854 );
not ( n56319 , n56318 );
not ( n56320 , n55853 );
not ( n56321 , n56320 );
or ( n56322 , n56319 , n56321 );
buf ( n56323 , n12481 );
not ( n56324 , n56323 );
buf ( n56325 , n56324 );
nand ( n56326 , C1 , n42854 );
nand ( n56327 , n56322 , n56326 );
not ( n56328 , n56327 );
and ( n56329 , n56317 , n56328 );
buf ( n56330 , n56316 );
buf ( n56331 , n56327 );
nand ( n56332 , n56330 , n56331 );
buf ( n56333 , n56332 );
buf ( n56334 , n48172 );
not ( n56335 , n56334 );
buf ( n56336 , n51804 );
not ( n56337 , n56336 );
or ( n56338 , n56335 , n56337 );
buf ( n56339 , n25159 );
buf ( n56340 , n28368 );
not ( n56341 , n56340 );
buf ( n56342 , n56341 );
buf ( n56343 , n56342 );
nand ( n56344 , n56339 , n56343 );
buf ( n56345 , n56344 );
buf ( n56346 , n56345 );
nand ( n56347 , n56338 , n56346 );
buf ( n56348 , n56347 );
buf ( n56349 , n56348 );
not ( n56350 , n56349 );
buf ( n56351 , n50128 );
not ( n56352 , n56351 );
or ( n56353 , n56350 , n56352 );
buf ( n56354 , n54133 );
not ( n56355 , n56354 );
buf ( n56356 , n42564 );
nand ( n56357 , n56355 , n56356 );
buf ( n56358 , n56357 );
buf ( n56359 , n56358 );
nand ( n56360 , n56353 , n56359 );
buf ( n56361 , n56360 );
buf ( n56362 , n56361 );
buf ( n56363 , n42504 );
not ( n56364 , n56363 );
buf ( n56365 , n42471 );
not ( n56366 , n56365 );
or ( n56367 , n56364 , n56366 );
buf ( n56368 , n42468 );
buf ( n56369 , n41721 );
nand ( n56370 , n56368 , n56369 );
buf ( n56371 , n56370 );
buf ( n56372 , n56371 );
nand ( n56373 , n56367 , n56372 );
buf ( n56374 , n56373 );
buf ( n56375 , n56374 );
not ( n56376 , n56375 );
buf ( n56377 , n47014 );
not ( n56378 , n56377 );
or ( n56379 , n56376 , n56378 );
buf ( n56380 , n38973 );
not ( n56381 , n56380 );
buf ( n56382 , n54040 );
nand ( n56383 , n56381 , n56382 );
buf ( n56384 , n56383 );
buf ( n56385 , n56384 );
nand ( n56386 , n56379 , n56385 );
buf ( n56387 , n56386 );
buf ( n56388 , n56387 );
xor ( n56389 , n56362 , n56388 );
buf ( n56390 , n50982 );
not ( n56391 , n56390 );
not ( n56392 , n41912 );
not ( n56393 , n41660 );
or ( n56394 , n56392 , n56393 );
nand ( n56395 , n47001 , n48390 );
nand ( n56396 , n56394 , n56395 );
buf ( n56397 , n56396 );
not ( n56398 , n56397 );
or ( n56399 , n56391 , n56398 );
buf ( n56400 , n56125 );
buf ( n56401 , n48671 );
nand ( n56402 , n56400 , n56401 );
buf ( n56403 , n56402 );
buf ( n56404 , n56403 );
nand ( n56405 , n56399 , n56404 );
buf ( n56406 , n56405 );
buf ( n56407 , n56406 );
and ( n56408 , n56389 , n56407 );
and ( n56409 , n56362 , n56388 );
or ( n56410 , n56408 , n56409 );
buf ( n56411 , n56410 );
and ( n56412 , n56333 , n56411 );
nor ( n56413 , n56329 , n56412 );
buf ( n56414 , n56413 );
not ( n56415 , n56414 );
or ( n56416 , n56288 , n56415 );
buf ( n56417 , n46117 );
not ( n56418 , n56417 );
buf ( n56419 , n44381 );
not ( n56420 , n56419 );
or ( n56421 , n56418 , n56420 );
buf ( n56422 , n41889 );
buf ( n56423 , n46126 );
nand ( n56424 , n56422 , n56423 );
buf ( n56425 , n56424 );
buf ( n56426 , n56425 );
nand ( n56427 , n56421 , n56426 );
buf ( n56428 , n56427 );
buf ( n56429 , n56428 );
not ( n56430 , n56429 );
buf ( n56431 , n41862 );
not ( n56432 , n56431 );
or ( n56433 , n56430 , n56432 );
nand ( n56434 , n45617 , n53988 );
buf ( n56435 , n56434 );
nand ( n56436 , n56433 , n56435 );
buf ( n56437 , n56436 );
not ( n56438 , n56437 );
and ( n56439 , n42847 , n41976 );
not ( n56440 , n42847 );
and ( n56441 , n56440 , n37472 );
nor ( n56442 , n56439 , n56441 );
buf ( n56443 , n56442 );
not ( n56444 , n56443 );
buf ( n56445 , n50671 );
not ( n56446 , n56445 );
or ( n56447 , n56444 , n56446 );
buf ( n56448 , n53970 );
buf ( n56449 , n41852 );
nand ( n56450 , n56448 , n56449 );
buf ( n56451 , n56450 );
buf ( n56452 , n56451 );
nand ( n56453 , n56447 , n56452 );
buf ( n56454 , n56453 );
not ( n56455 , n56454 );
or ( n56456 , n56438 , n56455 );
buf ( n56457 , n56437 );
buf ( n56458 , n56454 );
nor ( n56459 , n56457 , n56458 );
buf ( n56460 , n56459 );
buf ( n56461 , n42339 );
not ( n56462 , n56461 );
buf ( n56463 , n53897 );
not ( n56464 , n56463 );
or ( n56465 , n56462 , n56464 );
buf ( n56466 , n42343 );
not ( n56467 , n56466 );
buf ( n56468 , n41763 );
not ( n56469 , n56468 );
or ( n56470 , n56467 , n56469 );
buf ( n56471 , n41762 );
buf ( n56472 , n46855 );
nand ( n56473 , n56471 , n56472 );
buf ( n56474 , n56473 );
buf ( n56475 , n56474 );
nand ( n56476 , n56470 , n56475 );
buf ( n56477 , n56476 );
buf ( n56478 , n56477 );
buf ( n56479 , n42378 );
nand ( n56480 , n56478 , n56479 );
buf ( n56481 , n56480 );
buf ( n56482 , n56481 );
nand ( n56483 , n56465 , n56482 );
buf ( n56484 , n56483 );
buf ( n56485 , n56484 );
not ( n56486 , n56485 );
buf ( n56487 , n56486 );
or ( n56488 , n56460 , n56487 );
nand ( n56489 , n56456 , n56488 );
buf ( n56490 , n56489 );
nand ( n56491 , n56416 , n56490 );
buf ( n56492 , n56491 );
buf ( n56493 , n56492 );
buf ( n56494 , n56286 );
not ( n56495 , n56494 );
buf ( n56496 , n56413 );
not ( n56497 , n56496 );
buf ( n56498 , n56497 );
buf ( n56499 , n56498 );
nand ( n56500 , n56495 , n56499 );
buf ( n56501 , n56500 );
buf ( n56502 , n56501 );
nand ( n56503 , n56493 , n56502 );
buf ( n56504 , n56503 );
buf ( n56505 , n56504 );
xor ( n56506 , n56266 , n56505 );
buf ( n56507 , n54026 );
buf ( n56508 , n54074 );
xor ( n56509 , n56507 , n56508 );
buf ( n56510 , n54052 );
xnor ( n56511 , n56509 , n56510 );
buf ( n56512 , n56511 );
buf ( n56513 , n56512 );
buf ( n56514 , n42668 );
not ( n56515 , n56514 );
buf ( n56516 , n55692 );
not ( n56517 , n56516 );
or ( n56518 , n56515 , n56517 );
and ( n56519 , n29269 , n25227 );
not ( n56520 , n29269 );
and ( n56521 , n56520 , n25226 );
or ( n56522 , n56519 , n56521 );
buf ( n56523 , n56522 );
buf ( n56524 , n42712 );
nand ( n56525 , n56523 , n56524 );
buf ( n56526 , n56525 );
buf ( n56527 , n56526 );
nand ( n56528 , n56518 , n56527 );
buf ( n56529 , n56528 );
buf ( n56530 , n56529 );
not ( n56531 , n56530 );
buf ( n56532 , n56531 );
buf ( n56533 , n56532 );
nand ( n56534 , n56513 , n56533 );
buf ( n56535 , n56534 );
buf ( n56536 , n56535 );
not ( n56537 , n56536 );
xor ( n56538 , n55161 , n55191 );
xor ( n56539 , n56538 , n55264 );
buf ( n56540 , n56539 );
buf ( n56541 , n56540 );
not ( n56542 , n56541 );
buf ( n56543 , n29754 );
not ( n56544 , n56543 );
buf ( n56545 , n56544 );
buf ( n56546 , n56545 );
not ( n56547 , n56546 );
buf ( n56548 , n56547 );
buf ( n56549 , n56548 );
not ( n56550 , n56549 );
buf ( n56551 , n52670 );
not ( n56552 , n56551 );
or ( n56553 , n56550 , n56552 );
buf ( n56554 , n29754 );
not ( n56555 , n56554 );
buf ( n56556 , n25159 );
nand ( n56557 , n56555 , n56556 );
buf ( n56558 , n56557 );
buf ( n56559 , n56558 );
nand ( n56560 , n56553 , n56559 );
buf ( n56561 , n56560 );
buf ( n56562 , n56561 );
not ( n56563 , n56562 );
buf ( n56564 , n50128 );
not ( n56565 , n56564 );
or ( n56566 , n56563 , n56565 );
not ( n56567 , n42563 );
buf ( n56568 , n56567 );
buf ( n56569 , n56348 );
nand ( n56570 , n56568 , n56569 );
buf ( n56571 , n56570 );
buf ( n56572 , n56571 );
nand ( n56573 , n56566 , n56572 );
buf ( n56574 , n56573 );
buf ( n56575 , n56574 );
not ( n56576 , n56575 );
buf ( n56577 , n56576 );
buf ( n56578 , n56577 );
not ( n56579 , n56578 );
or ( n56580 , n56542 , n56579 );
nand ( n56581 , n54269 , n55241 );
xnor ( n56582 , n56581 , n55144 );
buf ( n56583 , n56582 );
not ( n56584 , n56583 );
buf ( n56585 , n56584 );
buf ( n56586 , n56585 );
buf ( n56587 , n55132 );
not ( n56588 , n56587 );
buf ( n56589 , n56588 );
buf ( n56590 , n56589 );
or ( n56591 , n56586 , n56590 );
buf ( n56592 , n55249 );
not ( n56593 , n56592 );
buf ( n56594 , n56593 );
buf ( n56595 , n56594 );
buf ( n56596 , n55156 );
not ( n56597 , n56596 );
buf ( n56598 , n56597 );
buf ( n56599 , n56598 );
or ( n56600 , n56595 , n56599 );
nand ( n56601 , n56591 , n56600 );
buf ( n56602 , n56601 );
not ( n56603 , n5221 );
not ( n56604 , n5240 );
or ( n56605 , n56603 , n56604 );
nand ( n56606 , n56605 , n5245 );
not ( n56607 , n56606 );
not ( n56608 , n7201 );
or ( n56609 , n56607 , n56608 );
or ( n56610 , n7201 , n56606 );
nand ( n56611 , n56609 , n56610 );
buf ( n56612 , n56611 );
not ( n56613 , n56612 );
buf ( n56614 , n56613 );
buf ( n56615 , n56614 );
buf ( n56616 , n16469 );
buf ( n56617 , n7201 );
and ( n56618 , n56616 , n56617 );
buf ( n56619 , n16472 );
buf ( n56620 , n7124 );
and ( n56621 , n56619 , n56620 );
nor ( n56622 , n56618 , n56621 );
buf ( n56623 , n56622 );
buf ( n56624 , n56623 );
nand ( n56625 , n56615 , n56624 );
buf ( n56626 , n56625 );
buf ( n56627 , n56626 );
not ( n56628 , n56627 );
buf ( n56629 , n56628 );
buf ( n56630 , n56629 );
not ( n56631 , n16469 );
buf ( n56632 , n56631 );
nand ( n56633 , n56630 , n56632 );
buf ( n56634 , n56633 );
buf ( n56635 , n56634 );
not ( n56636 , n56635 );
buf ( n56637 , n56611 );
not ( n56638 , n56637 );
buf ( n56639 , n56638 );
buf ( n56640 , n56639 );
not ( n56641 , n56631 );
buf ( n56642 , n56641 );
nor ( n56643 , n56640 , n56642 );
buf ( n56644 , n56643 );
buf ( n56645 , n56644 );
nor ( n56646 , n56636 , n56645 );
buf ( n56647 , n56646 );
xor ( n56648 , n56602 , n56647 );
buf ( n56649 , n55113 );
buf ( n56650 , n55201 );
not ( n56651 , n56650 );
buf ( n56652 , n56651 );
buf ( n56653 , n56652 );
and ( n56654 , n56649 , n56653 );
not ( n56655 , n55113 );
buf ( n56656 , n56655 );
buf ( n56657 , n55201 );
and ( n56658 , n56656 , n56657 );
nor ( n56659 , n56654 , n56658 );
buf ( n56660 , n56659 );
buf ( n56661 , n56660 );
buf ( n56662 , n55180 );
not ( n56663 , n56662 );
buf ( n56664 , n56663 );
buf ( n56665 , n56664 );
or ( n56666 , n56661 , n56665 );
buf ( n56667 , n55212 );
buf ( n56668 , n55166 );
not ( n56669 , n56668 );
buf ( n56670 , n56669 );
buf ( n56671 , n56670 );
not ( n56672 , n56671 );
buf ( n56673 , n56672 );
buf ( n56674 , n56673 );
or ( n56675 , n56667 , n56674 );
nand ( n56676 , n56666 , n56675 );
buf ( n56677 , n56676 );
and ( n56678 , n56648 , n56677 );
and ( n56679 , n56602 , n56647 );
or ( n56680 , n56678 , n56679 );
buf ( n56681 , n56680 );
buf ( n56682 , n55221 );
buf ( n56683 , n55257 );
or ( n56684 , n56682 , n56683 );
buf ( n56685 , n55260 );
nand ( n56686 , n56684 , n56685 );
buf ( n56687 , n56686 );
buf ( n56688 , n56687 );
xor ( n56689 , n56681 , n56688 );
buf ( n56690 , n56641 );
buf ( n56691 , n55152 );
and ( n56692 , n56690 , n56691 );
not ( n56693 , n56690 );
buf ( n56694 , n55205 );
and ( n56695 , n56693 , n56694 );
nor ( n56696 , n56692 , n56695 );
buf ( n56697 , n56696 );
buf ( n56698 , n56697 );
not ( n56699 , n56698 );
buf ( n56700 , n56699 );
buf ( n56701 , n56700 );
buf ( n56702 , n56629 );
and ( n56703 , n56701 , n56702 );
buf ( n56704 , n56644 );
nor ( n56705 , n56703 , n56704 );
buf ( n56706 , n56705 );
buf ( n56707 , n56706 );
and ( n56708 , n54469 , n54235 , n54288 );
not ( n56709 , n56708 );
not ( n56710 , n55230 );
or ( n56711 , n56709 , n56710 );
and ( n56712 , n55236 , n54288 );
nor ( n56713 , n56712 , n55095 );
nand ( n56714 , n56711 , n56713 );
not ( n56715 , n55099 );
nand ( n56716 , n56715 , n54258 );
nor ( n56717 , n56714 , n56716 );
not ( n56718 , n56717 );
nand ( n56719 , n56714 , n56716 );
nand ( n56720 , n56718 , n56719 );
buf ( n56721 , n56720 );
buf ( n56722 , n55132 );
and ( n56723 , n56721 , n56722 );
buf ( n56724 , n56582 );
buf ( n56725 , n55156 );
and ( n56726 , n56724 , n56725 );
nor ( n56727 , n56723 , n56726 );
buf ( n56728 , n56727 );
buf ( n56729 , n56728 );
nand ( n56730 , n56707 , n56729 );
buf ( n56731 , n56730 );
xor ( n56732 , n56602 , n56647 );
xor ( n56733 , n56732 , n56677 );
and ( n56734 , n56731 , n56733 );
buf ( n56735 , n56706 );
buf ( n56736 , n56728 );
or ( n56737 , n56735 , n56736 );
buf ( n56738 , n56731 );
nand ( n56739 , n56737 , n56738 );
buf ( n56740 , n56739 );
buf ( n56741 , n56740 );
buf ( n56742 , n56652 );
buf ( n56743 , n55249 );
and ( n56744 , n56742 , n56743 );
not ( n56745 , n56742 );
buf ( n56746 , n56594 );
and ( n56747 , n56745 , n56746 );
nor ( n56748 , n56744 , n56747 );
buf ( n56749 , n56748 );
buf ( n56750 , n56749 );
buf ( n56751 , n56664 );
or ( n56752 , n56750 , n56751 );
buf ( n56753 , n56660 );
buf ( n56754 , n56673 );
or ( n56755 , n56753 , n56754 );
nand ( n56756 , n56752 , n56755 );
buf ( n56757 , n56756 );
buf ( n56758 , n56757 );
xor ( n56759 , n56741 , n56758 );
buf ( n56760 , n55113 );
buf ( n56761 , n56641 );
and ( n56762 , n56760 , n56761 );
buf ( n56763 , n56655 );
buf ( n56764 , n56631 );
and ( n56765 , n56763 , n56764 );
nor ( n56766 , n56762 , n56765 );
buf ( n56767 , n56766 );
buf ( n56768 , n56767 );
buf ( n56769 , n56626 );
or ( n56770 , n56768 , n56769 );
buf ( n56771 , n56697 );
buf ( n56772 , n56639 );
or ( n56773 , n56771 , n56772 );
nand ( n56774 , n56770 , n56773 );
buf ( n56775 , n56774 );
buf ( n56776 , n56775 );
not ( n56777 , n56606 );
not ( n56778 , n56777 );
not ( n56779 , n6918 );
or ( n56780 , n56778 , n56779 );
buf ( n56781 , n3264 );
or ( n56782 , n56781 , n56777 );
nand ( n56783 , n56780 , n56782 );
buf ( n56784 , n56783 );
buf ( n56785 , n56781 );
buf ( n56786 , n6908 );
buf ( n56787 , n56786 );
not ( n56788 , n56787 );
buf ( n56789 , n56788 );
buf ( n56790 , n56789 );
and ( n56791 , n56785 , n56790 );
not ( n56792 , n56785 );
buf ( n56793 , n56786 );
and ( n56794 , n56792 , n56793 );
nor ( n56795 , n56791 , n56794 );
buf ( n56796 , n56795 );
buf ( n56797 , n56796 );
nand ( n56798 , n56784 , n56797 );
buf ( n56799 , n56798 );
not ( n56800 , n56799 );
buf ( n56801 , n56800 );
buf ( n56802 , n56777 );
not ( n56803 , n56802 );
buf ( n56804 , n56803 );
buf ( n56805 , n56804 );
nand ( n56806 , n56801 , n56805 );
buf ( n56807 , n56806 );
buf ( n56808 , n56807 );
buf ( n56809 , n56796 );
not ( n56810 , n56809 );
buf ( n56811 , n56810 );
buf ( n56812 , n56811 );
buf ( n56813 , n56804 );
nand ( n56814 , n56812 , n56813 );
buf ( n56815 , n56814 );
buf ( n56816 , n56815 );
and ( n56817 , n56808 , n56816 );
buf ( n56818 , n56817 );
buf ( n56819 , n56818 );
xor ( n56820 , n56776 , n56819 );
buf ( n56821 , n56582 );
buf ( n56822 , n56652 );
and ( n56823 , n56821 , n56822 );
buf ( n56824 , n56585 );
buf ( n56825 , n55201 );
and ( n56826 , n56824 , n56825 );
nor ( n56827 , n56823 , n56826 );
buf ( n56828 , n56827 );
buf ( n56829 , n56828 );
buf ( n56830 , n56664 );
or ( n56831 , n56829 , n56830 );
buf ( n56832 , n56749 );
buf ( n56833 , n56673 );
or ( n56834 , n56832 , n56833 );
nand ( n56835 , n56831 , n56834 );
buf ( n56836 , n56835 );
buf ( n56837 , n56836 );
and ( n56838 , n56820 , n56837 );
and ( n56839 , n56776 , n56819 );
or ( n56840 , n56838 , n56839 );
buf ( n56841 , n56840 );
buf ( n56842 , n56841 );
and ( n56843 , n56759 , n56842 );
and ( n56844 , n56741 , n56758 );
or ( n56845 , n56843 , n56844 );
buf ( n56846 , n56845 );
xor ( n56847 , n56602 , n56647 );
xor ( n56848 , n56847 , n56677 );
and ( n56849 , n56846 , n56848 );
and ( n56850 , n56731 , n56846 );
or ( n56851 , n56734 , n56849 , n56850 );
buf ( n56852 , n56851 );
and ( n56853 , n56689 , n56852 );
and ( n56854 , n56681 , n56688 );
or ( n56855 , n56853 , n56854 );
buf ( n56856 , n56855 );
buf ( n56857 , n56856 );
nand ( n56858 , n56580 , n56857 );
buf ( n56859 , n56858 );
buf ( n56860 , n56859 );
buf ( n56861 , n56540 );
not ( n56862 , n56861 );
buf ( n56863 , n56574 );
nand ( n56864 , n56862 , n56863 );
buf ( n56865 , n56864 );
buf ( n56866 , n56865 );
nand ( n56867 , n56860 , n56866 );
buf ( n56868 , n56867 );
buf ( n56869 , n56868 );
buf ( n56870 , n42378 );
not ( n56871 , n56870 );
buf ( n56872 , n42343 );
not ( n56873 , n56872 );
buf ( n56874 , n41835 );
not ( n56875 , n56874 );
or ( n56876 , n56873 , n56875 );
buf ( n56877 , n28305 );
buf ( n56878 , n46855 );
nand ( n56879 , n56877 , n56878 );
buf ( n56880 , n56879 );
buf ( n56881 , n56880 );
nand ( n56882 , n56876 , n56881 );
buf ( n56883 , n56882 );
buf ( n56884 , n56883 );
not ( n56885 , n56884 );
or ( n56886 , n56871 , n56885 );
buf ( n56887 , n56477 );
buf ( n56888 , n42339 );
nand ( n56889 , n56887 , n56888 );
buf ( n56890 , n56889 );
buf ( n56891 , n56890 );
nand ( n56892 , n56886 , n56891 );
buf ( n56893 , n56892 );
buf ( n56894 , n56893 );
xor ( n56895 , n56869 , n56894 );
buf ( n56896 , n41993 );
not ( n56897 , n56896 );
buf ( n56898 , n44054 );
not ( n56899 , n56898 );
or ( n56900 , n56897 , n56899 );
buf ( n56901 , n42411 );
buf ( n56902 , n43966 );
nand ( n56903 , n56901 , n56902 );
buf ( n56904 , n56903 );
buf ( n56905 , n56904 );
nand ( n56906 , n56900 , n56905 );
buf ( n56907 , n56906 );
buf ( n56908 , n56907 );
not ( n56909 , n56908 );
buf ( n56910 , n56909 );
or ( n56911 , n56910 , n44039 );
nand ( n56912 , n38382 , n55712 );
nand ( n56913 , n56911 , n56912 );
buf ( n56914 , n56913 );
and ( n56915 , n56895 , n56914 );
and ( n56916 , n56869 , n56894 );
or ( n56917 , n56915 , n56916 );
buf ( n56918 , n56917 );
buf ( n56919 , n56918 );
not ( n56920 , n56919 );
or ( n56921 , n56537 , n56920 );
buf ( n56922 , n56512 );
not ( n56923 , n56922 );
buf ( n56924 , n56923 );
buf ( n56925 , n56924 );
buf ( n56926 , n56529 );
nand ( n56927 , n56925 , n56926 );
buf ( n56928 , n56927 );
buf ( n56929 , n56928 );
nand ( n56930 , n56921 , n56929 );
buf ( n56931 , n56930 );
buf ( n56932 , n56931 );
buf ( n56933 , n44708 );
not ( n56934 , n56933 );
buf ( n56935 , n44533 );
not ( n56936 , n56935 );
buf ( n56937 , n37689 );
not ( n56938 , n56937 );
or ( n56939 , n56936 , n56938 );
buf ( n56940 , n43625 );
buf ( n56941 , n44530 );
nand ( n56942 , n56940 , n56941 );
buf ( n56943 , n56942 );
buf ( n56944 , n56943 );
nand ( n56945 , n56939 , n56944 );
buf ( n56946 , n56945 );
buf ( n56947 , n56946 );
not ( n56948 , n56947 );
or ( n56949 , n56934 , n56948 );
buf ( n56950 , n44533 );
not ( n56951 , n56950 );
buf ( n56952 , n43224 );
not ( n56953 , n56952 );
or ( n56954 , n56951 , n56953 );
buf ( n56955 , n37294 );
buf ( n56956 , n44530 );
nand ( n56957 , n56955 , n56956 );
buf ( n56958 , n56957 );
buf ( n56959 , n56958 );
nand ( n56960 , n56954 , n56959 );
buf ( n56961 , n56960 );
buf ( n56962 , n56961 );
buf ( n56963 , n44496 );
nand ( n56964 , n56962 , n56963 );
buf ( n56965 , n56964 );
buf ( n56966 , n56965 );
nand ( n56967 , n56949 , n56966 );
buf ( n56968 , n56967 );
buf ( n56969 , n56968 );
xor ( n56970 , n56932 , n56969 );
buf ( n56971 , n54080 );
buf ( n56972 , n53982 );
xor ( n56973 , n56971 , n56972 );
buf ( n56974 , n53996 );
xor ( n56975 , n56973 , n56974 );
buf ( n56976 , n56975 );
buf ( n56977 , n56976 );
and ( n56978 , n56970 , n56977 );
and ( n56979 , n56932 , n56969 );
or ( n56980 , n56978 , n56979 );
buf ( n56981 , n56980 );
buf ( n56982 , n56981 );
and ( n56983 , n56506 , n56982 );
and ( n56984 , n56266 , n56505 );
or ( n56985 , n56983 , n56984 );
buf ( n56986 , n56985 );
buf ( n56987 , n56986 );
and ( n56988 , n56262 , n56987 );
and ( n56989 , n56257 , n56261 );
or ( n56990 , n56988 , n56989 );
buf ( n56991 , n56990 );
not ( n56992 , n56991 );
or ( n56993 , n56100 , n56992 );
or ( n56994 , n56099 , n56991 );
xor ( n56995 , n55523 , n55580 );
xor ( n56996 , n56995 , n55584 );
buf ( n56997 , n56996 );
nand ( n56998 , n56994 , n56997 );
nand ( n56999 , n56993 , n56998 );
xor ( n57000 , n56096 , n56999 );
buf ( n57001 , n55518 );
buf ( n57002 , n55588 );
xor ( n57003 , n57001 , n57002 );
buf ( n57004 , n55515 );
xor ( n57005 , n57003 , n57004 );
buf ( n57006 , n57005 );
and ( n57007 , n57000 , n57006 );
and ( n57008 , n56096 , n56999 );
or ( n57009 , n57007 , n57008 );
buf ( n57010 , n57009 );
nand ( n57011 , n56093 , n57010 );
buf ( n57012 , n57011 );
buf ( n57013 , n57012 );
nand ( n57014 , n56082 , n57013 );
buf ( n57015 , n57014 );
buf ( n57016 , n57015 );
not ( n57017 , n57016 );
buf ( n57018 , n57017 );
buf ( n57019 , n57018 );
xor ( n57020 , n55600 , n57019 );
xor ( n57021 , n55476 , n55491 );
xor ( n57022 , n57021 , n55495 );
buf ( n57023 , n57022 );
buf ( n57024 , n57023 );
and ( n57025 , n57020 , n57024 );
and ( n57026 , n55600 , n57019 );
or ( n57027 , n57025 , n57026 );
buf ( n57028 , n57027 );
nand ( n57029 , n55500 , n57028 );
buf ( n57030 , n57029 );
xor ( n57031 , n52866 , n53356 );
xor ( n57032 , n57031 , n53369 );
buf ( n57033 , n57032 );
not ( n57034 , n57033 );
xor ( n57035 , n53461 , n53472 );
and ( n57036 , n57035 , n55499 );
and ( n57037 , n53461 , n53472 );
or ( n57038 , n57036 , n57037 );
nand ( n57039 , n57034 , n57038 );
buf ( n57040 , n57039 );
and ( n57041 , n57030 , n57040 );
buf ( n57042 , n57041 );
buf ( n57043 , n57042 );
xor ( n57044 , n55504 , n55508 );
xor ( n57045 , n57044 , n55595 );
buf ( n57046 , n57045 );
buf ( n57047 , n57046 );
buf ( n57048 , C0 );
buf ( n57049 , n57048 );
buf ( n57050 , n44496 );
not ( n57051 , n57050 );
buf ( n57052 , n55537 );
not ( n57053 , n57052 );
or ( n57054 , n57051 , n57053 );
buf ( n57055 , n56961 );
buf ( n57056 , n44708 );
nand ( n57057 , n57055 , n57056 );
buf ( n57058 , n57057 );
buf ( n57059 , n57058 );
nand ( n57060 , n57054 , n57059 );
buf ( n57061 , n57060 );
buf ( n57062 , n57061 );
xor ( n57063 , n57049 , n57062 );
buf ( n57064 , n46912 );
not ( n57065 , n57064 );
buf ( n57066 , n55568 );
not ( n57067 , n57066 );
or ( n57068 , n57065 , n57067 );
buf ( n57069 , n46875 );
not ( n57070 , n57069 );
buf ( n57071 , n49804 );
not ( n57072 , n57071 );
buf ( n57073 , n57072 );
buf ( n57074 , n57073 );
not ( n57075 , n57074 );
or ( n57076 , n57070 , n57075 );
buf ( n57077 , n42929 );
buf ( n57078 , n46887 );
nand ( n57079 , n57077 , n57078 );
buf ( n57080 , n57079 );
buf ( n57081 , n57080 );
nand ( n57082 , n57076 , n57081 );
buf ( n57083 , n57082 );
buf ( n57084 , n57083 );
buf ( n57085 , n47331 );
nand ( n57086 , n57084 , n57085 );
buf ( n57087 , n57086 );
buf ( n57088 , n57087 );
nand ( n57089 , n57068 , n57088 );
buf ( n57090 , n57089 );
buf ( n57091 , n57090 );
and ( n57092 , n57063 , n57091 );
or ( n57093 , n57092 , C0 );
buf ( n57094 , n57093 );
buf ( n57095 , n57094 );
buf ( n57096 , n54092 );
buf ( n57097 , n54112 );
not ( n57098 , n57097 );
buf ( n57099 , n55357 );
not ( n57100 , n57099 );
buf ( n57101 , n57100 );
buf ( n57102 , n57101 );
not ( n57103 , n57102 );
or ( n57104 , n57098 , n57103 );
buf ( n57105 , n55357 );
buf ( n57106 , n54109 );
nand ( n57107 , n57105 , n57106 );
buf ( n57108 , n57107 );
buf ( n57109 , n57108 );
nand ( n57110 , n57104 , n57109 );
buf ( n57111 , n57110 );
xnor ( n57112 , n57096 , n57111 );
buf ( n57113 , n57112 );
xor ( n57114 , n57095 , n57113 );
and ( n57115 , n55627 , n55619 );
not ( n57116 , n55627 );
and ( n57117 , n57116 , n55620 );
nor ( n57118 , n57115 , n57117 );
xor ( n57119 , n57118 , n55780 );
buf ( n57120 , n57119 );
and ( n57121 , n57114 , n57120 );
and ( n57122 , n57095 , n57113 );
or ( n57123 , n57121 , n57122 );
buf ( n57124 , n57123 );
buf ( n57125 , n57124 );
xor ( n57126 , n55609 , n55785 );
xor ( n57127 , n57126 , n55790 );
buf ( n57128 , n57127 );
buf ( n57129 , n57128 );
xor ( n57130 , n57125 , n57129 );
not ( n57131 , n46912 );
not ( n57132 , n57083 );
or ( n57133 , n57131 , n57132 );
buf ( n57134 , n46875 );
not ( n57135 , n57134 );
buf ( n57136 , n38218 );
not ( n57137 , n57136 );
or ( n57138 , n57135 , n57137 );
buf ( n57139 , n47969 );
buf ( n57140 , n46887 );
nand ( n57141 , n57139 , n57140 );
buf ( n57142 , n57141 );
buf ( n57143 , n57142 );
nand ( n57144 , n57138 , n57143 );
buf ( n57145 , n57144 );
nand ( n57146 , n57145 , n47331 );
nand ( n57147 , n57133 , n57146 );
or ( n57148 , C0 , n57147 );
not ( n57149 , n56232 );
not ( n57150 , n56225 );
or ( n57151 , n57149 , n57150 );
nand ( n57152 , n56224 , n56200 );
nand ( n57153 , n57151 , n57152 );
and ( n57154 , n57153 , n56177 );
not ( n57155 , n57153 );
buf ( n57156 , n56177 );
not ( n57157 , n57156 );
buf ( n57158 , n57157 );
and ( n57159 , n57155 , n57158 );
nor ( n57160 , n57154 , n57159 );
nand ( n57161 , n57148 , n57160 );
nand ( n57162 , C1 , n57161 );
not ( n57163 , n57162 );
buf ( n57164 , n51488 );
not ( n57165 , n57164 );
buf ( n57166 , n48836 );
not ( n57167 , n57166 );
buf ( n57168 , n40067 );
not ( n57169 , n57168 );
or ( n57170 , n57167 , n57169 );
buf ( n57171 , n36427 );
buf ( n57172 , n48836 );
not ( n57173 , n57172 );
buf ( n57174 , n57173 );
buf ( n57175 , n57174 );
nand ( n57176 , n57171 , n57175 );
buf ( n57177 , n57176 );
buf ( n57178 , n57177 );
nand ( n57179 , n57170 , n57178 );
buf ( n57180 , n57179 );
buf ( n57181 , n57180 );
not ( n57182 , n57181 );
or ( n57183 , n57165 , n57182 );
buf ( n57184 , n55617 );
buf ( n57185 , n52456 );
nand ( n57186 , n57184 , n57185 );
buf ( n57187 , n57186 );
buf ( n57188 , n57187 );
nand ( n57189 , n57183 , n57188 );
buf ( n57190 , n57189 );
buf ( n57191 , n57190 );
not ( n57192 , n57191 );
buf ( n57193 , n57192 );
nand ( n57194 , n57163 , n57193 );
not ( n57195 , n57194 );
buf ( n57196 , n55947 );
not ( n57197 , n57196 );
buf ( n57198 , n55931 );
not ( n57199 , n57198 );
or ( n57200 , n57197 , n57199 );
buf ( n57201 , n55928 );
buf ( n57202 , n55944 );
nand ( n57203 , n57201 , n57202 );
buf ( n57204 , n57203 );
buf ( n57205 , n57204 );
nand ( n57206 , n57200 , n57205 );
buf ( n57207 , n57206 );
not ( n57208 , n55923 );
and ( n57209 , n57207 , n57208 );
not ( n57210 , n57207 );
not ( n57211 , n57208 );
and ( n57212 , n57210 , n57211 );
nor ( n57213 , n57209 , n57212 );
not ( n57214 , n57213 );
or ( n57215 , n57195 , n57214 );
buf ( n57216 , n57193 );
not ( n57217 , n57216 );
buf ( n57218 , n57162 );
nand ( n57219 , n57217 , n57218 );
buf ( n57220 , n57219 );
nand ( n57221 , n57215 , n57220 );
buf ( n57222 , n57221 );
not ( n57223 , n57222 );
buf ( n57224 , n55959 );
buf ( n57225 , n55798 );
xor ( n57226 , n57224 , n57225 );
buf ( n57227 , n55827 );
xnor ( n57228 , n57226 , n57227 );
buf ( n57229 , n57228 );
not ( n57230 , n57229 );
buf ( n57231 , n57230 );
not ( n57232 , n57231 );
or ( n57233 , n57223 , n57232 );
buf ( n57234 , n57229 );
not ( n57235 , n57234 );
buf ( n57236 , n57221 );
not ( n57237 , n57236 );
buf ( n57238 , n57237 );
buf ( n57239 , n57238 );
not ( n57240 , n57239 );
or ( n57241 , n57235 , n57240 );
xor ( n57242 , n55653 , n55668 );
xor ( n57243 , n57242 , n55776 );
buf ( n57244 , n57243 );
buf ( n57245 , n48868 );
not ( n57246 , n57245 );
buf ( n57247 , n55820 );
not ( n57248 , n57247 );
or ( n57249 , n57246 , n57248 );
xor ( n57250 , n37072 , n48808 );
xnor ( n57251 , n57250 , n37071 );
buf ( n57252 , n57251 );
buf ( n57253 , n48855 );
nand ( n57254 , n57252 , n57253 );
buf ( n57255 , n57254 );
buf ( n57256 , n57255 );
nand ( n57257 , n57249 , n57256 );
buf ( n57258 , n57257 );
or ( n57259 , n57244 , n57258 );
xor ( n57260 , n55675 , n55697 );
xor ( n57261 , n57260 , n55773 );
buf ( n57262 , n57261 );
not ( n57263 , n57262 );
buf ( n57264 , n57263 );
buf ( n57265 , n57264 );
not ( n57266 , n57265 );
and ( n57267 , n55920 , n55891 );
not ( n57268 , n55920 );
and ( n57269 , n57268 , n55894 );
nor ( n57270 , n57267 , n57269 );
buf ( n57271 , n57270 );
buf ( n57272 , n55860 );
and ( n57273 , n57271 , n57272 );
not ( n57274 , n57271 );
buf ( n57275 , n55863 );
and ( n57276 , n57274 , n57275 );
nor ( n57277 , n57273 , n57276 );
buf ( n57278 , n57277 );
buf ( n57279 , n57278 );
not ( n57280 , n57279 );
buf ( n57281 , n57280 );
buf ( n57282 , n57281 );
not ( n57283 , n57282 );
buf ( n57284 , n57283 );
buf ( n57285 , n57284 );
not ( n57286 , n57285 );
or ( n57287 , n57266 , n57286 );
buf ( n57288 , n57261 );
not ( n57289 , n57288 );
buf ( n57290 , n57281 );
not ( n57291 , n57290 );
or ( n57292 , n57289 , n57291 );
not ( n57293 , n55881 );
buf ( n57294 , n47716 );
not ( n57295 , n57294 );
buf ( n57296 , n43371 );
not ( n57297 , n57296 );
or ( n57298 , n57295 , n57297 );
buf ( n57299 , n38108 );
buf ( n57300 , n47725 );
nand ( n57301 , n57299 , n57300 );
buf ( n57302 , n57301 );
buf ( n57303 , n57302 );
nand ( n57304 , n57298 , n57303 );
buf ( n57305 , n57304 );
not ( n57306 , n57305 );
or ( n57307 , n57293 , n57306 );
not ( n57308 , n55876 );
or ( n57309 , n57308 , n38057 );
nand ( n57310 , n57307 , n57309 );
buf ( n57311 , n57310 );
not ( n57312 , n57311 );
buf ( n57313 , n50060 );
not ( n57314 , n57313 );
buf ( n57315 , n42082 );
not ( n57316 , n57315 );
or ( n57317 , n57314 , n57316 );
buf ( n57318 , n39136 );
buf ( n57319 , n50067 );
nand ( n57320 , n57318 , n57319 );
buf ( n57321 , n57320 );
buf ( n57322 , n57321 );
nand ( n57323 , n57317 , n57322 );
buf ( n57324 , n57323 );
buf ( n57325 , n57324 );
not ( n57326 , n57325 );
not ( n57327 , n44776 );
or ( n57328 , n57326 , n57327 );
nand ( n57329 , n36912 , n56212 );
nand ( n57330 , n57328 , n57329 );
buf ( n57331 , n57330 );
not ( n57332 , n57331 );
or ( n57333 , n57312 , n57332 );
or ( n57334 , n57330 , n57310 );
buf ( n57335 , n42865 );
not ( n57336 , n57335 );
buf ( n57337 , n41778 );
not ( n57338 , n57337 );
or ( n57339 , n57336 , n57338 );
buf ( n57340 , n37327 );
buf ( n57341 , n42862 );
nand ( n57342 , n57340 , n57341 );
buf ( n57343 , n57342 );
buf ( n57344 , n57343 );
nand ( n57345 , n57339 , n57344 );
buf ( n57346 , n57345 );
buf ( n57347 , n57346 );
not ( n57348 , n57347 );
buf ( n57349 , n37394 );
not ( n57350 , n57349 );
or ( n57351 , n57348 , n57350 );
buf ( n57352 , n56160 );
buf ( n57353 , n37410 );
nand ( n57354 , n57352 , n57353 );
buf ( n57355 , n57354 );
buf ( n57356 , n57355 );
nand ( n57357 , n57351 , n57356 );
buf ( n57358 , n57357 );
not ( n57359 , n57358 );
not ( n57360 , n42668 );
not ( n57361 , n56522 );
or ( n57362 , n57360 , n57361 );
buf ( n57363 , n29287 );
not ( n57364 , n57363 );
buf ( n57365 , n25227 );
not ( n57366 , n57365 );
and ( n57367 , n57364 , n57366 );
buf ( n57368 , n29287 );
buf ( n57369 , n25227 );
and ( n57370 , n57368 , n57369 );
nor ( n57371 , n57367 , n57370 );
buf ( n57372 , n57371 );
or ( n57373 , n57372 , n42711 );
nand ( n57374 , n57362 , n57373 );
not ( n57375 , n57374 );
or ( n57376 , n57359 , n57375 );
buf ( n57377 , n57358 );
buf ( n57378 , n57374 );
or ( n57379 , n57377 , n57378 );
xor ( n57380 , n55726 , n55739 );
xor ( n57381 , n57380 , n55765 );
buf ( n57382 , n57381 );
nand ( n57383 , n57379 , n57382 );
buf ( n57384 , n57383 );
nand ( n57385 , n57376 , n57384 );
nand ( n57386 , n57334 , n57385 );
buf ( n57387 , n57386 );
nand ( n57388 , n57333 , n57387 );
buf ( n57389 , n57388 );
buf ( n57390 , n57389 );
nand ( n57391 , n57292 , n57390 );
buf ( n57392 , n57391 );
buf ( n57393 , n57392 );
nand ( n57394 , n57287 , n57393 );
buf ( n57395 , n57394 );
and ( n57396 , n57259 , n57395 );
and ( n57397 , n57244 , n57258 );
nor ( n57398 , n57396 , n57397 );
buf ( n57399 , n57398 );
not ( n57400 , n57399 );
buf ( n57401 , n57400 );
buf ( n57402 , n57401 );
nand ( n57403 , n57241 , n57402 );
buf ( n57404 , n57403 );
buf ( n57405 , n57404 );
nand ( n57406 , n57233 , n57405 );
buf ( n57407 , n57406 );
buf ( n57408 , n57407 );
and ( n57409 , n57130 , n57408 );
and ( n57410 , n57125 , n57129 );
or ( n57411 , n57409 , n57410 );
buf ( n57412 , n57411 );
buf ( n57413 , n57412 );
not ( n57414 , n57413 );
buf ( n57415 , n57414 );
buf ( n57416 , n57415 );
not ( n57417 , n57416 );
xor ( n57418 , n55795 , n56070 );
xor ( n57419 , n57418 , n56075 );
buf ( n57420 , n57419 );
not ( n57421 , n57420 );
buf ( n57422 , n57421 );
not ( n57423 , n57422 );
or ( n57424 , n57417 , n57423 );
buf ( n57425 , n56063 );
buf ( n57426 , n55965 );
xor ( n57427 , n57425 , n57426 );
buf ( n57428 , n57427 );
buf ( n57429 , n55970 );
not ( n57430 , n57429 );
and ( n57431 , n57428 , n57430 );
not ( n57432 , n57428 );
and ( n57433 , n57432 , n57429 );
nor ( n57434 , n57431 , n57433 );
not ( n57435 , n57434 );
not ( n57436 , n57435 );
not ( n57437 , n55989 );
not ( n57438 , n55994 );
or ( n57439 , n57437 , n57438 );
nand ( n57440 , n55993 , n55986 );
nand ( n57441 , n57439 , n57440 );
and ( n57442 , n57441 , n56057 );
not ( n57443 , n57441 );
buf ( n57444 , n56057 );
not ( n57445 , n57444 );
buf ( n57446 , n57445 );
and ( n57447 , n57443 , n57446 );
nor ( n57448 , n57442 , n57447 );
buf ( n57449 , n57448 );
not ( n57450 , n57449 );
xor ( n57451 , n56115 , n56238 );
buf ( n57452 , n57451 );
buf ( n57453 , n57452 );
buf ( n57454 , n56247 );
and ( n57455 , n57453 , n57454 );
not ( n57456 , n57453 );
buf ( n57457 , n56244 );
and ( n57458 , n57456 , n57457 );
nor ( n57459 , n57455 , n57458 );
buf ( n57460 , n57459 );
buf ( n57461 , n57460 );
not ( n57462 , n57461 );
buf ( n57463 , n57462 );
not ( n57464 , n57463 );
xor ( n57465 , n56024 , n56048 );
xor ( n57466 , n57465 , n56051 );
not ( n57467 , n57466 );
not ( n57468 , n48855 );
buf ( n57469 , n48821 );
buf ( n57470 , n37147 );
and ( n57471 , n57469 , n57470 );
not ( n57472 , n57469 );
buf ( n57473 , n37146 );
and ( n57474 , n57472 , n57473 );
nor ( n57475 , n57471 , n57474 );
buf ( n57476 , n57475 );
not ( n57477 , n57476 );
or ( n57478 , n57468 , n57477 );
buf ( n57479 , n57251 );
buf ( n57480 , n48868 );
nand ( n57481 , n57479 , n57480 );
buf ( n57482 , n57481 );
nand ( n57483 , n57478 , n57482 );
not ( n57484 , n57483 );
nand ( n57485 , n57484 , C1 );
not ( n57486 , n57485 );
or ( n57487 , n57467 , n57486 );
nand ( n57488 , n57487 , C1 );
not ( n57489 , n57488 );
or ( n57490 , n57464 , n57489 );
buf ( n57491 , n57488 );
not ( n57492 , n57491 );
buf ( n57493 , n57492 );
not ( n57494 , n57493 );
not ( n57495 , n57460 );
or ( n57496 , n57494 , n57495 );
not ( n57497 , n42266 );
not ( n57498 , n42899 );
or ( n57499 , n57497 , n57498 );
buf ( n57500 , n38821 );
buf ( n57501 , n42263 );
nand ( n57502 , n57500 , n57501 );
buf ( n57503 , n57502 );
nand ( n57504 , n57499 , n57503 );
buf ( n57505 , n57504 );
not ( n57506 , n57505 );
buf ( n57507 , n57506 );
buf ( n57508 , n57507 );
not ( n57509 , n57508 );
buf ( n57510 , n42249 );
not ( n57511 , n57510 );
and ( n57512 , n57509 , n57511 );
buf ( n57513 , n56195 );
buf ( n57514 , n42315 );
and ( n57515 , n57513 , n57514 );
nor ( n57516 , n57512 , n57515 );
buf ( n57517 , n57516 );
buf ( n57518 , n36444 );
buf ( n57519 , n12481 );
nand ( n57520 , n57518 , n57519 );
buf ( n57521 , n57520 );
buf ( n57522 , n47489 );
not ( n57523 , n57522 );
buf ( n57524 , n44949 );
buf ( n57525 , n37472 );
and ( n57526 , n57524 , n57525 );
not ( n57527 , n57524 );
buf ( n57528 , n51901 );
and ( n57529 , n57527 , n57528 );
or ( n57530 , n57526 , n57529 );
buf ( n57531 , n57530 );
nor ( n57532 , n57523 , n57531 );
nand ( n57533 , n57532 , n41855 );
not ( n57534 , n37443 );
nand ( n57535 , n57534 , n56442 );
nand ( n57536 , n57521 , n57533 , n57535 );
buf ( n57537 , n41736 );
not ( n57538 , n57537 );
buf ( n57539 , n52551 );
not ( n57540 , n57539 );
or ( n57541 , n57538 , n57540 );
buf ( n57542 , n24092 );
buf ( n57543 , n41733 );
nand ( n57544 , n57542 , n57543 );
buf ( n57545 , n57544 );
buf ( n57546 , n57545 );
nand ( n57547 , n57541 , n57546 );
buf ( n57548 , n57547 );
buf ( n57549 , n57548 );
not ( n57550 , n57549 );
buf ( n57551 , n52537 );
not ( n57552 , n57551 );
or ( n57553 , n57550 , n57552 );
buf ( n57554 , n55753 );
buf ( n57555 , n39983 );
nand ( n57556 , n57554 , n57555 );
buf ( n57557 , n57556 );
buf ( n57558 , n57557 );
nand ( n57559 , n57553 , n57558 );
buf ( n57560 , n57559 );
not ( n57561 , n57560 );
buf ( n57562 , n42008 );
not ( n57563 , n57562 );
buf ( n57564 , n47031 );
not ( n57565 , n57564 );
or ( n57566 , n57563 , n57565 );
buf ( n57567 , n38979 );
buf ( n57568 , n42017 );
nand ( n57569 , n57567 , n57568 );
buf ( n57570 , n57569 );
buf ( n57571 , n57570 );
nand ( n57572 , n57566 , n57571 );
buf ( n57573 , n57572 );
buf ( n57574 , n57573 );
not ( n57575 , n57574 );
buf ( n57576 , n47050 );
not ( n57577 , n57576 );
or ( n57578 , n57575 , n57577 );
buf ( n57579 , n47019 );
not ( n57580 , n57579 );
buf ( n57581 , n56374 );
nand ( n57582 , n57580 , n57581 );
buf ( n57583 , n57582 );
buf ( n57584 , n57583 );
nand ( n57585 , n57578 , n57584 );
buf ( n57586 , n57585 );
not ( n57587 , n57586 );
or ( n57588 , n57561 , n57587 );
or ( n57589 , n57586 , n57560 );
buf ( n57590 , n55737 );
buf ( n57591 , n46294 );
and ( n57592 , n57590 , n57591 );
buf ( n57593 , n54068 );
not ( n57594 , n57593 );
buf ( n57595 , n43362 );
not ( n57596 , n57595 );
or ( n57597 , n57594 , n57596 );
buf ( n57598 , n50624 );
not ( n57599 , n42560 );
buf ( n57600 , n57599 );
nand ( n57601 , n57598 , n57600 );
buf ( n57602 , n57601 );
buf ( n57603 , n57602 );
nand ( n57604 , n57597 , n57603 );
buf ( n57605 , n57604 );
buf ( n57606 , n57605 );
buf ( n57607 , n43938 );
and ( n57608 , n57606 , n57607 );
buf ( n57609 , n57608 );
buf ( n57610 , n57609 );
nor ( n57611 , n57592 , n57610 );
buf ( n57612 , n57611 );
buf ( n57613 , n57612 );
not ( n57614 , n57613 );
buf ( n57615 , n57614 );
nand ( n57616 , n57589 , n57615 );
nand ( n57617 , n57588 , n57616 );
nand ( n57618 , n57536 , n57617 );
not ( n57619 , n41855 );
not ( n57620 , n57532 );
or ( n57621 , n57619 , n57620 );
nand ( n57622 , n57621 , n57535 );
not ( n57623 , n57521 );
nand ( n57624 , n57622 , n57623 );
nand ( n57625 , n57517 , n57618 , n57624 );
not ( n57626 , n57625 );
xor ( n57627 , n55707 , n55719 );
xor ( n57628 , n57627 , n55769 );
buf ( n57629 , n57628 );
not ( n57630 , n57629 );
or ( n57631 , n57626 , n57630 );
not ( n57632 , n57517 );
nand ( n57633 , n57618 , n57624 );
nand ( n57634 , n57632 , n57633 );
nand ( n57635 , n57631 , n57634 );
buf ( n57636 , n57635 );
buf ( n57637 , n46225 );
not ( n57638 , n57637 );
buf ( n57639 , n45753 );
not ( n57640 , n57639 );
buf ( n57641 , n52229 );
not ( n57642 , n57641 );
or ( n57643 , n57640 , n57642 );
buf ( n57644 , n50463 );
buf ( n57645 , n45750 );
nand ( n57646 , n57644 , n57645 );
buf ( n57647 , n57646 );
buf ( n57648 , n57647 );
nand ( n57649 , n57643 , n57648 );
buf ( n57650 , n57649 );
buf ( n57651 , n57650 );
not ( n57652 , n57651 );
or ( n57653 , n57638 , n57652 );
buf ( n57654 , n56107 );
buf ( n57655 , n46246 );
nand ( n57656 , n57654 , n57655 );
buf ( n57657 , n57656 );
buf ( n57658 , n57657 );
nand ( n57659 , n57653 , n57658 );
buf ( n57660 , n57659 );
buf ( n57661 , n57660 );
xor ( n57662 , n57636 , n57661 );
buf ( n57663 , n53539 );
not ( n57664 , n57663 );
buf ( n57665 , n41718 );
not ( n57666 , n57665 );
or ( n57667 , n57664 , n57666 );
buf ( n57668 , n41715 );
buf ( n57669 , n53548 );
nand ( n57670 , n57668 , n57669 );
buf ( n57671 , n57670 );
buf ( n57672 , n57671 );
nand ( n57673 , n57667 , n57672 );
buf ( n57674 , n57673 );
buf ( n57675 , n57674 );
not ( n57676 , n57675 );
buf ( n57677 , n39803 );
not ( n57678 , n57677 );
or ( n57679 , n57676 , n57678 );
buf ( n57680 , n44141 );
buf ( n57681 , n56036 );
nand ( n57682 , n57680 , n57681 );
buf ( n57683 , n57682 );
buf ( n57684 , n57683 );
nand ( n57685 , n57679 , n57684 );
buf ( n57686 , n57685 );
buf ( n57687 , n57686 );
xor ( n57688 , n56133 , n56147 );
xor ( n57689 , n57688 , n56173 );
buf ( n57690 , n57689 );
buf ( n57691 , n57690 );
xor ( n57692 , n57687 , n57691 );
not ( n57693 , n42252 );
buf ( n57694 , n42266 );
not ( n57695 , n57694 );
buf ( n57696 , n42485 );
not ( n57697 , n57696 );
or ( n57698 , n57695 , n57697 );
buf ( n57699 , n38848 );
buf ( n57700 , n42263 );
nand ( n57701 , n57699 , n57700 );
buf ( n57702 , n57701 );
buf ( n57703 , n57702 );
nand ( n57704 , n57698 , n57703 );
buf ( n57705 , n57704 );
not ( n57706 , n57705 );
or ( n57707 , n57693 , n57706 );
nand ( n57708 , n57504 , n42315 );
nand ( n57709 , n57707 , n57708 );
buf ( n57710 , n46390 );
not ( n57711 , n57710 );
buf ( n57712 , n41890 );
not ( n57713 , n57712 );
or ( n57714 , n57711 , n57713 );
buf ( n57715 , n41889 );
buf ( n57716 , n46393 );
nand ( n57717 , n57715 , n57716 );
buf ( n57718 , n57717 );
buf ( n57719 , n57718 );
nand ( n57720 , n57714 , n57719 );
buf ( n57721 , n57720 );
not ( n57722 , n57721 );
not ( n57723 , n37872 );
or ( n57724 , n57722 , n57723 );
buf ( n57725 , n42175 );
buf ( n57726 , n56428 );
nand ( n57727 , n57725 , n57726 );
buf ( n57728 , n57727 );
nand ( n57729 , n57724 , n57728 );
or ( n57730 , n57709 , n57729 );
buf ( n57731 , n52780 );
not ( n57732 , n57731 );
buf ( n57733 , n43259 );
not ( n57734 , n57733 );
or ( n57735 , n57732 , n57734 );
buf ( n57736 , n33077 );
buf ( n57737 , n52789 );
nand ( n57738 , n57736 , n57737 );
buf ( n57739 , n57738 );
buf ( n57740 , n57739 );
nand ( n57741 , n57735 , n57740 );
buf ( n57742 , n57741 );
buf ( n57743 , n57742 );
not ( n57744 , n57743 );
buf ( n57745 , n51937 );
not ( n57746 , n57745 );
or ( n57747 , n57744 , n57746 );
buf ( n57748 , n42530 );
buf ( n57749 , n56301 );
nand ( n57750 , n57748 , n57749 );
buf ( n57751 , n57750 );
buf ( n57752 , n57751 );
nand ( n57753 , n57747 , n57752 );
buf ( n57754 , n57753 );
nand ( n57755 , n57730 , n57754 );
buf ( n57756 , n57755 );
nand ( n57757 , n57709 , n57729 );
buf ( n57758 , n57757 );
nand ( n57759 , n57756 , n57758 );
buf ( n57760 , n57759 );
buf ( n57761 , n57760 );
and ( n57762 , n57692 , n57761 );
and ( n57763 , n57687 , n57691 );
or ( n57764 , n57762 , n57763 );
buf ( n57765 , n57764 );
buf ( n57766 , n57765 );
and ( n57767 , n57662 , n57766 );
and ( n57768 , n57636 , n57661 );
or ( n57769 , n57767 , n57768 );
buf ( n57770 , n57769 );
nand ( n57771 , n57496 , n57770 );
nand ( n57772 , n57490 , n57771 );
not ( n57773 , n57772 );
or ( n57774 , n57450 , n57773 );
buf ( n57775 , n57772 );
not ( n57776 , n57775 );
buf ( n57777 , n57776 );
not ( n57778 , n57777 );
not ( n57779 , n57449 );
not ( n57780 , n57779 );
or ( n57781 , n57778 , n57780 );
xor ( n57782 , n56004 , n56020 );
xor ( n57783 , n57782 , n56054 );
buf ( n57784 , n57783 );
xor ( n57785 , n57049 , n57062 );
xor ( n57786 , n57785 , n57091 );
buf ( n57787 , n57786 );
buf ( n57788 , n57787 );
xor ( n57789 , n57784 , n57788 );
buf ( n57790 , n51488 );
not ( n57791 , n57790 );
buf ( n57792 , n48836 );
not ( n57793 , n57792 );
buf ( n57794 , n39897 );
not ( n57795 , n57794 );
or ( n57796 , n57793 , n57795 );
buf ( n57797 , n36396 );
buf ( n57798 , n51493 );
nand ( n57799 , n57797 , n57798 );
buf ( n57800 , n57799 );
buf ( n57801 , n57800 );
nand ( n57802 , n57796 , n57801 );
buf ( n57803 , n57802 );
buf ( n57804 , n57803 );
not ( n57805 , n57804 );
or ( n57806 , n57791 , n57805 );
buf ( n57807 , n57180 );
buf ( n57808 , n52456 );
nand ( n57809 , n57807 , n57808 );
buf ( n57810 , n57809 );
buf ( n57811 , n57810 );
nand ( n57812 , n57806 , n57811 );
buf ( n57813 , n57812 );
buf ( n57814 , n43198 );
not ( n57815 , n57814 );
buf ( n57816 , n44530 );
not ( n57817 , n57816 );
and ( n57818 , n57815 , n57817 );
buf ( n57819 , n39522 );
buf ( n57820 , n44530 );
and ( n57821 , n57819 , n57820 );
nor ( n57822 , n57818 , n57821 );
buf ( n57823 , n57822 );
not ( n57824 , n57823 );
not ( n57825 , n44518 );
and ( n57826 , n57824 , n57825 );
and ( n57827 , n56946 , n44496 );
nor ( n57828 , n57826 , n57827 );
not ( n57829 , n57828 );
not ( n57830 , n57829 );
buf ( n57831 , n56276 );
not ( n57832 , n57831 );
buf ( n57833 , n57832 );
buf ( n57834 , n57833 );
buf ( n57835 , n43868 );
and ( n57836 , n57834 , n57835 );
buf ( n57837 , n41608 );
not ( n57838 , n57837 );
buf ( n57839 , n37589 );
not ( n57840 , n57839 );
or ( n57841 , n57838 , n57840 );
buf ( n57842 , n44163 );
buf ( n57843 , n41611 );
nand ( n57844 , n57842 , n57843 );
buf ( n57845 , n57844 );
buf ( n57846 , n57845 );
nand ( n57847 , n57841 , n57846 );
buf ( n57848 , n57847 );
buf ( n57849 , n57848 );
not ( n57850 , n57849 );
buf ( n57851 , n41599 );
nor ( n57852 , n57850 , n57851 );
buf ( n57853 , n57852 );
buf ( n57854 , n57853 );
nor ( n57855 , n57836 , n57854 );
buf ( n57856 , n57855 );
buf ( n57857 , n57856 );
not ( n57858 , n57857 );
buf ( n57859 , n57858 );
not ( n57860 , n57859 );
or ( n57861 , n57830 , n57860 );
not ( n57862 , n57856 );
not ( n57863 , n57828 );
or ( n57864 , n57862 , n57863 );
and ( n57865 , n56454 , n56487 );
not ( n57866 , n56454 );
and ( n57867 , n57866 , n56484 );
or ( n57868 , n57865 , n57867 );
buf ( n57869 , n56437 );
and ( n57870 , n57868 , n57869 );
not ( n57871 , n57868 );
not ( n57872 , n57869 );
and ( n57873 , n57871 , n57872 );
nor ( n57874 , n57870 , n57873 );
nand ( n57875 , n57864 , n57874 );
nand ( n57876 , n57861 , n57875 );
or ( n57877 , n57813 , n57876 );
xor ( n57878 , n56932 , n56969 );
xor ( n57879 , n57878 , n56977 );
buf ( n57880 , n57879 );
nand ( n57881 , n57877 , n57880 );
buf ( n57882 , n57881 );
nand ( n57883 , n57876 , n57813 );
buf ( n57884 , n57883 );
nand ( n57885 , n57882 , n57884 );
buf ( n57886 , n57885 );
buf ( n57887 , n57886 );
and ( n57888 , n57789 , n57887 );
and ( n57889 , n57784 , n57788 );
or ( n57890 , n57888 , n57889 );
buf ( n57891 , n57890 );
buf ( n57892 , n57891 );
nand ( n57893 , n57781 , n57892 );
nand ( n57894 , n57774 , n57893 );
not ( n57895 , n57894 );
or ( n57896 , n57436 , n57895 );
or ( n57897 , n57894 , n57435 );
xor ( n57898 , n56099 , n56991 );
xor ( n57899 , n57898 , n56997 );
nand ( n57900 , n57897 , n57899 );
nand ( n57901 , n57896 , n57900 );
buf ( n57902 , n57901 );
nand ( n57903 , n57424 , n57902 );
buf ( n57904 , n57903 );
buf ( n57905 , n57904 );
buf ( n57906 , n57420 );
buf ( n57907 , n57412 );
nand ( n57908 , n57906 , n57907 );
buf ( n57909 , n57908 );
buf ( n57910 , n57909 );
and ( n57911 , n57905 , n57910 );
buf ( n57912 , n57911 );
buf ( n57913 , n57912 );
xor ( n57914 , n57047 , n57913 );
buf ( n57915 , n56079 );
not ( n57916 , n57915 );
buf ( n57917 , n56090 );
not ( n57918 , n57917 );
or ( n57919 , n57916 , n57918 );
buf ( n57920 , n55603 );
buf ( n57921 , n56085 );
nand ( n57922 , n57920 , n57921 );
buf ( n57923 , n57922 );
buf ( n57924 , n57923 );
nand ( n57925 , n57919 , n57924 );
buf ( n57926 , n57925 );
buf ( n57927 , n57926 );
buf ( n57928 , n57009 );
not ( n57929 , n57928 );
buf ( n57930 , n57929 );
buf ( n57931 , n57930 );
and ( n57932 , n57927 , n57931 );
not ( n57933 , n57927 );
buf ( n57934 , n57009 );
and ( n57935 , n57933 , n57934 );
nor ( n57936 , n57932 , n57935 );
buf ( n57937 , n57936 );
buf ( n57938 , n57937 );
and ( n57939 , n57914 , n57938 );
and ( n57940 , n57047 , n57913 );
or ( n57941 , n57939 , n57940 );
buf ( n57942 , n57941 );
not ( n57943 , n57942 );
xor ( n57944 , n55600 , n57019 );
xor ( n57945 , n57944 , n57024 );
buf ( n57946 , n57945 );
not ( n57947 , n57946 );
or ( n57948 , n57943 , n57947 );
xor ( n57949 , n57047 , n57913 );
xor ( n57950 , n57949 , n57938 );
buf ( n57951 , n57950 );
buf ( n57952 , n57951 );
xor ( n57953 , n56257 , n56261 );
xor ( n57954 , n57953 , n56987 );
buf ( n57955 , n57954 );
buf ( n57956 , n57955 );
xor ( n57957 , n57095 , n57113 );
xor ( n57958 , n57957 , n57120 );
buf ( n57959 , n57958 );
buf ( n57960 , n57959 );
xor ( n57961 , n57956 , n57960 );
buf ( n57962 , n57244 );
buf ( n57963 , n57258 );
xor ( n57964 , n57962 , n57963 );
buf ( n57965 , n57395 );
xor ( n57966 , n57964 , n57965 );
buf ( n57967 , n57966 );
not ( n57968 , n57967 );
xor ( n57969 , n56266 , n56505 );
xor ( n57970 , n57969 , n56982 );
buf ( n57971 , n57970 );
not ( n57972 , n57971 );
or ( n57973 , n57968 , n57972 );
or ( n57974 , n57971 , n57967 );
xor ( n57975 , n56411 , n56313 );
xnor ( n57976 , n57975 , n56327 );
buf ( n57977 , n57976 );
not ( n57978 , n57977 );
buf ( n57979 , n56532 );
not ( n57980 , n57979 );
buf ( n57981 , n56924 );
not ( n57982 , n57981 );
or ( n57983 , n57980 , n57982 );
buf ( n57984 , n56512 );
buf ( n57985 , n56529 );
nand ( n57986 , n57984 , n57985 );
buf ( n57987 , n57986 );
buf ( n57988 , n57987 );
nand ( n57989 , n57983 , n57988 );
buf ( n57990 , n57989 );
buf ( n57991 , n57990 );
buf ( n57992 , n56918 );
not ( n57993 , n57992 );
buf ( n57994 , n57993 );
buf ( n57995 , n57994 );
and ( n57996 , n57991 , n57995 );
not ( n57997 , n57991 );
buf ( n57998 , n56918 );
and ( n57999 , n57997 , n57998 );
nor ( n58000 , n57996 , n57999 );
buf ( n58001 , n58000 );
buf ( n58002 , n58001 );
not ( n58003 , n58002 );
buf ( n58004 , n58003 );
buf ( n58005 , n58004 );
not ( n58006 , n58005 );
or ( n58007 , n57978 , n58006 );
not ( n58008 , n57976 );
nand ( n58009 , n58008 , n58001 );
buf ( n58010 , n48323 );
not ( n58011 , n58010 );
buf ( n58012 , n43371 );
not ( n58013 , n58012 );
or ( n58014 , n58011 , n58013 );
buf ( n58015 , n45376 );
buf ( n58016 , n48320 );
nand ( n58017 , n58015 , n58016 );
buf ( n58018 , n58017 );
buf ( n58019 , n58018 );
nand ( n58020 , n58014 , n58019 );
buf ( n58021 , n58020 );
buf ( n58022 , n58021 );
not ( n58023 , n58022 );
buf ( n58024 , n43386 );
not ( n58025 , n58024 );
or ( n58026 , n58023 , n58025 );
buf ( n58027 , n57305 );
buf ( n58028 , n45144 );
nand ( n58029 , n58027 , n58028 );
buf ( n58030 , n58029 );
buf ( n58031 , n58030 );
nand ( n58032 , n58026 , n58031 );
buf ( n58033 , n58032 );
buf ( n58034 , n58033 );
xor ( n58035 , n56869 , n56894 );
xor ( n58036 , n58035 , n56914 );
buf ( n58037 , n58036 );
buf ( n58038 , n58037 );
xor ( n58039 , n58034 , n58038 );
buf ( n58040 , n44267 );
not ( n58041 , n58040 );
buf ( n58042 , n41608 );
not ( n58043 , n58042 );
buf ( n58044 , n42891 );
not ( n58045 , n58044 );
or ( n58046 , n58043 , n58045 );
buf ( n58047 , n37641 );
buf ( n58048 , n41611 );
nand ( n58049 , n58047 , n58048 );
buf ( n58050 , n58049 );
buf ( n58051 , n58050 );
nand ( n58052 , n58046 , n58051 );
buf ( n58053 , n58052 );
buf ( n58054 , n58053 );
not ( n58055 , n58054 );
or ( n58056 , n58041 , n58055 );
buf ( n58057 , n57848 );
buf ( n58058 , n41574 );
nand ( n58059 , n58057 , n58058 );
buf ( n58060 , n58059 );
buf ( n58061 , n58060 );
nand ( n58062 , n58056 , n58061 );
buf ( n58063 , n58062 );
buf ( n58064 , n58063 );
and ( n58065 , n58039 , n58064 );
and ( n58066 , n58034 , n58038 );
or ( n58067 , n58065 , n58066 );
buf ( n58068 , n58067 );
nand ( n58069 , n58009 , n58068 );
buf ( n58070 , n58069 );
nand ( n58071 , n58007 , n58070 );
buf ( n58072 , n58071 );
not ( n58073 , n58072 );
or ( n58074 , n56286 , n56489 );
nand ( n58075 , n56489 , n56286 );
nand ( n58076 , n58074 , n58075 );
buf ( n58077 , n56413 );
and ( n58078 , n58076 , n58077 );
not ( n58079 , n58076 );
and ( n58080 , n58079 , n56498 );
nor ( n58081 , n58078 , n58080 );
buf ( n58082 , n58081 );
not ( n58083 , n58082 );
buf ( n58084 , n58083 );
not ( n58085 , n58084 );
or ( n58086 , n58073 , n58085 );
buf ( n58087 , n58072 );
not ( n58088 , n58087 );
buf ( n58089 , n58088 );
not ( n58090 , n58089 );
not ( n58091 , n58081 );
or ( n58092 , n58090 , n58091 );
xor ( n58093 , n56362 , n56388 );
xor ( n58094 , n58093 , n56407 );
buf ( n58095 , n58094 );
not ( n58096 , n58095 );
buf ( n58097 , n48671 );
not ( n58098 , n58097 );
buf ( n58099 , n56396 );
not ( n58100 , n58099 );
or ( n58101 , n58098 , n58100 );
nand ( n58102 , n48390 , n41873 );
not ( n58103 , n58102 );
buf ( n58104 , n50575 );
buf ( n58105 , n41698 );
not ( n58106 , n58105 );
buf ( n58107 , n58106 );
buf ( n58108 , n58107 );
nand ( n58109 , n58104 , n58108 );
buf ( n58110 , n58109 );
not ( n58111 , n58110 );
or ( n58112 , n58103 , n58111 );
nand ( n58113 , n58112 , n50982 );
buf ( n58114 , n58113 );
nand ( n58115 , n58101 , n58114 );
buf ( n58116 , n58115 );
buf ( n58117 , n58116 );
not ( n58118 , n58117 );
buf ( n58119 , n43063 );
not ( n58120 , n58119 );
buf ( n58121 , n44054 );
not ( n58122 , n58121 );
or ( n58123 , n58120 , n58122 );
buf ( n58124 , n42411 );
buf ( n58125 , n43064 );
nand ( n58126 , n58124 , n58125 );
buf ( n58127 , n58126 );
buf ( n58128 , n58127 );
nand ( n58129 , n58123 , n58128 );
buf ( n58130 , n58129 );
not ( n58131 , n58130 );
not ( n58132 , n46620 );
or ( n58133 , n58131 , n58132 );
buf ( n58134 , n56907 );
buf ( n58135 , n38380 );
nand ( n58136 , n58134 , n58135 );
buf ( n58137 , n58136 );
nand ( n58138 , n58133 , n58137 );
buf ( n58139 , n58138 );
not ( n58140 , n58139 );
or ( n58141 , n58118 , n58140 );
buf ( n58142 , n58138 );
buf ( n58143 , n58116 );
or ( n58144 , n58142 , n58143 );
buf ( n58145 , n42339 );
not ( n58146 , n58145 );
buf ( n58147 , n56883 );
not ( n58148 , n58147 );
or ( n58149 , n58146 , n58148 );
not ( n58150 , n42343 );
not ( n58151 , n51250 );
or ( n58152 , n58150 , n58151 );
buf ( n58153 , n41822 );
buf ( n58154 , n46855 );
nand ( n58155 , n58153 , n58154 );
buf ( n58156 , n58155 );
nand ( n58157 , n58152 , n58156 );
buf ( n58158 , n58157 );
buf ( n58159 , n42378 );
nand ( n58160 , n58158 , n58159 );
buf ( n58161 , n58160 );
buf ( n58162 , n58161 );
nand ( n58163 , n58149 , n58162 );
buf ( n58164 , n58163 );
buf ( n58165 , n58164 );
nand ( n58166 , n58144 , n58165 );
buf ( n58167 , n58166 );
buf ( n58168 , n58167 );
nand ( n58169 , n58141 , n58168 );
buf ( n58170 , n58169 );
not ( n58171 , n58170 );
nand ( n58172 , n58096 , n58171 );
not ( n58173 , n58172 );
xor ( n58174 , n56681 , n56688 );
xor ( n58175 , n58174 , n56852 );
buf ( n58176 , n58175 );
buf ( n58177 , n58176 );
buf ( n58178 , n43905 );
not ( n58179 , n58178 );
buf ( n58180 , n57605 );
not ( n58181 , n58180 );
or ( n58182 , n58179 , n58181 );
and ( n58183 , n28368 , n25181 );
not ( n58184 , n28368 );
buf ( n58185 , n25180 );
and ( n58186 , n58184 , n58185 );
or ( n58187 , n58183 , n58186 );
buf ( n58188 , n58187 );
buf ( n58189 , n43935 );
nand ( n58190 , n58188 , n58189 );
buf ( n58191 , n58190 );
buf ( n58192 , n58191 );
nand ( n58193 , n58182 , n58192 );
buf ( n58194 , n58193 );
buf ( n58195 , n58194 );
xor ( n58196 , n58177 , n58195 );
buf ( n58197 , n42504 );
not ( n58198 , n58197 );
buf ( n58199 , n47857 );
not ( n58200 , n58199 );
or ( n58201 , n58198 , n58200 );
buf ( n58202 , n24092 );
buf ( n58203 , n41721 );
nand ( n58204 , n58202 , n58203 );
buf ( n58205 , n58204 );
buf ( n58206 , n58205 );
nand ( n58207 , n58201 , n58206 );
buf ( n58208 , n58207 );
buf ( n58209 , n58208 );
not ( n58210 , n58209 );
buf ( n58211 , n39999 );
not ( n58212 , n58211 );
or ( n58213 , n58210 , n58212 );
buf ( n58214 , n57548 );
buf ( n58215 , n46633 );
nand ( n58216 , n58214 , n58215 );
buf ( n58217 , n58216 );
buf ( n58218 , n58217 );
nand ( n58219 , n58213 , n58218 );
buf ( n58220 , n58219 );
buf ( n58221 , n58220 );
and ( n58222 , n58196 , n58221 );
and ( n58223 , n58177 , n58195 );
or ( n58224 , n58222 , n58223 );
buf ( n58225 , n58224 );
buf ( n58226 , n58225 );
not ( n58227 , n58226 );
buf ( n58228 , n42668 );
not ( n58229 , n58228 );
buf ( n58230 , n57372 );
not ( n58231 , n58230 );
buf ( n58232 , n58231 );
buf ( n58233 , n58232 );
not ( n58234 , n58233 );
or ( n58235 , n58229 , n58234 );
buf ( n58236 , n25228 );
not ( n58237 , n58236 );
buf ( n58238 , n41781 );
not ( n58239 , n58238 );
or ( n58240 , n58237 , n58239 );
buf ( n58241 , n41762 );
buf ( n58242 , n25227 );
nand ( n58243 , n58241 , n58242 );
buf ( n58244 , n58243 );
buf ( n58245 , n58244 );
nand ( n58246 , n58240 , n58245 );
buf ( n58247 , n58246 );
buf ( n58248 , n58247 );
buf ( n58249 , n46047 );
buf ( n58250 , n58249 );
nand ( n58251 , n58248 , n58250 );
buf ( n58252 , n58251 );
buf ( n58253 , n58252 );
nand ( n58254 , n58235 , n58253 );
buf ( n58255 , n58254 );
buf ( n58256 , n58255 );
not ( n58257 , n58256 );
or ( n58258 , n58227 , n58257 );
buf ( n58259 , n58255 );
buf ( n58260 , n58225 );
or ( n58261 , n58259 , n58260 );
buf ( n58262 , n56561 );
not ( n58263 , n58262 );
buf ( n58264 , n50128 );
not ( n58265 , n58264 );
or ( n58266 , n58263 , n58265 );
buf ( n58267 , n56571 );
nand ( n58268 , n58266 , n58267 );
buf ( n58269 , n58268 );
buf ( n58270 , n58269 );
not ( n58271 , n58270 );
buf ( n58272 , n56856 );
not ( n58273 , n58272 );
buf ( n58274 , n56540 );
not ( n58275 , n58274 );
and ( n58276 , n58273 , n58275 );
buf ( n58277 , n56856 );
buf ( n58278 , n56540 );
and ( n58279 , n58277 , n58278 );
nor ( n58280 , n58276 , n58279 );
buf ( n58281 , n58280 );
buf ( n58282 , n58281 );
not ( n58283 , n58282 );
and ( n58284 , n58271 , n58283 );
buf ( n58285 , n58269 );
buf ( n58286 , n58281 );
and ( n58287 , n58285 , n58286 );
nor ( n58288 , n58284 , n58287 );
buf ( n58289 , n58288 );
buf ( n58290 , n58289 );
not ( n58291 , n58290 );
buf ( n58292 , n58291 );
buf ( n58293 , n58292 );
nand ( n58294 , n58261 , n58293 );
buf ( n58295 , n58294 );
buf ( n58296 , n58295 );
nand ( n58297 , n58258 , n58296 );
buf ( n58298 , n58297 );
not ( n58299 , n58298 );
or ( n58300 , n58173 , n58299 );
nand ( n58301 , n58170 , n58095 );
nand ( n58302 , n58300 , n58301 );
buf ( n58303 , n58302 );
buf ( n58304 , n46912 );
not ( n58305 , n58304 );
buf ( n58306 , n57145 );
not ( n58307 , n58306 );
or ( n58308 , n58305 , n58307 );
and ( n58309 , n46887 , n38247 );
not ( n58310 , n46887 );
and ( n58311 , n58310 , n43031 );
nor ( n58312 , n58309 , n58311 );
buf ( n58313 , n58312 );
not ( n58314 , n58313 );
buf ( n58315 , n47331 );
nand ( n58316 , n58314 , n58315 );
buf ( n58317 , n58316 );
buf ( n58318 , n58317 );
nand ( n58319 , n58308 , n58318 );
buf ( n58320 , n58319 );
buf ( n58321 , n58320 );
xor ( n58322 , n58303 , n58321 );
buf ( n58323 , n51004 );
not ( n58324 , n58323 );
buf ( n58325 , n49425 );
not ( n58326 , n58325 );
or ( n58327 , n58324 , n58326 );
buf ( n58328 , n39136 );
buf ( n58329 , n51001 );
nand ( n58330 , n58328 , n58329 );
buf ( n58331 , n58330 );
buf ( n58332 , n58331 );
nand ( n58333 , n58327 , n58332 );
buf ( n58334 , n58333 );
not ( n58335 , n58334 );
not ( n58336 , n45155 );
or ( n58337 , n58335 , n58336 );
buf ( n58338 , n57324 );
buf ( n58339 , n44676 );
nand ( n58340 , n58338 , n58339 );
buf ( n58341 , n58340 );
nand ( n58342 , n58337 , n58341 );
not ( n58343 , n58342 );
xor ( n58344 , n57358 , n57374 );
xnor ( n58345 , n58344 , n57381 );
not ( n58346 , n58345 );
not ( n58347 , n58346 );
or ( n58348 , n58343 , n58347 );
not ( n58349 , n58342 );
not ( n58350 , n58349 );
not ( n58351 , n58345 );
or ( n58352 , n58350 , n58351 );
buf ( n58353 , n55841 );
not ( n58354 , n58353 );
buf ( n58355 , n41718 );
not ( n58356 , n58355 );
or ( n58357 , n58354 , n58356 );
buf ( n58358 , n36527 );
buf ( n58359 , n55841 );
not ( n58360 , n58359 );
buf ( n58361 , n58360 );
buf ( n58362 , n58361 );
nand ( n58363 , n58358 , n58362 );
buf ( n58364 , n58363 );
buf ( n58365 , n58364 );
nand ( n58366 , n58357 , n58365 );
buf ( n58367 , n58366 );
buf ( n58368 , n58367 );
not ( n58369 , n58368 );
buf ( n58370 , n39806 );
not ( n58371 , n58370 );
or ( n58372 , n58369 , n58371 );
buf ( n58373 , n36643 );
buf ( n58374 , n57674 );
nand ( n58375 , n58373 , n58374 );
buf ( n58376 , n58375 );
buf ( n58377 , n58376 );
nand ( n58378 , n58372 , n58377 );
buf ( n58379 , n58378 );
nand ( n58380 , n58352 , n58379 );
nand ( n58381 , n58348 , n58380 );
buf ( n58382 , n58381 );
and ( n58383 , n58322 , n58382 );
and ( n58384 , n58303 , n58321 );
or ( n58385 , n58383 , n58384 );
buf ( n58386 , n58385 );
nand ( n58387 , n58092 , n58386 );
nand ( n58388 , n58086 , n58387 );
nand ( n58389 , n57974 , n58388 );
nand ( n58390 , n57973 , n58389 );
buf ( n58391 , n58390 );
and ( n58392 , n57961 , n58391 );
and ( n58393 , n57956 , n57960 );
or ( n58394 , n58392 , n58393 );
buf ( n58395 , n58394 );
buf ( n58396 , n58395 );
xor ( n58397 , n57125 , n57129 );
xor ( n58398 , n58397 , n57408 );
buf ( n58399 , n58398 );
buf ( n58400 , n58399 );
xor ( n58401 , n58396 , n58400 );
not ( n58402 , n57401 );
not ( n58403 , n57238 );
or ( n58404 , n58402 , n58403 );
buf ( n58405 , n57221 );
buf ( n58406 , n57398 );
nand ( n58407 , n58405 , n58406 );
buf ( n58408 , n58407 );
nand ( n58409 , n58404 , n58408 );
not ( n58410 , n57230 );
and ( n58411 , n58409 , n58410 );
not ( n58412 , n58409 );
and ( n58413 , n58412 , n57230 );
nor ( n58414 , n58411 , n58413 );
buf ( n58415 , n58414 );
not ( n58416 , n58415 );
xor ( n58417 , n57448 , n57777 );
xor ( n58418 , n58417 , n57891 );
buf ( n58419 , n58418 );
not ( n58420 , n58419 );
or ( n58421 , n58416 , n58420 );
xor ( n58422 , n57190 , n57162 );
xnor ( n58423 , n58422 , n57213 );
buf ( n58424 , n58423 );
not ( n58425 , n58424 );
buf ( n58426 , n58425 );
buf ( n58427 , n58426 );
not ( n58428 , n58427 );
xor ( n58429 , n57261 , n57278 );
xor ( n58430 , n58429 , n57389 );
not ( n58431 , n57310 );
xor ( n58432 , n57385 , n58431 );
buf ( n58433 , n57330 );
xnor ( n58434 , n58432 , n58433 );
not ( n58435 , n58434 );
or ( n58436 , n58435 , C1 );
xor ( n58437 , n58431 , n57385 );
xor ( n58438 , n58437 , n57330 );
not ( n58439 , n58438 );
or ( n58440 , n58439 , C0 );
xor ( n58441 , n57517 , n57629 );
xor ( n58442 , n58441 , n57633 );
buf ( n58443 , n58442 );
not ( n58444 , n58443 );
buf ( n58445 , n58444 );
nand ( n58446 , n58440 , n58445 );
nand ( n58447 , n58436 , n58446 );
buf ( n58448 , n58447 );
not ( n58449 , n58448 );
buf ( n58450 , n58449 );
xor ( n58451 , n58430 , n58450 );
not ( n58452 , n57147 );
not ( n58453 , n58452 );
not ( n58454 , n57160 );
or ( n58455 , n58453 , n58454 );
or ( n58456 , n58452 , n57160 );
nand ( n58457 , n58455 , n58456 );
buf ( n58458 , C1 );
and ( n58459 , n58457 , n58458 );
nor ( n58460 , n58459 , C0 );
and ( n58461 , n58451 , n58460 );
and ( n58462 , n58430 , n58450 );
or ( n58463 , n58461 , n58462 );
buf ( n58464 , n58463 );
not ( n58465 , n58464 );
buf ( n58466 , n58465 );
buf ( n58467 , n58466 );
not ( n58468 , n58467 );
or ( n58469 , n58428 , n58468 );
buf ( n58470 , n58423 );
not ( n58471 , n58470 );
buf ( n58472 , n58463 );
not ( n58473 , n58472 );
or ( n58474 , n58471 , n58473 );
not ( n58475 , n57484 );
or ( n58476 , C0 , n58475 );
nand ( n58477 , n58476 , C1 );
and ( n58478 , n58477 , n57466 );
not ( n58479 , n58477 );
not ( n58480 , n57466 );
and ( n58481 , n58479 , n58480 );
nor ( n58482 , n58478 , n58481 );
buf ( n58483 , n58482 );
not ( n58484 , n58483 );
buf ( n58485 , n58484 );
not ( n58486 , n58485 );
xor ( n58487 , n57636 , n57661 );
xor ( n58488 , n58487 , n57766 );
buf ( n58489 , n58488 );
not ( n58490 , n58489 );
or ( n58491 , n58486 , n58490 );
buf ( n58492 , n58489 );
not ( n58493 , n58492 );
buf ( n58494 , n58493 );
not ( n58495 , n58494 );
not ( n58496 , n58482 );
or ( n58497 , n58495 , n58496 );
buf ( n58498 , n46246 );
not ( n58499 , n58498 );
buf ( n58500 , n57650 );
not ( n58501 , n58500 );
or ( n58502 , n58499 , n58501 );
buf ( n58503 , n53492 );
not ( n58504 , n58503 );
buf ( n58505 , n49178 );
not ( n58506 , n58505 );
or ( n58507 , n58504 , n58506 );
buf ( n58508 , n37294 );
buf ( n58509 , n45750 );
nand ( n58510 , n58508 , n58509 );
buf ( n58511 , n58510 );
buf ( n58512 , n58511 );
nand ( n58513 , n58507 , n58512 );
buf ( n58514 , n58513 );
buf ( n58515 , n58514 );
buf ( n58516 , n46225 );
nand ( n58517 , n58515 , n58516 );
buf ( n58518 , n58517 );
buf ( n58519 , n58518 );
nand ( n58520 , n58502 , n58519 );
buf ( n58521 , n58520 );
buf ( n58522 , n58521 );
and ( n58523 , n57617 , n57521 );
not ( n58524 , n57617 );
and ( n58525 , n58524 , n57623 );
nor ( n58526 , n58523 , n58525 );
nand ( n58527 , n57533 , n57535 );
and ( n58528 , n58526 , n58527 );
not ( n58529 , n58526 );
not ( n58530 , n58527 );
and ( n58531 , n58529 , n58530 );
nor ( n58532 , n58528 , n58531 );
not ( n58533 , n58532 );
not ( n58534 , n58533 );
not ( n58535 , n45617 );
not ( n58536 , n57721 );
or ( n58537 , n58535 , n58536 );
not ( n58538 , n41865 );
not ( n58539 , n37881 );
not ( n58540 , n47725 );
or ( n58541 , n58539 , n58540 );
nand ( n58542 , n49879 , n47716 );
nand ( n58543 , n58541 , n58542 );
nand ( n58544 , n58538 , n58543 );
nand ( n58545 , n58537 , n58544 );
buf ( n58546 , n36490 );
and ( n58547 , n51030 , n58546 );
nor ( n58548 , n58547 , n38468 );
buf ( n58549 , n58548 );
buf ( n58550 , n51030 );
buf ( n58551 , n36490 );
or ( n58552 , n58550 , n58551 );
buf ( n58553 , n12481 );
nand ( n58554 , n58552 , n58553 );
buf ( n58555 , n58554 );
buf ( n58556 , n58555 );
nand ( n58557 , n58549 , n58556 );
buf ( n58558 , n58557 );
not ( n58559 , n58558 );
or ( n58560 , n58545 , n58559 );
buf ( n58561 , n57586 );
not ( n58562 , n58561 );
buf ( n58563 , n58562 );
buf ( n58564 , n58563 );
not ( n58565 , n58564 );
and ( n58566 , n57560 , n57612 );
not ( n58567 , n57560 );
and ( n58568 , n58567 , n57615 );
or ( n58569 , n58566 , n58568 );
buf ( n58570 , n58569 );
not ( n58571 , n58570 );
or ( n58572 , n58565 , n58571 );
buf ( n58573 , n58569 );
buf ( n58574 , n58563 );
or ( n58575 , n58573 , n58574 );
nand ( n58576 , n58572 , n58575 );
buf ( n58577 , n58576 );
nand ( n58578 , n58560 , n58577 );
buf ( n58579 , n58578 );
nand ( n58580 , n58545 , n58559 );
buf ( n58581 , n58580 );
and ( n58582 , n58579 , n58581 );
buf ( n58583 , n58582 );
buf ( n58584 , n58583 );
not ( n58585 , n58584 );
buf ( n58586 , n58585 );
not ( n58587 , n58586 );
or ( n58588 , n58534 , n58587 );
buf ( n58589 , n58532 );
not ( n58590 , n58589 );
buf ( n58591 , n58583 );
not ( n58592 , n58591 );
or ( n58593 , n58590 , n58592 );
and ( n58594 , n46126 , n37473 );
not ( n58595 , n46126 );
and ( n58596 , n58595 , n48207 );
nor ( n58597 , n58594 , n58596 );
or ( n58598 , n41969 , n58597 );
nor ( n58599 , n41855 , n57531 );
not ( n58600 , n58599 );
nand ( n58601 , n58598 , n58600 );
buf ( n58602 , n42847 );
not ( n58603 , n58602 );
buf ( n58604 , n41772 );
not ( n58605 , n58604 );
or ( n58606 , n58603 , n58605 );
buf ( n58607 , n41769 );
buf ( n58608 , n46691 );
nand ( n58609 , n58607 , n58608 );
buf ( n58610 , n58609 );
buf ( n58611 , n58610 );
nand ( n58612 , n58606 , n58611 );
buf ( n58613 , n58612 );
not ( n58614 , n58613 );
not ( n58615 , n37397 );
or ( n58616 , n58614 , n58615 );
buf ( n58617 , n57346 );
buf ( n58618 , n45108 );
nand ( n58619 , n58617 , n58618 );
buf ( n58620 , n58619 );
nand ( n58621 , n58616 , n58620 );
or ( n58622 , n58601 , n58621 );
not ( n58623 , n50128 );
buf ( n58624 , n13653 );
not ( n58625 , n58624 );
buf ( n58626 , n51804 );
not ( n58627 , n58626 );
or ( n58628 , n58625 , n58627 );
buf ( n58629 , n52673 );
buf ( n58630 , n13653 );
not ( n58631 , n58630 );
buf ( n58632 , n58631 );
buf ( n58633 , n58632 );
nand ( n58634 , n58629 , n58633 );
buf ( n58635 , n58634 );
buf ( n58636 , n58635 );
nand ( n58637 , n58628 , n58636 );
buf ( n58638 , n58637 );
not ( n58639 , n58638 );
or ( n58640 , n58623 , n58639 );
buf ( n58641 , n56561 );
buf ( n58642 , n56567 );
nand ( n58643 , n58641 , n58642 );
buf ( n58644 , n58643 );
nand ( n58645 , n58640 , n58644 );
not ( n58646 , n58645 );
not ( n58647 , n50982 );
and ( n58648 , n42149 , n58107 );
not ( n58649 , n42149 );
and ( n58650 , n58649 , n48390 );
or ( n58651 , n58648 , n58650 );
not ( n58652 , n58651 );
or ( n58653 , n58647 , n58652 );
not ( n58654 , n58102 );
not ( n58655 , n58110 );
or ( n58656 , n58654 , n58655 );
nand ( n58657 , n58656 , n48671 );
nand ( n58658 , n58653 , n58657 );
not ( n58659 , n58658 );
or ( n58660 , n58646 , n58659 );
or ( n58661 , n58645 , n58658 );
buf ( n58662 , n43905 );
not ( n58663 , n58662 );
buf ( n58664 , n58187 );
not ( n58665 , n58664 );
or ( n58666 , n58663 , n58665 );
buf ( n58667 , n42560 );
not ( n58668 , n58667 );
buf ( n58669 , n56545 );
not ( n58670 , n58669 );
or ( n58671 , n58668 , n58670 );
buf ( n58672 , n42559 );
buf ( n58673 , n29754 );
nand ( n58674 , n58672 , n58673 );
buf ( n58675 , n58674 );
buf ( n58676 , n58675 );
nand ( n58677 , n58671 , n58676 );
buf ( n58678 , n58677 );
buf ( n58679 , n58678 );
buf ( n58680 , n53628 );
nand ( n58681 , n58679 , n58680 );
buf ( n58682 , n58681 );
buf ( n58683 , n58682 );
nand ( n58684 , n58666 , n58683 );
buf ( n58685 , n58684 );
not ( n58686 , n58685 );
xor ( n58687 , n56602 , n56647 );
xor ( n58688 , n58687 , n56677 );
xor ( n58689 , n56731 , n56846 );
xor ( n58690 , n58688 , n58689 );
not ( n58691 , n58690 );
or ( n58692 , n58686 , n58691 );
nor ( n58693 , n58690 , n58685 );
xor ( n58694 , n56741 , n56758 );
xor ( n58695 , n58694 , n56842 );
buf ( n58696 , n58695 );
buf ( n58697 , n58696 );
not ( n58698 , n55246 );
nand ( n58699 , n58698 , n55248 );
buf ( n58700 , n58699 );
buf ( n58701 , n56641 );
and ( n58702 , n58700 , n58701 );
buf ( n58703 , n56594 );
buf ( n58704 , n56631 );
and ( n58705 , n58703 , n58704 );
nor ( n58706 , n58702 , n58705 );
buf ( n58707 , n58706 );
buf ( n58708 , n58707 );
buf ( n58709 , n56626 );
or ( n58710 , n58708 , n58709 );
buf ( n58711 , n56767 );
buf ( n58712 , n56639 );
or ( n58713 , n58711 , n58712 );
nand ( n58714 , n58710 , n58713 );
buf ( n58715 , n58714 );
buf ( n58716 , n58715 );
buf ( n58717 , n55152 );
buf ( n58718 , n56606 );
buf ( n58719 , n58718 );
not ( n58720 , n58719 );
buf ( n58721 , n58720 );
buf ( n58722 , n58721 );
and ( n58723 , n58717 , n58722 );
buf ( n58724 , n55205 );
buf ( n58725 , n58718 );
and ( n58726 , n58724 , n58725 );
nor ( n58727 , n58723 , n58726 );
buf ( n58728 , n58727 );
buf ( n58729 , n58728 );
buf ( n58730 , n56799 );
or ( n58731 , n58729 , n58730 );
buf ( n58732 , n56815 );
nand ( n58733 , n58731 , n58732 );
buf ( n58734 , n58733 );
buf ( n58735 , n58734 );
nor ( n58736 , n58716 , n58735 );
buf ( n58737 , n58736 );
buf ( n58738 , n58737 );
not ( n58739 , n54235 );
not ( n58740 , n55086 );
or ( n58741 , n58739 , n58740 );
nand ( n58742 , n58741 , n55092 );
nand ( n58743 , n54288 , n55096 );
nor ( n58744 , n58742 , n58743 );
not ( n58745 , n58744 );
nand ( n58746 , n58742 , n58743 );
nand ( n58747 , n58745 , n58746 );
buf ( n58748 , n58747 );
buf ( n58749 , n55132 );
and ( n58750 , n58748 , n58749 );
buf ( n58751 , n56720 );
buf ( n58752 , n55156 );
and ( n58753 , n58751 , n58752 );
nor ( n58754 , n58750 , n58753 );
buf ( n58755 , n58754 );
buf ( n58756 , n58755 );
or ( n58757 , n58738 , n58756 );
buf ( n58758 , n58755 );
not ( n58759 , n58758 );
buf ( n58760 , n58737 );
not ( n58761 , n58760 );
or ( n58762 , n58759 , n58761 );
xor ( n58763 , n56776 , n56819 );
xor ( n58764 , n58763 , n56837 );
buf ( n58765 , n58764 );
buf ( n58766 , n58765 );
nand ( n58767 , n58762 , n58766 );
buf ( n58768 , n58767 );
buf ( n58769 , n58768 );
nand ( n58770 , n58757 , n58769 );
buf ( n58771 , n58770 );
buf ( n58772 , n58771 );
and ( n58773 , n58697 , n58772 );
buf ( n58774 , n58696 );
not ( n58775 , n58774 );
buf ( n58776 , n58771 );
not ( n58777 , n58776 );
and ( n58778 , n58775 , n58777 );
buf ( n58779 , n58765 );
buf ( n58780 , n58737 );
buf ( n58781 , n58755 );
xor ( n58782 , n58780 , n58781 );
buf ( n58783 , n58782 );
buf ( n58784 , n58783 );
xnor ( n58785 , n58779 , n58784 );
buf ( n58786 , n58785 );
buf ( n58787 , n58786 );
not ( n58788 , n58787 );
buf ( n58789 , n56720 );
buf ( n58790 , n56652 );
and ( n58791 , n58789 , n58790 );
not ( n58792 , n56720 );
buf ( n58793 , n58792 );
buf ( n58794 , n55201 );
and ( n58795 , n58793 , n58794 );
nor ( n58796 , n58791 , n58795 );
buf ( n58797 , n58796 );
buf ( n58798 , n58797 );
not ( n58799 , n58798 );
buf ( n58800 , n58799 );
buf ( n58801 , n58800 );
buf ( n58802 , n55180 );
and ( n58803 , n58801 , n58802 );
buf ( n58804 , n56828 );
not ( n58805 , n58804 );
buf ( n58806 , n58805 );
buf ( n58807 , n58806 );
buf ( n58808 , n56670 );
and ( n58809 , n58807 , n58808 );
nor ( n58810 , n58803 , n58809 );
buf ( n58811 , n58810 );
buf ( n58812 , n58811 );
not ( n58813 , n54210 );
not ( n58814 , n55086 );
or ( n58815 , n58813 , n58814 );
not ( n58816 , n55089 );
nand ( n58817 , n58815 , n58816 );
not ( n58818 , n55091 );
nand ( n58819 , n58818 , n54234 );
nor ( n58820 , n58817 , n58819 );
not ( n58821 , n58820 );
nand ( n58822 , n58817 , n58819 );
nand ( n58823 , n58821 , n58822 );
buf ( n58824 , n58823 );
buf ( n58825 , n55132 );
and ( n58826 , n58824 , n58825 );
buf ( n58827 , n58747 );
buf ( n58828 , n55156 );
and ( n58829 , n58827 , n58828 );
nor ( n58830 , n58826 , n58829 );
buf ( n58831 , n58830 );
buf ( n58832 , n58831 );
xor ( n58833 , n58812 , n58832 );
not ( n58834 , n58744 );
nand ( n58835 , n58834 , n58746 );
buf ( n58836 , n58835 );
buf ( n58837 , n56652 );
and ( n58838 , n58836 , n58837 );
buf ( n58839 , n58747 );
not ( n58840 , n58839 );
buf ( n58841 , n58840 );
buf ( n58842 , n58841 );
buf ( n58843 , n55201 );
and ( n58844 , n58842 , n58843 );
nor ( n58845 , n58838 , n58844 );
buf ( n58846 , n58845 );
buf ( n58847 , n58846 );
buf ( n58848 , n56664 );
or ( n58849 , n58847 , n58848 );
buf ( n58850 , n58797 );
buf ( n58851 , n56673 );
or ( n58852 , n58850 , n58851 );
nand ( n58853 , n58849 , n58852 );
buf ( n58854 , n58853 );
buf ( n58855 , n58854 );
nand ( n58856 , n54210 , n58816 );
xnor ( n58857 , n55086 , n58856 );
not ( n58858 , n58857 );
buf ( n58859 , n58858 );
buf ( n58860 , n56589 );
or ( n58861 , n58859 , n58860 );
not ( n58862 , n58823 );
buf ( n58863 , n58862 );
buf ( n58864 , n56598 );
or ( n58865 , n58863 , n58864 );
nand ( n58866 , n58861 , n58865 );
buf ( n58867 , n58866 );
buf ( n58868 , n58867 );
and ( n58869 , n58855 , n58868 );
buf ( n58870 , n58854 );
not ( n58871 , n58870 );
buf ( n58872 , n58867 );
not ( n58873 , n58872 );
and ( n58874 , n58871 , n58873 );
not ( n58875 , n15117 );
buf ( n58876 , n58875 );
buf ( n58877 , n15265 );
and ( n58878 , n58876 , n58877 );
not ( n58879 , n58876 );
not ( n58880 , n15265 );
buf ( n58881 , n58880 );
and ( n58882 , n58879 , n58881 );
nor ( n58883 , n58878 , n58882 );
buf ( n58884 , n58883 );
buf ( n58885 , n58884 );
not ( n58886 , n58885 );
buf ( n58887 , n58886 );
buf ( n58888 , n58887 );
not ( n58889 , n58888 );
buf ( n58890 , n58889 );
buf ( n58891 , n58890 );
buf ( n58892 , n56789 );
not ( n58893 , n58892 );
buf ( n58894 , n58893 );
buf ( n58895 , n58894 );
not ( n58896 , n58895 );
buf ( n58897 , n58896 );
buf ( n58898 , n58897 );
nor ( n58899 , n58891 , n58898 );
buf ( n58900 , n58899 );
buf ( n58901 , n58900 );
not ( n58902 , n58901 );
buf ( n58903 , n56786 );
buf ( n58904 , n58875 );
or ( n58905 , n58903 , n58904 );
buf ( n58906 , n56786 );
buf ( n58907 , n58875 );
nand ( n58908 , n58906 , n58907 );
buf ( n58909 , n58908 );
buf ( n58910 , n58909 );
buf ( n58911 , n58884 );
nand ( n58912 , n58905 , n58910 , n58911 );
buf ( n58913 , n58912 );
buf ( n58914 , n58913 );
not ( n58915 , n58914 );
buf ( n58916 , n58915 );
buf ( n58917 , n58916 );
buf ( n58918 , n58894 );
nand ( n58919 , n58917 , n58918 );
buf ( n58920 , n58919 );
buf ( n58921 , n58920 );
nand ( n58922 , n58902 , n58921 );
buf ( n58923 , n58922 );
buf ( n58924 , n58923 );
nor ( n58925 , n58874 , n58924 );
buf ( n58926 , n58925 );
buf ( n58927 , n58926 );
nor ( n58928 , n58869 , n58927 );
buf ( n58929 , n58928 );
buf ( n58930 , n58929 );
and ( n58931 , n58833 , n58930 );
and ( n58932 , n58812 , n58832 );
or ( n58933 , n58931 , n58932 );
buf ( n58934 , n58933 );
buf ( n58935 , n58934 );
not ( n58936 , n58935 );
and ( n58937 , n58788 , n58936 );
buf ( n58938 , n58786 );
buf ( n58939 , n58934 );
and ( n58940 , n58938 , n58939 );
buf ( n58941 , n58715 );
buf ( n58942 , n58734 );
and ( n58943 , n58941 , n58942 );
buf ( n58944 , n58737 );
nor ( n58945 , n58943 , n58944 );
buf ( n58946 , n58945 );
buf ( n58947 , n58946 );
not ( n58948 , n58947 );
buf ( n58949 , n58948 );
buf ( n58950 , n58949 );
buf ( n58951 , n56582 );
buf ( n58952 , n56641 );
and ( n58953 , n58951 , n58952 );
buf ( n58954 , n56585 );
buf ( n58955 , n56631 );
and ( n58956 , n58954 , n58955 );
nor ( n58957 , n58953 , n58956 );
buf ( n58958 , n58957 );
buf ( n58959 , n58958 );
buf ( n58960 , n56626 );
or ( n58961 , n58959 , n58960 );
buf ( n58962 , n58707 );
buf ( n58963 , n56639 );
or ( n58964 , n58962 , n58963 );
nand ( n58965 , n58961 , n58964 );
buf ( n58966 , n58965 );
buf ( n58967 , n58966 );
buf ( n58968 , n55113 );
buf ( n58969 , n58721 );
and ( n58970 , n58968 , n58969 );
buf ( n58971 , n56655 );
buf ( n58972 , n58718 );
and ( n58973 , n58971 , n58972 );
nor ( n58974 , n58970 , n58973 );
buf ( n58975 , n58974 );
buf ( n58976 , n58975 );
buf ( n58977 , n56799 );
or ( n58978 , n58976 , n58977 );
buf ( n58979 , n58728 );
buf ( n58980 , n56811 );
not ( n58981 , n58980 );
buf ( n58982 , n58981 );
buf ( n58983 , n58982 );
or ( n58984 , n58979 , n58983 );
nand ( n58985 , n58978 , n58984 );
buf ( n58986 , n58985 );
buf ( n58987 , n58986 );
xor ( n58988 , n58967 , n58987 );
buf ( n58989 , n55152 );
buf ( n58990 , n58897 );
and ( n58991 , n58989 , n58990 );
buf ( n58992 , n55205 );
buf ( n58993 , n58894 );
and ( n58994 , n58992 , n58993 );
nor ( n58995 , n58991 , n58994 );
buf ( n58996 , n58995 );
buf ( n58997 , n58996 );
not ( n58998 , n58997 );
buf ( n58999 , n58998 );
buf ( n59000 , n58999 );
buf ( n59001 , n58916 );
and ( n59002 , n59000 , n59001 );
buf ( n59003 , n58900 );
nor ( n59004 , n59002 , n59003 );
buf ( n59005 , n59004 );
buf ( n59006 , n59005 );
not ( n59007 , n55084 );
nand ( n59008 , n59007 , n54469 );
xnor ( n59009 , n55230 , n59008 );
buf ( n59010 , n59009 );
buf ( n59011 , n55132 );
and ( n59012 , n59010 , n59011 );
buf ( n59013 , n58857 );
buf ( n59014 , n55156 );
and ( n59015 , n59013 , n59014 );
nor ( n59016 , n59012 , n59015 );
buf ( n59017 , n59016 );
buf ( n59018 , n59017 );
nand ( n59019 , n59006 , n59018 );
buf ( n59020 , n59019 );
buf ( n59021 , n59020 );
and ( n59022 , n58988 , n59021 );
and ( n59023 , n58967 , n58987 );
or ( n59024 , n59022 , n59023 );
buf ( n59025 , n59024 );
buf ( n59026 , n59025 );
and ( n59027 , n58950 , n59026 );
buf ( n59028 , n58949 );
not ( n59029 , n59028 );
buf ( n59030 , n59025 );
not ( n59031 , n59030 );
and ( n59032 , n59029 , n59031 );
xor ( n59033 , n58812 , n58832 );
xor ( n59034 , n59033 , n58930 );
buf ( n59035 , n59034 );
buf ( n59036 , n59035 );
nor ( n59037 , n59032 , n59036 );
buf ( n59038 , n59037 );
buf ( n59039 , n59038 );
nor ( n59040 , n59027 , n59039 );
buf ( n59041 , n59040 );
buf ( n59042 , n59041 );
nor ( n59043 , n58940 , n59042 );
buf ( n59044 , n59043 );
buf ( n59045 , n59044 );
nor ( n59046 , n58937 , n59045 );
buf ( n59047 , n59046 );
buf ( n59048 , n59047 );
nor ( n59049 , n58778 , n59048 );
buf ( n59050 , n59049 );
buf ( n59051 , n59050 );
nor ( n59052 , n58773 , n59051 );
buf ( n59053 , n59052 );
or ( n59054 , n58693 , n59053 );
nand ( n59055 , n58692 , n59054 );
nand ( n59056 , n58661 , n59055 );
nand ( n59057 , n58660 , n59056 );
nand ( n59058 , n58622 , n59057 );
nand ( n59059 , n58601 , n58621 );
nand ( n59060 , n59058 , n59059 );
buf ( n59061 , n59060 );
nand ( n59062 , n58593 , n59061 );
buf ( n59063 , n59062 );
nand ( n59064 , n58588 , n59063 );
buf ( n59065 , n59064 );
xor ( n59066 , n58522 , n59065 );
xor ( n59067 , n57687 , n57691 );
xor ( n59068 , n59067 , n57761 );
buf ( n59069 , n59068 );
buf ( n59070 , n59069 );
and ( n59071 , n59066 , n59070 );
and ( n59072 , n58522 , n59065 );
or ( n59073 , n59071 , n59072 );
buf ( n59074 , n59073 );
nand ( n59075 , n58497 , n59074 );
nand ( n59076 , n58491 , n59075 );
buf ( n59077 , n59076 );
nand ( n59078 , n58474 , n59077 );
buf ( n59079 , n59078 );
buf ( n59080 , n59079 );
nand ( n59081 , n58469 , n59080 );
buf ( n59082 , n59081 );
buf ( n59083 , n59082 );
nand ( n59084 , n58421 , n59083 );
buf ( n59085 , n59084 );
buf ( n59086 , n59085 );
buf ( n59087 , n58414 );
not ( n59088 , n59087 );
buf ( n59089 , n58418 );
not ( n59090 , n59089 );
buf ( n59091 , n59090 );
buf ( n59092 , n59091 );
nand ( n59093 , n59088 , n59092 );
buf ( n59094 , n59093 );
buf ( n59095 , n59094 );
nand ( n59096 , n59086 , n59095 );
buf ( n59097 , n59096 );
buf ( n59098 , n59097 );
and ( n59099 , n58401 , n59098 );
and ( n59100 , n58396 , n58400 );
or ( n59101 , n59099 , n59100 );
buf ( n59102 , n59101 );
buf ( n59103 , n59102 );
buf ( n59104 , n59103 );
buf ( n59105 , n59104 );
xor ( n59106 , n56096 , n56999 );
xor ( n59107 , n59106 , n57006 );
not ( n59108 , n59107 );
and ( n59109 , n57415 , n57420 );
not ( n59110 , n57415 );
and ( n59111 , n59110 , n57421 );
nor ( n59112 , n59109 , n59111 );
and ( n59113 , n59112 , n57901 );
not ( n59114 , n59112 );
not ( n59115 , n57901 );
and ( n59116 , n59114 , n59115 );
nor ( n59117 , n59113 , n59116 );
nand ( n59118 , n59108 , n59117 );
and ( n59119 , n59105 , n59118 );
not ( n59120 , n59107 );
nor ( n59121 , n59120 , n59117 );
nor ( n59122 , n59119 , n59121 );
buf ( n59123 , n59122 );
nand ( n59124 , n57952 , n59123 );
buf ( n59125 , n59124 );
nand ( n59126 , n57948 , n59125 );
not ( n59127 , n59126 );
buf ( n59128 , n59127 );
nand ( n59129 , n57043 , n59128 );
buf ( n59130 , n59129 );
buf ( n59131 , n59130 );
not ( n59132 , n59131 );
buf ( n59133 , n59132 );
not ( n59134 , n59082 );
not ( n59135 , n59134 );
not ( n59136 , n58414 );
not ( n59137 , n59136 );
or ( n59138 , n59135 , n59137 );
nand ( n59139 , n58414 , n59082 );
nand ( n59140 , n59138 , n59139 );
and ( n59141 , n59140 , n59091 );
not ( n59142 , n59140 );
buf ( n59143 , n59091 );
not ( n59144 , n59143 );
buf ( n59145 , n59144 );
and ( n59146 , n59142 , n59145 );
nor ( n59147 , n59141 , n59146 );
buf ( n59148 , n59076 );
buf ( n59149 , n58426 );
and ( n59150 , n59148 , n59149 );
not ( n59151 , n59148 );
buf ( n59152 , n58423 );
and ( n59153 , n59151 , n59152 );
nor ( n59154 , n59150 , n59153 );
buf ( n59155 , n59154 );
xnor ( n59156 , n58463 , n59155 );
buf ( n59157 , n59156 );
buf ( n59158 , n57488 );
buf ( n59159 , n57463 );
and ( n59160 , n59158 , n59159 );
not ( n59161 , n59158 );
buf ( n59162 , n57460 );
and ( n59163 , n59161 , n59162 );
nor ( n59164 , n59160 , n59163 );
buf ( n59165 , n59164 );
xor ( n59166 , n57770 , n59165 );
buf ( n59167 , n59166 );
xor ( n59168 , n57784 , n57788 );
xor ( n59169 , n59168 , n57887 );
buf ( n59170 , n59169 );
buf ( n59171 , n59170 );
xor ( n59172 , n59167 , n59171 );
buf ( n59173 , n48868 );
not ( n59174 , n59173 );
buf ( n59175 , n57476 );
not ( n59176 , n59175 );
or ( n59177 , n59174 , n59176 );
buf ( n59178 , n48808 );
not ( n59179 , n59178 );
buf ( n59180 , n39280 );
not ( n59181 , n59180 );
or ( n59182 , n59179 , n59181 );
buf ( n59183 , n42929 );
buf ( n59184 , n48821 );
nand ( n59185 , n59183 , n59184 );
buf ( n59186 , n59185 );
buf ( n59187 , n59186 );
nand ( n59188 , n59182 , n59187 );
buf ( n59189 , n59188 );
buf ( n59190 , n59189 );
buf ( n59191 , n48855 );
nand ( n59192 , n59190 , n59191 );
buf ( n59193 , n59192 );
buf ( n59194 , n59193 );
nand ( n59195 , n59177 , n59194 );
buf ( n59196 , n59195 );
not ( n59197 , n59196 );
not ( n59198 , n44708 );
not ( n59199 , n44533 );
not ( n59200 , n47626 );
or ( n59201 , n59199 , n59200 );
not ( n59202 , n37782 );
buf ( n59203 , n59202 );
buf ( n59204 , n59203 );
buf ( n59205 , n44530 );
nand ( n59206 , n59204 , n59205 );
buf ( n59207 , n59206 );
nand ( n59208 , n59201 , n59207 );
not ( n59209 , n59208 );
or ( n59210 , n59198 , n59209 );
not ( n59211 , n57823 );
nand ( n59212 , n59211 , n44496 );
nand ( n59213 , n59210 , n59212 );
not ( n59214 , n59213 );
not ( n59215 , n46225 );
not ( n59216 , n51872 );
not ( n59217 , n45750 );
or ( n59218 , n59216 , n59217 );
buf ( n59219 , n43625 );
not ( n59220 , n59219 );
buf ( n59221 , n59220 );
nand ( n59222 , n59221 , n53492 );
nand ( n59223 , n59218 , n59222 );
not ( n59224 , n59223 );
or ( n59225 , n59215 , n59224 );
nand ( n59226 , n58514 , n46246 );
nand ( n59227 , n59225 , n59226 );
not ( n59228 , n59227 );
or ( n59229 , n59214 , n59228 );
not ( n59230 , n59213 );
buf ( n59231 , n59230 );
not ( n59232 , n59231 );
not ( n59233 , n59227 );
buf ( n59234 , n59233 );
not ( n59235 , n59234 );
or ( n59236 , n59232 , n59235 );
not ( n59237 , n42315 );
not ( n59238 , n57705 );
or ( n59239 , n59237 , n59238 );
buf ( n59240 , n42260 );
not ( n59241 , n59240 );
buf ( n59242 , n59241 );
buf ( n59243 , n59242 );
not ( n59244 , n59243 );
buf ( n59245 , n42425 );
not ( n59246 , n59245 );
or ( n59247 , n59244 , n59246 );
buf ( n59248 , n43446 );
buf ( n59249 , n42263 );
nand ( n59250 , n59248 , n59249 );
buf ( n59251 , n59250 );
buf ( n59252 , n59251 );
nand ( n59253 , n59247 , n59252 );
buf ( n59254 , n59253 );
buf ( n59255 , n59254 );
buf ( n59256 , n42252 );
nand ( n59257 , n59255 , n59256 );
buf ( n59258 , n59257 );
nand ( n59259 , n59239 , n59258 );
not ( n59260 , n41993 );
not ( n59261 , n42471 );
or ( n59262 , n59260 , n59261 );
buf ( n59263 , n38979 );
buf ( n59264 , n43966 );
nand ( n59265 , n59263 , n59264 );
buf ( n59266 , n59265 );
nand ( n59267 , n59262 , n59266 );
buf ( n59268 , n59267 );
not ( n59269 , n59268 );
buf ( n59270 , n47050 );
not ( n59271 , n59270 );
or ( n59272 , n59269 , n59271 );
buf ( n59273 , n57573 );
buf ( n59274 , n52595 );
nand ( n59275 , n59273 , n59274 );
buf ( n59276 , n59275 );
buf ( n59277 , n59276 );
nand ( n59278 , n59272 , n59277 );
buf ( n59279 , n59278 );
not ( n59280 , n59279 );
not ( n59281 , n42339 );
not ( n59282 , n58157 );
or ( n59283 , n59281 , n59282 );
buf ( n59284 , n42343 );
not ( n59285 , n59284 );
buf ( n59286 , n41915 );
not ( n59287 , n59286 );
or ( n59288 , n59285 , n59287 );
buf ( n59289 , n47001 );
not ( n59290 , n59289 );
buf ( n59291 , n59290 );
buf ( n59292 , n59291 );
buf ( n59293 , n46855 );
nand ( n59294 , n59292 , n59293 );
buf ( n59295 , n59294 );
buf ( n59296 , n59295 );
nand ( n59297 , n59288 , n59296 );
buf ( n59298 , n59297 );
buf ( n59299 , n59298 );
buf ( n59300 , n42378 );
nand ( n59301 , n59299 , n59300 );
buf ( n59302 , n59301 );
nand ( n59303 , n59283 , n59302 );
not ( n59304 , n59303 );
or ( n59305 , n59280 , n59304 );
or ( n59306 , n59279 , n59303 );
xor ( n59307 , n58177 , n58195 );
xor ( n59308 , n59307 , n58221 );
buf ( n59309 , n59308 );
nand ( n59310 , n59306 , n59309 );
nand ( n59311 , n59305 , n59310 );
xor ( n59312 , n59259 , n59311 );
buf ( n59313 , n58247 );
buf ( n59314 , n42668 );
nand ( n59315 , n59313 , n59314 );
buf ( n59316 , n59315 );
buf ( n59317 , n25228 );
not ( n59318 , n59317 );
buf ( n59319 , n42119 );
not ( n59320 , n59319 );
or ( n59321 , n59318 , n59320 );
buf ( n59322 , n28305 );
buf ( n59323 , n25227 );
nand ( n59324 , n59322 , n59323 );
buf ( n59325 , n59324 );
buf ( n59326 , n59325 );
nand ( n59327 , n59321 , n59326 );
buf ( n59328 , n59327 );
nand ( n59329 , n59328 , n42712 );
nand ( n59330 , n59316 , n59329 );
not ( n59331 , n59330 );
not ( n59332 , n59331 );
not ( n59333 , n38404 );
and ( n59334 , n42865 , n47068 );
not ( n59335 , n42865 );
and ( n59336 , n59335 , n42414 );
nor ( n59337 , n59334 , n59336 );
not ( n59338 , n59337 );
or ( n59339 , n59333 , n59338 );
nand ( n59340 , n58130 , n38380 );
nand ( n59341 , n59339 , n59340 );
not ( n59342 , n59341 );
not ( n59343 , n59342 );
or ( n59344 , n59332 , n59343 );
buf ( n59345 , n41736 );
not ( n59346 , n59345 );
buf ( n59347 , n51804 );
not ( n59348 , n59347 );
or ( n59349 , n59346 , n59348 );
buf ( n59350 , n25159 );
buf ( n59351 , n41733 );
nand ( n59352 , n59350 , n59351 );
buf ( n59353 , n59352 );
buf ( n59354 , n59353 );
nand ( n59355 , n59349 , n59354 );
buf ( n59356 , n59355 );
buf ( n59357 , n59356 );
not ( n59358 , n59357 );
buf ( n59359 , n50128 );
not ( n59360 , n59359 );
or ( n59361 , n59358 , n59360 );
buf ( n59362 , n58638 );
buf ( n59363 , n42564 );
nand ( n59364 , n59362 , n59363 );
buf ( n59365 , n59364 );
buf ( n59366 , n59365 );
nand ( n59367 , n59361 , n59366 );
buf ( n59368 , n59367 );
buf ( n59369 , n59368 );
buf ( n59370 , n42008 );
not ( n59371 , n59370 );
buf ( n59372 , n47857 );
not ( n59373 , n59372 );
or ( n59374 , n59371 , n59373 );
buf ( n59375 , n24092 );
buf ( n59376 , n42017 );
nand ( n59377 , n59375 , n59376 );
buf ( n59378 , n59377 );
buf ( n59379 , n59378 );
nand ( n59380 , n59374 , n59379 );
buf ( n59381 , n59380 );
buf ( n59382 , n59381 );
not ( n59383 , n59382 );
buf ( n59384 , n50608 );
not ( n59385 , n59384 );
or ( n59386 , n59383 , n59385 );
buf ( n59387 , n58208 );
buf ( n59388 , n39983 );
nand ( n59389 , n59387 , n59388 );
buf ( n59390 , n59389 );
buf ( n59391 , n59390 );
nand ( n59392 , n59386 , n59391 );
buf ( n59393 , n59392 );
buf ( n59394 , n59393 );
xor ( n59395 , n59369 , n59394 );
buf ( n59396 , n48671 );
not ( n59397 , n59396 );
buf ( n59398 , n58651 );
not ( n59399 , n59398 );
or ( n59400 , n59397 , n59399 );
buf ( n59401 , n58107 );
not ( n59402 , n59401 );
buf ( n59403 , n59402 );
buf ( n59404 , n59403 );
not ( n59405 , n59404 );
buf ( n59406 , n43362 );
not ( n59407 , n59406 );
or ( n59408 , n59405 , n59407 );
buf ( n59409 , n50624 );
buf ( n59410 , n41660 );
nand ( n59411 , n59409 , n59410 );
buf ( n59412 , n59411 );
buf ( n59413 , n59412 );
nand ( n59414 , n59408 , n59413 );
buf ( n59415 , n59414 );
buf ( n59416 , n59415 );
buf ( n59417 , n50982 );
nand ( n59418 , n59416 , n59417 );
buf ( n59419 , n59418 );
buf ( n59420 , n59419 );
nand ( n59421 , n59400 , n59420 );
buf ( n59422 , n59421 );
buf ( n59423 , n59422 );
and ( n59424 , n59395 , n59423 );
and ( n59425 , n59369 , n59394 );
or ( n59426 , n59424 , n59425 );
buf ( n59427 , n59426 );
nand ( n59428 , n59344 , n59427 );
not ( n59429 , n59329 );
not ( n59430 , n59316 );
or ( n59431 , n59429 , n59430 );
nand ( n59432 , n59431 , n59341 );
nand ( n59433 , n59428 , n59432 );
and ( n59434 , n59312 , n59433 );
and ( n59435 , n59259 , n59311 );
or ( n59436 , n59434 , n59435 );
buf ( n59437 , n59436 );
nand ( n59438 , n59236 , n59437 );
buf ( n59439 , n59438 );
nand ( n59440 , n59229 , n59439 );
not ( n59441 , n59440 );
or ( n59442 , n59197 , n59441 );
or ( n59443 , n59440 , n59196 );
and ( n59444 , n58095 , n58171 );
not ( n59445 , n58095 );
and ( n59446 , n59445 , n58170 );
nor ( n59447 , n59444 , n59446 );
xor ( n59448 , n59447 , n58298 );
not ( n59449 , n59448 );
buf ( n59450 , n59449 );
not ( n59451 , n59450 );
xor ( n59452 , n57709 , n57729 );
xor ( n59453 , n59452 , n57754 );
buf ( n59454 , n59453 );
not ( n59455 , n59454 );
or ( n59456 , n59451 , n59455 );
buf ( n59457 , n59449 );
buf ( n59458 , n59453 );
or ( n59459 , n59457 , n59458 );
buf ( n59460 , n58289 );
buf ( n59461 , n58255 );
xor ( n59462 , n59460 , n59461 );
buf ( n59463 , n58225 );
xor ( n59464 , n59462 , n59463 );
buf ( n59465 , n59464 );
buf ( n59466 , n59465 );
not ( n59467 , n59466 );
buf ( n59468 , n59467 );
not ( n59469 , n59468 );
not ( n59470 , n55881 );
buf ( n59471 , n50060 );
not ( n59472 , n59471 );
buf ( n59473 , n43371 );
not ( n59474 , n59473 );
or ( n59475 , n59472 , n59474 );
buf ( n59476 , n43403 );
buf ( n59477 , n50067 );
nand ( n59478 , n59476 , n59477 );
buf ( n59479 , n59478 );
buf ( n59480 , n59479 );
nand ( n59481 , n59475 , n59480 );
buf ( n59482 , n59481 );
not ( n59483 , n59482 );
or ( n59484 , n59470 , n59483 );
buf ( n59485 , n58021 );
buf ( n59486 , n46172 );
nand ( n59487 , n59485 , n59486 );
buf ( n59488 , n59487 );
nand ( n59489 , n59484 , n59488 );
not ( n59490 , n59489 );
or ( n59491 , n59469 , n59490 );
not ( n59492 , n59465 );
not ( n59493 , n59489 );
not ( n59494 , n59493 );
or ( n59495 , n59492 , n59494 );
buf ( n59496 , n59254 );
buf ( n59497 , n42315 );
nand ( n59498 , n59496 , n59497 );
buf ( n59499 , n59498 );
buf ( n59500 , n59242 );
not ( n59501 , n59500 );
buf ( n59502 , n41799 );
not ( n59503 , n59502 );
or ( n59504 , n59501 , n59503 );
buf ( n59505 , n42398 );
buf ( n59506 , n42263 );
nand ( n59507 , n59505 , n59506 );
buf ( n59508 , n59507 );
buf ( n59509 , n59508 );
nand ( n59510 , n59504 , n59509 );
buf ( n59511 , n59510 );
nand ( n59512 , n59511 , n42252 );
nand ( n59513 , n59499 , n59512 );
buf ( n59514 , n44952 );
not ( n59515 , n59514 );
buf ( n59516 , n41805 );
not ( n59517 , n59516 );
or ( n59518 , n59515 , n59517 );
buf ( n59519 , n41769 );
buf ( n59520 , n44961 );
nand ( n59521 , n59519 , n59520 );
buf ( n59522 , n59521 );
buf ( n59523 , n59522 );
nand ( n59524 , n59518 , n59523 );
buf ( n59525 , n59524 );
not ( n59526 , n59525 );
not ( n59527 , n37397 );
or ( n59528 , n59526 , n59527 );
buf ( n59529 , n58613 );
buf ( n59530 , n42135 );
nand ( n59531 , n59529 , n59530 );
buf ( n59532 , n59531 );
nand ( n59533 , n59528 , n59532 );
nor ( n59534 , n59513 , n59533 );
buf ( n59535 , n58645 );
buf ( n59536 , n58658 );
xor ( n59537 , n59535 , n59536 );
buf ( n59538 , n59055 );
xnor ( n59539 , n59537 , n59538 );
buf ( n59540 , n59539 );
or ( n59541 , n59534 , n59540 );
not ( n59542 , n59512 );
not ( n59543 , n59499 );
or ( n59544 , n59542 , n59543 );
nand ( n59545 , n59544 , n59533 );
nand ( n59546 , n59541 , n59545 );
nand ( n59547 , n59495 , n59546 );
nand ( n59548 , n59491 , n59547 );
buf ( n59549 , n59548 );
nand ( n59550 , n59459 , n59549 );
buf ( n59551 , n59550 );
buf ( n59552 , n59551 );
nand ( n59553 , n59456 , n59552 );
buf ( n59554 , n59553 );
nand ( n59555 , n59443 , n59554 );
nand ( n59556 , n59442 , n59555 );
buf ( n59557 , n59556 );
buf ( n59558 , C0 );
buf ( n59559 , n59558 );
buf ( n59560 , n52456 );
not ( n59561 , n59560 );
buf ( n59562 , n57803 );
not ( n59563 , n59562 );
or ( n59564 , n59561 , n59563 );
buf ( n59565 , n48836 );
not ( n59566 , n59565 );
buf ( n59567 , n47813 );
not ( n59568 , n59567 );
or ( n59569 , n59566 , n59568 );
buf ( n59570 , n45839 );
not ( n59571 , n59570 );
buf ( n59572 , n57174 );
nand ( n59573 , n59571 , n59572 );
buf ( n59574 , n59573 );
buf ( n59575 , n59574 );
nand ( n59576 , n59569 , n59575 );
buf ( n59577 , n59576 );
buf ( n59578 , n59577 );
buf ( n59579 , n51488 );
nand ( n59580 , n59578 , n59579 );
buf ( n59581 , n59580 );
buf ( n59582 , n59581 );
nand ( n59583 , n59564 , n59582 );
buf ( n59584 , n59583 );
buf ( n59585 , n59584 );
xor ( n59586 , n59559 , n59585 );
not ( n59587 , n57874 );
not ( n59588 , n59587 );
not ( n59589 , n57859 );
or ( n59590 , n59588 , n59589 );
nand ( n59591 , n57874 , n57856 );
nand ( n59592 , n59590 , n59591 );
buf ( n59593 , n59592 );
buf ( n59594 , n57828 );
buf ( n59595 , n59594 );
buf ( n59596 , n59595 );
buf ( n59597 , n59596 );
not ( n59598 , n59597 );
buf ( n59599 , n59598 );
buf ( n59600 , n59599 );
and ( n59601 , n59593 , n59600 );
not ( n59602 , n59593 );
buf ( n59603 , n59596 );
and ( n59604 , n59602 , n59603 );
nor ( n59605 , n59601 , n59604 );
buf ( n59606 , n59605 );
buf ( n59607 , n59606 );
and ( n59608 , n59586 , n59607 );
or ( n59609 , n59608 , C0 );
buf ( n59610 , n59609 );
buf ( n59611 , n59610 );
xor ( n59612 , n59557 , n59611 );
xor ( n59613 , n58081 , n58072 );
xnor ( n59614 , n59613 , n58386 );
buf ( n59615 , n59614 );
and ( n59616 , n59612 , n59615 );
and ( n59617 , n59557 , n59611 );
or ( n59618 , n59616 , n59617 );
buf ( n59619 , n59618 );
buf ( n59620 , n59619 );
xor ( n59621 , n59172 , n59620 );
buf ( n59622 , n59621 );
buf ( n59623 , n59622 );
xor ( n59624 , n59157 , n59623 );
xor ( n59625 , n59557 , n59611 );
xor ( n59626 , n59625 , n59615 );
buf ( n59627 , n59626 );
buf ( n59628 , n59627 );
xor ( n59629 , n57876 , n57880 );
xnor ( n59630 , n59629 , n57813 );
buf ( n59631 , n41574 );
not ( n59632 , n59631 );
buf ( n59633 , n58053 );
not ( n59634 , n59633 );
or ( n59635 , n59632 , n59634 );
buf ( n59636 , n41611 );
buf ( n59637 , n42458 );
and ( n59638 , n59636 , n59637 );
not ( n59639 , n59636 );
buf ( n59640 , n42455 );
and ( n59641 , n59639 , n59640 );
nor ( n59642 , n59638 , n59641 );
buf ( n59643 , n59642 );
buf ( n59644 , n59643 );
not ( n59645 , n59644 );
buf ( n59646 , n44267 );
nand ( n59647 , n59645 , n59646 );
buf ( n59648 , n59647 );
buf ( n59649 , n59648 );
nand ( n59650 , n59635 , n59649 );
buf ( n59651 , n59650 );
not ( n59652 , n59651 );
buf ( n59653 , n53539 );
not ( n59654 , n59653 );
buf ( n59655 , n39493 );
not ( n59656 , n59655 );
or ( n59657 , n59654 , n59656 );
buf ( n59658 , n33077 );
buf ( n59659 , n53548 );
nand ( n59660 , n59658 , n59659 );
buf ( n59661 , n59660 );
buf ( n59662 , n59661 );
nand ( n59663 , n59657 , n59662 );
buf ( n59664 , n59663 );
buf ( n59665 , n59664 );
not ( n59666 , n59665 );
buf ( n59667 , n42521 );
not ( n59668 , n59667 );
or ( n59669 , n59666 , n59668 );
buf ( n59670 , n42530 );
buf ( n59671 , n57742 );
nand ( n59672 , n59670 , n59671 );
buf ( n59673 , n59672 );
buf ( n59674 , n59673 );
nand ( n59675 , n59669 , n59674 );
buf ( n59676 , n59675 );
not ( n59677 , n59676 );
or ( n59678 , n59652 , n59677 );
buf ( n59679 , n59651 );
buf ( n59680 , n59676 );
nor ( n59681 , n59679 , n59680 );
buf ( n59682 , n59681 );
buf ( n59683 , n58116 );
buf ( n59684 , n58138 );
xor ( n59685 , n59683 , n59684 );
buf ( n59686 , n58164 );
xnor ( n59687 , n59685 , n59686 );
buf ( n59688 , n59687 );
or ( n59689 , n59682 , n59688 );
nand ( n59690 , n59678 , n59689 );
buf ( n59691 , n59690 );
buf ( n59692 , n48855 );
not ( n59693 , n59692 );
buf ( n59694 , n48808 );
not ( n59695 , n59694 );
buf ( n59696 , n39407 );
not ( n59697 , n59696 );
or ( n59698 , n59695 , n59697 );
buf ( n59699 , n45227 );
buf ( n59700 , n48818 );
nand ( n59701 , n59699 , n59700 );
buf ( n59702 , n59701 );
buf ( n59703 , n59702 );
nand ( n59704 , n59698 , n59703 );
buf ( n59705 , n59704 );
buf ( n59706 , n59705 );
not ( n59707 , n59706 );
or ( n59708 , n59693 , n59707 );
buf ( n59709 , n59189 );
buf ( n59710 , n48868 );
nand ( n59711 , n59709 , n59710 );
buf ( n59712 , n59711 );
buf ( n59713 , n59712 );
nand ( n59714 , n59708 , n59713 );
buf ( n59715 , n59714 );
buf ( n59716 , n59715 );
xor ( n59717 , n59691 , n59716 );
xor ( n59718 , n58034 , n58038 );
xor ( n59719 , n59718 , n58064 );
buf ( n59720 , n59719 );
buf ( n59721 , n59720 );
and ( n59722 , n59717 , n59721 );
and ( n59723 , n59691 , n59716 );
or ( n59724 , n59722 , n59723 );
buf ( n59725 , n59724 );
not ( n59726 , n59725 );
buf ( n59727 , n57976 );
buf ( n59728 , n58004 );
xor ( n59729 , n59727 , n59728 );
buf ( n59730 , n58068 );
xnor ( n59731 , n59729 , n59730 );
buf ( n59732 , n59731 );
nand ( n59733 , n59726 , n59732 );
not ( n59734 , n59733 );
xor ( n59735 , n58303 , n58321 );
xor ( n59736 , n59735 , n58382 );
buf ( n59737 , n59736 );
not ( n59738 , n59737 );
or ( n59739 , n59734 , n59738 );
buf ( n59740 , n59732 );
not ( n59741 , n59740 );
buf ( n59742 , n59741 );
nand ( n59743 , n59742 , n59725 );
nand ( n59744 , n59739 , n59743 );
and ( n59745 , n59630 , n59744 );
not ( n59746 , n59630 );
not ( n59747 , n59744 );
and ( n59748 , n59746 , n59747 );
nor ( n59749 , n59745 , n59748 );
xor ( n59750 , n58430 , n58450 );
xor ( n59751 , n59750 , n58460 );
and ( n59752 , n59749 , n59751 );
not ( n59753 , n59749 );
not ( n59754 , n59751 );
and ( n59755 , n59753 , n59754 );
nor ( n59756 , n59752 , n59755 );
buf ( n59757 , n59756 );
or ( n59758 , n59628 , n59757 );
xor ( n59759 , n59559 , n59585 );
xor ( n59760 , n59759 , n59607 );
buf ( n59761 , n59760 );
not ( n59762 , n59060 );
and ( n59763 , n59762 , n58532 );
not ( n59764 , n59762 );
and ( n59765 , n59764 , n58533 );
nor ( n59766 , n59763 , n59765 );
buf ( n59767 , n59766 );
buf ( n59768 , n58586 );
and ( n59769 , n59767 , n59768 );
not ( n59770 , n59767 );
buf ( n59771 , n58583 );
and ( n59772 , n59770 , n59771 );
nor ( n59773 , n59769 , n59772 );
buf ( n59774 , n59773 );
buf ( n59775 , n59774 );
not ( n59776 , n59775 );
buf ( n59777 , n59776 );
buf ( n59778 , n59777 );
not ( n59779 , n59778 );
not ( n59780 , n59436 );
not ( n59781 , n59230 );
not ( n59782 , n59227 );
or ( n59783 , n59781 , n59782 );
or ( n59784 , n59227 , n59230 );
nand ( n59785 , n59783 , n59784 );
not ( n59786 , n59785 );
or ( n59787 , n59780 , n59786 );
or ( n59788 , n59785 , n59436 );
nand ( n59789 , n59787 , n59788 );
buf ( n59790 , n59789 );
not ( n59791 , n59790 );
or ( n59792 , n59779 , n59791 );
buf ( n59793 , n46912 );
not ( n59794 , n59793 );
buf ( n59795 , n46875 );
not ( n59796 , n59795 );
buf ( n59797 , n43879 );
not ( n59798 , n59797 );
or ( n59799 , n59796 , n59798 );
buf ( n59800 , n37264 );
buf ( n59801 , n46887 );
nand ( n59802 , n59800 , n59801 );
buf ( n59803 , n59802 );
buf ( n59804 , n59803 );
nand ( n59805 , n59799 , n59804 );
buf ( n59806 , n59805 );
buf ( n59807 , n59806 );
not ( n59808 , n59807 );
or ( n59809 , n59794 , n59808 );
buf ( n59810 , n46875 );
not ( n59811 , n59810 );
buf ( n59812 , n43224 );
not ( n59813 , n59812 );
or ( n59814 , n59811 , n59813 );
buf ( n59815 , n43224 );
buf ( n59816 , n46875 );
or ( n59817 , n59815 , n59816 );
buf ( n59818 , n59817 );
buf ( n59819 , n59818 );
nand ( n59820 , n59814 , n59819 );
buf ( n59821 , n59820 );
buf ( n59822 , n59821 );
buf ( n59823 , n47331 );
nand ( n59824 , n59822 , n59823 );
buf ( n59825 , n59824 );
buf ( n59826 , n59825 );
nand ( n59827 , n59809 , n59826 );
buf ( n59828 , n59827 );
not ( n59829 , n59468 );
not ( n59830 , n59493 );
or ( n59831 , n59829 , n59830 );
buf ( n59832 , n59465 );
buf ( n59833 , n59489 );
nand ( n59834 , n59832 , n59833 );
buf ( n59835 , n59834 );
nand ( n59836 , n59831 , n59835 );
xor ( n59837 , n59836 , n59546 );
xor ( n59838 , n59828 , n59837 );
not ( n59839 , n36085 );
buf ( n59840 , n59839 );
not ( n59841 , n59840 );
buf ( n59842 , n36920 );
not ( n59843 , n59842 );
or ( n59844 , n59841 , n59843 );
buf ( n59845 , n39475 );
nand ( n59846 , n59844 , n59845 );
buf ( n59847 , n59846 );
buf ( n59848 , n59847 );
not ( n59849 , n59848 );
buf ( n59850 , n36085 );
not ( n59851 , n59850 );
buf ( n59852 , n36923 );
not ( n59853 , n59852 );
or ( n59854 , n59851 , n59853 );
buf ( n59855 , n12481 );
nand ( n59856 , n59854 , n59855 );
buf ( n59857 , n59856 );
buf ( n59858 , n59857 );
nand ( n59859 , n59849 , n59858 );
buf ( n59860 , n59859 );
not ( n59861 , n59860 );
xor ( n59862 , n59369 , n59394 );
xor ( n59863 , n59862 , n59423 );
buf ( n59864 , n59863 );
buf ( n59865 , n59864 );
not ( n59866 , n59865 );
buf ( n59867 , n59866 );
not ( n59868 , n59867 );
or ( n59869 , n59861 , n59868 );
buf ( n59870 , n58696 );
buf ( n59871 , n58771 );
xor ( n59872 , n59870 , n59871 );
buf ( n59873 , n59872 );
buf ( n59874 , n59873 );
not ( n59875 , n59874 );
buf ( n59876 , n59047 );
not ( n59877 , n59876 );
or ( n59878 , n59875 , n59877 );
buf ( n59879 , n59047 );
buf ( n59880 , n59873 );
or ( n59881 , n59879 , n59880 );
nand ( n59882 , n59878 , n59881 );
buf ( n59883 , n59882 );
buf ( n59884 , n59883 );
buf ( n59885 , n13653 );
not ( n59886 , n59885 );
buf ( n59887 , n54067 );
not ( n59888 , n59887 );
or ( n59889 , n59886 , n59888 );
buf ( n59890 , n58632 );
buf ( n59891 , n58185 );
nand ( n59892 , n59890 , n59891 );
buf ( n59893 , n59892 );
buf ( n59894 , n59893 );
nand ( n59895 , n59889 , n59894 );
buf ( n59896 , n59895 );
buf ( n59897 , n59896 );
not ( n59898 , n59897 );
buf ( n59899 , n43935 );
not ( n59900 , n59899 );
or ( n59901 , n59898 , n59900 );
buf ( n59902 , n58678 );
buf ( n59903 , n53649 );
nand ( n59904 , n59902 , n59903 );
buf ( n59905 , n59904 );
buf ( n59906 , n59905 );
nand ( n59907 , n59901 , n59906 );
buf ( n59908 , n59907 );
buf ( n59909 , n59908 );
xor ( n59910 , n59884 , n59909 );
buf ( n59911 , n48671 );
not ( n59912 , n59911 );
buf ( n59913 , n59415 );
not ( n59914 , n59913 );
or ( n59915 , n59912 , n59914 );
not ( n59916 , n42072 );
not ( n59917 , n59403 );
or ( n59918 , n59916 , n59917 );
buf ( n59919 , n56342 );
not ( n59920 , n59919 );
buf ( n59921 , n41660 );
nand ( n59922 , n59920 , n59921 );
buf ( n59923 , n59922 );
nand ( n59924 , n59918 , n59923 );
buf ( n59925 , n59924 );
buf ( n59926 , n50979 );
not ( n59927 , n59926 );
buf ( n59928 , n59927 );
buf ( n59929 , n59928 );
nand ( n59930 , n59925 , n59929 );
buf ( n59931 , n59930 );
buf ( n59932 , n59931 );
nand ( n59933 , n59915 , n59932 );
buf ( n59934 , n59933 );
buf ( n59935 , n59934 );
xor ( n59936 , n59910 , n59935 );
buf ( n59937 , n59936 );
not ( n59938 , n59937 );
buf ( n59939 , n59041 );
not ( n59940 , n59939 );
buf ( n59941 , n58786 );
buf ( n59942 , n58934 );
xor ( n59943 , n59941 , n59942 );
buf ( n59944 , n59943 );
buf ( n59945 , n59944 );
not ( n59946 , n59945 );
or ( n59947 , n59940 , n59946 );
buf ( n59948 , n59944 );
buf ( n59949 , n59041 );
or ( n59950 , n59948 , n59949 );
nand ( n59951 , n59947 , n59950 );
buf ( n59952 , n59951 );
buf ( n59953 , n59952 );
buf ( n59954 , n59035 );
not ( n59955 , n59954 );
buf ( n59956 , n59025 );
buf ( n59957 , n58949 );
and ( n59958 , n59956 , n59957 );
not ( n59959 , n59956 );
buf ( n59960 , n58946 );
and ( n59961 , n59959 , n59960 );
nor ( n59962 , n59958 , n59961 );
buf ( n59963 , n59962 );
buf ( n59964 , n59963 );
not ( n59965 , n59964 );
or ( n59966 , n59955 , n59965 );
buf ( n59967 , n59963 );
buf ( n59968 , n59035 );
or ( n59969 , n59967 , n59968 );
nand ( n59970 , n59966 , n59969 );
buf ( n59971 , n59970 );
buf ( n59972 , n59971 );
buf ( n59973 , n56720 );
buf ( n59974 , n56641 );
and ( n59975 , n59973 , n59974 );
buf ( n59976 , n58792 );
buf ( n59977 , n56631 );
and ( n59978 , n59976 , n59977 );
nor ( n59979 , n59975 , n59978 );
buf ( n59980 , n59979 );
buf ( n59981 , n59980 );
buf ( n59982 , n56626 );
or ( n59983 , n59981 , n59982 );
buf ( n59984 , n58958 );
buf ( n59985 , n56639 );
or ( n59986 , n59984 , n59985 );
nand ( n59987 , n59983 , n59986 );
buf ( n59988 , n59987 );
buf ( n59989 , n59988 );
buf ( n59990 , n58699 );
buf ( n59991 , n58721 );
and ( n59992 , n59990 , n59991 );
buf ( n59993 , n56594 );
buf ( n59994 , n58718 );
and ( n59995 , n59993 , n59994 );
nor ( n59996 , n59992 , n59995 );
buf ( n59997 , n59996 );
buf ( n59998 , n59997 );
buf ( n59999 , n56799 );
or ( n60000 , n59998 , n59999 );
buf ( n60001 , n58975 );
buf ( n60002 , n58982 );
or ( n60003 , n60001 , n60002 );
nand ( n60004 , n60000 , n60003 );
buf ( n60005 , n60004 );
buf ( n60006 , n60005 );
xor ( n60007 , n59989 , n60006 );
buf ( n60008 , n58823 );
buf ( n60009 , n56652 );
and ( n60010 , n60008 , n60009 );
buf ( n60011 , n58862 );
buf ( n60012 , n55201 );
and ( n60013 , n60011 , n60012 );
nor ( n60014 , n60010 , n60013 );
buf ( n60015 , n60014 );
buf ( n60016 , n60015 );
buf ( n60017 , n56664 );
or ( n60018 , n60016 , n60017 );
buf ( n60019 , n58846 );
buf ( n60020 , n56673 );
or ( n60021 , n60019 , n60020 );
nand ( n60022 , n60018 , n60021 );
buf ( n60023 , n60022 );
buf ( n60024 , n60023 );
and ( n60025 , n60007 , n60024 );
and ( n60026 , n59989 , n60006 );
or ( n60027 , n60025 , n60026 );
buf ( n60028 , n60027 );
buf ( n60029 , n58854 );
not ( n60030 , n60029 );
buf ( n60031 , n58867 );
not ( n60032 , n60031 );
buf ( n60033 , n58923 );
not ( n60034 , n60033 );
and ( n60035 , n60032 , n60034 );
buf ( n60036 , n58867 );
buf ( n60037 , n58923 );
and ( n60038 , n60036 , n60037 );
nor ( n60039 , n60035 , n60038 );
buf ( n60040 , n60039 );
buf ( n60041 , n60040 );
not ( n60042 , n60041 );
or ( n60043 , n60030 , n60042 );
buf ( n60044 , n60040 );
buf ( n60045 , n58854 );
or ( n60046 , n60044 , n60045 );
nand ( n60047 , n60043 , n60046 );
buf ( n60048 , n60047 );
xor ( n60049 , n60028 , n60048 );
xor ( n60050 , n58967 , n58987 );
xor ( n60051 , n60050 , n59021 );
buf ( n60052 , n60051 );
and ( n60053 , n60049 , n60052 );
and ( n60054 , n60028 , n60048 );
or ( n60055 , n60053 , n60054 );
buf ( n60056 , n60055 );
xor ( n60057 , n59972 , n60056 );
not ( n60058 , n54431 );
not ( n60059 , n55075 );
or ( n60060 , n60058 , n60059 );
not ( n60061 , n55078 );
nand ( n60062 , n60060 , n60061 );
not ( n60063 , n55080 );
nand ( n60064 , n60063 , n54457 );
nor ( n60065 , n60062 , n60064 );
not ( n60066 , n60065 );
nand ( n60067 , n60062 , n60064 );
nand ( n60068 , n60066 , n60067 );
buf ( n60069 , n60068 );
not ( n60070 , n60069 );
buf ( n60071 , n60070 );
buf ( n60072 , n60071 );
buf ( n60073 , n56589 );
or ( n60074 , n60072 , n60073 );
buf ( n60075 , n59009 );
not ( n60076 , n60075 );
buf ( n60077 , n60076 );
buf ( n60078 , n60077 );
buf ( n60079 , n56598 );
or ( n60080 , n60078 , n60079 );
nand ( n60081 , n60074 , n60080 );
buf ( n60082 , n60081 );
buf ( n60083 , n15265 );
buf ( n60084 , n2251 );
buf ( n60085 , n60084 );
not ( n60086 , n60085 );
buf ( n60087 , n60086 );
buf ( n60088 , n60087 );
and ( n60089 , n60083 , n60088 );
not ( n60090 , n15265 );
buf ( n60091 , n60090 );
buf ( n60092 , n60084 );
and ( n60093 , n60091 , n60092 );
nor ( n60094 , n60089 , n60093 );
buf ( n60095 , n60094 );
not ( n60096 , n14273 );
and ( n60097 , n60096 , n60087 );
not ( n60098 , n60096 );
and ( n60099 , n60098 , n60084 );
or ( n60100 , n60097 , n60099 );
and ( n60101 , n60095 , n60100 );
nand ( n60102 , n60101 , n58880 );
buf ( n60103 , n60102 );
not ( n60104 , n60100 );
buf ( n60105 , n60104 );
buf ( n60106 , n58880 );
nand ( n60107 , n60105 , n60106 );
buf ( n60108 , n60107 );
buf ( n60109 , n60108 );
and ( n60110 , n60103 , n60109 );
buf ( n60111 , n60110 );
xor ( n60112 , n60082 , n60111 );
buf ( n60113 , n56582 );
buf ( n60114 , n58721 );
and ( n60115 , n60113 , n60114 );
buf ( n60116 , n56585 );
buf ( n60117 , n58718 );
and ( n60118 , n60116 , n60117 );
nor ( n60119 , n60115 , n60118 );
buf ( n60120 , n60119 );
buf ( n60121 , n60120 );
buf ( n60122 , n56799 );
or ( n60123 , n60121 , n60122 );
buf ( n60124 , n59997 );
buf ( n60125 , n58982 );
or ( n60126 , n60124 , n60125 );
nand ( n60127 , n60123 , n60126 );
buf ( n60128 , n60127 );
and ( n60129 , n60112 , n60128 );
and ( n60130 , n60082 , n60111 );
or ( n60131 , n60129 , n60130 );
buf ( n60132 , n60131 );
buf ( n60133 , n59005 );
buf ( n60134 , n59017 );
or ( n60135 , n60133 , n60134 );
buf ( n60136 , n59020 );
nand ( n60137 , n60135 , n60136 );
buf ( n60138 , n60137 );
buf ( n60139 , n60138 );
xor ( n60140 , n60132 , n60139 );
buf ( n60141 , n58835 );
buf ( n60142 , n56641 );
and ( n60143 , n60141 , n60142 );
buf ( n60144 , n58841 );
buf ( n60145 , n56631 );
and ( n60146 , n60144 , n60145 );
nor ( n60147 , n60143 , n60146 );
buf ( n60148 , n60147 );
buf ( n60149 , n60148 );
buf ( n60150 , n56626 );
or ( n60151 , n60149 , n60150 );
buf ( n60152 , n59980 );
buf ( n60153 , n56639 );
or ( n60154 , n60152 , n60153 );
nand ( n60155 , n60151 , n60154 );
buf ( n60156 , n60155 );
buf ( n60157 , n60156 );
buf ( n60158 , n55113 );
buf ( n60159 , n58897 );
and ( n60160 , n60158 , n60159 );
buf ( n60161 , n56655 );
buf ( n60162 , n58894 );
and ( n60163 , n60161 , n60162 );
nor ( n60164 , n60160 , n60163 );
buf ( n60165 , n60164 );
buf ( n60166 , n60165 );
buf ( n60167 , n58913 );
or ( n60168 , n60166 , n60167 );
buf ( n60169 , n58996 );
buf ( n60170 , n58890 );
or ( n60171 , n60169 , n60170 );
nand ( n60172 , n60168 , n60171 );
buf ( n60173 , n60172 );
buf ( n60174 , n60173 );
xor ( n60175 , n60157 , n60174 );
buf ( n60176 , n58857 );
buf ( n60177 , n56652 );
and ( n60178 , n60176 , n60177 );
buf ( n60179 , n58858 );
buf ( n60180 , n55201 );
and ( n60181 , n60179 , n60180 );
nor ( n60182 , n60178 , n60181 );
buf ( n60183 , n60182 );
buf ( n60184 , n60183 );
buf ( n60185 , n56664 );
or ( n60186 , n60184 , n60185 );
buf ( n60187 , n60015 );
buf ( n60188 , n56673 );
or ( n60189 , n60187 , n60188 );
nand ( n60190 , n60186 , n60189 );
buf ( n60191 , n60190 );
buf ( n60192 , n60191 );
and ( n60193 , n60175 , n60192 );
and ( n60194 , n60157 , n60174 );
or ( n60195 , n60193 , n60194 );
buf ( n60196 , n60195 );
buf ( n60197 , n60196 );
and ( n60198 , n60140 , n60197 );
and ( n60199 , n60132 , n60139 );
or ( n60200 , n60198 , n60199 );
buf ( n60201 , n60200 );
xor ( n60202 , n60028 , n60048 );
xor ( n60203 , n60202 , n60052 );
and ( n60204 , n60201 , n60203 );
buf ( n60205 , n59009 );
buf ( n60206 , n56652 );
and ( n60207 , n60205 , n60206 );
buf ( n60208 , n60077 );
buf ( n60209 , n55201 );
and ( n60210 , n60208 , n60209 );
nor ( n60211 , n60207 , n60210 );
buf ( n60212 , n60211 );
buf ( n60213 , n60212 );
not ( n60214 , n60213 );
buf ( n60215 , n60214 );
buf ( n60216 , n60215 );
buf ( n60217 , n55180 );
and ( n60218 , n60216 , n60217 );
buf ( n60219 , n60183 );
not ( n60220 , n60219 );
buf ( n60221 , n60220 );
buf ( n60222 , n60221 );
buf ( n60223 , n56670 );
and ( n60224 , n60222 , n60223 );
nor ( n60225 , n60218 , n60224 );
buf ( n60226 , n60225 );
buf ( n60227 , n60226 );
nand ( n60228 , n60061 , n54431 );
xnor ( n60229 , n60228 , n55075 );
buf ( n60230 , n60229 );
buf ( n60231 , n55132 );
and ( n60232 , n60230 , n60231 );
buf ( n60233 , n60068 );
buf ( n60234 , n55156 );
and ( n60235 , n60233 , n60234 );
nor ( n60236 , n60232 , n60235 );
buf ( n60237 , n60236 );
buf ( n60238 , n60237 );
nand ( n60239 , n60227 , n60238 );
buf ( n60240 , n60239 );
xor ( n60241 , n60082 , n60111 );
xor ( n60242 , n60241 , n60128 );
and ( n60243 , n60240 , n60242 );
buf ( n60244 , n58699 );
buf ( n60245 , n58897 );
and ( n60246 , n60244 , n60245 );
buf ( n60247 , n56594 );
buf ( n60248 , n58894 );
and ( n60249 , n60247 , n60248 );
nor ( n60250 , n60246 , n60249 );
buf ( n60251 , n60250 );
buf ( n60252 , n60251 );
buf ( n60253 , n58913 );
or ( n60254 , n60252 , n60253 );
buf ( n60255 , n60165 );
buf ( n60256 , n58890 );
or ( n60257 , n60255 , n60256 );
nand ( n60258 , n60254 , n60257 );
buf ( n60259 , n60258 );
buf ( n60260 , n55152 );
not ( n60261 , n60090 );
buf ( n60262 , n60261 );
and ( n60263 , n60260 , n60262 );
buf ( n60264 , n55205 );
buf ( n60265 , n60090 );
and ( n60266 , n60264 , n60265 );
nor ( n60267 , n60263 , n60266 );
buf ( n60268 , n60267 );
buf ( n60269 , n60268 );
not ( n60270 , n60101 );
buf ( n60271 , n60270 );
or ( n60272 , n60269 , n60271 );
buf ( n60273 , n60108 );
nand ( n60274 , n60272 , n60273 );
buf ( n60275 , n60274 );
xor ( n60276 , n60259 , n60275 );
buf ( n60277 , n56720 );
buf ( n60278 , n58721 );
and ( n60279 , n60277 , n60278 );
buf ( n60280 , n58792 );
buf ( n60281 , n58718 );
and ( n60282 , n60280 , n60281 );
nor ( n60283 , n60279 , n60282 );
buf ( n60284 , n60283 );
buf ( n60285 , n60284 );
buf ( n60286 , n56799 );
or ( n60287 , n60285 , n60286 );
buf ( n60288 , n60120 );
buf ( n60289 , n58982 );
or ( n60290 , n60288 , n60289 );
nand ( n60291 , n60287 , n60290 );
buf ( n60292 , n60291 );
and ( n60293 , n60276 , n60292 );
and ( n60294 , n60259 , n60275 );
or ( n60295 , n60293 , n60294 );
xor ( n60296 , n60082 , n60111 );
xor ( n60297 , n60296 , n60128 );
and ( n60298 , n60295 , n60297 );
and ( n60299 , n60240 , n60295 );
or ( n60300 , n60243 , n60298 , n60299 );
xor ( n60301 , n59989 , n60006 );
xor ( n60302 , n60301 , n60024 );
buf ( n60303 , n60302 );
xor ( n60304 , n60300 , n60303 );
xor ( n60305 , n60132 , n60139 );
xor ( n60306 , n60305 , n60197 );
buf ( n60307 , n60306 );
and ( n60308 , n60304 , n60307 );
and ( n60309 , n60300 , n60303 );
or ( n60310 , n60308 , n60309 );
xor ( n60311 , n60028 , n60048 );
xor ( n60312 , n60311 , n60052 );
and ( n60313 , n60310 , n60312 );
and ( n60314 , n60201 , n60310 );
or ( n60315 , n60204 , n60313 , n60314 );
buf ( n60316 , n60315 );
and ( n60317 , n60057 , n60316 );
and ( n60318 , n59972 , n60056 );
or ( n60319 , n60317 , n60318 );
buf ( n60320 , n60319 );
buf ( n60321 , n60320 );
xor ( n60322 , n59953 , n60321 );
buf ( n60323 , n25180 );
not ( n60324 , n60323 );
buf ( n60325 , n28344 );
buf ( n60326 , n60325 );
buf ( n60327 , n60326 );
buf ( n60328 , n60327 );
not ( n60329 , n60328 );
buf ( n60330 , n60329 );
buf ( n60331 , n60330 );
not ( n60332 , n60331 );
and ( n60333 , n60324 , n60332 );
buf ( n60334 , n54068 );
buf ( n60335 , n41733 );
and ( n60336 , n60334 , n60335 );
nor ( n60337 , n60333 , n60336 );
buf ( n60338 , n60337 );
not ( n60339 , n60338 );
buf ( n60340 , n60339 );
not ( n60341 , n60340 );
buf ( n60342 , n43935 );
not ( n60343 , n60342 );
or ( n60344 , n60341 , n60343 );
buf ( n60345 , n59896 );
buf ( n60346 , n43905 );
nand ( n60347 , n60345 , n60346 );
buf ( n60348 , n60347 );
buf ( n60349 , n60348 );
nand ( n60350 , n60344 , n60349 );
buf ( n60351 , n60350 );
buf ( n60352 , n60351 );
and ( n60353 , n60322 , n60352 );
and ( n60354 , n59953 , n60321 );
or ( n60355 , n60353 , n60354 );
buf ( n60356 , n60355 );
not ( n60357 , n60356 );
nand ( n60358 , n59938 , n60357 );
not ( n60359 , n60358 );
buf ( n60360 , n42712 );
not ( n60361 , n60360 );
buf ( n60362 , n25226 );
not ( n60363 , n60362 );
buf ( n60364 , n42195 );
not ( n60365 , n60364 );
or ( n60366 , n60363 , n60365 );
buf ( n60367 , n29360 );
buf ( n60368 , n25227 );
nand ( n60369 , n60367 , n60368 );
buf ( n60370 , n60369 );
buf ( n60371 , n60370 );
nand ( n60372 , n60366 , n60371 );
buf ( n60373 , n60372 );
buf ( n60374 , n60373 );
not ( n60375 , n60374 );
or ( n60376 , n60361 , n60375 );
buf ( n60377 , n25228 );
not ( n60378 , n60377 );
buf ( n60379 , n51250 );
not ( n60380 , n60379 );
or ( n60381 , n60378 , n60380 );
buf ( n60382 , n41822 );
buf ( n60383 , n25227 );
nand ( n60384 , n60382 , n60383 );
buf ( n60385 , n60384 );
buf ( n60386 , n60385 );
nand ( n60387 , n60381 , n60386 );
buf ( n60388 , n60387 );
buf ( n60389 , n60388 );
buf ( n60390 , n42668 );
nand ( n60391 , n60389 , n60390 );
buf ( n60392 , n60391 );
buf ( n60393 , n60392 );
nand ( n60394 , n60376 , n60393 );
buf ( n60395 , n60394 );
not ( n60396 , n60395 );
or ( n60397 , n60359 , n60396 );
nand ( n60398 , n59937 , n60356 );
nand ( n60399 , n60397 , n60398 );
nand ( n60400 , n59869 , n60399 );
buf ( n60401 , n60400 );
buf ( n60402 , n59860 );
not ( n60403 , n60402 );
buf ( n60404 , n59864 );
nand ( n60405 , n60403 , n60404 );
buf ( n60406 , n60405 );
buf ( n60407 , n60406 );
nand ( n60408 , n60401 , n60407 );
buf ( n60409 , n60408 );
buf ( n60410 , n60409 );
xor ( n60411 , n59533 , n59540 );
xnor ( n60412 , n60411 , n59513 );
buf ( n60413 , n60412 );
xor ( n60414 , n60410 , n60413 );
buf ( n60415 , n44670 );
and ( n60416 , n52780 , n49425 );
not ( n60417 , n52780 );
and ( n60418 , n60417 , n43095 );
or ( n60419 , n60416 , n60418 );
buf ( n60420 , n60419 );
not ( n60421 , n60420 );
buf ( n60422 , n60421 );
buf ( n60423 , n60422 );
or ( n60424 , n60415 , n60423 );
buf ( n60425 , n36909 );
buf ( n60426 , n53946 );
buf ( n60427 , n44689 );
and ( n60428 , n60426 , n60427 );
not ( n60429 , n60426 );
buf ( n60430 , n36929 );
and ( n60431 , n60429 , n60430 );
nor ( n60432 , n60428 , n60431 );
buf ( n60433 , n60432 );
buf ( n60434 , n60433 );
or ( n60435 , n60425 , n60434 );
nand ( n60436 , n60424 , n60435 );
buf ( n60437 , n60436 );
buf ( n60438 , n60437 );
and ( n60439 , n60414 , n60438 );
and ( n60440 , n60410 , n60413 );
or ( n60441 , n60439 , n60440 );
buf ( n60442 , n60441 );
and ( n60443 , n59838 , n60442 );
and ( n60444 , n59828 , n59837 );
or ( n60445 , n60443 , n60444 );
buf ( n60446 , n60445 );
nand ( n60447 , n59792 , n60446 );
buf ( n60448 , n60447 );
buf ( n60449 , n60448 );
buf ( n60450 , n59789 );
not ( n60451 , n60450 );
buf ( n60452 , n60451 );
buf ( n60453 , n60452 );
buf ( n60454 , n59774 );
nand ( n60455 , n60453 , n60454 );
buf ( n60456 , n60455 );
buf ( n60457 , n60456 );
nand ( n60458 , n60449 , n60457 );
buf ( n60459 , n60458 );
xor ( n60460 , n59761 , n60459 );
buf ( n60461 , n59725 );
buf ( n60462 , n59737 );
xor ( n60463 , n60461 , n60462 );
buf ( n60464 , n59742 );
xor ( n60465 , n60463 , n60464 );
buf ( n60466 , n60465 );
and ( n60467 , n60460 , n60466 );
and ( n60468 , n59761 , n60459 );
or ( n60469 , n60467 , n60468 );
buf ( n60470 , n60469 );
nand ( n60471 , n59758 , n60470 );
buf ( n60472 , n60471 );
buf ( n60473 , n60472 );
buf ( n60474 , n59756 );
buf ( n60475 , n59627 );
nand ( n60476 , n60474 , n60475 );
buf ( n60477 , n60476 );
buf ( n60478 , n60477 );
nand ( n60479 , n60473 , n60478 );
buf ( n60480 , n60479 );
buf ( n60481 , n60480 );
and ( n60482 , n59624 , n60481 );
and ( n60483 , n59157 , n59623 );
or ( n60484 , n60482 , n60483 );
buf ( n60485 , n60484 );
xor ( n60486 , n59147 , n60485 );
xor ( n60487 , n59167 , n59171 );
and ( n60488 , n60487 , n59620 );
and ( n60489 , n59167 , n59171 );
or ( n60490 , n60488 , n60489 );
buf ( n60491 , n60490 );
xor ( n60492 , n57956 , n57960 );
xor ( n60493 , n60492 , n58391 );
buf ( n60494 , n60493 );
xor ( n60495 , n60491 , n60494 );
not ( n60496 , n59751 );
not ( n60497 , n59630 );
and ( n60498 , n60496 , n60497 );
nand ( n60499 , n59630 , n59751 );
buf ( n60500 , n59744 );
and ( n60501 , n60499 , n60500 );
nor ( n60502 , n60498 , n60501 );
not ( n60503 , n60502 );
not ( n60504 , n60503 );
and ( n60505 , n57971 , n58388 );
not ( n60506 , n57971 );
not ( n60507 , n58388 );
and ( n60508 , n60506 , n60507 );
nor ( n60509 , n60505 , n60508 );
xnor ( n60510 , n60509 , n57967 );
not ( n60511 , n60510 );
not ( n60512 , n60511 );
or ( n60513 , n60504 , n60512 );
not ( n60514 , n60510 );
not ( n60515 , n60502 );
or ( n60516 , n60514 , n60515 );
not ( n60517 , n58445 );
or ( n60518 , C0 , n60517 );
buf ( n60519 , C1 );
nand ( n60520 , n60518 , n60519 );
not ( n60521 , n58434 );
and ( n60522 , n60520 , n60521 );
not ( n60523 , n60520 );
not ( n60524 , n58438 );
and ( n60525 , n60523 , n60524 );
nor ( n60526 , n60522 , n60525 );
not ( n60527 , n60526 );
not ( n60528 , n60527 );
buf ( n60529 , n57174 );
not ( n60530 , n60529 );
buf ( n60531 , n50876 );
not ( n60532 , n60531 );
or ( n60533 , n60530 , n60532 );
buf ( n60534 , n42360 );
buf ( n60535 , n51496 );
nand ( n60536 , n60534 , n60535 );
buf ( n60537 , n60536 );
buf ( n60538 , n60537 );
nand ( n60539 , n60533 , n60538 );
buf ( n60540 , n60539 );
buf ( n60541 , n60540 );
buf ( n60542 , n51488 );
and ( n60543 , n60541 , n60542 );
buf ( n60544 , n59577 );
buf ( n60545 , n52456 );
buf ( n60546 , n60545 );
and ( n60547 , n60544 , n60546 );
nor ( n60548 , n60543 , n60547 );
buf ( n60549 , n60548 );
buf ( n60550 , n60549 );
not ( n60551 , n60550 );
or ( n60552 , n60551 , C0 );
buf ( n60553 , n59208 );
buf ( n60554 , n44496 );
and ( n60555 , n60553 , n60554 );
buf ( n60556 , n44533 );
not ( n60557 , n60556 );
buf ( n60558 , n44157 );
not ( n60559 , n60558 );
or ( n60560 , n60557 , n60559 );
buf ( n60561 , n39489 );
buf ( n60562 , n44530 );
nand ( n60563 , n60561 , n60562 );
buf ( n60564 , n60563 );
buf ( n60565 , n60564 );
nand ( n60566 , n60560 , n60565 );
buf ( n60567 , n60566 );
buf ( n60568 , n60567 );
not ( n60569 , n60568 );
buf ( n60570 , n44518 );
nor ( n60571 , n60569 , n60570 );
buf ( n60572 , n60571 );
buf ( n60573 , n60572 );
nor ( n60574 , n60555 , n60573 );
buf ( n60575 , n60574 );
not ( n60576 , n60575 );
buf ( n60577 , n36520 );
not ( n60578 , n60577 );
buf ( n60579 , n56325 );
buf ( n60580 , n36527 );
and ( n60581 , n60579 , n60580 );
not ( n60582 , n60579 );
buf ( n60583 , n38468 );
buf ( n60584 , n60583 );
and ( n60585 , n60582 , n60584 );
nor ( n60586 , n60581 , n60585 );
buf ( n60587 , n60586 );
buf ( n60588 , n60587 );
not ( n60589 , n60588 );
and ( n60590 , n60578 , n60589 );
buf ( n60591 , n58367 );
not ( n60592 , n60591 );
buf ( n60593 , n39813 );
nor ( n60594 , n60592 , n60593 );
buf ( n60595 , n60594 );
buf ( n60596 , n60595 );
nor ( n60597 , n60590 , n60596 );
buf ( n60598 , n60597 );
not ( n60599 , n60598 );
or ( n60600 , n60576 , n60599 );
xor ( n60601 , n58558 , n58577 );
xnor ( n60602 , n60601 , n58545 );
nand ( n60603 , n60600 , n60602 );
buf ( n60604 , n60603 );
buf ( n60605 , n60575 );
not ( n60606 , n60605 );
buf ( n60607 , n60598 );
not ( n60608 , n60607 );
buf ( n60609 , n60608 );
buf ( n60610 , n60609 );
nand ( n60611 , n60606 , n60610 );
buf ( n60612 , n60611 );
buf ( n60613 , n60612 );
nand ( n60614 , n60604 , n60613 );
buf ( n60615 , n60614 );
buf ( n60616 , n60615 );
nand ( n60617 , n60552 , n60616 );
buf ( n60618 , n60617 );
buf ( n60619 , n60618 );
buf ( n60620 , n60549 );
not ( n60621 , n60620 );
buf ( n60622 , n60621 );
buf ( n60623 , C1 );
buf ( n60624 , n60623 );
nand ( n60625 , n60619 , n60624 );
buf ( n60626 , n60625 );
not ( n60627 , n60626 );
or ( n60628 , n60528 , n60627 );
buf ( n60629 , n58312 );
not ( n60630 , n60629 );
buf ( n60631 , n46915 );
not ( n60632 , n60631 );
and ( n60633 , n60630 , n60632 );
buf ( n60634 , n59806 );
buf ( n60635 , n47331 );
and ( n60636 , n60634 , n60635 );
nor ( n60637 , n60633 , n60636 );
buf ( n60638 , n60637 );
buf ( n60639 , n60638 );
buf ( n60640 , n60639 );
not ( n60641 , n60640 );
and ( n60642 , n58342 , n58345 );
not ( n60643 , n58342 );
and ( n60644 , n60643 , n58346 );
nor ( n60645 , n60642 , n60644 );
and ( n60646 , n60645 , n58379 );
not ( n60647 , n60645 );
buf ( n60648 , n58379 );
not ( n60649 , n60648 );
buf ( n60650 , n60649 );
and ( n60651 , n60647 , n60650 );
nor ( n60652 , n60646 , n60651 );
buf ( n60653 , n60652 );
not ( n60654 , n60653 );
or ( n60655 , n60641 , n60654 );
buf ( n60656 , n36982 );
buf ( n60657 , n60433 );
or ( n60658 , n60656 , n60657 );
buf ( n60659 , n58334 );
not ( n60660 , n60659 );
buf ( n60661 , n60660 );
buf ( n60662 , n60661 );
buf ( n60663 , n36909 );
or ( n60664 , n60662 , n60663 );
nand ( n60665 , n60658 , n60664 );
buf ( n60666 , n60665 );
buf ( n60667 , n60666 );
not ( n60668 , n60667 );
xor ( n60669 , n58621 , n59057 );
not ( n60670 , n60669 );
not ( n60671 , n60670 );
not ( n60672 , n58601 );
or ( n60673 , n60671 , n60672 );
not ( n60674 , n58601 );
nand ( n60675 , n60674 , n60669 );
nand ( n60676 , n60673 , n60675 );
buf ( n60677 , n60676 );
not ( n60678 , n60677 );
or ( n60679 , n60668 , n60678 );
or ( n60680 , n60666 , n60676 );
buf ( n60681 , n59053 );
not ( n60682 , n60681 );
buf ( n60683 , n58690 );
not ( n60684 , n60683 );
and ( n60685 , n60682 , n60684 );
buf ( n60686 , n59053 );
buf ( n60687 , n58690 );
and ( n60688 , n60686 , n60687 );
nor ( n60689 , n60685 , n60688 );
buf ( n60690 , n60689 );
buf ( n60691 , n60690 );
not ( n60692 , n60691 );
buf ( n60693 , n58685 );
not ( n60694 , n60693 );
or ( n60695 , n60692 , n60694 );
buf ( n60696 , n58685 );
buf ( n60697 , n60690 );
or ( n60698 , n60696 , n60697 );
nand ( n60699 , n60695 , n60698 );
buf ( n60700 , n60699 );
buf ( n60701 , n60700 );
not ( n60702 , n47014 );
buf ( n60703 , n43063 );
not ( n60704 , n60703 );
buf ( n60705 , n42471 );
not ( n60706 , n60705 );
or ( n60707 , n60704 , n60706 );
buf ( n60708 , n42468 );
buf ( n60709 , n43064 );
nand ( n60710 , n60708 , n60709 );
buf ( n60711 , n60710 );
buf ( n60712 , n60711 );
nand ( n60713 , n60707 , n60712 );
buf ( n60714 , n60713 );
not ( n60715 , n60714 );
or ( n60716 , n60702 , n60715 );
nand ( n60717 , n52595 , n59267 );
nand ( n60718 , n60716 , n60717 );
buf ( n60719 , n60718 );
xor ( n60720 , n60701 , n60719 );
not ( n60721 , n42336 );
not ( n60722 , n59298 );
or ( n60723 , n60721 , n60722 );
not ( n60724 , n42343 );
not ( n60725 , n41879 );
or ( n60726 , n60724 , n60725 );
nand ( n60727 , n41876 , n46855 );
nand ( n60728 , n60726 , n60727 );
nand ( n60729 , n60728 , n42378 );
nand ( n60730 , n60723 , n60729 );
buf ( n60731 , n60730 );
and ( n60732 , n60720 , n60731 );
and ( n60733 , n60701 , n60719 );
or ( n60734 , n60732 , n60733 );
buf ( n60735 , n60734 );
buf ( n60736 , n60735 );
buf ( n60737 , n58597 );
buf ( n60738 , n37443 );
or ( n60739 , n60737 , n60738 );
buf ( n60740 , n46390 );
buf ( n60741 , n51901 );
and ( n60742 , n60740 , n60741 );
not ( n60743 , n60740 );
buf ( n60744 , n37472 );
and ( n60745 , n60743 , n60744 );
nor ( n60746 , n60742 , n60745 );
buf ( n60747 , n60746 );
nand ( n60748 , n60747 , n37443 , n57522 );
buf ( n60749 , n60748 );
nand ( n60750 , n60739 , n60749 );
buf ( n60751 , n60750 );
buf ( n60752 , n60751 );
xor ( n60753 , n60736 , n60752 );
buf ( n60754 , n48323 );
not ( n60755 , n60754 );
buf ( n60756 , n37880 );
not ( n60757 , n60756 );
or ( n60758 , n60755 , n60757 );
nand ( n60759 , n37881 , n48320 );
buf ( n60760 , n60759 );
nand ( n60761 , n60758 , n60760 );
buf ( n60762 , n60761 );
buf ( n60763 , n60762 );
not ( n60764 , n60763 );
buf ( n60765 , n41862 );
not ( n60766 , n60765 );
or ( n60767 , n60764 , n60766 );
buf ( n60768 , n41905 );
buf ( n60769 , n58543 );
nand ( n60770 , n60768 , n60769 );
buf ( n60771 , n60770 );
buf ( n60772 , n60771 );
nand ( n60773 , n60767 , n60772 );
buf ( n60774 , n60773 );
buf ( n60775 , n60774 );
and ( n60776 , n60753 , n60775 );
and ( n60777 , n60736 , n60752 );
or ( n60778 , n60776 , n60777 );
buf ( n60779 , n60778 );
nand ( n60780 , n60680 , n60779 );
buf ( n60781 , n60780 );
nand ( n60782 , n60679 , n60781 );
buf ( n60783 , n60782 );
buf ( n60784 , n60783 );
nand ( n60785 , n60655 , n60784 );
buf ( n60786 , n60785 );
not ( n60787 , n60786 );
not ( n60788 , n60652 );
buf ( n60789 , n60788 );
not ( n60790 , n60638 );
buf ( n60791 , n60790 );
nand ( n60792 , n60789 , n60791 );
buf ( n60793 , n60792 );
not ( n60794 , n60793 );
or ( n60795 , n60787 , n60794 );
not ( n60796 , n60626 );
nand ( n60797 , n60796 , n60526 );
nand ( n60798 , n60795 , n60797 );
nand ( n60799 , n60628 , n60798 );
buf ( n60800 , n58494 );
not ( n60801 , n60800 );
buf ( n60802 , n58485 );
not ( n60803 , n60802 );
or ( n60804 , n60801 , n60803 );
buf ( n60805 , n58482 );
buf ( n60806 , n58489 );
nand ( n60807 , n60805 , n60806 );
buf ( n60808 , n60807 );
buf ( n60809 , n60808 );
nand ( n60810 , n60804 , n60809 );
buf ( n60811 , n60810 );
buf ( n60812 , n60811 );
buf ( n60813 , n59074 );
and ( n60814 , n60812 , n60813 );
not ( n60815 , n60812 );
buf ( n60816 , n59074 );
not ( n60817 , n60816 );
buf ( n60818 , n60817 );
buf ( n60819 , n60818 );
and ( n60820 , n60815 , n60819 );
nor ( n60821 , n60814 , n60820 );
buf ( n60822 , n60821 );
xor ( n60823 , n60799 , n60822 );
xor ( n60824 , n59196 , n59554 );
xnor ( n60825 , n60824 , n59440 );
buf ( n60826 , n60825 );
not ( n60827 , n60826 );
buf ( n60828 , n60827 );
not ( n60829 , n60828 );
xor ( n60830 , n58522 , n59065 );
xor ( n60831 , n60830 , n59070 );
buf ( n60832 , n60831 );
not ( n60833 , n60832 );
or ( n60834 , n60829 , n60833 );
buf ( n60835 , n60832 );
not ( n60836 , n60835 );
buf ( n60837 , n60836 );
not ( n60838 , n60837 );
not ( n60839 , n60825 );
or ( n60840 , n60838 , n60839 );
buf ( n60841 , C1 );
buf ( n60842 , n48868 );
not ( n60843 , n60842 );
buf ( n60844 , n59705 );
not ( n60845 , n60844 );
or ( n60846 , n60843 , n60845 );
buf ( n60847 , n48855 );
and ( n60848 , n48808 , n43031 );
not ( n60849 , n48808 );
and ( n60850 , n60849 , n38244 );
or ( n60851 , n60848 , n60850 );
buf ( n60852 , n60851 );
nand ( n60853 , n60847 , n60852 );
buf ( n60854 , n60853 );
buf ( n60855 , n60854 );
nand ( n60856 , n60846 , n60855 );
buf ( n60857 , n60856 );
buf ( n60858 , n60857 );
xor ( n60859 , n59259 , n59311 );
xor ( n60860 , n60859 , n59433 );
buf ( n60861 , n60860 );
xor ( n60862 , n60858 , n60861 );
xor ( n60863 , n59279 , n59303 );
xor ( n60864 , n60863 , n59309 );
buf ( n60865 , n60864 );
buf ( n60866 , n43250 );
not ( n60867 , n60866 );
buf ( n60868 , n55841 );
not ( n60869 , n60868 );
buf ( n60870 , n36500 );
not ( n60871 , n60870 );
or ( n60872 , n60869 , n60871 );
buf ( n60873 , n43503 );
buf ( n60874 , n55840 );
nand ( n60875 , n60873 , n60874 );
buf ( n60876 , n60875 );
buf ( n60877 , n60876 );
nand ( n60878 , n60872 , n60877 );
buf ( n60879 , n60878 );
buf ( n60880 , n60879 );
not ( n60881 , n60880 );
or ( n60882 , n60867 , n60881 );
buf ( n60883 , n32969 );
buf ( n60884 , n59664 );
nand ( n60885 , n60883 , n60884 );
buf ( n60886 , n60885 );
buf ( n60887 , n60886 );
nand ( n60888 , n60882 , n60887 );
buf ( n60889 , n60888 );
buf ( n60890 , n60889 );
xor ( n60891 , n60865 , n60890 );
nand ( n60892 , n59330 , n59341 , n59427 );
not ( n60893 , n59427 );
nand ( n60894 , n59341 , n59331 , n60893 );
nand ( n60895 , n59342 , n59331 , n59427 );
nand ( n60896 , n59342 , n59330 , n60893 );
nand ( n60897 , n60892 , n60894 , n60895 , n60896 );
buf ( n60898 , n60897 );
and ( n60899 , n60891 , n60898 );
and ( n60900 , n60865 , n60890 );
or ( n60901 , n60899 , n60900 );
buf ( n60902 , n60901 );
buf ( n60903 , n60902 );
and ( n60904 , n60862 , n60903 );
and ( n60905 , n60858 , n60861 );
or ( n60906 , n60904 , n60905 );
buf ( n60907 , n60906 );
buf ( n60908 , n60907 );
not ( n60909 , n60908 );
buf ( n60910 , n60909 );
not ( n60911 , n60910 );
or ( n60912 , C0 , n60911 );
buf ( n60913 , n59643 );
not ( n60914 , n60913 );
buf ( n60915 , n41577 );
not ( n60916 , n60915 );
and ( n60917 , n60914 , n60916 );
buf ( n60918 , n41608 );
not ( n60919 , n60918 );
buf ( n60920 , n43311 );
not ( n60921 , n60920 );
or ( n60922 , n60919 , n60921 );
buf ( n60923 , n44992 );
buf ( n60924 , n41611 );
nand ( n60925 , n60923 , n60924 );
buf ( n60926 , n60925 );
buf ( n60927 , n60926 );
nand ( n60928 , n60922 , n60927 );
buf ( n60929 , n60928 );
buf ( n60930 , n60929 );
buf ( n60931 , n44267 );
and ( n60932 , n60930 , n60931 );
nor ( n60933 , n60917 , n60932 );
buf ( n60934 , n60933 );
nand ( n60935 , n44141 , n12481 );
or ( n60936 , n60934 , n60935 );
buf ( n60937 , n60935 );
not ( n60938 , n60937 );
buf ( n60939 , n60934 );
not ( n60940 , n60939 );
or ( n60941 , n60938 , n60940 );
xor ( n60942 , n59884 , n59909 );
and ( n60943 , n60942 , n59935 );
and ( n60944 , n59884 , n59909 );
or ( n60945 , n60943 , n60944 );
buf ( n60946 , n60945 );
buf ( n60947 , n60946 );
buf ( n60948 , n41993 );
not ( n60949 , n60948 );
buf ( n60950 , n52551 );
not ( n60951 , n60950 );
or ( n60952 , n60949 , n60951 );
buf ( n60953 , n24092 );
buf ( n60954 , n43966 );
nand ( n60955 , n60953 , n60954 );
buf ( n60956 , n60955 );
buf ( n60957 , n60956 );
nand ( n60958 , n60952 , n60957 );
buf ( n60959 , n60958 );
buf ( n60960 , n60959 );
not ( n60961 , n60960 );
buf ( n60962 , n50608 );
not ( n60963 , n60962 );
or ( n60964 , n60961 , n60963 );
buf ( n60965 , n59381 );
buf ( n60966 , n46633 );
nand ( n60967 , n60965 , n60966 );
buf ( n60968 , n60967 );
buf ( n60969 , n60968 );
nand ( n60970 , n60964 , n60969 );
buf ( n60971 , n60970 );
not ( n60972 , n60971 );
not ( n60973 , n50128 );
buf ( n60974 , n42504 );
not ( n60975 , n60974 );
buf ( n60976 , n51804 );
not ( n60977 , n60976 );
or ( n60978 , n60975 , n60977 );
buf ( n60979 , n25159 );
buf ( n60980 , n41721 );
nand ( n60981 , n60979 , n60980 );
buf ( n60982 , n60981 );
buf ( n60983 , n60982 );
nand ( n60984 , n60978 , n60983 );
buf ( n60985 , n60984 );
not ( n60986 , n60985 );
or ( n60987 , n60973 , n60986 );
nand ( n60988 , n56567 , n59356 );
nand ( n60989 , n60987 , n60988 );
not ( n60990 , n60989 );
nand ( n60991 , n60972 , n60990 );
not ( n60992 , n60991 );
not ( n60993 , n42378 );
buf ( n60994 , n42343 );
not ( n60995 , n60994 );
buf ( n60996 , n47836 );
not ( n60997 , n60996 );
or ( n60998 , n60995 , n60997 );
buf ( n60999 , n42149 );
buf ( n61000 , n46855 );
nand ( n61001 , n60999 , n61000 );
buf ( n61002 , n61001 );
buf ( n61003 , n61002 );
nand ( n61004 , n60998 , n61003 );
buf ( n61005 , n61004 );
not ( n61006 , n61005 );
or ( n61007 , n60993 , n61006 );
buf ( n61008 , n60728 );
buf ( n61009 , n42336 );
nand ( n61010 , n61008 , n61009 );
buf ( n61011 , n61010 );
nand ( n61012 , n61007 , n61011 );
not ( n61013 , n61012 );
or ( n61014 , n60992 , n61013 );
nand ( n61015 , n60989 , n60971 );
nand ( n61016 , n61014 , n61015 );
buf ( n61017 , n61016 );
xor ( n61018 , n60947 , n61017 );
and ( n61019 , n42847 , n44054 );
not ( n61020 , n42847 );
and ( n61021 , n61020 , n47068 );
or ( n61022 , n61019 , n61021 );
not ( n61023 , n61022 );
not ( n61024 , n44042 );
or ( n61025 , n61023 , n61024 );
not ( n61026 , n38379 );
nand ( n61027 , n61026 , n59337 );
nand ( n61028 , n61025 , n61027 );
buf ( n61029 , n61028 );
and ( n61030 , n61018 , n61029 );
and ( n61031 , n60947 , n61017 );
or ( n61032 , n61030 , n61031 );
buf ( n61033 , n61032 );
buf ( n61034 , n61033 );
nand ( n61035 , n60941 , n61034 );
buf ( n61036 , n61035 );
nand ( n61037 , n60936 , n61036 );
buf ( n61038 , n61037 );
buf ( n61039 , n46246 );
not ( n61040 , n61039 );
buf ( n61041 , n59223 );
not ( n61042 , n61041 );
or ( n61043 , n61040 , n61042 );
buf ( n61044 , n45753 );
not ( n61045 , n61044 );
buf ( n61046 , n44316 );
not ( n61047 , n61046 );
or ( n61048 , n61045 , n61047 );
buf ( n61049 , n39522 );
buf ( n61050 , n45750 );
nand ( n61051 , n61049 , n61050 );
buf ( n61052 , n61051 );
buf ( n61053 , n61052 );
nand ( n61054 , n61048 , n61053 );
buf ( n61055 , n61054 );
buf ( n61056 , n61055 );
buf ( n61057 , n46225 );
nand ( n61058 , n61056 , n61057 );
buf ( n61059 , n61058 );
buf ( n61060 , n61059 );
nand ( n61061 , n61043 , n61060 );
buf ( n61062 , n61061 );
buf ( n61063 , n61062 );
xor ( n61064 , n61038 , n61063 );
and ( n61065 , n51004 , n44635 );
not ( n61066 , n51004 );
and ( n61067 , n61066 , n49391 );
or ( n61068 , n61065 , n61067 );
buf ( n61069 , n61068 );
not ( n61070 , n61069 );
buf ( n61071 , n47101 );
not ( n61072 , n61071 );
or ( n61073 , n61070 , n61072 );
buf ( n61074 , n59482 );
buf ( n61075 , n47108 );
nand ( n61076 , n61074 , n61075 );
buf ( n61077 , n61076 );
buf ( n61078 , n61077 );
nand ( n61079 , n61073 , n61078 );
buf ( n61080 , n61079 );
buf ( n61081 , n61080 );
not ( n61082 , n61081 );
buf ( n61083 , n44708 );
not ( n61084 , n61083 );
not ( n61085 , n44533 );
not ( n61086 , n45394 );
or ( n61087 , n61085 , n61086 );
not ( n61088 , n42891 );
nand ( n61089 , n61088 , n44530 );
nand ( n61090 , n61087 , n61089 );
buf ( n61091 , n61090 );
not ( n61092 , n61091 );
or ( n61093 , n61084 , n61092 );
buf ( n61094 , n60567 );
buf ( n61095 , n44496 );
nand ( n61096 , n61094 , n61095 );
buf ( n61097 , n61096 );
buf ( n61098 , n61097 );
nand ( n61099 , n61093 , n61098 );
buf ( n61100 , n61099 );
buf ( n61101 , n61100 );
not ( n61102 , n61101 );
or ( n61103 , n61082 , n61102 );
buf ( n61104 , n61080 );
not ( n61105 , n61104 );
buf ( n61106 , n61105 );
buf ( n61107 , n61106 );
not ( n61108 , n61107 );
buf ( n61109 , n61100 );
not ( n61110 , n61109 );
buf ( n61111 , n61110 );
buf ( n61112 , n61111 );
not ( n61113 , n61112 );
or ( n61114 , n61108 , n61113 );
buf ( n61115 , n42668 );
not ( n61116 , n61115 );
buf ( n61117 , n59328 );
not ( n61118 , n61117 );
or ( n61119 , n61116 , n61118 );
buf ( n61120 , n60388 );
buf ( n61121 , n58249 );
nand ( n61122 , n61120 , n61121 );
buf ( n61123 , n61122 );
buf ( n61124 , n61123 );
nand ( n61125 , n61119 , n61124 );
buf ( n61126 , n61125 );
buf ( n61127 , n46117 );
not ( n61128 , n61127 );
buf ( n61129 , n41805 );
not ( n61130 , n61129 );
or ( n61131 , n61128 , n61130 );
buf ( n61132 , n41769 );
buf ( n61133 , n46126 );
nand ( n61134 , n61132 , n61133 );
buf ( n61135 , n61134 );
buf ( n61136 , n61135 );
nand ( n61137 , n61131 , n61136 );
buf ( n61138 , n61137 );
buf ( n61139 , n61138 );
not ( n61140 , n61139 );
buf ( n61141 , n37397 );
not ( n61142 , n61141 );
or ( n61143 , n61140 , n61142 );
buf ( n61144 , n59525 );
buf ( n61145 , n42135 );
nand ( n61146 , n61144 , n61145 );
buf ( n61147 , n61146 );
buf ( n61148 , n61147 );
nand ( n61149 , n61143 , n61148 );
buf ( n61150 , n61149 );
or ( n61151 , n61126 , n61150 );
buf ( n61152 , n42315 );
not ( n61153 , n61152 );
buf ( n61154 , n59511 );
not ( n61155 , n61154 );
or ( n61156 , n61153 , n61155 );
buf ( n61157 , n59242 );
not ( n61158 , n61157 );
buf ( n61159 , n41763 );
not ( n61160 , n61159 );
or ( n61161 , n61158 , n61160 );
buf ( n61162 , n41762 );
buf ( n61163 , n42263 );
nand ( n61164 , n61162 , n61163 );
buf ( n61165 , n61164 );
buf ( n61166 , n61165 );
nand ( n61167 , n61161 , n61166 );
buf ( n61168 , n61167 );
buf ( n61169 , n61168 );
buf ( n61170 , n42252 );
nand ( n61171 , n61169 , n61170 );
buf ( n61172 , n61171 );
buf ( n61173 , n61172 );
nand ( n61174 , n61156 , n61173 );
buf ( n61175 , n61174 );
nand ( n61176 , n61151 , n61175 );
buf ( n61177 , n61176 );
buf ( n61178 , n61150 );
buf ( n61179 , n61126 );
nand ( n61180 , n61178 , n61179 );
buf ( n61181 , n61180 );
buf ( n61182 , n61181 );
nand ( n61183 , n61177 , n61182 );
buf ( n61184 , n61183 );
buf ( n61185 , n61184 );
nand ( n61186 , n61114 , n61185 );
buf ( n61187 , n61186 );
buf ( n61188 , n61187 );
nand ( n61189 , n61103 , n61188 );
buf ( n61190 , n61189 );
buf ( n61191 , n61190 );
and ( n61192 , n61064 , n61191 );
and ( n61193 , n61038 , n61063 );
or ( n61194 , n61192 , n61193 );
buf ( n61195 , n61194 );
buf ( n61196 , n61195 );
nand ( n61197 , n60912 , n61196 );
buf ( n61198 , C1 );
nand ( n61199 , n61197 , n61198 );
nand ( n61200 , n60840 , n61199 );
nand ( n61201 , n60834 , n61200 );
and ( n61202 , n60823 , n61201 );
and ( n61203 , n60799 , n60822 );
or ( n61204 , n61202 , n61203 );
nand ( n61205 , n60516 , n61204 );
nand ( n61206 , n60513 , n61205 );
xor ( n61207 , n60495 , n61206 );
xor ( n61208 , n60486 , n61207 );
not ( n61209 , n61208 );
not ( n61210 , n60503 );
not ( n61211 , n60511 );
and ( n61212 , n61210 , n61211 );
and ( n61213 , n60503 , n60511 );
nor ( n61214 , n61212 , n61213 );
buf ( n61215 , n61204 );
not ( n61216 , n61215 );
buf ( n61217 , n61216 );
not ( n61218 , n61217 );
and ( n61219 , n61214 , n61218 );
not ( n61220 , n61214 );
and ( n61221 , n61220 , n61217 );
nor ( n61222 , n61219 , n61221 );
buf ( n61223 , n61222 );
buf ( n61224 , n60786 );
buf ( n61225 , n60793 );
nand ( n61226 , n61224 , n61225 );
buf ( n61227 , n61226 );
buf ( n61228 , n61227 );
not ( n61229 , n61228 );
buf ( n61230 , n60626 );
not ( n61231 , n61230 );
buf ( n61232 , n61231 );
buf ( n61233 , n61232 );
not ( n61234 , n61233 );
or ( n61235 , n61229 , n61234 );
buf ( n61236 , n61227 );
not ( n61237 , n61236 );
buf ( n61238 , n61237 );
buf ( n61239 , n61238 );
buf ( n61240 , n60626 );
nand ( n61241 , n61239 , n61240 );
buf ( n61242 , n61241 );
buf ( n61243 , n61242 );
nand ( n61244 , n61235 , n61243 );
buf ( n61245 , n61244 );
not ( n61246 , n60527 );
and ( n61247 , n61245 , n61246 );
not ( n61248 , n61245 );
and ( n61249 , n61248 , n60527 );
nor ( n61250 , n61247 , n61249 );
buf ( n61251 , n61250 );
not ( n61252 , n61251 );
xor ( n61253 , n60666 , n60676 );
or ( n61254 , n60779 , n61253 );
nand ( n61255 , n61253 , n60779 );
nand ( n61256 , n61254 , n61255 );
buf ( n61257 , n61256 );
buf ( n61258 , n59651 );
buf ( n61259 , n59688 );
xor ( n61260 , n61258 , n61259 );
buf ( n61261 , n61260 );
xnor ( n61262 , n59676 , n61261 );
buf ( n61263 , n61262 );
not ( n61264 , n61263 );
buf ( n61265 , n61264 );
buf ( n61266 , n61265 );
nand ( n61267 , n61257 , n61266 );
buf ( n61268 , n61267 );
xor ( n61269 , n60736 , n60752 );
xor ( n61270 , n61269 , n60775 );
buf ( n61271 , n61270 );
buf ( n61272 , n61271 );
buf ( n61273 , n46225 );
not ( n61274 , n61273 );
buf ( n61275 , n45750 );
not ( n61276 , n61275 );
buf ( n61277 , n43684 );
not ( n61278 , n61277 );
or ( n61279 , n61276 , n61278 );
buf ( n61280 , n59202 );
not ( n61281 , n61280 );
buf ( n61282 , n53492 );
nand ( n61283 , n61281 , n61282 );
buf ( n61284 , n61283 );
buf ( n61285 , n61284 );
nand ( n61286 , n61279 , n61285 );
buf ( n61287 , n61286 );
buf ( n61288 , n61287 );
not ( n61289 , n61288 );
or ( n61290 , n61274 , n61289 );
buf ( n61291 , n61055 );
buf ( n61292 , n46246 );
nand ( n61293 , n61291 , n61292 );
buf ( n61294 , n61293 );
buf ( n61295 , n61294 );
nand ( n61296 , n61290 , n61295 );
buf ( n61297 , n61296 );
buf ( n61298 , n61297 );
xor ( n61299 , n61272 , n61298 );
buf ( n61300 , n43868 );
not ( n61301 , n61300 );
buf ( n61302 , n60929 );
not ( n61303 , n61302 );
or ( n61304 , n61301 , n61303 );
buf ( n61305 , n41608 );
not ( n61306 , n61305 );
buf ( n61307 , n42425 );
not ( n61308 , n61307 );
or ( n61309 , n61306 , n61308 );
buf ( n61310 , n50043 );
buf ( n61311 , n41611 );
nand ( n61312 , n61310 , n61311 );
buf ( n61313 , n61312 );
buf ( n61314 , n61313 );
nand ( n61315 , n61309 , n61314 );
buf ( n61316 , n61315 );
buf ( n61317 , n61316 );
buf ( n61318 , n44267 );
nand ( n61319 , n61317 , n61318 );
buf ( n61320 , n61319 );
buf ( n61321 , n61320 );
nand ( n61322 , n61304 , n61321 );
buf ( n61323 , n61322 );
buf ( n61324 , n61323 );
and ( n61325 , n12481 , n39481 );
not ( n61326 , n12481 );
and ( n61327 , n61326 , n33080 );
nor ( n61328 , n61325 , n61327 );
buf ( n61329 , n61328 );
not ( n61330 , n61329 );
buf ( n61331 , n42521 );
not ( n61332 , n61331 );
or ( n61333 , n61330 , n61332 );
buf ( n61334 , n42834 );
buf ( n61335 , n60879 );
nand ( n61336 , n61334 , n61335 );
buf ( n61337 , n61336 );
buf ( n61338 , n61337 );
nand ( n61339 , n61333 , n61338 );
buf ( n61340 , n61339 );
buf ( n61341 , n61340 );
xor ( n61342 , n61324 , n61341 );
buf ( n61343 , n42865 );
not ( n61344 , n61343 );
buf ( n61345 , n42471 );
not ( n61346 , n61345 );
or ( n61347 , n61344 , n61346 );
buf ( n61348 , n42468 );
buf ( n61349 , n42862 );
nand ( n61350 , n61348 , n61349 );
buf ( n61351 , n61350 );
buf ( n61352 , n61351 );
nand ( n61353 , n61347 , n61352 );
buf ( n61354 , n61353 );
buf ( n61355 , n61354 );
not ( n61356 , n61355 );
buf ( n61357 , n45059 );
not ( n61358 , n61357 );
or ( n61359 , n61356 , n61358 );
buf ( n61360 , n60714 );
buf ( n61361 , n50104 );
nand ( n61362 , n61360 , n61361 );
buf ( n61363 , n61362 );
buf ( n61364 , n61363 );
nand ( n61365 , n61359 , n61364 );
buf ( n61366 , n61365 );
buf ( n61367 , n61366 );
buf ( n61368 , n43063 );
not ( n61369 , n61368 );
buf ( n61370 , n52551 );
not ( n61371 , n61370 );
or ( n61372 , n61369 , n61371 );
buf ( n61373 , n50591 );
buf ( n61374 , n43064 );
nand ( n61375 , n61373 , n61374 );
buf ( n61376 , n61375 );
buf ( n61377 , n61376 );
nand ( n61378 , n61372 , n61377 );
buf ( n61379 , n61378 );
buf ( n61380 , n61379 );
not ( n61381 , n61380 );
buf ( n61382 , n50608 );
not ( n61383 , n61382 );
or ( n61384 , n61381 , n61383 );
buf ( n61385 , n60959 );
buf ( n61386 , n39983 );
nand ( n61387 , n61385 , n61386 );
buf ( n61388 , n61387 );
buf ( n61389 , n61388 );
nand ( n61390 , n61384 , n61389 );
buf ( n61391 , n61390 );
buf ( n61392 , n61391 );
not ( n61393 , n61392 );
buf ( n61394 , n42336 );
not ( n61395 , n61394 );
buf ( n61396 , n61005 );
not ( n61397 , n61396 );
or ( n61398 , n61395 , n61397 );
buf ( n61399 , n42343 );
not ( n61400 , n61399 );
buf ( n61401 , n47436 );
not ( n61402 , n61401 );
or ( n61403 , n61400 , n61402 );
buf ( n61404 , n50624 );
buf ( n61405 , n46855 );
nand ( n61406 , n61404 , n61405 );
buf ( n61407 , n61406 );
buf ( n61408 , n61407 );
nand ( n61409 , n61403 , n61408 );
buf ( n61410 , n61409 );
buf ( n61411 , n61410 );
buf ( n61412 , n42378 );
nand ( n61413 , n61411 , n61412 );
buf ( n61414 , n61413 );
buf ( n61415 , n61414 );
nand ( n61416 , n61398 , n61415 );
buf ( n61417 , n61416 );
buf ( n61418 , n61417 );
not ( n61419 , n61418 );
or ( n61420 , n61393 , n61419 );
buf ( n61421 , n61391 );
buf ( n61422 , n61417 );
or ( n61423 , n61421 , n61422 );
xor ( n61424 , n59972 , n60056 );
xor ( n61425 , n61424 , n60316 );
buf ( n61426 , n61425 );
not ( n61427 , n61426 );
buf ( n61428 , n48671 );
not ( n61429 , n61428 );
and ( n61430 , n29754 , n41657 );
not ( n61431 , n29754 );
buf ( n61432 , n41656 );
not ( n61433 , n61432 );
buf ( n61434 , n61433 );
and ( n61435 , n61431 , n61434 );
or ( n61436 , n61430 , n61435 );
buf ( n61437 , n61436 );
not ( n61438 , n61437 );
or ( n61439 , n61429 , n61438 );
buf ( n61440 , n41655 );
buf ( n61441 , n61440 );
buf ( n61442 , n61441 );
not ( n61443 , n61442 );
buf ( n61444 , n13653 );
not ( n61445 , n61444 );
buf ( n61446 , n61445 );
not ( n61447 , n61446 );
or ( n61448 , n61443 , n61447 );
buf ( n61449 , n13653 );
buf ( n61450 , n41657 );
nand ( n61451 , n61449 , n61450 );
buf ( n61452 , n61451 );
nand ( n61453 , n61448 , n61452 );
not ( n61454 , n50979 );
nand ( n61455 , n61453 , n61454 );
buf ( n61456 , n61455 );
nand ( n61457 , n61439 , n61456 );
buf ( n61458 , n61457 );
not ( n61459 , n61458 );
or ( n61460 , n61427 , n61459 );
or ( n61461 , n61458 , n61426 );
not ( n61462 , n42556 );
and ( n61463 , n41721 , n61462 );
not ( n61464 , n41721 );
and ( n61465 , n61464 , n54067 );
or ( n61466 , n61463 , n61465 );
buf ( n61467 , n61466 );
not ( n61468 , n61467 );
buf ( n61469 , n61468 );
not ( n61470 , n61469 );
not ( n61471 , n43932 );
and ( n61472 , n61470 , n61471 );
and ( n61473 , n60339 , n43905 );
nor ( n61474 , n61472 , n61473 );
not ( n61475 , n61474 );
nand ( n61476 , n61461 , n61475 );
nand ( n61477 , n61460 , n61476 );
buf ( n61478 , n61477 );
nand ( n61479 , n61423 , n61478 );
buf ( n61480 , n61479 );
buf ( n61481 , n61480 );
nand ( n61482 , n61420 , n61481 );
buf ( n61483 , n61482 );
buf ( n61484 , n61483 );
xor ( n61485 , n61367 , n61484 );
not ( n61486 , n44042 );
buf ( n61487 , n44949 );
buf ( n61488 , n38411 );
and ( n61489 , n61487 , n61488 );
not ( n61490 , n61487 );
buf ( n61491 , n42411 );
and ( n61492 , n61490 , n61491 );
or ( n61493 , n61489 , n61492 );
buf ( n61494 , n61493 );
not ( n61495 , n61494 );
not ( n61496 , n61495 );
or ( n61497 , n61486 , n61496 );
nand ( n61498 , n61022 , n38382 );
nand ( n61499 , n61497 , n61498 );
buf ( n61500 , n61499 );
and ( n61501 , n61485 , n61500 );
and ( n61502 , n61367 , n61484 );
or ( n61503 , n61501 , n61502 );
buf ( n61504 , n61503 );
buf ( n61505 , n61504 );
and ( n61506 , n61342 , n61505 );
and ( n61507 , n61324 , n61341 );
or ( n61508 , n61506 , n61507 );
buf ( n61509 , n61508 );
buf ( n61510 , n61509 );
and ( n61511 , n61299 , n61510 );
and ( n61512 , n61272 , n61298 );
or ( n61513 , n61511 , n61512 );
buf ( n61514 , n61513 );
and ( n61515 , n61268 , n61514 );
nor ( n61516 , n61256 , n61265 );
nor ( n61517 , n61515 , n61516 );
not ( n61518 , n61517 );
and ( n61519 , n60615 , C1 );
or ( n61520 , n61519 , C0 );
buf ( n61521 , n61520 );
buf ( n61522 , n60622 );
xnor ( n61523 , n61521 , n61522 );
buf ( n61524 , n61523 );
not ( n61525 , n61524 );
or ( n61526 , n61518 , n61525 );
or ( n61527 , n61524 , n61517 );
buf ( n61528 , n60540 );
buf ( n61529 , n52456 );
and ( n61530 , n61528 , n61529 );
buf ( n61531 , n48836 );
not ( n61532 , n61531 );
buf ( n61533 , n39280 );
not ( n61534 , n61533 );
or ( n61535 , n61532 , n61534 );
buf ( n61536 , n39277 );
buf ( n61537 , n51493 );
nand ( n61538 , n61536 , n61537 );
buf ( n61539 , n61538 );
buf ( n61540 , n61539 );
nand ( n61541 , n61535 , n61540 );
buf ( n61542 , n61541 );
buf ( n61543 , n61542 );
not ( n61544 , n61543 );
buf ( n61545 , n51489 );
nor ( n61546 , n61544 , n61545 );
buf ( n61547 , n61546 );
buf ( n61548 , n61547 );
nor ( n61549 , n61530 , n61548 );
buf ( n61550 , n61549 );
buf ( n61551 , n61550 );
buf ( n61552 , C1 );
buf ( n61553 , n61552 );
buf ( n61554 , C1 );
buf ( n61555 , n61554 );
buf ( n61556 , C1 );
nand ( n61557 , n61527 , n61556 );
nand ( n61558 , n61526 , n61557 );
buf ( n61559 , n61558 );
not ( n61560 , n61559 );
or ( n61561 , n61252 , n61560 );
xor ( n61562 , n59691 , n59716 );
xor ( n61563 , n61562 , n59721 );
buf ( n61564 , n61563 );
not ( n61565 , n61564 );
not ( n61566 , n59548 );
not ( n61567 , n61566 );
not ( n61568 , n59449 );
or ( n61569 , n61567 , n61568 );
nand ( n61570 , n59448 , n59548 );
nand ( n61571 , n61569 , n61570 );
not ( n61572 , n59453 );
not ( n61573 , n61572 );
and ( n61574 , n61571 , n61573 );
not ( n61575 , n61571 );
and ( n61576 , n61575 , n61572 );
nor ( n61577 , n61574 , n61576 );
not ( n61578 , n61577 );
nand ( n61579 , n61565 , n61578 );
not ( n61580 , n61579 );
xor ( n61581 , n60790 , n60783 );
xnor ( n61582 , n61581 , n60652 );
not ( n61583 , n61582 );
or ( n61584 , n61580 , n61583 );
nand ( n61585 , n61564 , n61577 );
nand ( n61586 , n61584 , n61585 );
buf ( n61587 , n61586 );
nand ( n61588 , n61561 , n61587 );
buf ( n61589 , n61588 );
not ( n61590 , n61250 );
not ( n61591 , n61558 );
nand ( n61592 , n61590 , n61591 );
nand ( n61593 , n61589 , n61592 );
buf ( n61594 , n61593 );
not ( n61595 , n61594 );
xor ( n61596 , n60799 , n60822 );
xor ( n61597 , n61596 , n61201 );
buf ( n61598 , n61597 );
not ( n61599 , n61598 );
or ( n61600 , n61595 , n61599 );
not ( n61601 , n61597 );
buf ( n61602 , n61601 );
not ( n61603 , n61602 );
not ( n61604 , n61593 );
buf ( n61605 , n61604 );
not ( n61606 , n61605 );
or ( n61607 , n61603 , n61606 );
xor ( n61608 , n60832 , n60828 );
xnor ( n61609 , n61608 , n61199 );
not ( n61610 , n61609 );
not ( n61611 , n61610 );
and ( n61612 , n61195 , n60841 );
or ( n61613 , n61612 , C0 );
and ( n61614 , n61613 , n60910 );
not ( n61615 , n61613 );
and ( n61616 , n61615 , n60907 );
nor ( n61617 , n61614 , n61616 );
not ( n61618 , n61617 );
buf ( n61619 , n59777 );
not ( n61620 , n61619 );
buf ( n61621 , n60452 );
not ( n61622 , n61621 );
or ( n61623 , n61620 , n61622 );
buf ( n61624 , n59789 );
buf ( n61625 , n59774 );
nand ( n61626 , n61624 , n61625 );
buf ( n61627 , n61626 );
buf ( n61628 , n61627 );
nand ( n61629 , n61623 , n61628 );
buf ( n61630 , n61629 );
buf ( n61631 , n61630 );
buf ( n61632 , n60445 );
not ( n61633 , n61632 );
buf ( n61634 , n61633 );
buf ( n61635 , n61634 );
and ( n61636 , n61631 , n61635 );
not ( n61637 , n61631 );
buf ( n61638 , n60445 );
and ( n61639 , n61637 , n61638 );
nor ( n61640 , n61636 , n61639 );
buf ( n61641 , n61640 );
not ( n61642 , n61641 );
and ( n61643 , n61618 , n61642 );
not ( n61644 , n37514 );
and ( n61645 , n47725 , n41828 );
not ( n61646 , n47725 );
and ( n61647 , n61646 , n41977 );
nor ( n61648 , n61645 , n61647 );
not ( n61649 , n61648 );
and ( n61650 , n61644 , n61649 );
buf ( n61651 , n60747 );
not ( n61652 , n61651 );
buf ( n61653 , n41973 );
nor ( n61654 , n61652 , n61653 );
buf ( n61655 , n61654 );
nor ( n61656 , n61650 , n61655 );
buf ( n61657 , n61656 );
not ( n61658 , n61657 );
buf ( n61659 , n50060 );
not ( n61660 , n61659 );
buf ( n61661 , n41925 );
not ( n61662 , n61661 );
or ( n61663 , n61660 , n61662 );
buf ( n61664 , n41947 );
buf ( n61665 , n50067 );
nand ( n61666 , n61664 , n61665 );
buf ( n61667 , n61666 );
buf ( n61668 , n61667 );
nand ( n61669 , n61663 , n61668 );
buf ( n61670 , n61669 );
buf ( n61671 , n61670 );
not ( n61672 , n61671 );
buf ( n61673 , n37872 );
not ( n61674 , n61673 );
or ( n61675 , n61672 , n61674 );
buf ( n61676 , n45617 );
buf ( n61677 , n60762 );
nand ( n61678 , n61676 , n61677 );
buf ( n61679 , n61678 );
buf ( n61680 , n61679 );
nand ( n61681 , n61675 , n61680 );
buf ( n61682 , n61681 );
buf ( n61683 , n61682 );
not ( n61684 , n61683 );
buf ( n61685 , n61684 );
buf ( n61686 , n61685 );
not ( n61687 , n61686 );
or ( n61688 , n61658 , n61687 );
xor ( n61689 , n60701 , n60719 );
xor ( n61690 , n61689 , n60731 );
buf ( n61691 , n61690 );
buf ( n61692 , n61691 );
nand ( n61693 , n61688 , n61692 );
buf ( n61694 , n61693 );
buf ( n61695 , n61694 );
buf ( n61696 , n61656 );
not ( n61697 , n61696 );
buf ( n61698 , n61697 );
buf ( n61699 , n61698 );
buf ( n61700 , n61682 );
nand ( n61701 , n61699 , n61700 );
buf ( n61702 , n61701 );
buf ( n61703 , n61702 );
nand ( n61704 , n61695 , n61703 );
buf ( n61705 , n61704 );
buf ( n61706 , n61705 );
buf ( n61707 , n47331 );
not ( n61708 , n61707 );
buf ( n61709 , n51622 );
not ( n61710 , n61709 );
buf ( n61711 , n39240 );
not ( n61712 , n61711 );
or ( n61713 , n61710 , n61712 );
buf ( n61714 , n44300 );
buf ( n61715 , n46875 );
or ( n61716 , n61714 , n61715 );
buf ( n61717 , n61716 );
buf ( n61718 , n61717 );
nand ( n61719 , n61713 , n61718 );
buf ( n61720 , n61719 );
buf ( n61721 , n61720 );
not ( n61722 , n61721 );
or ( n61723 , n61708 , n61722 );
buf ( n61724 , n59821 );
buf ( n61725 , n46912 );
nand ( n61726 , n61724 , n61725 );
buf ( n61727 , n61726 );
buf ( n61728 , n61727 );
nand ( n61729 , n61723 , n61728 );
buf ( n61730 , n61729 );
buf ( n61731 , n61730 );
xor ( n61732 , n61706 , n61731 );
xor ( n61733 , n60947 , n61017 );
xor ( n61734 , n61733 , n61029 );
buf ( n61735 , n61734 );
buf ( n61736 , n61735 );
buf ( n61737 , n37397 );
not ( n61738 , n61737 );
buf ( n61739 , n61738 );
buf ( n61740 , n61739 );
not ( n61741 , n61740 );
buf ( n61742 , n46393 );
buf ( n61743 , n41779 );
and ( n61744 , n61742 , n61743 );
not ( n61745 , n61742 );
buf ( n61746 , n43442 );
and ( n61747 , n61745 , n61746 );
nor ( n61748 , n61744 , n61747 );
buf ( n61749 , n61748 );
buf ( n61750 , n61749 );
not ( n61751 , n61750 );
and ( n61752 , n61741 , n61751 );
buf ( n61753 , n61138 );
not ( n61754 , n61753 );
buf ( n61755 , n37416 );
nor ( n61756 , n61754 , n61755 );
buf ( n61757 , n61756 );
buf ( n61758 , n61757 );
nor ( n61759 , n61752 , n61758 );
buf ( n61760 , n61759 );
buf ( n61761 , n61760 );
not ( n61762 , n61761 );
buf ( n61763 , n61762 );
not ( n61764 , n61763 );
not ( n61765 , n44267 );
not ( n61766 , n41608 );
buf ( n61767 , n29290 );
not ( n61768 , n61767 );
buf ( n61769 , n61768 );
not ( n61770 , n61769 );
or ( n61771 , n61766 , n61770 );
buf ( n61772 , n39653 );
buf ( n61773 , n41611 );
nand ( n61774 , n61772 , n61773 );
buf ( n61775 , n61774 );
nand ( n61776 , n61771 , n61775 );
not ( n61777 , n61776 );
or ( n61778 , n61765 , n61777 );
nand ( n61779 , n61316 , n43868 );
nand ( n61780 , n61778 , n61779 );
not ( n61781 , n61780 );
or ( n61782 , n61764 , n61781 );
not ( n61783 , n61780 );
not ( n61784 , n61783 );
not ( n61785 , n61760 );
or ( n61786 , n61784 , n61785 );
not ( n61787 , n61012 );
not ( n61788 , n60971 );
not ( n61789 , n60990 );
and ( n61790 , n61788 , n61789 );
and ( n61791 , n60971 , n60990 );
nor ( n61792 , n61790 , n61791 );
not ( n61793 , n61792 );
or ( n61794 , n61787 , n61793 );
or ( n61795 , n61012 , n61792 );
nand ( n61796 , n61794 , n61795 );
buf ( n61797 , n61796 );
nand ( n61798 , n61786 , n61797 );
nand ( n61799 , n61782 , n61798 );
buf ( n61800 , n61799 );
xor ( n61801 , n61736 , n61800 );
buf ( n61802 , n53946 );
not ( n61803 , n61802 );
buf ( n61804 , n38068 );
not ( n61805 , n61804 );
or ( n61806 , n61803 , n61805 );
buf ( n61807 , n49391 );
buf ( n61808 , n52094 );
nand ( n61809 , n61807 , n61808 );
buf ( n61810 , n61809 );
buf ( n61811 , n61810 );
nand ( n61812 , n61806 , n61811 );
buf ( n61813 , n61812 );
buf ( n61814 , n61813 );
not ( n61815 , n61814 );
buf ( n61816 , n38130 );
not ( n61817 , n61816 );
or ( n61818 , n61815 , n61817 );
buf ( n61819 , n61068 );
buf ( n61820 , n38060 );
nand ( n61821 , n61819 , n61820 );
buf ( n61822 , n61821 );
buf ( n61823 , n61822 );
nand ( n61824 , n61818 , n61823 );
buf ( n61825 , n61824 );
buf ( n61826 , n61825 );
and ( n61827 , n61801 , n61826 );
and ( n61828 , n61736 , n61800 );
or ( n61829 , n61827 , n61828 );
buf ( n61830 , n61829 );
buf ( n61831 , n61830 );
and ( n61832 , n61732 , n61831 );
and ( n61833 , n61706 , n61731 );
or ( n61834 , n61832 , n61833 );
buf ( n61835 , n61834 );
buf ( n61836 , n61835 );
xor ( n61837 , n61038 , n61063 );
xor ( n61838 , n61837 , n61191 );
buf ( n61839 , n61838 );
buf ( n61840 , n61839 );
xor ( n61841 , n61836 , n61840 );
buf ( n61842 , n52456 );
not ( n61843 , n61842 );
buf ( n61844 , n61542 );
not ( n61845 , n61844 );
or ( n61846 , n61843 , n61845 );
not ( n61847 , n48836 );
buf ( n61848 , n61847 );
buf ( n61849 , n61848 );
buf ( n61850 , n61849 );
buf ( n61851 , n61850 );
not ( n61852 , n61851 );
buf ( n61853 , n61852 );
buf ( n61854 , n61853 );
not ( n61855 , n61854 );
buf ( n61856 , n38218 );
not ( n61857 , n61856 );
or ( n61858 , n61855 , n61857 );
buf ( n61859 , n47969 );
buf ( n61860 , n61850 );
nand ( n61861 , n61859 , n61860 );
buf ( n61862 , n61861 );
buf ( n61863 , n61862 );
nand ( n61864 , n61858 , n61863 );
buf ( n61865 , n61864 );
buf ( n61866 , n61865 );
buf ( n61867 , n51488 );
nand ( n61868 , n61866 , n61867 );
buf ( n61869 , n61868 );
buf ( n61870 , n61869 );
nand ( n61871 , n61846 , n61870 );
buf ( n61872 , n61871 );
xor ( n61873 , n60865 , n60890 );
xor ( n61874 , n61873 , n60898 );
buf ( n61875 , n61874 );
xor ( n61876 , n61872 , n61875 );
buf ( n61877 , n44496 );
not ( n61878 , n61877 );
buf ( n61879 , n61090 );
not ( n61880 , n61879 );
or ( n61881 , n61878 , n61880 );
buf ( n61882 , n44533 );
not ( n61883 , n61882 );
buf ( n61884 , n42461 );
not ( n61885 , n61884 );
or ( n61886 , n61883 , n61885 );
nand ( n61887 , n38821 , n44530 );
buf ( n61888 , n61887 );
nand ( n61889 , n61886 , n61888 );
buf ( n61890 , n61889 );
buf ( n61891 , n61890 );
buf ( n61892 , n44708 );
nand ( n61893 , n61891 , n61892 );
buf ( n61894 , n61893 );
buf ( n61895 , n61894 );
nand ( n61896 , n61881 , n61895 );
buf ( n61897 , n61896 );
buf ( n61898 , n61897 );
buf ( n61899 , n53539 );
not ( n61900 , n61899 );
buf ( n61901 , n43104 );
not ( n61902 , n61901 );
or ( n61903 , n61900 , n61902 );
buf ( n61904 , n43095 );
buf ( n61905 , n53548 );
nand ( n61906 , n61904 , n61905 );
buf ( n61907 , n61906 );
buf ( n61908 , n61907 );
nand ( n61909 , n61903 , n61908 );
buf ( n61910 , n61909 );
buf ( n61911 , n61910 );
not ( n61912 , n61911 );
buf ( n61913 , n45423 );
not ( n61914 , n61913 );
or ( n61915 , n61912 , n61914 );
buf ( n61916 , n44679 );
buf ( n61917 , n60419 );
nand ( n61918 , n61916 , n61917 );
buf ( n61919 , n61918 );
buf ( n61920 , n61919 );
nand ( n61921 , n61915 , n61920 );
buf ( n61922 , n61921 );
buf ( n61923 , n61922 );
xor ( n61924 , n61898 , n61923 );
buf ( n61925 , n48671 );
not ( n61926 , n61925 );
buf ( n61927 , n59924 );
not ( n61928 , n61927 );
or ( n61929 , n61926 , n61928 );
buf ( n61930 , n61436 );
buf ( n61931 , n50982 );
nand ( n61932 , n61930 , n61931 );
buf ( n61933 , n61932 );
buf ( n61934 , n61933 );
nand ( n61935 , n61929 , n61934 );
buf ( n61936 , n61935 );
buf ( n61937 , n61936 );
buf ( n61938 , n42008 );
not ( n61939 , n61938 );
buf ( n61940 , n52670 );
not ( n61941 , n61940 );
or ( n61942 , n61939 , n61941 );
buf ( n61943 , n52673 );
buf ( n61944 , n55708 );
nand ( n61945 , n61943 , n61944 );
buf ( n61946 , n61945 );
buf ( n61947 , n61946 );
nand ( n61948 , n61942 , n61947 );
buf ( n61949 , n61948 );
buf ( n61950 , n61949 );
not ( n61951 , n61950 );
buf ( n61952 , n42628 );
not ( n61953 , n61952 );
or ( n61954 , n61951 , n61953 );
buf ( n61955 , n60985 );
buf ( n61956 , n47872 );
nand ( n61957 , n61955 , n61956 );
buf ( n61958 , n61957 );
buf ( n61959 , n61958 );
nand ( n61960 , n61954 , n61959 );
buf ( n61961 , n61960 );
buf ( n61962 , n61961 );
xor ( n61963 , n61937 , n61962 );
xor ( n61964 , n59953 , n60321 );
xor ( n61965 , n61964 , n60352 );
buf ( n61966 , n61965 );
buf ( n61967 , n61966 );
and ( n61968 , n61963 , n61967 );
and ( n61969 , n61937 , n61962 );
or ( n61970 , n61968 , n61969 );
buf ( n61971 , n61970 );
buf ( n61972 , n61971 );
not ( n61973 , n42252 );
and ( n61974 , n42119 , n59242 );
not ( n61975 , n42119 );
and ( n61976 , n61975 , n42263 );
or ( n61977 , n61974 , n61976 );
not ( n61978 , n61977 );
or ( n61979 , n61973 , n61978 );
buf ( n61980 , n61168 );
buf ( n61981 , n42315 );
nand ( n61982 , n61980 , n61981 );
buf ( n61983 , n61982 );
nand ( n61984 , n61979 , n61983 );
buf ( n61985 , n61984 );
xor ( n61986 , n61972 , n61985 );
buf ( n61987 , n39715 );
buf ( n61988 , n12481 );
and ( n61989 , n61987 , n61988 );
buf ( n61990 , n61989 );
buf ( n61991 , n61990 );
and ( n61992 , n61986 , n61991 );
and ( n61993 , n61972 , n61985 );
or ( n61994 , n61992 , n61993 );
buf ( n61995 , n61994 );
buf ( n61996 , n61995 );
and ( n61997 , n61924 , n61996 );
and ( n61998 , n61898 , n61923 );
or ( n61999 , n61997 , n61998 );
buf ( n62000 , n61999 );
and ( n62001 , n61876 , n62000 );
and ( n62002 , n61872 , n61875 );
or ( n62003 , n62001 , n62002 );
buf ( n62004 , n62003 );
and ( n62005 , n61841 , n62004 );
and ( n62006 , n61836 , n61840 );
or ( n62007 , n62005 , n62006 );
buf ( n62008 , n62007 );
buf ( n62009 , n61617 );
buf ( n62010 , n61641 );
nand ( n62011 , n62009 , n62010 );
buf ( n62012 , n62011 );
and ( n62013 , n62008 , n62012 );
nor ( n62014 , n61643 , n62013 );
not ( n62015 , n62014 );
not ( n62016 , n62015 );
or ( n62017 , n61611 , n62016 );
buf ( n62018 , n61609 );
not ( n62019 , n62018 );
buf ( n62020 , n62014 );
not ( n62021 , n62020 );
or ( n62022 , n62019 , n62021 );
xor ( n62023 , n59761 , n60459 );
xor ( n62024 , n62023 , n60466 );
buf ( n62025 , n62024 );
nand ( n62026 , n62022 , n62025 );
buf ( n62027 , n62026 );
nand ( n62028 , n62017 , n62027 );
buf ( n62029 , n62028 );
nand ( n62030 , n61607 , n62029 );
buf ( n62031 , n62030 );
buf ( n62032 , n62031 );
nand ( n62033 , n61600 , n62032 );
buf ( n62034 , n62033 );
buf ( n62035 , n62034 );
xor ( n62036 , n61223 , n62035 );
xor ( n62037 , n59157 , n59623 );
xor ( n62038 , n62037 , n60481 );
buf ( n62039 , n62038 );
buf ( n62040 , n62039 );
and ( n62041 , n62036 , n62040 );
and ( n62042 , n61223 , n62035 );
or ( n62043 , n62041 , n62042 );
buf ( n62044 , n62043 );
buf ( n62045 , n62044 );
not ( n62046 , n62045 );
buf ( n62047 , n62046 );
nand ( n62048 , n61209 , n62047 );
buf ( n62049 , n62048 );
xor ( n62050 , n61223 , n62035 );
xor ( n62051 , n62050 , n62040 );
buf ( n62052 , n62051 );
buf ( n62053 , n62052 );
not ( n62054 , n62053 );
buf ( n62055 , n62054 );
not ( n62056 , n62028 );
not ( n62057 , n61593 );
not ( n62058 , n61601 );
or ( n62059 , n62057 , n62058 );
or ( n62060 , n61601 , n61593 );
nand ( n62061 , n62059 , n62060 );
not ( n62062 , n62061 );
or ( n62063 , n62056 , n62062 );
not ( n62064 , n61593 );
not ( n62065 , n61601 );
or ( n62066 , n62064 , n62065 );
or ( n62067 , n61601 , n61593 );
nand ( n62068 , n62066 , n62067 );
or ( n62069 , n62068 , n62028 );
nand ( n62070 , n62063 , n62069 );
buf ( n62071 , n62070 );
not ( n62072 , n62071 );
buf ( n62073 , n62072 );
not ( n62074 , n62073 );
buf ( n62075 , n59756 );
buf ( n62076 , n59627 );
and ( n62077 , n62075 , n62076 );
not ( n62078 , n62075 );
buf ( n62079 , n59627 );
not ( n62080 , n62079 );
buf ( n62081 , n62080 );
buf ( n62082 , n62081 );
and ( n62083 , n62078 , n62082 );
nor ( n62084 , n62077 , n62083 );
buf ( n62085 , n62084 );
buf ( n62086 , n62085 );
buf ( n62087 , n60469 );
and ( n62088 , n62086 , n62087 );
not ( n62089 , n62086 );
buf ( n62090 , n60469 );
not ( n62091 , n62090 );
buf ( n62092 , n62091 );
buf ( n62093 , n62092 );
and ( n62094 , n62089 , n62093 );
nor ( n62095 , n62088 , n62094 );
buf ( n62096 , n62095 );
not ( n62097 , n62096 );
or ( n62098 , n62074 , n62097 );
buf ( n62099 , n62096 );
not ( n62100 , n62099 );
buf ( n62101 , n62100 );
not ( n62102 , n62101 );
not ( n62103 , n62070 );
or ( n62104 , n62102 , n62103 );
xor ( n62105 , n61586 , n61250 );
xnor ( n62106 , n62105 , n61591 );
buf ( n62107 , n62106 );
not ( n62108 , n62107 );
buf ( n62109 , n62108 );
buf ( n62110 , n62109 );
not ( n62111 , n62110 );
xor ( n62112 , n61836 , n61840 );
xor ( n62113 , n62112 , n62004 );
buf ( n62114 , n62113 );
not ( n62115 , n62114 );
buf ( n62116 , n61262 );
buf ( n62117 , n61514 );
xor ( n62118 , n62116 , n62117 );
buf ( n62119 , n61256 );
xnor ( n62120 , n62118 , n62119 );
buf ( n62121 , n62120 );
buf ( n62122 , n62121 );
not ( n62123 , n62122 );
buf ( n62124 , n61865 );
not ( n62125 , n51473 );
buf ( n62126 , n62125 );
and ( n62127 , n62124 , n62126 );
and ( n62128 , n38244 , n51493 );
not ( n62129 , n38244 );
and ( n62130 , n62129 , n48836 );
or ( n62131 , n62128 , n62130 );
buf ( n62132 , n62131 );
buf ( n62133 , n51488 );
and ( n62134 , n62132 , n62133 );
buf ( n62135 , n62134 );
buf ( n62136 , n62135 );
nor ( n62137 , n62127 , n62136 );
buf ( n62138 , n62137 );
buf ( n62139 , n62138 );
not ( n62140 , n62139 );
buf ( n62141 , n62140 );
buf ( n62142 , n62141 );
not ( n62143 , n62142 );
buf ( n62144 , n48868 );
not ( n62145 , n62144 );
and ( n62146 , n48808 , n43879 );
not ( n62147 , n48808 );
and ( n62148 , n62147 , n37265 );
or ( n62149 , n62146 , n62148 );
buf ( n62150 , n62149 );
not ( n62151 , n62150 );
or ( n62152 , n62145 , n62151 );
buf ( n62153 , n48821 );
not ( n62154 , n62153 );
buf ( n62155 , n62154 );
buf ( n62156 , n62155 );
not ( n62157 , n62156 );
buf ( n62158 , n43224 );
not ( n62159 , n62158 );
or ( n62160 , n62157 , n62159 );
buf ( n62161 , n37293 );
buf ( n62162 , n48821 );
nand ( n62163 , n62161 , n62162 );
buf ( n62164 , n62163 );
buf ( n62165 , n62164 );
nand ( n62166 , n62160 , n62165 );
buf ( n62167 , n62166 );
buf ( n62168 , n62167 );
buf ( n62169 , n48855 );
nand ( n62170 , n62168 , n62169 );
buf ( n62171 , n62170 );
buf ( n62172 , n62171 );
nand ( n62173 , n62152 , n62172 );
buf ( n62174 , n62173 );
buf ( n62175 , n62174 );
not ( n62176 , n62175 );
or ( n62177 , n62143 , n62176 );
buf ( n62178 , n62174 );
not ( n62179 , n62178 );
buf ( n62180 , n62179 );
buf ( n62181 , n62180 );
not ( n62182 , n62181 );
buf ( n62183 , n62138 );
not ( n62184 , n62183 );
or ( n62185 , n62182 , n62184 );
buf ( n62186 , n52780 );
not ( n62187 , n62186 );
buf ( n62188 , n38068 );
not ( n62189 , n62188 );
or ( n62190 , n62187 , n62189 );
buf ( n62191 , n49391 );
buf ( n62192 , n52789 );
nand ( n62193 , n62191 , n62192 );
buf ( n62194 , n62193 );
buf ( n62195 , n62194 );
nand ( n62196 , n62190 , n62195 );
buf ( n62197 , n62196 );
buf ( n62198 , n62197 );
not ( n62199 , n62198 );
buf ( n62200 , n46165 );
not ( n62201 , n62200 );
or ( n62202 , n62199 , n62201 );
buf ( n62203 , n61813 );
buf ( n62204 , n47108 );
nand ( n62205 , n62203 , n62204 );
buf ( n62206 , n62205 );
buf ( n62207 , n62206 );
nand ( n62208 , n62202 , n62207 );
buf ( n62209 , n62208 );
buf ( n62210 , n62209 );
buf ( n62211 , n46225 );
not ( n62212 , n62211 );
buf ( n62213 , n53492 );
not ( n62214 , n62213 );
buf ( n62215 , n39701 );
not ( n62216 , n62215 );
or ( n62217 , n62214 , n62216 );
not ( n62218 , n39203 );
not ( n62219 , n37639 );
or ( n62220 , n62218 , n62219 );
nand ( n62221 , n62220 , n45747 );
buf ( n62222 , n62221 );
nand ( n62223 , n62217 , n62222 );
buf ( n62224 , n62223 );
buf ( n62225 , n62224 );
not ( n62226 , n62225 );
or ( n62227 , n62212 , n62226 );
buf ( n62228 , n53492 );
not ( n62229 , n62228 );
buf ( n62230 , n37589 );
not ( n62231 , n62230 );
or ( n62232 , n62229 , n62231 );
buf ( n62233 , n39489 );
buf ( n62234 , n45747 );
nand ( n62235 , n62233 , n62234 );
buf ( n62236 , n62235 );
buf ( n62237 , n62236 );
nand ( n62238 , n62232 , n62237 );
buf ( n62239 , n62238 );
buf ( n62240 , n62239 );
buf ( n62241 , n46246 );
nand ( n62242 , n62240 , n62241 );
buf ( n62243 , n62242 );
buf ( n62244 , n62243 );
nand ( n62245 , n62227 , n62244 );
buf ( n62246 , n62245 );
buf ( n62247 , n62246 );
xor ( n62248 , n62210 , n62247 );
buf ( n62249 , n55841 );
not ( n62250 , n62249 );
buf ( n62251 , n44689 );
not ( n62252 , n62251 );
or ( n62253 , n62250 , n62252 );
buf ( n62254 , n39136 );
buf ( n62255 , n58361 );
nand ( n62256 , n62254 , n62255 );
buf ( n62257 , n62256 );
buf ( n62258 , n62257 );
nand ( n62259 , n62253 , n62258 );
buf ( n62260 , n62259 );
buf ( n62261 , n62260 );
not ( n62262 , n62261 );
buf ( n62263 , n45423 );
not ( n62264 , n62263 );
or ( n62265 , n62262 , n62264 );
buf ( n62266 , n44679 );
buf ( n62267 , n61910 );
nand ( n62268 , n62266 , n62267 );
buf ( n62269 , n62268 );
buf ( n62270 , n62269 );
nand ( n62271 , n62265 , n62270 );
buf ( n62272 , n62271 );
buf ( n62273 , n62272 );
and ( n62274 , n62248 , n62273 );
and ( n62275 , n62210 , n62247 );
or ( n62276 , n62274 , n62275 );
buf ( n62277 , n62276 );
buf ( n62278 , n62277 );
nand ( n62279 , n62185 , n62278 );
buf ( n62280 , n62279 );
buf ( n62281 , n62280 );
nand ( n62282 , n62177 , n62281 );
buf ( n62283 , n62282 );
buf ( n62284 , n62283 );
xor ( n62285 , n61272 , n61298 );
xor ( n62286 , n62285 , n61510 );
buf ( n62287 , n62286 );
buf ( n62288 , n62287 );
xor ( n62289 , n62284 , n62288 );
xor ( n62290 , n61706 , n61731 );
xor ( n62291 , n62290 , n61831 );
buf ( n62292 , n62291 );
buf ( n62293 , n62292 );
and ( n62294 , n62289 , n62293 );
and ( n62295 , n62284 , n62288 );
or ( n62296 , n62294 , n62295 );
buf ( n62297 , n62296 );
buf ( n62298 , n62297 );
not ( n62299 , n62298 );
buf ( n62300 , n62299 );
buf ( n62301 , n62300 );
nand ( n62302 , n62123 , n62301 );
buf ( n62303 , n62302 );
not ( n62304 , n62303 );
or ( n62305 , n62115 , n62304 );
buf ( n62306 , n62121 );
not ( n62307 , n62306 );
buf ( n62308 , n62300 );
nor ( n62309 , n62307 , n62308 );
buf ( n62310 , n62309 );
not ( n62311 , n62310 );
nand ( n62312 , n62305 , n62311 );
not ( n62313 , n62312 );
and ( n62314 , n61268 , n61514 );
nor ( n62315 , n62314 , n61516 );
not ( n62316 , n62315 );
not ( n62317 , n62316 );
or ( n62318 , C0 , n62317 );
nand ( n62319 , C0 , n62315 );
nand ( n62320 , n62318 , n62319 );
and ( n62321 , n62320 , n61524 );
not ( n62322 , n62320 );
not ( n62323 , n61524 );
and ( n62324 , n62322 , n62323 );
nor ( n62325 , n62321 , n62324 );
not ( n62326 , n62325 );
not ( n62327 , n62326 );
or ( n62328 , n62313 , n62327 );
not ( n62329 , n62114 );
not ( n62330 , n62303 );
or ( n62331 , n62329 , n62330 );
nand ( n62332 , n62331 , n62311 );
not ( n62333 , n62325 );
or ( n62334 , n62332 , n62333 );
not ( n62335 , n62008 );
not ( n62336 , n62335 );
not ( n62337 , n61617 );
or ( n62338 , n62336 , n62337 );
not ( n62339 , n61617 );
nand ( n62340 , n62339 , n62008 );
nand ( n62341 , n62338 , n62340 );
buf ( n62342 , n61641 );
and ( n62343 , n62341 , n62342 );
not ( n62344 , n62341 );
not ( n62345 , n62342 );
and ( n62346 , n62344 , n62345 );
nor ( n62347 , n62343 , n62346 );
nand ( n62348 , n62334 , n62347 );
nand ( n62349 , n62328 , n62348 );
not ( n62350 , n62349 );
buf ( n62351 , n62350 );
not ( n62352 , n62351 );
or ( n62353 , n62111 , n62352 );
xor ( n62354 , n59828 , n59837 );
xor ( n62355 , n62354 , n60442 );
buf ( n62356 , n61691 );
buf ( n62357 , n61682 );
xor ( n62358 , n62356 , n62357 );
buf ( n62359 , n61698 );
xnor ( n62360 , n62358 , n62359 );
buf ( n62361 , n62360 );
buf ( n62362 , n62361 );
not ( n62363 , n62362 );
or ( n62364 , n44316 , n46890 );
or ( n62365 , n42596 , n51622 );
nand ( n62366 , n62364 , n62365 );
buf ( n62367 , n62366 );
not ( n62368 , n62367 );
buf ( n62369 , n46910 );
not ( n62370 , n62369 );
and ( n62371 , n62368 , n62370 );
buf ( n62372 , n61720 );
buf ( n62373 , n46912 );
and ( n62374 , n62372 , n62373 );
nor ( n62375 , n62371 , n62374 );
buf ( n62376 , n62375 );
buf ( n62377 , n62376 );
not ( n62378 , n62377 );
or ( n62379 , n62363 , n62378 );
not ( n62380 , n43798 );
buf ( n62381 , n51001 );
buf ( n62382 , n49228 );
and ( n62383 , n62381 , n62382 );
not ( n62384 , n62381 );
buf ( n62385 , n49879 );
and ( n62386 , n62384 , n62385 );
nor ( n62387 , n62383 , n62386 );
buf ( n62388 , n62387 );
not ( n62389 , n62388 );
and ( n62390 , n62380 , n62389 );
and ( n62391 , n45617 , n61670 );
nor ( n62392 , n62390 , n62391 );
not ( n62393 , n62392 );
buf ( n62394 , n37514 );
not ( n62395 , n62394 );
buf ( n62396 , n48320 );
buf ( n62397 , n37474 );
and ( n62398 , n62396 , n62397 );
not ( n62399 , n62396 );
buf ( n62400 , n41839 );
and ( n62401 , n62399 , n62400 );
nor ( n62402 , n62398 , n62401 );
buf ( n62403 , n62402 );
buf ( n62404 , n62403 );
not ( n62405 , n62404 );
and ( n62406 , n62395 , n62405 );
buf ( n62407 , n47725 );
buf ( n62408 , n41839 );
and ( n62409 , n62407 , n62408 );
not ( n62410 , n62407 );
buf ( n62411 , n41978 );
and ( n62412 , n62410 , n62411 );
or ( n62413 , n62409 , n62412 );
buf ( n62414 , n62413 );
buf ( n62415 , n62414 );
buf ( n62416 , n37449 );
nor ( n62417 , n62415 , n62416 );
buf ( n62418 , n62417 );
buf ( n62419 , n62418 );
nor ( n62420 , n62406 , n62419 );
buf ( n62421 , n62420 );
not ( n62422 , n62421 );
or ( n62423 , n62393 , n62422 );
xor ( n62424 , n60357 , n59937 );
xnor ( n62425 , n62424 , n60395 );
nand ( n62426 , n62423 , n62425 );
buf ( n62427 , n62426 );
buf ( n62428 , n62421 );
not ( n62429 , n62428 );
buf ( n62430 , n62392 );
not ( n62431 , n62430 );
buf ( n62432 , n62431 );
buf ( n62433 , n62432 );
nand ( n62434 , n62429 , n62433 );
buf ( n62435 , n62434 );
buf ( n62436 , n62435 );
nand ( n62437 , n62427 , n62436 );
buf ( n62438 , n62437 );
buf ( n62439 , n62438 );
nand ( n62440 , n62379 , n62439 );
buf ( n62441 , n62440 );
buf ( n62442 , n62441 );
buf ( n62443 , n62376 );
not ( n62444 , n62443 );
buf ( n62445 , n62361 );
not ( n62446 , n62445 );
buf ( n62447 , n62446 );
buf ( n62448 , n62447 );
nand ( n62449 , n62444 , n62448 );
buf ( n62450 , n62449 );
buf ( n62451 , n62450 );
nand ( n62452 , n62442 , n62451 );
buf ( n62453 , n62452 );
buf ( n62454 , n62453 );
buf ( n62455 , C0 );
or ( n62456 , n62454 , n62455 );
buf ( n62457 , n61287 );
buf ( n62458 , n46246 );
and ( n62459 , n62457 , n62458 );
buf ( n62460 , n62239 );
not ( n62461 , n62460 );
buf ( n62462 , n45742 );
nor ( n62463 , n62461 , n62462 );
buf ( n62464 , n62463 );
buf ( n62465 , n62464 );
nor ( n62466 , n62459 , n62465 );
buf ( n62467 , n62466 );
not ( n62468 , n62467 );
not ( n62469 , n62468 );
xor ( n62470 , n61126 , n61175 );
xnor ( n62471 , n62470 , n61150 );
not ( n62472 , n62471 );
not ( n62473 , n62472 );
or ( n62474 , n62469 , n62473 );
not ( n62475 , n62467 );
not ( n62476 , n62471 );
or ( n62477 , n62475 , n62476 );
not ( n62478 , n59864 );
not ( n62479 , n59860 );
not ( n62480 , n62479 );
or ( n62481 , n62478 , n62480 );
not ( n62482 , n59864 );
nand ( n62483 , n62482 , n59860 );
nand ( n62484 , n62481 , n62483 );
xor ( n62485 , n62484 , n60399 );
not ( n62486 , n62485 );
nand ( n62487 , n62477 , n62486 );
nand ( n62488 , n62474 , n62487 );
buf ( n62489 , n62488 );
nand ( n62490 , n62456 , n62489 );
buf ( n62491 , n62490 );
nand ( n62492 , C1 , n62491 );
xor ( n62493 , n62355 , n62492 );
xor ( n62494 , n60410 , n60413 );
xor ( n62495 , n62494 , n60438 );
buf ( n62496 , n62495 );
buf ( n62497 , C0 );
buf ( n62498 , n62496 );
buf ( n62499 , n62497 );
or ( n62500 , n62498 , n62499 );
buf ( n62501 , n60373 );
buf ( n62502 , n42668 );
and ( n62503 , n62501 , n62502 );
buf ( n62504 , n47072 );
not ( n62505 , n62504 );
buf ( n62506 , n25226 );
not ( n62507 , n62506 );
or ( n62508 , n62505 , n62507 );
buf ( n62509 , n50575 );
not ( n62510 , n25226 );
buf ( n62511 , n62510 );
nand ( n62512 , n62509 , n62511 );
buf ( n62513 , n62512 );
buf ( n62514 , n62513 );
nand ( n62515 , n62508 , n62514 );
buf ( n62516 , n62515 );
buf ( n62517 , n62516 );
not ( n62518 , n62517 );
buf ( n62519 , n42711 );
nor ( n62520 , n62518 , n62519 );
buf ( n62521 , n62520 );
buf ( n62522 , n62521 );
nor ( n62523 , n62503 , n62522 );
buf ( n62524 , n62523 );
buf ( n62525 , n62524 );
not ( n62526 , n62525 );
buf ( n62527 , n42847 );
not ( n62528 , n62527 );
buf ( n62529 , n38994 );
not ( n62530 , n62529 );
or ( n62531 , n62528 , n62530 );
buf ( n62532 , n42468 );
buf ( n62533 , n46691 );
nand ( n62534 , n62532 , n62533 );
buf ( n62535 , n62534 );
buf ( n62536 , n62535 );
nand ( n62537 , n62531 , n62536 );
buf ( n62538 , n62537 );
buf ( n62539 , n62538 );
not ( n62540 , n62539 );
buf ( n62541 , n47050 );
not ( n62542 , n62541 );
or ( n62543 , n62540 , n62542 );
buf ( n62544 , n61354 );
buf ( n62545 , n52595 );
nand ( n62546 , n62544 , n62545 );
buf ( n62547 , n62546 );
buf ( n62548 , n62547 );
nand ( n62549 , n62543 , n62548 );
buf ( n62550 , n62549 );
buf ( n62551 , n62550 );
not ( n62552 , n62551 );
buf ( n62553 , n62552 );
buf ( n62554 , n62553 );
not ( n62555 , n62554 );
or ( n62556 , n62526 , n62555 );
buf ( n62557 , n42336 );
not ( n62558 , n62557 );
buf ( n62559 , n61410 );
not ( n62560 , n62559 );
or ( n62561 , n62558 , n62560 );
and ( n62562 , n28368 , n46855 );
not ( n62563 , n28368 );
and ( n62564 , n62563 , n42343 );
or ( n62565 , n62562 , n62564 );
buf ( n62566 , n62565 );
buf ( n62567 , n42378 );
nand ( n62568 , n62566 , n62567 );
buf ( n62569 , n62568 );
buf ( n62570 , n62569 );
nand ( n62571 , n62561 , n62570 );
buf ( n62572 , n62571 );
buf ( n62573 , n62572 );
xor ( n62574 , n60028 , n60048 );
xor ( n62575 , n62574 , n60052 );
xor ( n62576 , n60201 , n60310 );
xor ( n62577 , n62575 , n62576 );
buf ( n62578 , n62577 );
not ( n62579 , n41642 );
buf ( n62580 , n62579 );
not ( n62581 , n62580 );
buf ( n62582 , n62581 );
not ( n62583 , n62582 );
not ( n62584 , n61453 );
or ( n62585 , n62583 , n62584 );
buf ( n62586 , n50979 );
not ( n62587 , n62586 );
buf ( n62588 , n62587 );
buf ( n62589 , n62588 );
buf ( n62590 , n61442 );
not ( n62591 , n62590 );
buf ( n62592 , n60330 );
not ( n62593 , n62592 );
or ( n62594 , n62591 , n62593 );
buf ( n62595 , n41736 );
buf ( n62596 , n61442 );
not ( n62597 , n62596 );
buf ( n62598 , n62597 );
buf ( n62599 , n62598 );
nand ( n62600 , n62595 , n62599 );
buf ( n62601 , n62600 );
buf ( n62602 , n62601 );
nand ( n62603 , n62594 , n62602 );
buf ( n62604 , n62603 );
buf ( n62605 , n62604 );
nand ( n62606 , n62589 , n62605 );
buf ( n62607 , n62606 );
nand ( n62608 , n62585 , n62607 );
buf ( n62609 , n62608 );
or ( n62610 , n62578 , n62609 );
buf ( n62611 , n60226 );
buf ( n62612 , n60237 );
or ( n62613 , n62611 , n62612 );
buf ( n62614 , n60240 );
nand ( n62615 , n62613 , n62614 );
buf ( n62616 , n62615 );
buf ( n62617 , n62616 );
buf ( n62618 , n58823 );
buf ( n62619 , n56641 );
and ( n62620 , n62618 , n62619 );
buf ( n62621 , n58862 );
buf ( n62622 , n56631 );
and ( n62623 , n62621 , n62622 );
nor ( n62624 , n62620 , n62623 );
buf ( n62625 , n62624 );
buf ( n62626 , n62625 );
buf ( n62627 , n56626 );
or ( n62628 , n62626 , n62627 );
buf ( n62629 , n60148 );
buf ( n62630 , n56639 );
or ( n62631 , n62629 , n62630 );
nand ( n62632 , n62628 , n62631 );
buf ( n62633 , n62632 );
buf ( n62634 , n62633 );
xor ( n62635 , n62617 , n62634 );
not ( n62636 , n54574 );
not ( n62637 , n55068 );
or ( n62638 , n62636 , n62637 );
not ( n62639 , n55071 );
nand ( n62640 , n62638 , n62639 );
not ( n62641 , n55073 );
nand ( n62642 , n62641 , n54526 );
xnor ( n62643 , n62640 , n62642 );
buf ( n62644 , n62643 );
not ( n62645 , n62644 );
buf ( n62646 , n62645 );
buf ( n62647 , n62646 );
buf ( n62648 , n56589 );
or ( n62649 , n62647 , n62648 );
buf ( n62650 , n60229 );
not ( n62651 , n62650 );
buf ( n62652 , n62651 );
buf ( n62653 , n62652 );
buf ( n62654 , n56598 );
or ( n62655 , n62653 , n62654 );
nand ( n62656 , n62649 , n62655 );
buf ( n62657 , n62656 );
buf ( n62658 , n62657 );
buf ( n62659 , n10265 );
buf ( n62660 , n62659 );
not ( n62661 , n62660 );
buf ( n62662 , n62661 );
not ( n62663 , n60096 );
or ( n62664 , n62662 , n62663 );
or ( n62665 , n62659 , n60096 );
nand ( n62666 , n62664 , n62665 );
buf ( n62667 , n62666 );
buf ( n62668 , n3049 );
buf ( n62669 , n62668 );
buf ( n62670 , n62662 );
and ( n62671 , n62669 , n62670 );
not ( n62672 , n62669 );
buf ( n62673 , n62659 );
and ( n62674 , n62672 , n62673 );
or ( n62675 , n62671 , n62674 );
buf ( n62676 , n62675 );
buf ( n62677 , n62676 );
and ( n62678 , n62667 , n62677 );
buf ( n62679 , n62678 );
buf ( n62680 , n62679 );
buf ( n62681 , n60096 );
buf ( n62682 , n62681 );
not ( n62683 , n62682 );
buf ( n62684 , n62683 );
buf ( n62685 , n62684 );
nand ( n62686 , n62680 , n62685 );
buf ( n62687 , n62686 );
buf ( n62688 , n62687 );
buf ( n62689 , n62676 );
not ( n62690 , n62689 );
buf ( n62691 , n62690 );
buf ( n62692 , n62691 );
buf ( n62693 , n62663 );
nand ( n62694 , n62692 , n62693 );
buf ( n62695 , n62694 );
buf ( n62696 , n62695 );
and ( n62697 , n62688 , n62696 );
buf ( n62698 , n62697 );
buf ( n62699 , n62698 );
xor ( n62700 , n62658 , n62699 );
buf ( n62701 , n60068 );
buf ( n62702 , n56652 );
and ( n62703 , n62701 , n62702 );
buf ( n62704 , n60071 );
buf ( n62705 , n55201 );
and ( n62706 , n62704 , n62705 );
nor ( n62707 , n62703 , n62706 );
buf ( n62708 , n62707 );
buf ( n62709 , n62708 );
buf ( n62710 , n56664 );
or ( n62711 , n62709 , n62710 );
buf ( n62712 , n60212 );
buf ( n62713 , n56673 );
or ( n62714 , n62712 , n62713 );
nand ( n62715 , n62711 , n62714 );
buf ( n62716 , n62715 );
buf ( n62717 , n62716 );
and ( n62718 , n62700 , n62717 );
and ( n62719 , n62658 , n62699 );
or ( n62720 , n62718 , n62719 );
buf ( n62721 , n62720 );
buf ( n62722 , n62721 );
and ( n62723 , n62635 , n62722 );
and ( n62724 , n62617 , n62634 );
or ( n62725 , n62723 , n62724 );
buf ( n62726 , n62725 );
xor ( n62727 , n60157 , n60174 );
xor ( n62728 , n62727 , n60192 );
buf ( n62729 , n62728 );
xor ( n62730 , n62726 , n62729 );
xor ( n62731 , n60082 , n60111 );
xor ( n62732 , n62731 , n60128 );
xor ( n62733 , n60240 , n60295 );
xor ( n62734 , n62732 , n62733 );
and ( n62735 , n62730 , n62734 );
and ( n62736 , n62726 , n62729 );
or ( n62737 , n62735 , n62736 );
xor ( n62738 , n60300 , n60303 );
xor ( n62739 , n62738 , n60307 );
and ( n62740 , n62737 , n62739 );
buf ( n62741 , n55113 );
buf ( n62742 , n60261 );
and ( n62743 , n62741 , n62742 );
buf ( n62744 , n56655 );
buf ( n62745 , n60090 );
and ( n62746 , n62744 , n62745 );
nor ( n62747 , n62743 , n62746 );
buf ( n62748 , n62747 );
buf ( n62749 , n62748 );
buf ( n62750 , n60270 );
or ( n62751 , n62749 , n62750 );
buf ( n62752 , n60268 );
buf ( n62753 , n60100 );
or ( n62754 , n62752 , n62753 );
nand ( n62755 , n62751 , n62754 );
buf ( n62756 , n62755 );
buf ( n62757 , n62756 );
buf ( n62758 , n60229 );
buf ( n62759 , n56652 );
and ( n62760 , n62758 , n62759 );
buf ( n62761 , n62652 );
buf ( n62762 , n55201 );
and ( n62763 , n62761 , n62762 );
nor ( n62764 , n62760 , n62763 );
buf ( n62765 , n62764 );
buf ( n62766 , n62765 );
not ( n62767 , n62766 );
buf ( n62768 , n62767 );
buf ( n62769 , n62768 );
buf ( n62770 , n55180 );
and ( n62771 , n62769 , n62770 );
buf ( n62772 , n62708 );
not ( n62773 , n62772 );
buf ( n62774 , n62773 );
buf ( n62775 , n62774 );
buf ( n62776 , n56670 );
and ( n62777 , n62775 , n62776 );
nor ( n62778 , n62771 , n62777 );
buf ( n62779 , n62778 );
buf ( n62780 , n62779 );
nand ( n62781 , n62639 , n54574 );
xnor ( n62782 , n55068 , n62781 );
buf ( n62783 , n62782 );
buf ( n62784 , n55132 );
and ( n62785 , n62783 , n62784 );
buf ( n62786 , n62643 );
buf ( n62787 , n55156 );
and ( n62788 , n62786 , n62787 );
nor ( n62789 , n62785 , n62788 );
buf ( n62790 , n62789 );
buf ( n62791 , n62790 );
nand ( n62792 , n62780 , n62791 );
buf ( n62793 , n62792 );
buf ( n62794 , n62793 );
xor ( n62795 , n62757 , n62794 );
buf ( n62796 , n56582 );
buf ( n62797 , n58897 );
and ( n62798 , n62796 , n62797 );
buf ( n62799 , n56585 );
buf ( n62800 , n58894 );
and ( n62801 , n62799 , n62800 );
nor ( n62802 , n62798 , n62801 );
buf ( n62803 , n62802 );
buf ( n62804 , n62803 );
buf ( n62805 , n58913 );
or ( n62806 , n62804 , n62805 );
buf ( n62807 , n60251 );
buf ( n62808 , n58890 );
or ( n62809 , n62807 , n62808 );
nand ( n62810 , n62806 , n62809 );
buf ( n62811 , n62810 );
buf ( n62812 , n62811 );
and ( n62813 , n62795 , n62812 );
and ( n62814 , n62757 , n62794 );
or ( n62815 , n62813 , n62814 );
buf ( n62816 , n62815 );
xor ( n62817 , n60259 , n60275 );
xor ( n62818 , n62817 , n60292 );
and ( n62819 , n62816 , n62818 );
buf ( n62820 , n56631 );
buf ( n62821 , n58858 );
and ( n62822 , n62820 , n62821 );
not ( n62823 , n62820 );
buf ( n62824 , n58857 );
and ( n62825 , n62823 , n62824 );
nor ( n62826 , n62822 , n62825 );
buf ( n62827 , n62826 );
buf ( n62828 , n62827 );
buf ( n62829 , n56626 );
or ( n62830 , n62828 , n62829 );
buf ( n62831 , n62625 );
buf ( n62832 , n56639 );
or ( n62833 , n62831 , n62832 );
nand ( n62834 , n62830 , n62833 );
buf ( n62835 , n62834 );
buf ( n62836 , n62835 );
buf ( n62837 , n58747 );
buf ( n62838 , n58721 );
and ( n62839 , n62837 , n62838 );
buf ( n62840 , n58841 );
buf ( n62841 , n58718 );
and ( n62842 , n62840 , n62841 );
nor ( n62843 , n62839 , n62842 );
buf ( n62844 , n62843 );
buf ( n62845 , n62844 );
buf ( n62846 , n56799 );
or ( n62847 , n62845 , n62846 );
buf ( n62848 , n60284 );
buf ( n62849 , n58982 );
or ( n62850 , n62848 , n62849 );
nand ( n62851 , n62847 , n62850 );
buf ( n62852 , n62851 );
buf ( n62853 , n62852 );
xor ( n62854 , n62836 , n62853 );
xor ( n62855 , n62658 , n62699 );
xor ( n62856 , n62855 , n62717 );
buf ( n62857 , n62856 );
buf ( n62858 , n62857 );
and ( n62859 , n62854 , n62858 );
and ( n62860 , n62836 , n62853 );
or ( n62861 , n62859 , n62860 );
buf ( n62862 , n62861 );
xor ( n62863 , n60259 , n60275 );
xor ( n62864 , n62863 , n60292 );
and ( n62865 , n62862 , n62864 );
and ( n62866 , n62816 , n62862 );
or ( n62867 , n62819 , n62865 , n62866 );
xor ( n62868 , n62726 , n62729 );
xor ( n62869 , n62868 , n62734 );
and ( n62870 , n62867 , n62869 );
buf ( n62871 , n56720 );
buf ( n62872 , n58897 );
and ( n62873 , n62871 , n62872 );
buf ( n62874 , n58792 );
buf ( n62875 , n58894 );
and ( n62876 , n62874 , n62875 );
nor ( n62877 , n62873 , n62876 );
buf ( n62878 , n62877 );
buf ( n62879 , n62878 );
buf ( n62880 , n58913 );
or ( n62881 , n62879 , n62880 );
buf ( n62882 , n62803 );
buf ( n62883 , n58890 );
or ( n62884 , n62882 , n62883 );
nand ( n62885 , n62881 , n62884 );
buf ( n62886 , n62885 );
buf ( n62887 , n55249 );
buf ( n62888 , n60261 );
and ( n62889 , n62887 , n62888 );
buf ( n62890 , n56594 );
buf ( n62891 , n60090 );
and ( n62892 , n62890 , n62891 );
nor ( n62893 , n62889 , n62892 );
buf ( n62894 , n62893 );
buf ( n62895 , n62894 );
buf ( n62896 , n60270 );
or ( n62897 , n62895 , n62896 );
buf ( n62898 , n62748 );
buf ( n62899 , n60100 );
or ( n62900 , n62898 , n62899 );
nand ( n62901 , n62897 , n62900 );
buf ( n62902 , n62901 );
xor ( n62903 , n62886 , n62902 );
buf ( n62904 , n58823 );
buf ( n62905 , n58721 );
and ( n62906 , n62904 , n62905 );
buf ( n62907 , n58862 );
buf ( n62908 , n58718 );
and ( n62909 , n62907 , n62908 );
nor ( n62910 , n62906 , n62909 );
buf ( n62911 , n62910 );
buf ( n62912 , n62911 );
buf ( n62913 , n56799 );
or ( n62914 , n62912 , n62913 );
buf ( n62915 , n62844 );
buf ( n62916 , n58982 );
or ( n62917 , n62915 , n62916 );
nand ( n62918 , n62914 , n62917 );
buf ( n62919 , n62918 );
and ( n62920 , n62903 , n62919 );
and ( n62921 , n62886 , n62902 );
or ( n62922 , n62920 , n62921 );
buf ( n62923 , n62922 );
buf ( n62924 , n55152 );
buf ( n62925 , n62681 );
and ( n62926 , n62924 , n62925 );
buf ( n62927 , n55205 );
buf ( n62928 , n62663 );
and ( n62929 , n62927 , n62928 );
nor ( n62930 , n62926 , n62929 );
buf ( n62931 , n62930 );
buf ( n62932 , n62931 );
buf ( n62933 , n62679 );
not ( n62934 , n62933 );
buf ( n62935 , n62934 );
buf ( n62936 , n62935 );
or ( n62937 , n62932 , n62936 );
buf ( n62938 , n62695 );
nand ( n62939 , n62937 , n62938 );
buf ( n62940 , n62939 );
buf ( n62941 , n62940 );
buf ( n62942 , n59009 );
buf ( n62943 , n56641 );
and ( n62944 , n62942 , n62943 );
buf ( n62945 , n60077 );
buf ( n62946 , n56631 );
and ( n62947 , n62945 , n62946 );
nor ( n62948 , n62944 , n62947 );
buf ( n62949 , n62948 );
buf ( n62950 , n62949 );
buf ( n62951 , n56626 );
or ( n62952 , n62950 , n62951 );
buf ( n62953 , n62827 );
buf ( n62954 , n56639 );
or ( n62955 , n62953 , n62954 );
nand ( n62956 , n62952 , n62955 );
buf ( n62957 , n62956 );
buf ( n62958 , n62957 );
xor ( n62959 , n62941 , n62958 );
not ( n62960 , n55066 );
nand ( n62961 , n62960 , n54733 );
not ( n62962 , n62961 );
nand ( n62963 , n55056 , n54711 );
not ( n62964 , n54726 );
or ( n62965 , n62963 , n62964 );
not ( n62966 , n55064 );
nand ( n62967 , n62965 , n62966 );
not ( n62968 , n62967 );
or ( n62969 , n62962 , n62968 );
or ( n62970 , n62961 , n62967 );
nand ( n62971 , n62969 , n62970 );
buf ( n62972 , n62971 );
not ( n62973 , n62972 );
buf ( n62974 , n62973 );
buf ( n62975 , n62974 );
buf ( n62976 , n56589 );
or ( n62977 , n62975 , n62976 );
buf ( n62978 , n62782 );
not ( n62979 , n62978 );
buf ( n62980 , n62979 );
buf ( n62981 , n62980 );
buf ( n62982 , n56598 );
or ( n62983 , n62981 , n62982 );
nand ( n62984 , n62977 , n62983 );
buf ( n62985 , n62984 );
buf ( n62986 , n62985 );
buf ( n62987 , n62668 );
buf ( n62988 , n6932 );
not ( n62989 , n62988 );
buf ( n62990 , n62989 );
buf ( n62991 , n62990 );
and ( n62992 , n62987 , n62991 );
not ( n62993 , n62987 );
buf ( n62994 , n6932 );
and ( n62995 , n62993 , n62994 );
nor ( n62996 , n62992 , n62995 );
buf ( n62997 , n62996 );
buf ( n62998 , n62997 );
not ( n62999 , n1854 );
not ( n63000 , n62999 );
nand ( n63001 , n62990 , n63000 );
buf ( n63002 , n63001 );
buf ( n63003 , n62999 );
buf ( n63004 , n63003 );
buf ( n63005 , n6932 );
nand ( n63006 , n63004 , n63005 );
buf ( n63007 , n63006 );
buf ( n63008 , n63007 );
and ( n63009 , n63002 , n63008 );
buf ( n63010 , n63009 );
buf ( n63011 , n63010 );
and ( n63012 , n62998 , n63011 );
buf ( n63013 , n63012 );
buf ( n63014 , n63013 );
not ( n63015 , n62668 );
buf ( n63016 , n63015 );
nand ( n63017 , n63014 , n63016 );
buf ( n63018 , n63017 );
buf ( n63019 , n63018 );
buf ( n63020 , n63010 );
not ( n63021 , n63020 );
buf ( n63022 , n63021 );
buf ( n63023 , n63022 );
buf ( n63024 , n63015 );
nand ( n63025 , n63023 , n63024 );
buf ( n63026 , n63025 );
buf ( n63027 , n63026 );
and ( n63028 , n63019 , n63027 );
buf ( n63029 , n63028 );
buf ( n63030 , n63029 );
xor ( n63031 , n62986 , n63030 );
buf ( n63032 , n62643 );
buf ( n63033 , n56652 );
and ( n63034 , n63032 , n63033 );
buf ( n63035 , n62646 );
buf ( n63036 , n55201 );
and ( n63037 , n63035 , n63036 );
nor ( n63038 , n63034 , n63037 );
buf ( n63039 , n63038 );
buf ( n63040 , n63039 );
buf ( n63041 , n56664 );
or ( n63042 , n63040 , n63041 );
buf ( n63043 , n62765 );
buf ( n63044 , n56673 );
or ( n63045 , n63043 , n63044 );
nand ( n63046 , n63042 , n63045 );
buf ( n63047 , n63046 );
buf ( n63048 , n63047 );
and ( n63049 , n63031 , n63048 );
and ( n63050 , n62986 , n63030 );
or ( n63051 , n63049 , n63050 );
buf ( n63052 , n63051 );
buf ( n63053 , n63052 );
and ( n63054 , n62959 , n63053 );
and ( n63055 , n62941 , n62958 );
or ( n63056 , n63054 , n63055 );
buf ( n63057 , n63056 );
buf ( n63058 , n63057 );
xor ( n63059 , n62923 , n63058 );
xor ( n63060 , n62757 , n62794 );
xor ( n63061 , n63060 , n62812 );
buf ( n63062 , n63061 );
buf ( n63063 , n63062 );
and ( n63064 , n63059 , n63063 );
and ( n63065 , n62923 , n63058 );
or ( n63066 , n63064 , n63065 );
buf ( n63067 , n63066 );
xor ( n63068 , n62617 , n62634 );
xor ( n63069 , n63068 , n62722 );
buf ( n63070 , n63069 );
xor ( n63071 , n63067 , n63070 );
xor ( n63072 , n60259 , n60275 );
xor ( n63073 , n63072 , n60292 );
xor ( n63074 , n62816 , n62862 );
xor ( n63075 , n63073 , n63074 );
and ( n63076 , n63071 , n63075 );
and ( n63077 , n63067 , n63070 );
or ( n63078 , n63076 , n63077 );
xor ( n63079 , n62726 , n62729 );
xor ( n63080 , n63079 , n62734 );
and ( n63081 , n63078 , n63080 );
and ( n63082 , n62867 , n63078 );
or ( n63083 , n62870 , n63081 , n63082 );
xor ( n63084 , n60300 , n60303 );
xor ( n63085 , n63084 , n60307 );
and ( n63086 , n63083 , n63085 );
and ( n63087 , n62737 , n63083 );
or ( n63088 , n62740 , n63086 , n63087 );
buf ( n63089 , n63088 );
nand ( n63090 , n62610 , n63089 );
buf ( n63091 , n63090 );
buf ( n63092 , n63091 );
buf ( n63093 , n62608 );
buf ( n63094 , n62577 );
nand ( n63095 , n63093 , n63094 );
buf ( n63096 , n63095 );
buf ( n63097 , n63096 );
nand ( n63098 , n63092 , n63097 );
buf ( n63099 , n63098 );
buf ( n63100 , n63099 );
xor ( n63101 , n62573 , n63100 );
xor ( n63102 , n61426 , n61474 );
xnor ( n63103 , n63102 , n61458 );
buf ( n63104 , n63103 );
and ( n63105 , n63101 , n63104 );
and ( n63106 , n62573 , n63100 );
or ( n63107 , n63105 , n63106 );
buf ( n63108 , n63107 );
buf ( n63109 , n63108 );
nand ( n63110 , n62556 , n63109 );
buf ( n63111 , n63110 );
buf ( n63112 , n63111 );
buf ( n63113 , n62550 );
buf ( n63114 , n62524 );
not ( n63115 , n63114 );
buf ( n63116 , n63115 );
buf ( n63117 , n63116 );
nand ( n63118 , n63113 , n63117 );
buf ( n63119 , n63118 );
buf ( n63120 , n63119 );
nand ( n63121 , n63112 , n63120 );
buf ( n63122 , n63121 );
buf ( n63123 , n63122 );
buf ( n63124 , n44517 );
not ( n63125 , n63124 );
buf ( n63126 , n44533 );
not ( n63127 , n63126 );
buf ( n63128 , n43311 );
not ( n63129 , n63128 );
or ( n63130 , n63127 , n63129 );
buf ( n63131 , n38848 );
buf ( n63132 , n44530 );
nand ( n63133 , n63131 , n63132 );
buf ( n63134 , n63133 );
buf ( n63135 , n63134 );
nand ( n63136 , n63130 , n63135 );
buf ( n63137 , n63136 );
buf ( n63138 , n63137 );
not ( n63139 , n63138 );
or ( n63140 , n63125 , n63139 );
buf ( n63141 , n61890 );
buf ( n63142 , n44496 );
nand ( n63143 , n63141 , n63142 );
buf ( n63144 , n63143 );
buf ( n63145 , n63144 );
nand ( n63146 , n63140 , n63145 );
buf ( n63147 , n63146 );
buf ( n63148 , n63147 );
xor ( n63149 , n63123 , n63148 );
buf ( n63150 , n61977 );
buf ( n63151 , n42315 );
and ( n63152 , n63150 , n63151 );
buf ( n63153 , n59242 );
not ( n63154 , n63153 );
buf ( n63155 , n29325 );
not ( n63156 , n63155 );
or ( n63157 , n63154 , n63156 );
buf ( n63158 , n29328 );
buf ( n63159 , n42260 );
nand ( n63160 , n63158 , n63159 );
buf ( n63161 , n63160 );
buf ( n63162 , n63161 );
nand ( n63163 , n63157 , n63162 );
buf ( n63164 , n63163 );
buf ( n63165 , n63164 );
not ( n63166 , n63165 );
buf ( n63167 , n42249 );
nor ( n63168 , n63166 , n63167 );
buf ( n63169 , n63168 );
buf ( n63170 , n63169 );
nor ( n63171 , n63152 , n63170 );
buf ( n63172 , n63171 );
buf ( n63173 , n63172 );
not ( n63174 , n63173 );
buf ( n63175 , n44039 );
not ( n63176 , n63175 );
buf ( n63177 , n47068 );
not ( n63178 , n63177 );
buf ( n63179 , n46126 );
not ( n63180 , n63179 );
and ( n63181 , n63178 , n63180 );
buf ( n63182 , n46623 );
buf ( n63183 , n46126 );
and ( n63184 , n63182 , n63183 );
nor ( n63185 , n63181 , n63184 );
buf ( n63186 , n63185 );
buf ( n63187 , n63186 );
not ( n63188 , n63187 );
and ( n63189 , n63176 , n63188 );
buf ( n63190 , n61494 );
buf ( n63191 , n52171 );
nor ( n63192 , n63190 , n63191 );
buf ( n63193 , n63192 );
buf ( n63194 , n63193 );
nor ( n63195 , n63189 , n63194 );
buf ( n63196 , n63195 );
buf ( n63197 , n63196 );
not ( n63198 , n63197 );
or ( n63199 , n63174 , n63198 );
buf ( n63200 , n41993 );
not ( n63201 , n63200 );
buf ( n63202 , n52670 );
not ( n63203 , n63202 );
or ( n63204 , n63201 , n63203 );
buf ( n63205 , n25159 );
buf ( n63206 , n43966 );
nand ( n63207 , n63205 , n63206 );
buf ( n63208 , n63207 );
buf ( n63209 , n63208 );
nand ( n63210 , n63204 , n63209 );
buf ( n63211 , n63210 );
buf ( n63212 , n63211 );
not ( n63213 , n63212 );
buf ( n63214 , n50128 );
not ( n63215 , n63214 );
or ( n63216 , n63213 , n63215 );
buf ( n63217 , n61949 );
buf ( n63218 , n56567 );
nand ( n63219 , n63217 , n63218 );
buf ( n63220 , n63219 );
buf ( n63221 , n63220 );
nand ( n63222 , n63216 , n63221 );
buf ( n63223 , n63222 );
buf ( n63224 , n63223 );
not ( n63225 , n63224 );
buf ( n63226 , n42865 );
not ( n63227 , n63226 );
buf ( n63228 , n46073 );
not ( n63229 , n63228 );
or ( n63230 , n63227 , n63229 );
buf ( n63231 , n24092 );
buf ( n63232 , n42862 );
nand ( n63233 , n63231 , n63232 );
buf ( n63234 , n63233 );
buf ( n63235 , n63234 );
nand ( n63236 , n63230 , n63235 );
buf ( n63237 , n63236 );
buf ( n63238 , n63237 );
not ( n63239 , n63238 );
buf ( n63240 , n52537 );
not ( n63241 , n63240 );
or ( n63242 , n63239 , n63241 );
buf ( n63243 , n61379 );
buf ( n63244 , n48975 );
nand ( n63245 , n63243 , n63244 );
buf ( n63246 , n63245 );
buf ( n63247 , n63246 );
nand ( n63248 , n63242 , n63247 );
buf ( n63249 , n63248 );
buf ( n63250 , n63249 );
not ( n63251 , n63250 );
or ( n63252 , n63225 , n63251 );
buf ( n63253 , n63249 );
buf ( n63254 , n63223 );
or ( n63255 , n63253 , n63254 );
buf ( n63256 , n58249 );
not ( n63257 , n63256 );
buf ( n63258 , n25226 );
not ( n63259 , n63258 );
buf ( n63260 , n46657 );
not ( n63261 , n63260 );
or ( n63262 , n63259 , n63261 );
buf ( n63263 , n42149 );
buf ( n63264 , n62510 );
nand ( n63265 , n63263 , n63264 );
buf ( n63266 , n63265 );
buf ( n63267 , n63266 );
nand ( n63268 , n63262 , n63267 );
buf ( n63269 , n63268 );
buf ( n63270 , n63269 );
not ( n63271 , n63270 );
or ( n63272 , n63257 , n63271 );
buf ( n63273 , n42668 );
buf ( n63274 , n62516 );
nand ( n63275 , n63273 , n63274 );
buf ( n63276 , n63275 );
buf ( n63277 , n63276 );
nand ( n63278 , n63272 , n63277 );
buf ( n63279 , n63278 );
buf ( n63280 , n63279 );
nand ( n63281 , n63255 , n63280 );
buf ( n63282 , n63281 );
buf ( n63283 , n63282 );
nand ( n63284 , n63252 , n63283 );
buf ( n63285 , n63284 );
buf ( n63286 , n63285 );
nand ( n63287 , n63199 , n63286 );
buf ( n63288 , n63287 );
buf ( n63289 , n63288 );
or ( n63290 , n63196 , n63172 );
buf ( n63291 , n63290 );
nand ( n63292 , n63289 , n63291 );
buf ( n63293 , n63292 );
buf ( n63294 , n63293 );
and ( n63295 , n63149 , n63294 );
and ( n63296 , n63123 , n63148 );
or ( n63297 , n63295 , n63296 );
buf ( n63298 , n63297 );
buf ( n63299 , n63298 );
xor ( n63300 , n61324 , n61341 );
xor ( n63301 , n63300 , n61505 );
buf ( n63302 , n63301 );
buf ( n63303 , n63302 );
xor ( n63304 , n63299 , n63303 );
xor ( n63305 , n61367 , n61484 );
xor ( n63306 , n63305 , n61500 );
buf ( n63307 , n63306 );
buf ( n63308 , n63307 );
xor ( n63309 , n61937 , n61962 );
xor ( n63310 , n63309 , n61967 );
buf ( n63311 , n63310 );
buf ( n63312 , n63311 );
xor ( n63313 , n61477 , n61391 );
xor ( n63314 , n63313 , n61417 );
buf ( n63315 , n63314 );
xor ( n63316 , n63312 , n63315 );
buf ( n63317 , n47716 );
not ( n63318 , n63317 );
buf ( n63319 , n41805 );
not ( n63320 , n63319 );
or ( n63321 , n63318 , n63320 );
buf ( n63322 , n53861 );
buf ( n63323 , n47725 );
nand ( n63324 , n63322 , n63323 );
buf ( n63325 , n63324 );
buf ( n63326 , n63325 );
nand ( n63327 , n63321 , n63326 );
buf ( n63328 , n63327 );
buf ( n63329 , n63328 );
not ( n63330 , n63329 );
buf ( n63331 , n37397 );
not ( n63332 , n63331 );
or ( n63333 , n63330 , n63332 );
buf ( n63334 , n61749 );
not ( n63335 , n63334 );
buf ( n63336 , n42135 );
nand ( n63337 , n63335 , n63336 );
buf ( n63338 , n63337 );
buf ( n63339 , n63338 );
nand ( n63340 , n63333 , n63339 );
buf ( n63341 , n63340 );
buf ( n63342 , n63341 );
and ( n63343 , n63316 , n63342 );
and ( n63344 , n63312 , n63315 );
or ( n63345 , n63343 , n63344 );
buf ( n63346 , n63345 );
buf ( n63347 , n63346 );
xor ( n63348 , n63308 , n63347 );
xor ( n63349 , n61972 , n61985 );
xor ( n63350 , n63349 , n61991 );
buf ( n63351 , n63350 );
buf ( n63352 , n63351 );
and ( n63353 , n63348 , n63352 );
and ( n63354 , n63308 , n63347 );
or ( n63355 , n63353 , n63354 );
buf ( n63356 , n63355 );
buf ( n63357 , n63356 );
and ( n63358 , n63304 , n63357 );
and ( n63359 , n63299 , n63303 );
or ( n63360 , n63358 , n63359 );
buf ( n63361 , n63360 );
buf ( n63362 , n63361 );
nand ( n63363 , n62500 , n63362 );
buf ( n63364 , n63363 );
nand ( n63365 , C1 , n63364 );
and ( n63366 , n62493 , n63365 );
and ( n63367 , n62355 , n62492 );
or ( n63368 , n63366 , n63367 );
buf ( n63369 , n63368 );
not ( n63370 , n63369 );
buf ( n63371 , n60575 );
buf ( n63372 , n60598 );
and ( n63373 , n63371 , n63372 );
not ( n63374 , n63371 );
buf ( n63375 , n60609 );
and ( n63376 , n63374 , n63375 );
nor ( n63377 , n63373 , n63376 );
buf ( n63378 , n63377 );
and ( n63379 , n63378 , n60602 );
not ( n63380 , n63378 );
not ( n63381 , n60602 );
and ( n63382 , n63380 , n63381 );
nor ( n63383 , n63379 , n63382 );
buf ( n63384 , n63383 );
xor ( n63385 , n60858 , n60861 );
xor ( n63386 , n63385 , n60903 );
buf ( n63387 , n63386 );
buf ( n63388 , n63387 );
xor ( n63389 , n63384 , n63388 );
buf ( n63390 , n48855 );
not ( n63391 , n63390 );
buf ( n63392 , n62149 );
not ( n63393 , n63392 );
or ( n63394 , n63391 , n63393 );
nand ( n63395 , n60851 , n48868 );
buf ( n63396 , n63395 );
nand ( n63397 , n63394 , n63396 );
buf ( n63398 , n63397 );
buf ( n63399 , n63398 );
not ( n63400 , n60934 );
xor ( n63401 , n60935 , n63400 );
xnor ( n63402 , n63401 , n61033 );
buf ( n63403 , n63402 );
xor ( n63404 , n63399 , n63403 );
buf ( n63405 , n61080 );
not ( n63406 , n63405 );
buf ( n63407 , n61111 );
not ( n63408 , n63407 );
or ( n63409 , n63406 , n63408 );
buf ( n63410 , n61100 );
buf ( n63411 , n61106 );
nand ( n63412 , n63410 , n63411 );
buf ( n63413 , n63412 );
buf ( n63414 , n63413 );
nand ( n63415 , n63409 , n63414 );
buf ( n63416 , n63415 );
buf ( n63417 , n63416 );
buf ( n63418 , n61184 );
and ( n63419 , n63417 , n63418 );
not ( n63420 , n63417 );
buf ( n63421 , n61184 );
not ( n63422 , n63421 );
buf ( n63423 , n63422 );
buf ( n63424 , n63423 );
and ( n63425 , n63420 , n63424 );
nor ( n63426 , n63419 , n63425 );
buf ( n63427 , n63426 );
buf ( n63428 , n63427 );
and ( n63429 , n63404 , n63428 );
and ( n63430 , n63399 , n63403 );
or ( n63431 , n63429 , n63430 );
buf ( n63432 , n63431 );
buf ( n63433 , n63432 );
and ( n63434 , n63389 , n63433 );
and ( n63435 , n63384 , n63388 );
or ( n63436 , n63434 , n63435 );
buf ( n63437 , n63436 );
buf ( n63438 , n63437 );
not ( n63439 , n63438 );
and ( n63440 , n61564 , n61577 );
not ( n63441 , n61564 );
and ( n63442 , n63441 , n61578 );
nor ( n63443 , n63440 , n63442 );
and ( n63444 , n63443 , n61582 );
not ( n63445 , n63443 );
not ( n63446 , n61582 );
and ( n63447 , n63445 , n63446 );
nor ( n63448 , n63444 , n63447 );
buf ( n63449 , n63448 );
not ( n63450 , n63449 );
buf ( n63451 , n63450 );
buf ( n63452 , n63451 );
nand ( n63453 , n63439 , n63452 );
buf ( n63454 , n63453 );
buf ( n63455 , n63454 );
not ( n63456 , n63455 );
or ( n63457 , n63370 , n63456 );
buf ( n63458 , n63437 );
buf ( n63459 , n63448 );
nand ( n63460 , n63458 , n63459 );
buf ( n63461 , n63460 );
buf ( n63462 , n63461 );
nand ( n63463 , n63457 , n63462 );
buf ( n63464 , n63463 );
buf ( n63465 , n63464 );
nand ( n63466 , n62353 , n63465 );
buf ( n63467 , n63466 );
nand ( n63468 , n62349 , n62106 );
nand ( n63469 , n63467 , n63468 );
nand ( n63470 , n62104 , n63469 );
nand ( n63471 , n62098 , n63470 );
not ( n63472 , n63471 );
nand ( n63473 , n62055 , n63472 );
buf ( n63474 , n63473 );
and ( n63475 , n62049 , n63474 );
buf ( n63476 , n63475 );
xor ( n63477 , n57434 , n57894 );
xnor ( n63478 , n63477 , n57899 );
buf ( n63479 , n63478 );
xor ( n63480 , n60491 , n60494 );
and ( n63481 , n63480 , n61206 );
and ( n63482 , n60491 , n60494 );
or ( n63483 , n63481 , n63482 );
buf ( n63484 , n63483 );
xor ( n63485 , n63479 , n63484 );
xor ( n63486 , n58396 , n58400 );
xor ( n63487 , n63486 , n59098 );
buf ( n63488 , n63487 );
buf ( n63489 , n63488 );
xor ( n63490 , n63485 , n63489 );
buf ( n63491 , n63490 );
buf ( n63492 , n63491 );
not ( n63493 , n63492 );
buf ( n63494 , n63493 );
xor ( n63495 , n59147 , n60485 );
and ( n63496 , n63495 , n61207 );
and ( n63497 , n59147 , n60485 );
or ( n63498 , n63496 , n63497 );
buf ( n63499 , n63498 );
not ( n63500 , n63499 );
buf ( n63501 , n63500 );
nand ( n63502 , n63494 , n63501 );
buf ( n63503 , n63502 );
buf ( n63504 , n63503 );
buf ( n63505 , n63504 );
xor ( n63506 , n59107 , n59102 );
xnor ( n63507 , n63506 , n59117 );
buf ( n63508 , n63507 );
not ( n63509 , n63508 );
buf ( n63510 , n63509 );
buf ( n63511 , n63510 );
xor ( n63512 , n63479 , n63484 );
and ( n63513 , n63512 , n63489 );
and ( n63514 , n63479 , n63484 );
or ( n63515 , n63513 , n63514 );
buf ( n63516 , n63515 );
buf ( n63517 , n63516 );
not ( n63518 , n63517 );
buf ( n63519 , n63518 );
buf ( n63520 , n63519 );
nand ( n63521 , n63511 , n63520 );
buf ( n63522 , n63521 );
and ( n63523 , n63476 , n63505 , n63522 );
xor ( n63524 , n63399 , n63403 );
xor ( n63525 , n63524 , n63428 );
buf ( n63526 , n63525 );
xor ( n63527 , n61898 , n61923 );
xor ( n63528 , n63527 , n61996 );
buf ( n63529 , n63528 );
not ( n63530 , n63529 );
xor ( n63531 , n61736 , n61800 );
xor ( n63532 , n63531 , n61826 );
buf ( n63533 , n63532 );
not ( n63534 , n63533 );
or ( n63535 , n63530 , n63534 );
buf ( n63536 , n63529 );
buf ( n63537 , n63533 );
or ( n63538 , n63536 , n63537 );
buf ( n63539 , n61796 );
buf ( n63540 , n61780 );
xor ( n63541 , n63539 , n63540 );
buf ( n63542 , n61763 );
xor ( n63543 , n63541 , n63542 );
buf ( n63544 , n63543 );
buf ( n63545 , n63544 );
buf ( n63546 , n47331 );
not ( n63547 , n63546 );
buf ( n63548 , n46875 );
not ( n63549 , n63548 );
buf ( n63550 , n42973 );
not ( n63551 , n63550 );
or ( n63552 , n63549 , n63551 );
buf ( n63553 , n38480 );
buf ( n63554 , n46890 );
nand ( n63555 , n63553 , n63554 );
buf ( n63556 , n63555 );
buf ( n63557 , n63556 );
nand ( n63558 , n63552 , n63557 );
buf ( n63559 , n63558 );
buf ( n63560 , n63559 );
not ( n63561 , n63560 );
or ( n63562 , n63547 , n63561 );
buf ( n63563 , n62366 );
not ( n63564 , n63563 );
buf ( n63565 , n46912 );
nand ( n63566 , n63564 , n63565 );
buf ( n63567 , n63566 );
buf ( n63568 , n63567 );
nand ( n63569 , n63562 , n63568 );
buf ( n63570 , n63569 );
buf ( n63571 , n63570 );
xor ( n63572 , n63545 , n63571 );
buf ( n63573 , n61776 );
not ( n63574 , n63573 );
buf ( n63575 , n43868 );
not ( n63576 , n63575 );
or ( n63577 , n63574 , n63576 );
buf ( n63578 , n41608 );
not ( n63579 , n63578 );
buf ( n63580 , n41781 );
not ( n63581 , n63580 );
or ( n63582 , n63579 , n63581 );
buf ( n63583 , n41762 );
buf ( n63584 , n41604 );
nand ( n63585 , n63583 , n63584 );
buf ( n63586 , n63585 );
buf ( n63587 , n63586 );
nand ( n63588 , n63582 , n63587 );
buf ( n63589 , n63588 );
buf ( n63590 , n63589 );
buf ( n63591 , n44267 );
nand ( n63592 , n63590 , n63591 );
buf ( n63593 , n63592 );
buf ( n63594 , n63593 );
nand ( n63595 , n63577 , n63594 );
buf ( n63596 , n63595 );
not ( n63597 , n63596 );
buf ( n63598 , n63597 );
not ( n63599 , n63598 );
buf ( n63600 , n37514 );
not ( n63601 , n63600 );
buf ( n63602 , n41843 );
not ( n63603 , n63602 );
buf ( n63604 , n50067 );
not ( n63605 , n63604 );
and ( n63606 , n63603 , n63605 );
buf ( n63607 , n41844 );
buf ( n63608 , n50067 );
and ( n63609 , n63607 , n63608 );
nor ( n63610 , n63606 , n63609 );
buf ( n63611 , n63610 );
buf ( n63612 , n63611 );
not ( n63613 , n63612 );
and ( n63614 , n63601 , n63613 );
buf ( n63615 , n62403 );
buf ( n63616 , n37449 );
nor ( n63617 , n63615 , n63616 );
buf ( n63618 , n63617 );
buf ( n63619 , n63618 );
nor ( n63620 , n63614 , n63619 );
buf ( n63621 , n63620 );
buf ( n63622 , n63621 );
not ( n63623 , n63622 );
or ( n63624 , n63599 , n63623 );
buf ( n63625 , n42008 );
not ( n63626 , n63625 );
buf ( n63627 , n52725 );
not ( n63628 , n63627 );
or ( n63629 , n63626 , n63628 );
buf ( n63630 , n25180 );
buf ( n63631 , n42008 );
not ( n63632 , n63631 );
buf ( n63633 , n63632 );
buf ( n63634 , n63633 );
nand ( n63635 , n63630 , n63634 );
buf ( n63636 , n63635 );
buf ( n63637 , n63636 );
nand ( n63638 , n63629 , n63637 );
buf ( n63639 , n63638 );
buf ( n63640 , n63639 );
not ( n63641 , n63640 );
buf ( n63642 , n53628 );
not ( n63643 , n63642 );
or ( n63644 , n63641 , n63643 );
buf ( n63645 , n61466 );
buf ( n63646 , n53649 );
nand ( n63647 , n63645 , n63646 );
buf ( n63648 , n63647 );
buf ( n63649 , n63648 );
nand ( n63650 , n63644 , n63649 );
buf ( n63651 , n63650 );
buf ( n63652 , n63651 );
buf ( n63653 , n42336 );
not ( n63654 , n63653 );
buf ( n63655 , n62565 );
not ( n63656 , n63655 );
or ( n63657 , n63654 , n63656 );
and ( n63658 , n29754 , n46855 );
not ( n63659 , n29754 );
and ( n63660 , n63659 , n42343 );
or ( n63661 , n63658 , n63660 );
buf ( n63662 , n63661 );
buf ( n63663 , n42378 );
nand ( n63664 , n63662 , n63663 );
buf ( n63665 , n63664 );
buf ( n63666 , n63665 );
nand ( n63667 , n63657 , n63666 );
buf ( n63668 , n63667 );
buf ( n63669 , n63668 );
xor ( n63670 , n63652 , n63669 );
buf ( n63671 , n63088 );
buf ( n63672 , n62577 );
xnor ( n63673 , n63671 , n63672 );
buf ( n63674 , n63673 );
buf ( n63675 , n63674 );
not ( n63676 , n63675 );
buf ( n63677 , n62608 );
not ( n63678 , n63677 );
or ( n63679 , n63676 , n63678 );
buf ( n63680 , n62608 );
buf ( n63681 , n63674 );
or ( n63682 , n63680 , n63681 );
nand ( n63683 , n63679 , n63682 );
buf ( n63684 , n63683 );
buf ( n63685 , n63684 );
and ( n63686 , n63670 , n63685 );
and ( n63687 , n63652 , n63669 );
or ( n63688 , n63686 , n63687 );
buf ( n63689 , n63688 );
buf ( n63690 , n63689 );
buf ( n63691 , n42315 );
not ( n63692 , n63691 );
buf ( n63693 , n63164 );
not ( n63694 , n63693 );
or ( n63695 , n63692 , n63694 );
buf ( n63696 , n59242 );
not ( n63697 , n63696 );
buf ( n63698 , n41915 );
not ( n63699 , n63698 );
or ( n63700 , n63697 , n63699 );
buf ( n63701 , n41912 );
buf ( n63702 , n42260 );
nand ( n63703 , n63701 , n63702 );
buf ( n63704 , n63703 );
buf ( n63705 , n63704 );
nand ( n63706 , n63700 , n63705 );
buf ( n63707 , n63706 );
buf ( n63708 , n63707 );
buf ( n63709 , n42252 );
nand ( n63710 , n63708 , n63709 );
buf ( n63711 , n63710 );
buf ( n63712 , n63711 );
nand ( n63713 , n63695 , n63712 );
buf ( n63714 , n63713 );
buf ( n63715 , n63714 );
xor ( n63716 , n63690 , n63715 );
buf ( n63717 , n38979 );
not ( n63718 , n63717 );
buf ( n63719 , n44949 );
not ( n63720 , n63719 );
and ( n63721 , n63718 , n63720 );
buf ( n63722 , n38979 );
buf ( n63723 , n44949 );
and ( n63724 , n63722 , n63723 );
nor ( n63725 , n63721 , n63724 );
buf ( n63726 , n63725 );
buf ( n63727 , n63726 );
not ( n63728 , n63727 );
buf ( n63729 , n63728 );
buf ( n63730 , n63729 );
not ( n63731 , n63730 );
buf ( n63732 , n47050 );
not ( n63733 , n63732 );
or ( n63734 , n63731 , n63733 );
buf ( n63735 , n62538 );
buf ( n63736 , n50104 );
nand ( n63737 , n63735 , n63736 );
buf ( n63738 , n63737 );
buf ( n63739 , n63738 );
nand ( n63740 , n63734 , n63739 );
buf ( n63741 , n63740 );
buf ( n63742 , n63741 );
and ( n63743 , n63716 , n63742 );
and ( n63744 , n63690 , n63715 );
or ( n63745 , n63743 , n63744 );
buf ( n63746 , n63745 );
buf ( n63747 , n63746 );
nand ( n63748 , n63624 , n63747 );
buf ( n63749 , n63748 );
buf ( n63750 , n63749 );
buf ( n63751 , n63621 );
not ( n63752 , n63751 );
buf ( n63753 , n63596 );
nand ( n63754 , n63752 , n63753 );
buf ( n63755 , n63754 );
buf ( n63756 , n63755 );
nand ( n63757 , n63750 , n63756 );
buf ( n63758 , n63757 );
buf ( n63759 , n63758 );
and ( n63760 , n63572 , n63759 );
and ( n63761 , n63545 , n63571 );
or ( n63762 , n63760 , n63761 );
buf ( n63763 , n63762 );
buf ( n63764 , n63763 );
nand ( n63765 , n63538 , n63764 );
buf ( n63766 , n63765 );
nand ( n63767 , n63535 , n63766 );
xor ( n63768 , n63526 , n63767 );
xor ( n63769 , n61872 , n61875 );
xor ( n63770 , n63769 , n62000 );
xor ( n63771 , n63768 , n63770 );
buf ( n63772 , n63771 );
xor ( n63773 , n63308 , n63347 );
xor ( n63774 , n63773 , n63352 );
buf ( n63775 , n63774 );
buf ( n63776 , n63775 );
xor ( n63777 , n63312 , n63315 );
xor ( n63778 , n63777 , n63342 );
buf ( n63779 , n63778 );
buf ( n63780 , n63779 );
buf ( n63781 , n12481 );
buf ( n63782 , n39235 );
and ( n63783 , n63781 , n63782 );
not ( n63784 , n63781 );
buf ( n63785 , n36932 );
and ( n63786 , n63784 , n63785 );
nor ( n63787 , n63783 , n63786 );
buf ( n63788 , n63787 );
buf ( n63789 , n63788 );
not ( n63790 , n63789 );
buf ( n63791 , n45423 );
not ( n63792 , n63791 );
or ( n63793 , n63790 , n63792 );
buf ( n63794 , n47409 );
buf ( n63795 , n62260 );
nand ( n63796 , n63794 , n63795 );
buf ( n63797 , n63796 );
buf ( n63798 , n63797 );
nand ( n63799 , n63793 , n63798 );
buf ( n63800 , n63799 );
buf ( n63801 , n63800 );
xor ( n63802 , n63780 , n63801 );
buf ( n63803 , n48323 );
not ( n63804 , n63803 );
buf ( n63805 , n41805 );
not ( n63806 , n63805 );
or ( n63807 , n63804 , n63806 );
buf ( n63808 , n42114 );
buf ( n63809 , n48320 );
nand ( n63810 , n63808 , n63809 );
buf ( n63811 , n63810 );
buf ( n63812 , n63811 );
nand ( n63813 , n63807 , n63812 );
buf ( n63814 , n63813 );
buf ( n63815 , n63814 );
not ( n63816 , n63815 );
buf ( n63817 , n37400 );
not ( n63818 , n63817 );
or ( n63819 , n63816 , n63818 );
buf ( n63820 , n63328 );
buf ( n63821 , n37413 );
nand ( n63822 , n63820 , n63821 );
buf ( n63823 , n63822 );
buf ( n63824 , n63823 );
nand ( n63825 , n63819 , n63824 );
buf ( n63826 , n63825 );
buf ( n63827 , n63826 );
not ( n63828 , n42668 );
not ( n63829 , n63269 );
or ( n63830 , n63828 , n63829 );
not ( n63831 , n42711 );
buf ( n63832 , n43362 );
not ( n63833 , n63832 );
buf ( n63834 , n25226 );
not ( n63835 , n63834 );
or ( n63836 , n63833 , n63835 );
buf ( n63837 , n50624 );
buf ( n63838 , n62510 );
nand ( n63839 , n63837 , n63838 );
buf ( n63840 , n63839 );
buf ( n63841 , n63840 );
nand ( n63842 , n63836 , n63841 );
buf ( n63843 , n63842 );
nand ( n63844 , n63831 , n63843 );
nand ( n63845 , n63830 , n63844 );
not ( n63846 , n63845 );
buf ( n63847 , n63846 );
not ( n63848 , n63847 );
not ( n63849 , n47020 );
not ( n63850 , n63726 );
and ( n63851 , n63849 , n63850 );
buf ( n63852 , n46117 );
not ( n63853 , n63852 );
buf ( n63854 , n42471 );
not ( n63855 , n63854 );
or ( n63856 , n63853 , n63855 );
buf ( n63857 , n38979 );
buf ( n63858 , n46126 );
nand ( n63859 , n63857 , n63858 );
buf ( n63860 , n63859 );
buf ( n63861 , n63860 );
nand ( n63862 , n63856 , n63861 );
buf ( n63863 , n63862 );
not ( n63864 , n63863 );
nor ( n63865 , n63864 , n45056 );
nor ( n63866 , n63851 , n63865 );
buf ( n63867 , n63866 );
not ( n63868 , n63867 );
or ( n63869 , n63848 , n63868 );
xor ( n63870 , n60300 , n60303 );
xor ( n63871 , n63870 , n60307 );
xor ( n63872 , n62737 , n63083 );
xor ( n63873 , n63871 , n63872 );
buf ( n63874 , n63873 );
buf ( n63875 , n13662 );
buf ( n63876 , n41698 );
and ( n63877 , n63875 , n63876 );
not ( n63878 , n63875 );
buf ( n63879 , n62598 );
and ( n63880 , n63878 , n63879 );
nor ( n63881 , n63877 , n63880 );
buf ( n63882 , n63881 );
buf ( n63883 , n63882 );
not ( n63884 , n63883 );
buf ( n63885 , n61454 );
not ( n63886 , n63885 );
or ( n63887 , n63884 , n63886 );
buf ( n63888 , n62604 );
buf ( n63889 , n48671 );
nand ( n63890 , n63888 , n63889 );
buf ( n63891 , n63890 );
buf ( n63892 , n63891 );
nand ( n63893 , n63887 , n63892 );
buf ( n63894 , n63893 );
buf ( n63895 , n63894 );
xor ( n63896 , n63874 , n63895 );
buf ( n63897 , n42336 );
not ( n63898 , n63897 );
buf ( n63899 , n63661 );
not ( n63900 , n63899 );
or ( n63901 , n63898 , n63900 );
buf ( n63902 , n42343 );
not ( n63903 , n63902 );
buf ( n63904 , n13653 );
not ( n63905 , n63904 );
buf ( n63906 , n63905 );
buf ( n63907 , n63906 );
not ( n63908 , n63907 );
or ( n63909 , n63903 , n63908 );
buf ( n63910 , n13653 );
buf ( n63911 , n24950 );
buf ( n63912 , n63911 );
buf ( n63913 , n63912 );
buf ( n63914 , n63913 );
nand ( n63915 , n63910 , n63914 );
buf ( n63916 , n63915 );
buf ( n63917 , n63916 );
nand ( n63918 , n63909 , n63917 );
buf ( n63919 , n63918 );
nand ( n63920 , n63919 , n42374 );
buf ( n63921 , n63920 );
nand ( n63922 , n63901 , n63921 );
buf ( n63923 , n63922 );
buf ( n63924 , n63923 );
xor ( n63925 , n63896 , n63924 );
buf ( n63926 , n63925 );
not ( n63927 , n63926 );
buf ( n63928 , n41993 );
not ( n63929 , n63928 );
buf ( n63930 , n52725 );
not ( n63931 , n63930 );
or ( n63932 , n63929 , n63931 );
buf ( n63933 , n42560 );
buf ( n63934 , n43966 );
nand ( n63935 , n63933 , n63934 );
buf ( n63936 , n63935 );
buf ( n63937 , n63936 );
nand ( n63938 , n63932 , n63937 );
buf ( n63939 , n63938 );
buf ( n63940 , n63939 );
not ( n63941 , n63940 );
buf ( n63942 , n43935 );
not ( n63943 , n63942 );
or ( n63944 , n63941 , n63943 );
buf ( n63945 , n63639 );
buf ( n63946 , n53649 );
nand ( n63947 , n63945 , n63946 );
buf ( n63948 , n63947 );
buf ( n63949 , n63948 );
nand ( n63950 , n63944 , n63949 );
buf ( n63951 , n63950 );
buf ( n63952 , n63951 );
not ( n63953 , n63952 );
xor ( n63954 , n62726 , n62729 );
xor ( n63955 , n63954 , n62734 );
xor ( n63956 , n62867 , n63078 );
xor ( n63957 , n63955 , n63956 );
buf ( n63958 , n63957 );
buf ( n63959 , n58857 );
buf ( n63960 , n58721 );
and ( n63961 , n63959 , n63960 );
buf ( n63962 , n58858 );
buf ( n63963 , n58718 );
and ( n63964 , n63962 , n63963 );
nor ( n63965 , n63961 , n63964 );
buf ( n63966 , n63965 );
buf ( n63967 , n63966 );
buf ( n63968 , n56799 );
or ( n63969 , n63967 , n63968 );
buf ( n63970 , n62911 );
buf ( n63971 , n58982 );
or ( n63972 , n63970 , n63971 );
nand ( n63973 , n63969 , n63972 );
buf ( n63974 , n63973 );
buf ( n63975 , n55113 );
buf ( n63976 , n62681 );
and ( n63977 , n63975 , n63976 );
buf ( n63978 , n56655 );
buf ( n63979 , n62663 );
and ( n63980 , n63978 , n63979 );
nor ( n63981 , n63977 , n63980 );
buf ( n63982 , n63981 );
buf ( n63983 , n63982 );
buf ( n63984 , n62935 );
or ( n63985 , n63983 , n63984 );
buf ( n63986 , n62931 );
buf ( n63987 , n62676 );
or ( n63988 , n63986 , n63987 );
nand ( n63989 , n63985 , n63988 );
buf ( n63990 , n63989 );
xor ( n63991 , n63974 , n63990 );
buf ( n63992 , n56582 );
buf ( n63993 , n60261 );
and ( n63994 , n63992 , n63993 );
buf ( n63995 , n56585 );
buf ( n63996 , n60090 );
and ( n63997 , n63995 , n63996 );
nor ( n63998 , n63994 , n63997 );
buf ( n63999 , n63998 );
buf ( n64000 , n63999 );
buf ( n64001 , n60270 );
or ( n64002 , n64000 , n64001 );
buf ( n64003 , n62894 );
buf ( n64004 , n60100 );
or ( n64005 , n64003 , n64004 );
nand ( n64006 , n64002 , n64005 );
buf ( n64007 , n64006 );
and ( n64008 , n63991 , n64007 );
and ( n64009 , n63974 , n63990 );
or ( n64010 , n64008 , n64009 );
buf ( n64011 , n64010 );
buf ( n64012 , n62779 );
buf ( n64013 , n62790 );
or ( n64014 , n64012 , n64013 );
buf ( n64015 , n62793 );
nand ( n64016 , n64014 , n64015 );
buf ( n64017 , n64016 );
buf ( n64018 , n64017 );
xor ( n64019 , n64011 , n64018 );
buf ( n64020 , n60068 );
buf ( n64021 , n56641 );
and ( n64022 , n64020 , n64021 );
buf ( n64023 , n60071 );
buf ( n64024 , n56631 );
and ( n64025 , n64023 , n64024 );
nor ( n64026 , n64022 , n64025 );
buf ( n64027 , n64026 );
buf ( n64028 , n64027 );
buf ( n64029 , n56626 );
or ( n64030 , n64028 , n64029 );
buf ( n64031 , n62949 );
buf ( n64032 , n56639 );
or ( n64033 , n64031 , n64032 );
nand ( n64034 , n64030 , n64033 );
buf ( n64035 , n64034 );
buf ( n64036 , n64035 );
buf ( n64037 , n62782 );
buf ( n64038 , n56652 );
and ( n64039 , n64037 , n64038 );
buf ( n64040 , n62980 );
buf ( n64041 , n55201 );
and ( n64042 , n64040 , n64041 );
nor ( n64043 , n64039 , n64042 );
buf ( n64044 , n64043 );
buf ( n64045 , n64044 );
not ( n64046 , n64045 );
buf ( n64047 , n64046 );
buf ( n64048 , n64047 );
buf ( n64049 , n55180 );
and ( n64050 , n64048 , n64049 );
buf ( n64051 , n63039 );
not ( n64052 , n64051 );
buf ( n64053 , n64052 );
buf ( n64054 , n64053 );
buf ( n64055 , n56670 );
and ( n64056 , n64054 , n64055 );
nor ( n64057 , n64050 , n64056 );
buf ( n64058 , n64057 );
buf ( n64059 , n64058 );
nand ( n64060 , n55063 , n54726 );
not ( n64061 , n64060 );
not ( n64062 , n55060 );
nand ( n64063 , n62963 , n64062 );
not ( n64064 , n64063 );
or ( n64065 , n64061 , n64064 );
not ( n64066 , n64060 );
nand ( n64067 , n64066 , n62963 , n64062 );
nand ( n64068 , n64065 , n64067 );
buf ( n64069 , n64068 );
buf ( n64070 , n55132 );
and ( n64071 , n64069 , n64070 );
buf ( n64072 , n62971 );
buf ( n64073 , n64072 );
buf ( n64074 , n55156 );
and ( n64075 , n64073 , n64074 );
nor ( n64076 , n64071 , n64075 );
buf ( n64077 , n64076 );
buf ( n64078 , n64077 );
nand ( n64079 , n64059 , n64078 );
buf ( n64080 , n64079 );
buf ( n64081 , n64080 );
xor ( n64082 , n64036 , n64081 );
buf ( n64083 , n58835 );
buf ( n64084 , n58897 );
and ( n64085 , n64083 , n64084 );
buf ( n64086 , n58841 );
buf ( n64087 , n58894 );
and ( n64088 , n64086 , n64087 );
nor ( n64089 , n64085 , n64088 );
buf ( n64090 , n64089 );
buf ( n64091 , n64090 );
buf ( n64092 , n58913 );
or ( n64093 , n64091 , n64092 );
buf ( n64094 , n62878 );
buf ( n64095 , n58890 );
or ( n64096 , n64094 , n64095 );
nand ( n64097 , n64093 , n64096 );
buf ( n64098 , n64097 );
buf ( n64099 , n64098 );
and ( n64100 , n64082 , n64099 );
and ( n64101 , n64036 , n64081 );
or ( n64102 , n64100 , n64101 );
buf ( n64103 , n64102 );
buf ( n64104 , n64103 );
and ( n64105 , n64019 , n64104 );
and ( n64106 , n64011 , n64018 );
or ( n64107 , n64105 , n64106 );
buf ( n64108 , n64107 );
xor ( n64109 , n62836 , n62853 );
xor ( n64110 , n64109 , n62858 );
buf ( n64111 , n64110 );
xor ( n64112 , n64108 , n64111 );
xor ( n64113 , n62923 , n63058 );
xor ( n64114 , n64113 , n63063 );
buf ( n64115 , n64114 );
and ( n64116 , n64112 , n64115 );
and ( n64117 , n64108 , n64111 );
or ( n64118 , n64116 , n64117 );
xor ( n64119 , n63067 , n63070 );
xor ( n64120 , n64119 , n63075 );
and ( n64121 , n64118 , n64120 );
xor ( n64122 , n62941 , n62958 );
xor ( n64123 , n64122 , n63053 );
buf ( n64124 , n64123 );
xor ( n64125 , n62886 , n62902 );
xor ( n64126 , n64125 , n62919 );
and ( n64127 , n64124 , n64126 );
buf ( n64128 , n55152 );
not ( n64129 , n63015 );
buf ( n64130 , n64129 );
and ( n64131 , n64128 , n64130 );
buf ( n64132 , n55205 );
not ( n64133 , n64129 );
buf ( n64134 , n64133 );
and ( n64135 , n64132 , n64134 );
nor ( n64136 , n64131 , n64135 );
buf ( n64137 , n64136 );
buf ( n64138 , n64137 );
buf ( n64139 , n63013 );
not ( n64140 , n64139 );
buf ( n64141 , n64140 );
buf ( n64142 , n64141 );
or ( n64143 , n64138 , n64142 );
buf ( n64144 , n63026 );
nand ( n64145 , n64143 , n64144 );
buf ( n64146 , n64145 );
buf ( n64147 , n64146 );
buf ( n64148 , n60229 );
buf ( n64149 , n56641 );
and ( n64150 , n64148 , n64149 );
buf ( n64151 , n62652 );
buf ( n64152 , n56631 );
and ( n64153 , n64151 , n64152 );
nor ( n64154 , n64150 , n64153 );
buf ( n64155 , n64154 );
buf ( n64156 , n64155 );
buf ( n64157 , n56626 );
or ( n64158 , n64156 , n64157 );
buf ( n64159 , n64027 );
buf ( n64160 , n56639 );
or ( n64161 , n64159 , n64160 );
nand ( n64162 , n64158 , n64161 );
buf ( n64163 , n64162 );
buf ( n64164 , n64163 );
xor ( n64165 , n64147 , n64164 );
buf ( n64166 , n59009 );
buf ( n64167 , n58721 );
and ( n64168 , n64166 , n64167 );
buf ( n64169 , n60077 );
buf ( n64170 , n58718 );
and ( n64171 , n64169 , n64170 );
nor ( n64172 , n64168 , n64171 );
buf ( n64173 , n64172 );
buf ( n64174 , n64173 );
buf ( n64175 , n56799 );
or ( n64176 , n64174 , n64175 );
buf ( n64177 , n63966 );
buf ( n64178 , n58982 );
or ( n64179 , n64177 , n64178 );
nand ( n64180 , n64176 , n64179 );
buf ( n64181 , n64180 );
buf ( n64182 , n64181 );
and ( n64183 , n64165 , n64182 );
and ( n64184 , n64147 , n64164 );
or ( n64185 , n64183 , n64184 );
buf ( n64186 , n64185 );
buf ( n64187 , n64186 );
xor ( n64188 , n62986 , n63030 );
xor ( n64189 , n64188 , n63048 );
buf ( n64190 , n64189 );
buf ( n64191 , n64190 );
xor ( n64192 , n64187 , n64191 );
buf ( n64193 , n58699 );
buf ( n64194 , n62681 );
and ( n64195 , n64193 , n64194 );
buf ( n64196 , n56594 );
buf ( n64197 , n62663 );
and ( n64198 , n64196 , n64197 );
nor ( n64199 , n64195 , n64198 );
buf ( n64200 , n64199 );
buf ( n64201 , n64200 );
buf ( n64202 , n62935 );
or ( n64203 , n64201 , n64202 );
buf ( n64204 , n63982 );
buf ( n64205 , n62676 );
or ( n64206 , n64204 , n64205 );
nand ( n64207 , n64203 , n64206 );
buf ( n64208 , n64207 );
buf ( n64209 , n64208 );
nand ( n64210 , n64062 , n54711 );
xnor ( n64211 , n55056 , n64210 );
buf ( n64212 , n64211 );
buf ( n64213 , n55132 );
and ( n64214 , n64212 , n64213 );
buf ( n64215 , n64068 );
buf ( n64216 , n55156 );
and ( n64217 , n64215 , n64216 );
nor ( n64218 , n64214 , n64217 );
buf ( n64219 , n64218 );
buf ( n64220 , n64219 );
buf ( n64221 , n62999 );
not ( n64222 , n64221 );
buf ( n64223 , n64222 );
buf ( n64224 , n64223 );
buf ( n64225 , n1664 );
not ( n64226 , n64225 );
buf ( n64227 , n64226 );
buf ( n64228 , n64227 );
nand ( n64229 , n64224 , n64228 );
buf ( n64230 , n64229 );
buf ( n64231 , n64230 );
buf ( n64232 , n64223 );
buf ( n64233 , n1664 );
nand ( n64234 , n64232 , n64233 );
buf ( n64235 , n64234 );
buf ( n64236 , n64235 );
nand ( n64237 , n64231 , n64236 );
buf ( n64238 , n64237 );
buf ( n64239 , n64238 );
nand ( n64240 , n64220 , n64239 );
buf ( n64241 , n64240 );
buf ( n64242 , n64241 );
xor ( n64243 , n64209 , n64242 );
buf ( n64244 , n58894 );
buf ( n64245 , n58862 );
and ( n64246 , n64244 , n64245 );
not ( n64247 , n64244 );
buf ( n64248 , n58823 );
and ( n64249 , n64247 , n64248 );
nor ( n64250 , n64246 , n64249 );
buf ( n64251 , n64250 );
buf ( n64252 , n64251 );
buf ( n64253 , n58913 );
or ( n64254 , n64252 , n64253 );
buf ( n64255 , n64090 );
buf ( n64256 , n58890 );
or ( n64257 , n64255 , n64256 );
nand ( n64258 , n64254 , n64257 );
buf ( n64259 , n64258 );
buf ( n64260 , n64259 );
and ( n64261 , n64243 , n64260 );
and ( n64262 , n64209 , n64242 );
or ( n64263 , n64261 , n64262 );
buf ( n64264 , n64263 );
buf ( n64265 , n64264 );
and ( n64266 , n64192 , n64265 );
and ( n64267 , n64187 , n64191 );
or ( n64268 , n64266 , n64267 );
buf ( n64269 , n64268 );
xor ( n64270 , n62886 , n62902 );
xor ( n64271 , n64270 , n62919 );
and ( n64272 , n64269 , n64271 );
and ( n64273 , n64124 , n64269 );
or ( n64274 , n64127 , n64272 , n64273 );
xor ( n64275 , n64108 , n64111 );
xor ( n64276 , n64275 , n64115 );
and ( n64277 , n64274 , n64276 );
xor ( n64278 , n64036 , n64081 );
xor ( n64279 , n64278 , n64099 );
buf ( n64280 , n64279 );
xor ( n64281 , n63974 , n63990 );
xor ( n64282 , n64281 , n64007 );
and ( n64283 , n64280 , n64282 );
buf ( n64284 , n56720 );
buf ( n64285 , n60261 );
and ( n64286 , n64284 , n64285 );
buf ( n64287 , n58792 );
buf ( n64288 , n60090 );
and ( n64289 , n64287 , n64288 );
nor ( n64290 , n64286 , n64289 );
buf ( n64291 , n64290 );
buf ( n64292 , n64291 );
buf ( n64293 , n60270 );
or ( n64294 , n64292 , n64293 );
buf ( n64295 , n63999 );
buf ( n64296 , n60100 );
or ( n64297 , n64295 , n64296 );
nand ( n64298 , n64294 , n64297 );
buf ( n64299 , n64298 );
buf ( n64300 , n64058 );
buf ( n64301 , n64077 );
or ( n64302 , n64300 , n64301 );
buf ( n64303 , n64080 );
nand ( n64304 , n64302 , n64303 );
buf ( n64305 , n64304 );
xor ( n64306 , n64299 , n64305 );
buf ( n64307 , n56631 );
buf ( n64308 , n62646 );
and ( n64309 , n64307 , n64308 );
not ( n64310 , n64307 );
buf ( n64311 , n62643 );
and ( n64312 , n64310 , n64311 );
nor ( n64313 , n64309 , n64312 );
buf ( n64314 , n64313 );
buf ( n64315 , n64314 );
buf ( n64316 , n56626 );
or ( n64317 , n64315 , n64316 );
buf ( n64318 , n64155 );
buf ( n64319 , n56639 );
or ( n64320 , n64318 , n64319 );
nand ( n64321 , n64317 , n64320 );
buf ( n64322 , n64321 );
buf ( n64323 , n64322 );
buf ( n64324 , n62971 );
buf ( n64325 , n56652 );
and ( n64326 , n64324 , n64325 );
buf ( n64327 , n62974 );
buf ( n64328 , n55201 );
and ( n64329 , n64327 , n64328 );
nor ( n64330 , n64326 , n64329 );
buf ( n64331 , n64330 );
buf ( n64332 , n64331 );
buf ( n64333 , n56664 );
or ( n64334 , n64332 , n64333 );
buf ( n64335 , n64044 );
buf ( n64336 , n56673 );
or ( n64337 , n64335 , n64336 );
nand ( n64338 , n64334 , n64337 );
buf ( n64339 , n64338 );
buf ( n64340 , n64339 );
xor ( n64341 , n64323 , n64340 );
buf ( n64342 , n60068 );
buf ( n64343 , n58721 );
and ( n64344 , n64342 , n64343 );
buf ( n64345 , n60071 );
buf ( n64346 , n58718 );
and ( n64347 , n64345 , n64346 );
nor ( n64348 , n64344 , n64347 );
buf ( n64349 , n64348 );
buf ( n64350 , n64349 );
buf ( n64351 , n56799 );
or ( n64352 , n64350 , n64351 );
buf ( n64353 , n64173 );
buf ( n64354 , n58982 );
or ( n64355 , n64353 , n64354 );
nand ( n64356 , n64352 , n64355 );
buf ( n64357 , n64356 );
buf ( n64358 , n64357 );
and ( n64359 , n64341 , n64358 );
and ( n64360 , n64323 , n64340 );
or ( n64361 , n64359 , n64360 );
buf ( n64362 , n64361 );
and ( n64363 , n64306 , n64362 );
and ( n64364 , n64299 , n64305 );
or ( n64365 , n64363 , n64364 );
xor ( n64366 , n63974 , n63990 );
xor ( n64367 , n64366 , n64007 );
and ( n64368 , n64365 , n64367 );
and ( n64369 , n64280 , n64365 );
or ( n64370 , n64283 , n64368 , n64369 );
xor ( n64371 , n64011 , n64018 );
xor ( n64372 , n64371 , n64104 );
buf ( n64373 , n64372 );
or ( n64374 , n64370 , n64373 );
not ( n64375 , n64374 );
xor ( n64376 , n62886 , n62902 );
xor ( n64377 , n64376 , n62919 );
xor ( n64378 , n64124 , n64269 );
xor ( n64379 , n64377 , n64378 );
not ( n64380 , n64379 );
or ( n64381 , n64375 , n64380 );
nand ( n64382 , n64373 , n64370 );
nand ( n64383 , n64381 , n64382 );
xor ( n64384 , n64108 , n64111 );
xor ( n64385 , n64384 , n64115 );
and ( n64386 , n64383 , n64385 );
and ( n64387 , n64274 , n64383 );
or ( n64388 , n64277 , n64386 , n64387 );
xor ( n64389 , n63067 , n63070 );
xor ( n64390 , n64389 , n63075 );
and ( n64391 , n64388 , n64390 );
and ( n64392 , n64118 , n64388 );
or ( n64393 , n64121 , n64391 , n64392 );
buf ( n64394 , n64393 );
xor ( n64395 , n63958 , n64394 );
buf ( n64396 , n42008 );
not ( n64397 , n64396 );
buf ( n64398 , n41657 );
not ( n64399 , n64398 );
or ( n64400 , n64397 , n64399 );
buf ( n64401 , n61434 );
buf ( n64402 , n63633 );
nand ( n64403 , n64401 , n64402 );
buf ( n64404 , n64403 );
buf ( n64405 , n64404 );
nand ( n64406 , n64400 , n64405 );
buf ( n64407 , n64406 );
buf ( n64408 , n64407 );
not ( n64409 , n64408 );
nand ( n64410 , n62579 , n41699 , n41702 );
buf ( n64411 , n64410 );
not ( n64412 , n64411 );
buf ( n64413 , n64412 );
buf ( n64414 , n64413 );
not ( n64415 , n64414 );
or ( n64416 , n64409 , n64415 );
buf ( n64417 , n63882 );
buf ( n64418 , n62582 );
nand ( n64419 , n64417 , n64418 );
buf ( n64420 , n64419 );
buf ( n64421 , n64420 );
nand ( n64422 , n64416 , n64421 );
buf ( n64423 , n64422 );
buf ( n64424 , n64423 );
and ( n64425 , n64395 , n64424 );
and ( n64426 , n63958 , n64394 );
or ( n64427 , n64425 , n64426 );
buf ( n64428 , n64427 );
buf ( n64429 , n64428 );
not ( n64430 , n64429 );
buf ( n64431 , n64430 );
buf ( n64432 , n64431 );
nand ( n64433 , n63953 , n64432 );
buf ( n64434 , n64433 );
not ( n64435 , n64434 );
or ( n64436 , n63927 , n64435 );
buf ( n64437 , n64428 );
buf ( n64438 , n63951 );
nand ( n64439 , n64437 , n64438 );
buf ( n64440 , n64439 );
nand ( n64441 , n64436 , n64440 );
buf ( n64442 , n64441 );
nand ( n64443 , n63869 , n64442 );
buf ( n64444 , n64443 );
buf ( n64445 , n64444 );
buf ( n64446 , n63866 );
not ( n64447 , n64446 );
buf ( n64448 , n63845 );
nand ( n64449 , n64447 , n64448 );
buf ( n64450 , n64449 );
buf ( n64451 , n64450 );
nand ( n64452 , n64445 , n64451 );
buf ( n64453 , n64452 );
buf ( n64454 , n64453 );
xor ( n64455 , n63827 , n64454 );
buf ( n64456 , n41947 );
not ( n64457 , n64456 );
buf ( n64458 , n52789 );
not ( n64459 , n64458 );
and ( n64460 , n64457 , n64459 );
buf ( n64461 , n41947 );
buf ( n64462 , n52789 );
and ( n64463 , n64461 , n64462 );
nor ( n64464 , n64460 , n64463 );
buf ( n64465 , n64464 );
buf ( n64466 , n64465 );
not ( n64467 , n64466 );
buf ( n64468 , n64467 );
buf ( n64469 , n64468 );
not ( n64470 , n64469 );
buf ( n64471 , n37872 );
not ( n64472 , n64471 );
or ( n64473 , n64470 , n64472 );
buf ( n64474 , n42175 );
buf ( n64475 , n53946 );
not ( n64476 , n64475 );
buf ( n64477 , n41925 );
not ( n64478 , n64477 );
or ( n64479 , n64476 , n64478 );
buf ( n64480 , n43813 );
buf ( n64481 , n52094 );
nand ( n64482 , n64480 , n64481 );
buf ( n64483 , n64482 );
buf ( n64484 , n64483 );
nand ( n64485 , n64479 , n64484 );
buf ( n64486 , n64485 );
buf ( n64487 , n64486 );
nand ( n64488 , n64474 , n64487 );
buf ( n64489 , n64488 );
buf ( n64490 , n64489 );
nand ( n64491 , n64473 , n64490 );
buf ( n64492 , n64491 );
buf ( n64493 , n64492 );
and ( n64494 , n64455 , n64493 );
and ( n64495 , n63827 , n64454 );
or ( n64496 , n64494 , n64495 );
buf ( n64497 , n64496 );
buf ( n64498 , n64497 );
and ( n64499 , n63802 , n64498 );
and ( n64500 , n63780 , n63801 );
or ( n64501 , n64499 , n64500 );
buf ( n64502 , n64501 );
buf ( n64503 , n64502 );
xor ( n64504 , n63776 , n64503 );
not ( n64505 , n43371 );
buf ( n64506 , n36901 );
buf ( n64507 , n64506 );
buf ( n64508 , n64507 );
nor ( n64509 , n64505 , n64508 );
not ( n64510 , n64509 );
not ( n64511 , n56325 );
and ( n64512 , n64510 , n64511 );
buf ( n64513 , n64508 );
not ( n64514 , n64513 );
buf ( n64515 , n49391 );
not ( n64516 , n64515 );
or ( n64517 , n64514 , n64516 );
buf ( n64518 , n43095 );
nand ( n64519 , n64517 , n64518 );
buf ( n64520 , n64519 );
nor ( n64521 , n64512 , n64520 );
not ( n64522 , n64486 );
not ( n64523 , n37872 );
or ( n64524 , n64522 , n64523 );
buf ( n64525 , n62388 );
not ( n64526 , n64525 );
buf ( n64527 , n37919 );
nand ( n64528 , n64526 , n64527 );
buf ( n64529 , n64528 );
nand ( n64530 , n64524 , n64529 );
xor ( n64531 , n64521 , n64530 );
not ( n64532 , n63108 );
not ( n64533 , n64532 );
buf ( n64534 , n63116 );
not ( n64535 , n64534 );
buf ( n64536 , n62553 );
not ( n64537 , n64536 );
or ( n64538 , n64535 , n64537 );
buf ( n64539 , n62553 );
buf ( n64540 , n63116 );
or ( n64541 , n64539 , n64540 );
nand ( n64542 , n64538 , n64541 );
buf ( n64543 , n64542 );
not ( n64544 , n64543 );
or ( n64545 , n64533 , n64544 );
or ( n64546 , n64543 , n64532 );
nand ( n64547 , n64545 , n64546 );
xor ( n64548 , n64531 , n64547 );
buf ( n64549 , n64548 );
not ( n64550 , n64549 );
not ( n64551 , n48868 );
not ( n64552 , n48808 );
not ( n64553 , n37717 );
or ( n64554 , n64552 , n64553 );
not ( n64555 , n42573 );
nand ( n64556 , n64555 , n48821 );
nand ( n64557 , n64554 , n64556 );
not ( n64558 , n64557 );
or ( n64559 , n64551 , n64558 );
not ( n64560 , n48818 );
not ( n64561 , n43198 );
or ( n64562 , n64560 , n64561 );
or ( n64563 , n39522 , n48821 );
nand ( n64564 , n64562 , n64563 );
buf ( n64565 , n64564 );
buf ( n64566 , n48855 );
nand ( n64567 , n64565 , n64566 );
buf ( n64568 , n64567 );
nand ( n64569 , n64559 , n64568 );
buf ( n64570 , n64569 );
not ( n64571 , n64570 );
or ( n64572 , n64550 , n64571 );
buf ( n64573 , n64548 );
buf ( n64574 , n64569 );
or ( n64575 , n64573 , n64574 );
xor ( n64576 , n63690 , n63715 );
xor ( n64577 , n64576 , n63742 );
buf ( n64578 , n64577 );
buf ( n64579 , n64578 );
not ( n64580 , n44253 );
not ( n64581 , n63611 );
not ( n64582 , n64581 );
or ( n64583 , n64580 , n64582 );
or ( n64584 , n41828 , n51004 );
nand ( n64585 , n41981 , n51004 );
nand ( n64586 , n64584 , n64585 );
not ( n64587 , n64586 );
nand ( n64588 , n64587 , n41966 );
nand ( n64589 , n64583 , n64588 );
buf ( n64590 , n64589 );
xor ( n64591 , n64579 , n64590 );
buf ( n64592 , n44679 );
buf ( n64593 , n12481 );
and ( n64594 , n64592 , n64593 );
buf ( n64595 , n64594 );
buf ( n64596 , n64595 );
and ( n64597 , n64591 , n64596 );
and ( n64598 , n64579 , n64590 );
or ( n64599 , n64597 , n64598 );
buf ( n64600 , n64599 );
buf ( n64601 , n64600 );
nand ( n64602 , n64575 , n64601 );
buf ( n64603 , n64602 );
buf ( n64604 , n64603 );
nand ( n64605 , n64572 , n64604 );
buf ( n64606 , n64605 );
buf ( n64607 , n64606 );
and ( n64608 , n64504 , n64607 );
and ( n64609 , n63776 , n64503 );
or ( n64610 , n64608 , n64609 );
buf ( n64611 , n64610 );
buf ( n64612 , n64611 );
buf ( n64613 , C0 );
buf ( n64614 , n64613 );
not ( n64615 , n46246 );
not ( n64616 , n45747 );
buf ( n64617 , n64616 );
not ( n64618 , n64617 );
buf ( n64619 , n42461 );
not ( n64620 , n64619 );
or ( n64621 , n64618 , n64620 );
buf ( n64622 , n38821 );
buf ( n64623 , n45747 );
nand ( n64624 , n64622 , n64623 );
buf ( n64625 , n64624 );
buf ( n64626 , n64625 );
nand ( n64627 , n64621 , n64626 );
buf ( n64628 , n64627 );
not ( n64629 , n64628 );
or ( n64630 , n64615 , n64629 );
and ( n64631 , n64616 , n44989 );
not ( n64632 , n64616 );
and ( n64633 , n64632 , n38848 );
or ( n64634 , n64631 , n64633 );
nand ( n64635 , n64634 , n46225 );
nand ( n64636 , n64630 , n64635 );
not ( n64637 , n64636 );
buf ( n64638 , n64637 );
not ( n64639 , n64638 );
buf ( n64640 , n43868 );
not ( n64641 , n64640 );
buf ( n64642 , n41608 );
not ( n64643 , n64642 );
buf ( n64644 , n44025 );
not ( n64645 , n64644 );
or ( n64646 , n64643 , n64645 );
buf ( n64647 , n28306 );
buf ( n64648 , n41604 );
nand ( n64649 , n64647 , n64648 );
buf ( n64650 , n64649 );
buf ( n64651 , n64650 );
nand ( n64652 , n64646 , n64651 );
buf ( n64653 , n64652 );
buf ( n64654 , n64653 );
not ( n64655 , n64654 );
or ( n64656 , n64641 , n64655 );
buf ( n64657 , n41608 );
not ( n64658 , n64657 );
buf ( n64659 , n45075 );
not ( n64660 , n64659 );
or ( n64661 , n64658 , n64660 );
buf ( n64662 , n41822 );
buf ( n64663 , n41604 );
nand ( n64664 , n64662 , n64663 );
buf ( n64665 , n64664 );
buf ( n64666 , n64665 );
nand ( n64667 , n64661 , n64666 );
buf ( n64668 , n64667 );
buf ( n64669 , n64668 );
buf ( n64670 , n44267 );
nand ( n64671 , n64669 , n64670 );
buf ( n64672 , n64671 );
buf ( n64673 , n64672 );
nand ( n64674 , n64656 , n64673 );
buf ( n64675 , n64674 );
buf ( n64676 , n64675 );
not ( n64677 , n45069 );
not ( n64678 , n47725 );
and ( n64679 , n64677 , n64678 );
not ( n64680 , n47068 );
and ( n64681 , n64680 , n47725 );
nor ( n64682 , n64679 , n64681 );
not ( n64683 , n64682 );
not ( n64684 , n46620 );
or ( n64685 , n64683 , n64684 );
buf ( n64686 , n46390 );
not ( n64687 , n64686 );
buf ( n64688 , n42403 );
not ( n64689 , n64688 );
or ( n64690 , n64687 , n64689 );
buf ( n64691 , n46623 );
buf ( n64692 , n46393 );
nand ( n64693 , n64691 , n64692 );
buf ( n64694 , n64693 );
buf ( n64695 , n64694 );
nand ( n64696 , n64690 , n64695 );
buf ( n64697 , n64696 );
buf ( n64698 , n64697 );
buf ( n64699 , n38380 );
nand ( n64700 , n64698 , n64699 );
buf ( n64701 , n64700 );
nand ( n64702 , n64685 , n64701 );
buf ( n64703 , n64702 );
or ( n64704 , n64676 , n64703 );
buf ( n64705 , n64704 );
buf ( n64706 , n42865 );
not ( n64707 , n64706 );
buf ( n64708 , n52670 );
not ( n64709 , n64708 );
or ( n64710 , n64707 , n64709 );
buf ( n64711 , n25159 );
buf ( n64712 , n42862 );
nand ( n64713 , n64711 , n64712 );
buf ( n64714 , n64713 );
buf ( n64715 , n64714 );
nand ( n64716 , n64710 , n64715 );
buf ( n64717 , n64716 );
buf ( n64718 , n64717 );
not ( n64719 , n64718 );
buf ( n64720 , n50128 );
not ( n64721 , n64720 );
or ( n64722 , n64719 , n64721 );
buf ( n64723 , n47872 );
buf ( n64724 , n43063 );
not ( n64725 , n64724 );
buf ( n64726 , n52670 );
not ( n64727 , n64726 );
or ( n64728 , n64725 , n64727 );
buf ( n64729 , n25159 );
buf ( n64730 , n43064 );
nand ( n64731 , n64729 , n64730 );
buf ( n64732 , n64731 );
buf ( n64733 , n64732 );
nand ( n64734 , n64728 , n64733 );
buf ( n64735 , n64734 );
buf ( n64736 , n64735 );
nand ( n64737 , n64723 , n64736 );
buf ( n64738 , n64737 );
buf ( n64739 , n64738 );
nand ( n64740 , n64722 , n64739 );
buf ( n64741 , n64740 );
not ( n64742 , n64741 );
buf ( n64743 , n42668 );
not ( n64744 , n64743 );
buf ( n64745 , n63843 );
not ( n64746 , n64745 );
or ( n64747 , n64744 , n64746 );
buf ( n64748 , n25226 );
not ( n64749 , n64748 );
not ( n64750 , n48169 );
or ( n64751 , n64749 , n64750 );
buf ( n64752 , n28368 );
not ( n64753 , n64748 );
buf ( n64754 , n64753 );
nand ( n64755 , n64752 , n64754 );
buf ( n64756 , n64755 );
nand ( n64757 , n64751 , n64756 );
nand ( n64758 , n64757 , n58249 );
buf ( n64759 , n64758 );
nand ( n64760 , n64747 , n64759 );
buf ( n64761 , n64760 );
not ( n64762 , n64761 );
or ( n64763 , n64742 , n64762 );
not ( n64764 , n64741 );
not ( n64765 , n64764 );
not ( n64766 , n64761 );
not ( n64767 , n64766 );
or ( n64768 , n64765 , n64767 );
not ( n64769 , n24092 );
not ( n64770 , n44949 );
or ( n64771 , n64769 , n64770 );
nand ( n64772 , n47857 , n44952 );
nand ( n64773 , n64771 , n64772 );
not ( n64774 , n64773 );
buf ( n64775 , n48970 );
not ( n64776 , n64775 );
buf ( n64777 , n64776 );
not ( n64778 , n64777 );
or ( n64779 , n64774 , n64778 );
buf ( n64780 , n42847 );
buf ( n64781 , n55743 );
and ( n64782 , n64780 , n64781 );
not ( n64783 , n64780 );
buf ( n64784 , n24092 );
and ( n64785 , n64783 , n64784 );
nor ( n64786 , n64782 , n64785 );
buf ( n64787 , n64786 );
or ( n64788 , n39980 , n64787 );
nand ( n64789 , n64779 , n64788 );
nand ( n64790 , n64768 , n64789 );
nand ( n64791 , n64763 , n64790 );
and ( n64792 , n64705 , n64791 );
buf ( n64793 , n64675 );
buf ( n64794 , n64702 );
and ( n64795 , n64793 , n64794 );
buf ( n64796 , n64795 );
nor ( n64797 , n64792 , n64796 );
buf ( n64798 , n64797 );
not ( n64799 , n64798 );
or ( n64800 , n64639 , n64799 );
xor ( n64801 , n63652 , n63669 );
xor ( n64802 , n64801 , n63685 );
buf ( n64803 , n64802 );
not ( n64804 , n64803 );
buf ( n64805 , n42315 );
not ( n64806 , n64805 );
buf ( n64807 , n63707 );
not ( n64808 , n64807 );
or ( n64809 , n64806 , n64808 );
nand ( n64810 , n59242 , n41873 );
not ( n64811 , n64810 );
buf ( n64812 , n50575 );
buf ( n64813 , n42260 );
nand ( n64814 , n64812 , n64813 );
buf ( n64815 , n64814 );
not ( n64816 , n64815 );
or ( n64817 , n64811 , n64816 );
nand ( n64818 , n64817 , n42252 );
buf ( n64819 , n64818 );
nand ( n64820 , n64809 , n64819 );
buf ( n64821 , n64820 );
not ( n64822 , n64821 );
nand ( n64823 , n64804 , n64822 );
not ( n64824 , n64823 );
buf ( n64825 , n45376 );
buf ( n64826 , n37880 );
buf ( n64827 , n38120 );
nand ( n64828 , n64826 , n64827 );
buf ( n64829 , n64828 );
buf ( n64830 , n64829 );
buf ( n64831 , n12481 );
and ( n64832 , n64830 , n64831 );
buf ( n64833 , n37881 );
buf ( n64834 , n38112 );
and ( n64835 , n64833 , n64834 );
nor ( n64836 , n64832 , n64835 );
buf ( n64837 , n64836 );
buf ( n64838 , n64837 );
and ( n64839 , n64825 , n64838 );
buf ( n64840 , n64839 );
not ( n64841 , n64840 );
or ( n64842 , n64824 , n64841 );
nand ( n64843 , n64821 , n64803 );
nand ( n64844 , n64842 , n64843 );
buf ( n64845 , n64844 );
nand ( n64846 , n64800 , n64845 );
buf ( n64847 , n64846 );
buf ( n64848 , n64797 );
not ( n64849 , n64848 );
buf ( n64850 , n64849 );
buf ( n64851 , n64850 );
buf ( n64852 , n64636 );
nand ( n64853 , n64851 , n64852 );
buf ( n64854 , n64853 );
nand ( n64855 , n64847 , n64854 );
buf ( n64856 , n64855 );
not ( n64857 , n64856 );
buf ( n64858 , n46912 );
not ( n64859 , n64858 );
buf ( n64860 , n63559 );
not ( n64861 , n64860 );
or ( n64862 , n64859 , n64861 );
and ( n64863 , n44157 , n46875 );
not ( n64864 , n44157 );
and ( n64865 , n64864 , n46887 );
or ( n64866 , n64863 , n64865 );
buf ( n64867 , n64866 );
buf ( n64868 , n47331 );
nand ( n64869 , n64867 , n64868 );
buf ( n64870 , n64869 );
buf ( n64871 , n64870 );
nand ( n64872 , n64862 , n64871 );
buf ( n64873 , n64872 );
buf ( n64874 , n64873 );
not ( n64875 , n64874 );
or ( n64876 , n64857 , n64875 );
buf ( n64877 , n63746 );
not ( n64878 , n64877 );
buf ( n64879 , n64878 );
and ( n64880 , n63597 , n64879 );
not ( n64881 , n63597 );
and ( n64882 , n64881 , n63746 );
nor ( n64883 , n64880 , n64882 );
not ( n64884 , n63621 );
and ( n64885 , n64883 , n64884 );
not ( n64886 , n64883 );
and ( n64887 , n64886 , n63621 );
nor ( n64888 , n64885 , n64887 );
not ( n64889 , n64873 );
nand ( n64890 , n64889 , n64847 , n64854 );
nand ( n64891 , n64888 , n64890 );
buf ( n64892 , n64891 );
nand ( n64893 , n64876 , n64892 );
buf ( n64894 , n64893 );
buf ( n64895 , n64894 );
xor ( n64896 , n64614 , n64895 );
xor ( n64897 , n63545 , n63571 );
xor ( n64898 , n64897 , n63759 );
buf ( n64899 , n64898 );
buf ( n64900 , n64899 );
and ( n64901 , n64896 , n64900 );
or ( n64902 , n64901 , C0 );
buf ( n64903 , n64902 );
buf ( n64904 , n64903 );
xor ( n64905 , n64612 , n64904 );
buf ( n64906 , n63533 );
buf ( n64907 , n63529 );
xor ( n64908 , n64906 , n64907 );
buf ( n64909 , n63763 );
xor ( n64910 , n64908 , n64909 );
buf ( n64911 , n64910 );
buf ( n64912 , n64911 );
and ( n64913 , n64905 , n64912 );
and ( n64914 , n64612 , n64904 );
or ( n64915 , n64913 , n64914 );
buf ( n64916 , n64915 );
buf ( n64917 , n64916 );
xor ( n64918 , n63772 , n64917 );
and ( n64919 , n62485 , n62471 );
not ( n64920 , n62485 );
and ( n64921 , n64920 , n62472 );
nor ( n64922 , n64919 , n64921 );
and ( n64923 , n64922 , n62468 );
not ( n64924 , n64922 );
and ( n64925 , n64924 , n62467 );
nor ( n64926 , n64923 , n64925 );
buf ( n64927 , n64926 );
buf ( n64928 , C0 );
buf ( n64929 , n64928 );
xor ( n64930 , n64927 , n64929 );
xor ( n64931 , n64521 , n64530 );
and ( n64932 , n64931 , n64547 );
and ( n64933 , n64521 , n64530 );
or ( n64934 , n64932 , n64933 );
buf ( n64935 , n64934 );
not ( n64936 , n62421 );
xor ( n64937 , n62425 , n64936 );
xor ( n64938 , n64937 , n62432 );
buf ( n64939 , n64938 );
xor ( n64940 , n64935 , n64939 );
buf ( n64941 , n48855 );
not ( n64942 , n64941 );
buf ( n64943 , n64557 );
not ( n64944 , n64943 );
or ( n64945 , n64942 , n64944 );
buf ( n64946 , n62167 );
buf ( n64947 , n48868 );
nand ( n64948 , n64946 , n64947 );
buf ( n64949 , n64948 );
buf ( n64950 , n64949 );
nand ( n64951 , n64945 , n64950 );
buf ( n64952 , n64951 );
buf ( n64953 , n64952 );
and ( n64954 , n64940 , n64953 );
and ( n64955 , n64935 , n64939 );
or ( n64956 , n64954 , n64955 );
buf ( n64957 , n64956 );
buf ( n64958 , n64957 );
xor ( n64959 , n64930 , n64958 );
buf ( n64960 , n64959 );
buf ( n64961 , n64960 );
not ( n64962 , n43991 );
buf ( n64963 , n53539 );
not ( n64964 , n64963 );
buf ( n64965 , n44635 );
not ( n64966 , n64965 );
or ( n64967 , n64964 , n64966 );
buf ( n64968 , n43403 );
buf ( n64969 , n53548 );
nand ( n64970 , n64968 , n64969 );
buf ( n64971 , n64970 );
buf ( n64972 , n64971 );
nand ( n64973 , n64967 , n64972 );
buf ( n64974 , n64973 );
not ( n64975 , n64974 );
or ( n64976 , n64962 , n64975 );
buf ( n64977 , n62197 );
buf ( n64978 , n45144 );
nand ( n64979 , n64977 , n64978 );
buf ( n64980 , n64979 );
nand ( n64981 , n64976 , n64980 );
buf ( n64982 , n63223 );
buf ( n64983 , n63279 );
xor ( n64984 , n64982 , n64983 );
buf ( n64985 , n63249 );
xnor ( n64986 , n64984 , n64985 );
buf ( n64987 , n64986 );
buf ( n64988 , n64987 );
not ( n64989 , n64988 );
buf ( n64990 , n64989 );
not ( n64991 , n64990 );
buf ( n64992 , n44267 );
not ( n64993 , n64992 );
buf ( n64994 , n64653 );
not ( n64995 , n64994 );
or ( n64996 , n64993 , n64995 );
buf ( n64997 , n43868 );
buf ( n64998 , n63589 );
nand ( n64999 , n64997 , n64998 );
buf ( n65000 , n64999 );
buf ( n65001 , n65000 );
nand ( n65002 , n64996 , n65001 );
buf ( n65003 , n65002 );
buf ( n65004 , n65003 );
not ( n65005 , n65004 );
buf ( n65006 , n44517 );
not ( n65007 , n65006 );
buf ( n65008 , n44530 );
not ( n65009 , n65008 );
buf ( n65010 , n65009 );
buf ( n65011 , n65010 );
not ( n65012 , n65011 );
buf ( n65013 , n39656 );
not ( n65014 , n65013 );
or ( n65015 , n65012 , n65014 );
buf ( n65016 , n39653 );
buf ( n65017 , n44530 );
nand ( n65018 , n65016 , n65017 );
buf ( n65019 , n65018 );
buf ( n65020 , n65019 );
nand ( n65021 , n65015 , n65020 );
buf ( n65022 , n65021 );
buf ( n65023 , n65022 );
not ( n65024 , n65023 );
or ( n65025 , n65007 , n65024 );
buf ( n65026 , n65010 );
not ( n65027 , n65026 );
buf ( n65028 , n42425 );
not ( n65029 , n65028 );
or ( n65030 , n65027 , n65029 );
buf ( n65031 , n50043 );
buf ( n65032 , n44530 );
nand ( n65033 , n65031 , n65032 );
buf ( n65034 , n65033 );
buf ( n65035 , n65034 );
nand ( n65036 , n65030 , n65035 );
buf ( n65037 , n65036 );
buf ( n65038 , n65037 );
buf ( n65039 , n44496 );
nand ( n65040 , n65038 , n65039 );
buf ( n65041 , n65040 );
buf ( n65042 , n65041 );
nand ( n65043 , n65025 , n65042 );
buf ( n65044 , n65043 );
buf ( n65045 , n65044 );
not ( n65046 , n65045 );
buf ( n65047 , n65046 );
buf ( n65048 , n65047 );
nand ( n65049 , n65005 , n65048 );
buf ( n65050 , n65049 );
not ( n65051 , n65050 );
or ( n65052 , n64991 , n65051 );
nand ( n65053 , n65044 , n65003 );
nand ( n65054 , n65052 , n65053 );
xor ( n65055 , n64981 , n65054 );
xor ( n65056 , n63285 , n63172 );
xnor ( n65057 , n65056 , n63196 );
not ( n65058 , n65057 );
xnor ( n65059 , n65055 , n65058 );
buf ( n65060 , n65059 );
not ( n65061 , n65060 );
not ( n65062 , n48836 );
not ( n65063 , n43143 );
or ( n65064 , n65062 , n65063 );
buf ( n65065 , n50463 );
buf ( n65066 , n51493 );
nand ( n65067 , n65065 , n65066 );
buf ( n65068 , n65067 );
nand ( n65069 , n65064 , n65068 );
buf ( n65070 , n65069 );
buf ( n65071 , n52456 );
and ( n65072 , n65070 , n65071 );
and ( n65073 , n37293 , n51496 );
not ( n65074 , n37293 );
and ( n65075 , n65074 , n51493 );
nor ( n65076 , n65073 , n65075 );
not ( n65077 , n65076 );
nor ( n65078 , n65077 , n51489 );
buf ( n65079 , n65078 );
nor ( n65080 , n65072 , n65079 );
buf ( n65081 , n65080 );
buf ( n65082 , n65081 );
not ( n65083 , n65082 );
or ( n65084 , n65061 , n65083 );
buf ( n65085 , n65003 );
not ( n65086 , n65085 );
buf ( n65087 , n64987 );
not ( n65088 , n65087 );
or ( n65089 , n65086 , n65088 );
buf ( n65090 , n65003 );
buf ( n65091 , n64987 );
or ( n65092 , n65090 , n65091 );
nand ( n65093 , n65089 , n65092 );
buf ( n65094 , n65093 );
buf ( n65095 , n65094 );
buf ( n65096 , n65044 );
and ( n65097 , n65095 , n65096 );
not ( n65098 , n65095 );
buf ( n65099 , n65047 );
and ( n65100 , n65098 , n65099 );
nor ( n65101 , n65097 , n65100 );
buf ( n65102 , n65101 );
buf ( n65103 , n65102 );
not ( n65104 , n65103 );
buf ( n65105 , n65104 );
buf ( n65106 , n65105 );
not ( n65107 , n44496 );
not ( n65108 , n65022 );
or ( n65109 , n65107 , n65108 );
buf ( n65110 , n65010 );
not ( n65111 , n65110 );
buf ( n65112 , n41975 );
not ( n65113 , n65112 );
or ( n65114 , n65111 , n65113 );
buf ( n65115 , n28723 );
buf ( n65116 , n44530 );
nand ( n65117 , n65115 , n65116 );
buf ( n65118 , n65117 );
buf ( n65119 , n65118 );
nand ( n65120 , n65114 , n65119 );
buf ( n65121 , n65120 );
buf ( n65122 , n65121 );
buf ( n65123 , n44517 );
nand ( n65124 , n65122 , n65123 );
buf ( n65125 , n65124 );
nand ( n65126 , n65109 , n65125 );
buf ( n65127 , n65126 );
not ( n65128 , n65127 );
buf ( n65129 , n50060 );
not ( n65130 , n65129 );
buf ( n65131 , n45270 );
not ( n65132 , n65131 );
or ( n65133 , n65130 , n65132 );
buf ( n65134 , n41769 );
buf ( n65135 , n50067 );
nand ( n65136 , n65134 , n65135 );
buf ( n65137 , n65136 );
buf ( n65138 , n65137 );
nand ( n65139 , n65133 , n65138 );
buf ( n65140 , n65139 );
not ( n65141 , n65140 );
not ( n65142 , n37400 );
or ( n65143 , n65141 , n65142 );
buf ( n65144 , n63814 );
buf ( n65145 , n42135 );
nand ( n65146 , n65144 , n65145 );
buf ( n65147 , n65146 );
nand ( n65148 , n65143 , n65147 );
buf ( n65149 , n65148 );
not ( n65150 , n65149 );
or ( n65151 , n65128 , n65150 );
buf ( n65152 , n65126 );
buf ( n65153 , n65148 );
or ( n65154 , n65152 , n65153 );
buf ( n65155 , n42628 );
buf ( n65156 , n64735 );
and ( n65157 , n65155 , n65156 );
buf ( n65158 , n63211 );
not ( n65159 , n65158 );
buf ( n65160 , n42563 );
nor ( n65161 , n65159 , n65160 );
buf ( n65162 , n65161 );
buf ( n65163 , n65162 );
nor ( n65164 , n65157 , n65163 );
buf ( n65165 , n65164 );
not ( n65166 , n65165 );
xor ( n65167 , n63874 , n63895 );
and ( n65168 , n65167 , n63924 );
and ( n65169 , n63874 , n63895 );
or ( n65170 , n65168 , n65169 );
buf ( n65171 , n65170 );
not ( n65172 , n65171 );
or ( n65173 , n65166 , n65172 );
not ( n65174 , n65165 );
buf ( n65175 , n65171 );
not ( n65176 , n65175 );
buf ( n65177 , n65176 );
nand ( n65178 , n65174 , n65177 );
nand ( n65179 , n65173 , n65178 );
buf ( n65180 , n39998 );
not ( n65181 , n65180 );
buf ( n65182 , n64787 );
not ( n65183 , n65182 );
and ( n65184 , n65181 , n65183 );
buf ( n65185 , n63237 );
not ( n65186 , n65185 );
buf ( n65187 , n39980 );
nor ( n65188 , n65186 , n65187 );
buf ( n65189 , n65188 );
buf ( n65190 , n65189 );
nor ( n65191 , n65184 , n65190 );
buf ( n65192 , n65191 );
xnor ( n65193 , n65179 , n65192 );
buf ( n65194 , n65193 );
nand ( n65195 , n65154 , n65194 );
buf ( n65196 , n65195 );
buf ( n65197 , n65196 );
nand ( n65198 , n65151 , n65197 );
buf ( n65199 , n65198 );
buf ( n65200 , n65199 );
not ( n65201 , n65200 );
buf ( n65202 , n65201 );
buf ( n65203 , n65202 );
nand ( n65204 , n65106 , n65203 );
buf ( n65205 , n65204 );
buf ( n65206 , n65205 );
not ( n65207 , n65206 );
buf ( n65208 , n42252 );
not ( n65209 , n65208 );
buf ( n65210 , n59242 );
not ( n65211 , n65210 );
buf ( n65212 , n47836 );
not ( n65213 , n65212 );
or ( n65214 , n65211 , n65213 );
buf ( n65215 , n28411 );
buf ( n65216 , n42260 );
nand ( n65217 , n65215 , n65216 );
buf ( n65218 , n65217 );
buf ( n65219 , n65218 );
nand ( n65220 , n65214 , n65219 );
buf ( n65221 , n65220 );
buf ( n65222 , n65221 );
not ( n65223 , n65222 );
or ( n65224 , n65209 , n65223 );
not ( n65225 , n64810 );
not ( n65226 , n64815 );
or ( n65227 , n65225 , n65226 );
nand ( n65228 , n65227 , n42315 );
buf ( n65229 , n65228 );
nand ( n65230 , n65224 , n65229 );
buf ( n65231 , n65230 );
buf ( n65232 , n65231 );
not ( n65233 , n42374 );
and ( n65234 , n60327 , n63913 );
not ( n65235 , n60327 );
not ( n65236 , n42342 );
and ( n65237 , n65235 , n65236 );
or ( n65238 , n65234 , n65237 );
not ( n65239 , n65238 );
or ( n65240 , n65233 , n65239 );
nand ( n65241 , n63919 , n42336 );
nand ( n65242 , n65240 , n65241 );
buf ( n65243 , n65242 );
and ( n65244 , n29500 , n42556 );
not ( n65245 , n29500 );
and ( n65246 , n65245 , n42560 );
or ( n65247 , n65244 , n65246 );
buf ( n65248 , n65247 );
not ( n65249 , n65248 );
buf ( n65250 , n43935 );
not ( n65251 , n65250 );
or ( n65252 , n65249 , n65251 );
buf ( n65253 , n63939 );
buf ( n65254 , n43905 );
nand ( n65255 , n65253 , n65254 );
buf ( n65256 , n65255 );
buf ( n65257 , n65256 );
nand ( n65258 , n65252 , n65257 );
buf ( n65259 , n65258 );
buf ( n65260 , n65259 );
xor ( n65261 , n65243 , n65260 );
not ( n65262 , n42668 );
not ( n65263 , n64757 );
or ( n65264 , n65262 , n65263 );
and ( n65265 , n29754 , n64753 );
not ( n65266 , n29754 );
and ( n65267 , n65266 , n64748 );
or ( n65268 , n65265 , n65267 );
buf ( n65269 , n65268 );
buf ( n65270 , n58249 );
nand ( n65271 , n65269 , n65270 );
buf ( n65272 , n65271 );
nand ( n65273 , n65264 , n65272 );
buf ( n65274 , n65273 );
and ( n65275 , n65261 , n65274 );
and ( n65276 , n65243 , n65260 );
or ( n65277 , n65275 , n65276 );
buf ( n65278 , n65277 );
buf ( n65279 , n65278 );
or ( n65280 , n65232 , n65279 );
xor ( n65281 , n63951 , n64431 );
xnor ( n65282 , n65281 , n63926 );
buf ( n65283 , n65282 );
nand ( n65284 , n65280 , n65283 );
buf ( n65285 , n65284 );
buf ( n65286 , n65285 );
buf ( n65287 , n65231 );
buf ( n65288 , n65278 );
nand ( n65289 , n65287 , n65288 );
buf ( n65290 , n65289 );
buf ( n65291 , n65290 );
nand ( n65292 , n65286 , n65291 );
buf ( n65293 , n65292 );
buf ( n65294 , n65293 );
buf ( n65295 , n51901 );
not ( n65296 , n65295 );
buf ( n65297 , n52094 );
not ( n65298 , n65297 );
and ( n65299 , n65296 , n65298 );
buf ( n65300 , n51901 );
buf ( n65301 , n52094 );
and ( n65302 , n65300 , n65301 );
nor ( n65303 , n65299 , n65302 );
buf ( n65304 , n65303 );
not ( n65305 , n65304 );
not ( n65306 , n65305 );
not ( n65307 , n37511 );
not ( n65308 , n65307 );
or ( n65309 , n65306 , n65308 );
or ( n65310 , n64586 , n41973 );
nand ( n65311 , n65309 , n65310 );
buf ( n65312 , n65311 );
xor ( n65313 , n65294 , n65312 );
buf ( n65314 , n43798 );
buf ( n65315 , n53548 );
buf ( n65316 , n41947 );
and ( n65317 , n65315 , n65316 );
not ( n65318 , n65315 );
buf ( n65319 , n49879 );
and ( n65320 , n65318 , n65319 );
nor ( n65321 , n65317 , n65320 );
buf ( n65322 , n65321 );
buf ( n65323 , n65322 );
or ( n65324 , n65314 , n65323 );
buf ( n65325 , n37916 );
buf ( n65326 , n64465 );
or ( n65327 , n65325 , n65326 );
nand ( n65328 , n65324 , n65327 );
buf ( n65329 , n65328 );
buf ( n65330 , n65329 );
and ( n65331 , n65313 , n65330 );
and ( n65332 , n65294 , n65312 );
or ( n65333 , n65331 , n65332 );
buf ( n65334 , n65333 );
buf ( n65335 , n65334 );
not ( n65336 , n65335 );
or ( n65337 , n65207 , n65336 );
buf ( n65338 , n65102 );
buf ( n65339 , n65199 );
nand ( n65340 , n65338 , n65339 );
buf ( n65341 , n65340 );
buf ( n65342 , n65341 );
nand ( n65343 , n65337 , n65342 );
buf ( n65344 , n65343 );
buf ( n65345 , n65344 );
nand ( n65346 , n65084 , n65345 );
buf ( n65347 , n65346 );
buf ( n65348 , n65081 );
not ( n65349 , n65348 );
buf ( n65350 , n65059 );
not ( n65351 , n65350 );
buf ( n65352 , n65351 );
buf ( n65353 , n65352 );
nand ( n65354 , n65349 , n65353 );
buf ( n65355 , n65354 );
nand ( n65356 , n65347 , n65355 );
buf ( n65357 , n65356 );
not ( n65358 , n65357 );
xor ( n65359 , n64935 , n64939 );
xor ( n65360 , n65359 , n64953 );
buf ( n65361 , n65360 );
buf ( n65362 , n65361 );
not ( n65363 , n65362 );
or ( n65364 , n65358 , n65363 );
not ( n65365 , n65361 );
nand ( n65366 , n65365 , n65347 , n65355 );
buf ( n65367 , C1 );
buf ( n65368 , n44496 );
not ( n65369 , n65368 );
buf ( n65370 , n63137 );
not ( n65371 , n65370 );
or ( n65372 , n65369 , n65371 );
buf ( n65373 , n65037 );
buf ( n65374 , n44517 );
nand ( n65375 , n65373 , n65374 );
buf ( n65376 , n65375 );
buf ( n65377 , n65376 );
nand ( n65378 , n65372 , n65377 );
buf ( n65379 , n65378 );
not ( n65380 , n65165 );
not ( n65381 , n65177 );
or ( n65382 , n65380 , n65381 );
not ( n65383 , n65174 );
not ( n65384 , n65171 );
or ( n65385 , n65383 , n65384 );
nand ( n65386 , n65385 , n65192 );
nand ( n65387 , n65382 , n65386 );
buf ( n65388 , n65387 );
not ( n65389 , n65388 );
buf ( n65390 , n65389 );
buf ( n65391 , n65390 );
not ( n65392 , n65391 );
buf ( n65393 , n44039 );
not ( n65394 , n65393 );
buf ( n65395 , n64697 );
not ( n65396 , n65395 );
buf ( n65397 , n65396 );
buf ( n65398 , n65397 );
not ( n65399 , n65398 );
and ( n65400 , n65394 , n65399 );
buf ( n65401 , n63186 );
buf ( n65402 , n38381 );
nor ( n65403 , n65401 , n65402 );
buf ( n65404 , n65403 );
buf ( n65405 , n65404 );
nor ( n65406 , n65400 , n65405 );
buf ( n65407 , n65406 );
buf ( n65408 , n65407 );
not ( n65409 , n65408 );
buf ( n65410 , n65409 );
buf ( n65411 , n65410 );
not ( n65412 , n65411 );
or ( n65413 , n65392 , n65412 );
buf ( n65414 , n65387 );
not ( n65415 , n65414 );
buf ( n65416 , n65407 );
not ( n65417 , n65416 );
or ( n65418 , n65415 , n65417 );
xor ( n65419 , n62573 , n63100 );
xor ( n65420 , n65419 , n63104 );
buf ( n65421 , n65420 );
buf ( n65422 , n65421 );
nand ( n65423 , n65418 , n65422 );
buf ( n65424 , n65423 );
buf ( n65425 , n65424 );
nand ( n65426 , n65413 , n65425 );
buf ( n65427 , n65426 );
xor ( n65428 , n65379 , n65427 );
buf ( n65429 , n64628 );
not ( n65430 , n65429 );
buf ( n65431 , n45742 );
nor ( n65432 , n65430 , n65431 );
buf ( n65433 , n65432 );
not ( n65434 , n65433 );
nand ( n65435 , n62224 , n46246 );
nand ( n65436 , n65434 , n65435 );
xnor ( n65437 , n65428 , n65436 );
not ( n65438 , n65437 );
or ( n65439 , n65438 , C0 );
buf ( n65440 , n46912 );
not ( n65441 , n65440 );
buf ( n65442 , n64866 );
not ( n65443 , n65442 );
or ( n65444 , n65441 , n65443 );
buf ( n65445 , n51622 );
not ( n65446 , n65445 );
buf ( n65447 , n47119 );
not ( n65448 , n65447 );
or ( n65449 , n65446 , n65448 );
buf ( n65450 , n39205 );
buf ( n65451 , n46890 );
nand ( n65452 , n65450 , n65451 );
buf ( n65453 , n65452 );
buf ( n65454 , n65453 );
nand ( n65455 , n65449 , n65454 );
buf ( n65456 , n65455 );
buf ( n65457 , n65456 );
buf ( n65458 , n47331 );
nand ( n65459 , n65457 , n65458 );
buf ( n65460 , n65459 );
buf ( n65461 , n65460 );
nand ( n65462 , n65444 , n65461 );
buf ( n65463 , n65462 );
buf ( n65464 , n65463 );
buf ( n65465 , n55841 );
not ( n65466 , n65465 );
buf ( n65467 , n38068 );
not ( n65468 , n65467 );
or ( n65469 , n65466 , n65468 );
buf ( n65470 , n49391 );
buf ( n65471 , n58361 );
nand ( n65472 , n65470 , n65471 );
buf ( n65473 , n65472 );
buf ( n65474 , n65473 );
nand ( n65475 , n65469 , n65474 );
buf ( n65476 , n65475 );
buf ( n65477 , n65476 );
not ( n65478 , n65477 );
buf ( n65479 , n46165 );
not ( n65480 , n65479 );
or ( n65481 , n65478 , n65480 );
buf ( n65482 , n64974 );
buf ( n65483 , n43414 );
nand ( n65484 , n65482 , n65483 );
buf ( n65485 , n65484 );
buf ( n65486 , n65485 );
nand ( n65487 , n65481 , n65486 );
buf ( n65488 , n65487 );
buf ( n65489 , n65488 );
or ( n65490 , n65464 , n65489 );
buf ( n65491 , n65421 );
buf ( n65492 , n65390 );
xor ( n65493 , n65491 , n65492 );
buf ( n65494 , n65410 );
xor ( n65495 , n65493 , n65494 );
buf ( n65496 , n65495 );
buf ( n65497 , n65496 );
nand ( n65498 , n65490 , n65497 );
buf ( n65499 , n65498 );
buf ( n65500 , n65499 );
buf ( n65501 , n65463 );
buf ( n65502 , n65488 );
nand ( n65503 , n65501 , n65502 );
buf ( n65504 , n65503 );
buf ( n65505 , n65504 );
nand ( n65506 , n65500 , n65505 );
buf ( n65507 , n65506 );
nand ( n65508 , n65439 , n65507 );
nand ( n65509 , C1 , n65508 );
nand ( n65510 , n65366 , n65509 );
buf ( n65511 , n65510 );
nand ( n65512 , n65364 , n65511 );
buf ( n65513 , n65512 );
buf ( n65514 , n65513 );
xor ( n65515 , n64961 , n65514 );
xor ( n65516 , n63123 , n63148 );
xor ( n65517 , n65516 , n63294 );
buf ( n65518 , n65517 );
buf ( n65519 , n65518 );
not ( n65520 , n65379 );
not ( n65521 , n65427 );
or ( n65522 , n65520 , n65521 );
nor ( n65523 , n65427 , n65379 );
not ( n65524 , n65436 );
or ( n65525 , n65523 , n65524 );
nand ( n65526 , n65522 , n65525 );
buf ( n65527 , n65526 );
xor ( n65528 , n65519 , n65527 );
not ( n65529 , n64981 );
buf ( n65530 , n65529 );
not ( n65531 , n65530 );
buf ( n65532 , n65057 );
not ( n65533 , n65532 );
or ( n65534 , n65531 , n65533 );
not ( n65535 , n64990 );
not ( n65536 , n65050 );
or ( n65537 , n65535 , n65536 );
nand ( n65538 , n65537 , n65053 );
buf ( n65539 , n65538 );
nand ( n65540 , n65534 , n65539 );
buf ( n65541 , n65540 );
buf ( n65542 , n65541 );
buf ( n65543 , n65058 );
buf ( n65544 , n64981 );
nand ( n65545 , n65543 , n65544 );
buf ( n65546 , n65545 );
buf ( n65547 , n65546 );
nand ( n65548 , n65542 , n65547 );
buf ( n65549 , n65548 );
buf ( n65550 , n65549 );
and ( n65551 , n65528 , n65550 );
and ( n65552 , n65519 , n65527 );
or ( n65553 , n65551 , n65552 );
buf ( n65554 , n65553 );
buf ( n65555 , n65554 );
not ( n65556 , n65555 );
buf ( n65557 , C1 );
or ( n65558 , n65556 , C0 );
nand ( n65559 , n65558 , C1 );
buf ( n65560 , n65559 );
buf ( n65561 , n65560 );
xor ( n65562 , n62376 , n62438 );
and ( n65563 , n65562 , n62447 );
not ( n65564 , n65562 );
and ( n65565 , n65564 , n62361 );
nor ( n65566 , n65563 , n65565 );
buf ( n65567 , n65566 );
not ( n65568 , n65567 );
buf ( n65569 , n65568 );
buf ( n65570 , n65569 );
and ( n65571 , n65561 , n65570 );
not ( n65572 , n65561 );
buf ( n65573 , n65566 );
and ( n65574 , n65572 , n65573 );
nor ( n65575 , n65571 , n65574 );
buf ( n65576 , n65575 );
buf ( n65577 , n65576 );
and ( n65578 , n65515 , n65577 );
and ( n65579 , n64961 , n65514 );
or ( n65580 , n65578 , n65579 );
buf ( n65581 , n65580 );
buf ( n65582 , n65581 );
xor ( n65583 , n64918 , n65582 );
buf ( n65584 , n65583 );
buf ( n65585 , n65584 );
xor ( n65586 , n64612 , n64904 );
xor ( n65587 , n65586 , n64912 );
buf ( n65588 , n65587 );
buf ( n65589 , n65588 );
xor ( n65590 , n64961 , n65514 );
xor ( n65591 , n65590 , n65577 );
buf ( n65592 , n65591 );
buf ( n65593 , n65592 );
xor ( n65594 , n65589 , n65593 );
buf ( n65595 , n62174 );
buf ( n65596 , n62141 );
xor ( n65597 , n65595 , n65596 );
buf ( n65598 , n62277 );
xor ( n65599 , n65597 , n65598 );
buf ( n65600 , n65599 );
buf ( n65601 , n65600 );
buf ( n65602 , C0 );
buf ( n65603 , n51488 );
not ( n65604 , n65603 );
buf ( n65605 , n65069 );
not ( n65606 , n65605 );
or ( n65607 , n65604 , n65606 );
buf ( n65608 , n62131 );
buf ( n65609 , n62125 );
nand ( n65610 , n65608 , n65609 );
buf ( n65611 , n65610 );
buf ( n65612 , n65611 );
nand ( n65613 , n65607 , n65612 );
buf ( n65614 , n65613 );
buf ( n65615 , n65614 );
buf ( n65616 , n65602 );
or ( n65617 , n65615 , n65616 );
xor ( n65618 , n62210 , n62247 );
xor ( n65619 , n65618 , n62273 );
buf ( n65620 , n65619 );
buf ( n65621 , n65620 );
nand ( n65622 , n65617 , n65621 );
buf ( n65623 , n65622 );
buf ( n65624 , n65623 );
nand ( n65625 , C1 , n65624 );
buf ( n65626 , n65625 );
buf ( n65627 , n65626 );
xor ( n65628 , n65601 , n65627 );
buf ( n65629 , n65628 );
buf ( n65630 , n65629 );
xor ( n65631 , n63299 , n63303 );
xor ( n65632 , n65631 , n63357 );
buf ( n65633 , n65632 );
buf ( n65634 , n65633 );
xor ( n65635 , n65630 , n65634 );
buf ( n65636 , n65635 );
buf ( n65637 , n65636 );
xor ( n65638 , n65519 , n65527 );
xor ( n65639 , n65638 , n65550 );
buf ( n65640 , n65639 );
buf ( n65641 , n65640 );
buf ( n65642 , n51488 );
not ( n65643 , n65642 );
buf ( n65644 , n51493 );
buf ( n65645 , n37708 );
and ( n65646 , n65644 , n65645 );
not ( n65647 , n65644 );
buf ( n65648 , n37711 );
and ( n65649 , n65647 , n65648 );
nor ( n65650 , n65646 , n65649 );
buf ( n65651 , n65650 );
buf ( n65652 , n65651 );
not ( n65653 , n65652 );
or ( n65654 , n65643 , n65653 );
nand ( n65655 , n65076 , n52456 );
buf ( n65656 , n65655 );
nand ( n65657 , n65654 , n65656 );
buf ( n65658 , n65657 );
not ( n65659 , n65658 );
buf ( n65660 , n62155 );
buf ( n65661 , n37786 );
and ( n65662 , n65660 , n65661 );
not ( n65663 , n65660 );
buf ( n65664 , n59203 );
and ( n65665 , n65663 , n65664 );
nor ( n65666 , n65662 , n65665 );
buf ( n65667 , n65666 );
not ( n65668 , n65667 );
not ( n65669 , n48858 );
and ( n65670 , n65668 , n65669 );
and ( n65671 , n64564 , n48868 );
nor ( n65672 , n65670 , n65671 );
buf ( n65673 , n65672 );
not ( n65674 , n65673 );
buf ( n65675 , n65674 );
not ( n65676 , n65675 );
or ( n65677 , n65659 , n65676 );
buf ( n65678 , n65658 );
buf ( n65679 , n65675 );
nor ( n65680 , n65678 , n65679 );
buf ( n65681 , n65680 );
buf ( n65682 , n46246 );
not ( n65683 , n65682 );
buf ( n65684 , n64634 );
not ( n65685 , n65684 );
or ( n65686 , n65683 , n65685 );
buf ( n65687 , n64616 );
not ( n65688 , n65687 );
buf ( n65689 , n50040 );
not ( n65690 , n65689 );
or ( n65691 , n65688 , n65690 );
buf ( n65692 , n50043 );
buf ( n65693 , n45747 );
nand ( n65694 , n65692 , n65693 );
buf ( n65695 , n65694 );
buf ( n65696 , n65695 );
nand ( n65697 , n65691 , n65696 );
buf ( n65698 , n65697 );
buf ( n65699 , n65698 );
buf ( n65700 , n46225 );
nand ( n65701 , n65699 , n65700 );
buf ( n65702 , n65701 );
buf ( n65703 , n65702 );
nand ( n65704 , n65686 , n65703 );
buf ( n65705 , n65704 );
buf ( n65706 , n65705 );
not ( n65707 , n65706 );
buf ( n65708 , n65707 );
not ( n65709 , n65708 );
and ( n65710 , n64441 , n63846 );
not ( n65711 , n64441 );
and ( n65712 , n65711 , n63845 );
or ( n65713 , n65710 , n65712 );
xor ( n65714 , n63866 , n65713 );
not ( n65715 , n65714 );
and ( n65716 , n65709 , n65715 );
xor ( n65717 , n64803 , n64822 );
xnor ( n65718 , n65717 , n64840 );
buf ( n65719 , n65708 );
buf ( n65720 , n65714 );
nand ( n65721 , n65719 , n65720 );
buf ( n65722 , n65721 );
and ( n65723 , n65718 , n65722 );
nor ( n65724 , n65716 , n65723 );
or ( n65725 , n65681 , n65724 );
nand ( n65726 , n65677 , n65725 );
buf ( n65727 , n65726 );
xor ( n65728 , n63780 , n63801 );
xor ( n65729 , n65728 , n64498 );
buf ( n65730 , n65729 );
buf ( n65731 , n65730 );
buf ( n65732 , C0 );
buf ( n65733 , n65732 );
and ( n65734 , n65727 , n65731 );
or ( n65735 , C0 , n65734 );
buf ( n65736 , n65735 );
buf ( n65737 , n65736 );
xor ( n65738 , n65641 , n65737 );
xor ( n65739 , n63776 , n64503 );
xor ( n65740 , n65739 , n64607 );
buf ( n65741 , n65740 );
buf ( n65742 , n65741 );
and ( n65743 , n65738 , n65742 );
and ( n65744 , n65641 , n65737 );
or ( n65745 , n65743 , n65744 );
buf ( n65746 , n65745 );
buf ( n65747 , n65746 );
xor ( n65748 , n65637 , n65747 );
buf ( n65749 , n65620 );
not ( n65750 , n65749 );
buf ( n65751 , n65750 );
buf ( n65752 , n65751 );
not ( n65753 , n65752 );
xor ( n65754 , n65602 , n65614 );
buf ( n65755 , n65754 );
not ( n65756 , n65755 );
or ( n65757 , n65753 , n65756 );
buf ( n65758 , n65754 );
buf ( n65759 , n65751 );
or ( n65760 , n65758 , n65759 );
nand ( n65761 , n65757 , n65760 );
buf ( n65762 , n65761 );
buf ( n65763 , n65762 );
xor ( n65764 , n64614 , n64895 );
xor ( n65765 , n65764 , n64900 );
buf ( n65766 , n65765 );
buf ( n65767 , n65766 );
xor ( n65768 , n65763 , n65767 );
xor ( n65769 , n63827 , n64454 );
xor ( n65770 , n65769 , n64493 );
buf ( n65771 , n65770 );
not ( n65772 , n65771 );
buf ( n65773 , C0 );
xor ( n65774 , n64579 , n64590 );
xor ( n65775 , n65774 , n64596 );
buf ( n65776 , n65775 );
buf ( n65777 , n65776 );
or ( n65778 , n65773 , n65777 );
buf ( n65779 , n65778 );
not ( n65780 , n65779 );
or ( n65781 , n65772 , n65780 );
buf ( n65782 , C0 );
nand ( n65783 , n65781 , C1 );
not ( n65784 , n65783 );
or ( n65785 , n64569 , n64548 );
nand ( n65786 , n64548 , n64569 );
nand ( n65787 , n65785 , n65786 );
and ( n65788 , n65787 , n64600 );
not ( n65789 , n65787 );
not ( n65790 , n64600 );
and ( n65791 , n65789 , n65790 );
nor ( n65792 , n65788 , n65791 );
not ( n65793 , n65792 );
not ( n65794 , n65793 );
or ( n65795 , n65784 , n65794 );
not ( n65796 , n65792 );
and ( n65797 , n65779 , n65771 );
nor ( n65798 , n65797 , n65782 );
not ( n65799 , n65798 );
or ( n65800 , n65796 , n65799 );
not ( n65801 , n64873 );
not ( n65802 , n65801 );
and ( n65803 , n64888 , n65802 );
not ( n65804 , n64888 );
and ( n65805 , n65804 , n65801 );
nor ( n65806 , n65803 , n65805 );
buf ( n65807 , n64855 );
buf ( n65808 , n65807 );
buf ( n65809 , n65808 );
and ( n65810 , n65806 , n65809 );
not ( n65811 , n65806 );
not ( n65812 , n65809 );
and ( n65813 , n65811 , n65812 );
nor ( n65814 , n65810 , n65813 );
nand ( n65815 , n65800 , n65814 );
nand ( n65816 , n65795 , n65815 );
buf ( n65817 , n65816 );
and ( n65818 , n65768 , n65817 );
and ( n65819 , n65763 , n65767 );
or ( n65820 , n65818 , n65819 );
buf ( n65821 , n65820 );
buf ( n65822 , n65821 );
xor ( n65823 , n65748 , n65822 );
buf ( n65824 , n65823 );
buf ( n65825 , n65824 );
and ( n65826 , n65594 , n65825 );
and ( n65827 , n65589 , n65593 );
or ( n65828 , n65826 , n65827 );
buf ( n65829 , n65828 );
buf ( n65830 , n65829 );
xor ( n65831 , n65585 , n65830 );
buf ( n65832 , n62488 );
buf ( n65833 , C0 );
xor ( n65834 , n65832 , n65833 );
buf ( n65835 , n62453 );
xnor ( n65836 , n65834 , n65835 );
buf ( n65837 , n65836 );
buf ( n65838 , n65837 );
not ( n65839 , n65838 );
buf ( n65840 , n65839 );
not ( n65841 , n65840 );
xor ( n65842 , n64927 , n64929 );
and ( n65843 , n65842 , n64958 );
or ( n65844 , n65843 , C0 );
buf ( n65845 , n65844 );
not ( n65846 , n65845 );
not ( n65847 , n65846 );
or ( n65848 , n65841 , n65847 );
nand ( n65849 , n65845 , n65837 );
nand ( n65850 , n65848 , n65849 );
buf ( n65851 , n65557 );
buf ( n65852 , n65566 );
nand ( n65853 , n65851 , n65852 );
buf ( n65854 , n65853 );
and ( n65855 , n65854 , n65554 );
nor ( n65856 , C0 , n65855 );
buf ( n65857 , n65856 );
buf ( n65858 , n65857 );
buf ( n65859 , n65858 );
buf ( n65860 , n65859 );
not ( n65861 , n65860 );
buf ( n65862 , n65861 );
and ( n65863 , n65850 , n65862 );
not ( n65864 , n65850 );
and ( n65865 , n65864 , n65859 );
nor ( n65866 , n65863 , n65865 );
or ( n65867 , n65626 , n65600 );
and ( n65868 , n65867 , n65633 );
and ( n65869 , n65601 , n65627 );
buf ( n65870 , n65869 );
nor ( n65871 , n65868 , n65870 );
buf ( n65872 , n65871 );
not ( n65873 , n65872 );
xor ( n65874 , n62284 , n62288 );
xor ( n65875 , n65874 , n62293 );
buf ( n65876 , n65875 );
not ( n65877 , n65876 );
not ( n65878 , n65877 );
buf ( n65879 , n62496 );
buf ( n65880 , n62497 );
xor ( n65881 , n65879 , n65880 );
buf ( n65882 , n63361 );
xnor ( n65883 , n65881 , n65882 );
buf ( n65884 , n65883 );
buf ( n65885 , n65884 );
not ( n65886 , n65885 );
buf ( n65887 , n65886 );
not ( n65888 , n65887 );
or ( n65889 , n65878 , n65888 );
buf ( n65890 , n65876 );
buf ( n65891 , n65884 );
nand ( n65892 , n65890 , n65891 );
buf ( n65893 , n65892 );
nand ( n65894 , n65889 , n65893 );
not ( n65895 , n65894 );
or ( n65896 , n65873 , n65895 );
or ( n65897 , n65872 , n65894 );
nand ( n65898 , n65896 , n65897 );
xor ( n65899 , n65866 , n65898 );
xor ( n65900 , n65637 , n65747 );
and ( n65901 , n65900 , n65822 );
and ( n65902 , n65637 , n65747 );
or ( n65903 , n65901 , n65902 );
buf ( n65904 , n65903 );
xor ( n65905 , n65899 , n65904 );
buf ( n65906 , n65905 );
and ( n65907 , n65831 , n65906 );
and ( n65908 , n65585 , n65830 );
or ( n65909 , n65907 , n65908 );
buf ( n65910 , n65909 );
not ( n65911 , n65910 );
not ( n65912 , n65911 );
xor ( n65913 , n63772 , n64917 );
and ( n65914 , n65913 , n65582 );
and ( n65915 , n63772 , n64917 );
or ( n65916 , n65914 , n65915 );
buf ( n65917 , n65916 );
buf ( n65918 , n65917 );
xor ( n65919 , n65866 , n65898 );
and ( n65920 , n65919 , n65904 );
and ( n65921 , n65866 , n65898 );
or ( n65922 , n65920 , n65921 );
buf ( n65923 , n65922 );
xor ( n65924 , n65918 , n65923 );
xor ( n65925 , n62355 , n62492 );
xor ( n65926 , n65925 , n63365 );
buf ( n65927 , n65926 );
not ( n65928 , n65856 );
not ( n65929 , n65928 );
not ( n65930 , n65840 );
or ( n65931 , n65929 , n65930 );
not ( n65932 , n65837 );
not ( n65933 , n65856 );
or ( n65934 , n65932 , n65933 );
nand ( n65935 , n65934 , n65845 );
nand ( n65936 , n65931 , n65935 );
buf ( n65937 , n65936 );
and ( n65938 , n65927 , n65937 );
not ( n65939 , n65927 );
buf ( n65940 , n65936 );
not ( n65941 , n65940 );
buf ( n65942 , n65941 );
buf ( n65943 , n65942 );
and ( n65944 , n65939 , n65943 );
nor ( n65945 , n65938 , n65944 );
buf ( n65946 , n65945 );
buf ( n65947 , n65877 );
not ( n65948 , n65947 );
buf ( n65949 , n65871 );
not ( n65950 , n65949 );
or ( n65951 , n65948 , n65950 );
buf ( n65952 , n65887 );
nand ( n65953 , n65951 , n65952 );
buf ( n65954 , n65953 );
buf ( n65955 , n65871 );
not ( n65956 , n65955 );
not ( n65957 , n65877 );
buf ( n65958 , n65957 );
nand ( n65959 , n65956 , n65958 );
buf ( n65960 , n65959 );
nand ( n65961 , n65954 , n65960 );
xor ( n65962 , n65946 , n65961 );
buf ( n65963 , n62121 );
buf ( n65964 , n62300 );
xor ( n65965 , n65963 , n65964 );
buf ( n65966 , n62114 );
xnor ( n65967 , n65965 , n65966 );
buf ( n65968 , n65967 );
xor ( n65969 , n61551 , n61553 );
xor ( n65970 , n65969 , n61555 );
buf ( n65971 , n65970 );
buf ( n65972 , n65971 );
buf ( n65973 , n63526 );
not ( n65974 , n65973 );
buf ( n65975 , n63770 );
not ( n65976 , n65975 );
or ( n65977 , n65974 , n65976 );
buf ( n65978 , n63770 );
buf ( n65979 , n63526 );
or ( n65980 , n65978 , n65979 );
buf ( n65981 , n63767 );
nand ( n65982 , n65980 , n65981 );
buf ( n65983 , n65982 );
buf ( n65984 , n65983 );
nand ( n65985 , n65977 , n65984 );
buf ( n65986 , n65985 );
buf ( n65987 , n65986 );
xor ( n65988 , n65972 , n65987 );
xor ( n65989 , n63384 , n63388 );
xor ( n65990 , n65989 , n63433 );
buf ( n65991 , n65990 );
buf ( n65992 , n65991 );
xnor ( n65993 , n65988 , n65992 );
buf ( n65994 , n65993 );
buf ( n65995 , n65994 );
not ( n65996 , n65995 );
buf ( n65997 , n65996 );
and ( n65998 , n65968 , n65997 );
not ( n65999 , n65968 );
and ( n66000 , n65999 , n65994 );
or ( n66001 , n65998 , n66000 );
xor ( n66002 , n65962 , n66001 );
buf ( n66003 , n66002 );
xor ( n66004 , n65924 , n66003 );
buf ( n66005 , n66004 );
not ( n66006 , n66005 );
not ( n66007 , n66006 );
and ( n66008 , n65912 , n66007 );
not ( n66009 , n62326 );
not ( n66010 , n62332 );
not ( n66011 , n66010 );
or ( n66012 , n66009 , n66011 );
nand ( n66013 , n62312 , n62325 );
nand ( n66014 , n66012 , n66013 );
buf ( n66015 , n66014 );
buf ( n66016 , n62347 );
not ( n66017 , n66016 );
buf ( n66018 , n66017 );
buf ( n66019 , n66018 );
and ( n66020 , n66015 , n66019 );
not ( n66021 , n66015 );
buf ( n66022 , n62347 );
buf ( n66023 , n66022 );
and ( n66024 , n66021 , n66023 );
nor ( n66025 , n66020 , n66024 );
buf ( n66026 , n66025 );
buf ( n66027 , n66026 );
not ( n66028 , n65997 );
xor ( n66029 , n62121 , n62300 );
xor ( n66030 , n66029 , n62114 );
not ( n66031 , n66030 );
and ( n66032 , n66028 , n66031 );
buf ( n66033 , n65997 );
buf ( n66034 , n66030 );
nand ( n66035 , n66033 , n66034 );
buf ( n66036 , n66035 );
and ( n66037 , n66036 , n65962 );
nor ( n66038 , n66032 , n66037 );
buf ( n66039 , n66038 );
xor ( n66040 , n66027 , n66039 );
buf ( n66041 , n65971 );
not ( n66042 , n66041 );
buf ( n66043 , n65991 );
not ( n66044 , n66043 );
buf ( n66045 , n66044 );
buf ( n66046 , n66045 );
not ( n66047 , n66046 );
or ( n66048 , n66042 , n66047 );
buf ( n66049 , n65986 );
nand ( n66050 , n66048 , n66049 );
buf ( n66051 , n66050 );
buf ( n66052 , n66051 );
buf ( n66053 , n65971 );
not ( n66054 , n66053 );
buf ( n66055 , n65991 );
nand ( n66056 , n66054 , n66055 );
buf ( n66057 , n66056 );
buf ( n66058 , n66057 );
and ( n66059 , n66052 , n66058 );
buf ( n66060 , n66059 );
buf ( n66061 , n66060 );
and ( n66062 , n63437 , n63451 );
not ( n66063 , n63437 );
and ( n66064 , n66063 , n63448 );
nor ( n66065 , n66062 , n66064 );
xor ( n66066 , n63368 , n66065 );
buf ( n66067 , n66066 );
xor ( n66068 , n66061 , n66067 );
not ( n66069 , n65961 );
not ( n66070 , n66069 );
buf ( n66071 , n65942 );
buf ( n66072 , n66071 );
buf ( n66073 , n66072 );
not ( n66074 , n66073 );
and ( n66075 , n66070 , n66074 );
nand ( n66076 , n66073 , n66069 );
buf ( n66077 , n65926 );
buf ( n66078 , n66077 );
buf ( n66079 , n66078 );
and ( n66080 , n66076 , n66079 );
nor ( n66081 , n66075 , n66080 );
buf ( n66082 , n66081 );
xor ( n66083 , n66068 , n66082 );
buf ( n66084 , n66083 );
buf ( n66085 , n66084 );
xor ( n66086 , n66040 , n66085 );
buf ( n66087 , n66086 );
not ( n66088 , n66087 );
xor ( n66089 , n65918 , n65923 );
and ( n66090 , n66089 , n66003 );
and ( n66091 , n65918 , n65923 );
or ( n66092 , n66090 , n66091 );
buf ( n66093 , n66092 );
and ( n66094 , n66088 , n66093 );
nor ( n66095 , n66008 , n66094 );
not ( n66096 , n62015 );
not ( n66097 , n62024 );
not ( n66098 , n66097 );
or ( n66099 , n66096 , n66098 );
nand ( n66100 , n62024 , n62014 );
nand ( n66101 , n66099 , n66100 );
and ( n66102 , n66101 , n61609 );
not ( n66103 , n66101 );
and ( n66104 , n66103 , n61610 );
nor ( n66105 , n66102 , n66104 );
buf ( n66106 , n66105 );
xor ( n66107 , n66061 , n66067 );
and ( n66108 , n66107 , n66082 );
and ( n66109 , n66061 , n66067 );
or ( n66110 , n66108 , n66109 );
buf ( n66111 , n66110 );
buf ( n66112 , n66111 );
xor ( n66113 , n66106 , n66112 );
xor ( n66114 , n63464 , n62106 );
xnor ( n66115 , n66114 , n62349 );
buf ( n66116 , n66115 );
xor ( n66117 , n66113 , n66116 );
buf ( n66118 , n66117 );
buf ( n66119 , n66118 );
not ( n66120 , n66119 );
buf ( n66121 , n66120 );
xor ( n66122 , n66027 , n66039 );
and ( n66123 , n66122 , n66085 );
and ( n66124 , n66027 , n66039 );
or ( n66125 , n66123 , n66124 );
buf ( n66126 , n66125 );
buf ( n66127 , n66126 );
not ( n66128 , n66127 );
buf ( n66129 , n66128 );
nand ( n66130 , n66121 , n66129 );
xor ( n66131 , n65585 , n65830 );
xor ( n66132 , n66131 , n65906 );
buf ( n66133 , n66132 );
not ( n66134 , n42408 );
not ( n66135 , n48320 );
or ( n66136 , n66134 , n66135 );
nand ( n66137 , n42403 , n48323 );
nand ( n66138 , n66136 , n66137 );
not ( n66139 , n66138 );
and ( n66140 , n38402 , n38400 );
not ( n66141 , n66140 );
or ( n66142 , n66139 , n66141 );
not ( n66143 , n38402 );
nand ( n66144 , n66143 , n64682 );
nand ( n66145 , n66142 , n66144 );
buf ( n66146 , n66145 );
buf ( n66147 , n38051 );
buf ( n66148 , n56325 );
nor ( n66149 , n66147 , n66148 );
buf ( n66150 , n66149 );
buf ( n66151 , n66150 );
xor ( n66152 , n66146 , n66151 );
not ( n66153 , n44517 );
buf ( n66154 , n65010 );
not ( n66155 , n66154 );
buf ( n66156 , n42119 );
not ( n66157 , n66156 );
or ( n66158 , n66155 , n66157 );
buf ( n66159 , n28305 );
buf ( n66160 , n44530 );
nand ( n66161 , n66159 , n66160 );
buf ( n66162 , n66161 );
buf ( n66163 , n66162 );
nand ( n66164 , n66158 , n66163 );
buf ( n66165 , n66164 );
not ( n66166 , n66165 );
or ( n66167 , n66153 , n66166 );
nand ( n66168 , n65121 , n44496 );
nand ( n66169 , n66167 , n66168 );
buf ( n66170 , n66169 );
and ( n66171 , n66152 , n66170 );
and ( n66172 , n66146 , n66151 );
or ( n66173 , n66171 , n66172 );
buf ( n66174 , n66173 );
buf ( n66175 , n66174 );
buf ( n66176 , n46390 );
not ( n66177 , n66176 );
buf ( n66178 , n47031 );
not ( n66179 , n66178 );
or ( n66180 , n66177 , n66179 );
buf ( n66181 , n38979 );
buf ( n66182 , n46393 );
nand ( n66183 , n66181 , n66182 );
buf ( n66184 , n66183 );
buf ( n66185 , n66184 );
nand ( n66186 , n66180 , n66185 );
buf ( n66187 , n66186 );
buf ( n66188 , n66187 );
not ( n66189 , n66188 );
buf ( n66190 , n47050 );
not ( n66191 , n66190 );
or ( n66192 , n66189 , n66191 );
buf ( n66193 , n63863 );
buf ( n66194 , n42448 );
nand ( n66195 , n66193 , n66194 );
buf ( n66196 , n66195 );
buf ( n66197 , n66196 );
nand ( n66198 , n66192 , n66197 );
buf ( n66199 , n66198 );
buf ( n66200 , n66199 );
buf ( n66201 , n44267 );
not ( n66202 , n66201 );
buf ( n66203 , n41605 );
not ( n66204 , n66203 );
buf ( n66205 , n41915 );
not ( n66206 , n66205 );
or ( n66207 , n66204 , n66206 );
buf ( n66208 , n51798 );
not ( n66209 , n66208 );
buf ( n66210 , n41604 );
nand ( n66211 , n66209 , n66210 );
buf ( n66212 , n66211 );
buf ( n66213 , n66212 );
nand ( n66214 , n66207 , n66213 );
buf ( n66215 , n66214 );
buf ( n66216 , n66215 );
not ( n66217 , n66216 );
or ( n66218 , n66202 , n66217 );
buf ( n66219 , n64668 );
buf ( n66220 , n43868 );
nand ( n66221 , n66219 , n66220 );
buf ( n66222 , n66221 );
buf ( n66223 , n66222 );
nand ( n66224 , n66218 , n66223 );
buf ( n66225 , n66224 );
buf ( n66226 , n66225 );
xor ( n66227 , n66200 , n66226 );
buf ( n66228 , n42847 );
not ( n66229 , n66228 );
buf ( n66230 , n52670 );
not ( n66231 , n66230 );
or ( n66232 , n66229 , n66231 );
buf ( n66233 , n25159 );
buf ( n66234 , n46691 );
nand ( n66235 , n66233 , n66234 );
buf ( n66236 , n66235 );
buf ( n66237 , n66236 );
nand ( n66238 , n66232 , n66237 );
buf ( n66239 , n66238 );
buf ( n66240 , n66239 );
not ( n66241 , n66240 );
buf ( n66242 , n50128 );
not ( n66243 , n66242 );
or ( n66244 , n66241 , n66243 );
buf ( n66245 , n64717 );
buf ( n66246 , n42564 );
nand ( n66247 , n66245 , n66246 );
buf ( n66248 , n66247 );
buf ( n66249 , n66248 );
nand ( n66250 , n66244 , n66249 );
buf ( n66251 , n66250 );
buf ( n66252 , n66251 );
buf ( n66253 , n46117 );
not ( n66254 , n66253 );
buf ( n66255 , n50599 );
not ( n66256 , n66255 );
or ( n66257 , n66254 , n66256 );
buf ( n66258 , n50591 );
buf ( n66259 , n46126 );
nand ( n66260 , n66258 , n66259 );
buf ( n66261 , n66260 );
buf ( n66262 , n66261 );
nand ( n66263 , n66257 , n66262 );
buf ( n66264 , n66263 );
buf ( n66265 , n66264 );
not ( n66266 , n66265 );
buf ( n66267 , n52537 );
not ( n66268 , n66267 );
or ( n66269 , n66266 , n66268 );
nand ( n66270 , n64773 , n48975 );
buf ( n66271 , n66270 );
nand ( n66272 , n66269 , n66271 );
buf ( n66273 , n66272 );
buf ( n66274 , n66273 );
xor ( n66275 , n66252 , n66274 );
buf ( n66276 , n65221 );
not ( n66277 , n66276 );
buf ( n66278 , n66277 );
buf ( n66279 , n66278 );
buf ( n66280 , n42312 );
or ( n66281 , n66279 , n66280 );
buf ( n66282 , n59242 );
not ( n66283 , n66282 );
buf ( n66284 , n43362 );
not ( n66285 , n66284 );
or ( n66286 , n66283 , n66285 );
buf ( n66287 , n29407 );
buf ( n66288 , n42260 );
nand ( n66289 , n66287 , n66288 );
buf ( n66290 , n66289 );
buf ( n66291 , n66290 );
nand ( n66292 , n66286 , n66291 );
buf ( n66293 , n66292 );
buf ( n66294 , n66293 );
buf ( n66295 , n42252 );
nand ( n66296 , n66294 , n66295 );
buf ( n66297 , n66296 );
buf ( n66298 , n66297 );
nand ( n66299 , n66281 , n66298 );
buf ( n66300 , n66299 );
buf ( n66301 , n66300 );
and ( n66302 , n66275 , n66301 );
and ( n66303 , n66252 , n66274 );
or ( n66304 , n66302 , n66303 );
buf ( n66305 , n66304 );
buf ( n66306 , n66305 );
and ( n66307 , n66227 , n66306 );
and ( n66308 , n66200 , n66226 );
or ( n66309 , n66307 , n66308 );
buf ( n66310 , n66309 );
buf ( n66311 , n66310 );
xor ( n66312 , n66175 , n66311 );
buf ( n66313 , n46912 );
not ( n66314 , n66313 );
buf ( n66315 , n65456 );
not ( n66316 , n66315 );
or ( n66317 , n66314 , n66316 );
buf ( n66318 , n46875 );
not ( n66319 , n66318 );
buf ( n66320 , n42899 );
not ( n66321 , n66320 );
or ( n66322 , n66319 , n66321 );
buf ( n66323 , n42458 );
buf ( n66324 , n46887 );
nand ( n66325 , n66323 , n66324 );
buf ( n66326 , n66325 );
buf ( n66327 , n66326 );
nand ( n66328 , n66322 , n66327 );
buf ( n66329 , n66328 );
buf ( n66330 , n66329 );
buf ( n66331 , n47331 );
nand ( n66332 , n66330 , n66331 );
buf ( n66333 , n66332 );
buf ( n66334 , n66333 );
nand ( n66335 , n66317 , n66334 );
buf ( n66336 , n66335 );
buf ( n66337 , n66336 );
and ( n66338 , n66312 , n66337 );
and ( n66339 , n66175 , n66311 );
or ( n66340 , n66338 , n66339 );
buf ( n66341 , n66340 );
not ( n66342 , n64636 );
not ( n66343 , n64844 );
or ( n66344 , n66342 , n66343 );
or ( n66345 , n64844 , n64636 );
nand ( n66346 , n66344 , n66345 );
and ( n66347 , n66346 , n64850 );
not ( n66348 , n66346 );
and ( n66349 , n66348 , n64797 );
or ( n66350 , n66347 , n66349 );
xor ( n66351 , n66341 , n66350 );
buf ( n66352 , n12481 );
not ( n66353 , n66352 );
buf ( n66354 , n47898 );
not ( n66355 , n66354 );
or ( n66356 , n66353 , n66355 );
buf ( n66357 , n49391 );
buf ( n66358 , n56325 );
nand ( n66359 , n66357 , n66358 );
buf ( n66360 , n66359 );
buf ( n66361 , n66360 );
nand ( n66362 , n66356 , n66361 );
buf ( n66363 , n66362 );
buf ( n66364 , n66363 );
not ( n66365 , n66364 );
buf ( n66366 , n46165 );
not ( n66367 , n66366 );
or ( n66368 , n66365 , n66367 );
buf ( n66369 , n47108 );
buf ( n66370 , n65476 );
nand ( n66371 , n66369 , n66370 );
buf ( n66372 , n66371 );
buf ( n66373 , n66372 );
nand ( n66374 , n66368 , n66373 );
buf ( n66375 , n66374 );
buf ( n66376 , n66375 );
buf ( n66377 , n64702 );
buf ( n66378 , n64791 );
xor ( n66379 , n66377 , n66378 );
buf ( n66380 , n64675 );
xor ( n66381 , n66379 , n66380 );
buf ( n66382 , n66381 );
buf ( n66383 , n66382 );
xor ( n66384 , n66376 , n66383 );
xor ( n66385 , n63958 , n64394 );
xor ( n66386 , n66385 , n64424 );
buf ( n66387 , n66386 );
buf ( n66388 , n66387 );
not ( n66389 , n66388 );
xor ( n66390 , n63067 , n63070 );
xor ( n66391 , n66390 , n63075 );
xor ( n66392 , n64118 , n64388 );
xor ( n66393 , n66391 , n66392 );
not ( n66394 , n66393 );
buf ( n66395 , n66394 );
buf ( n66396 , n28430 );
not ( n66397 , n66396 );
buf ( n66398 , n66397 );
not ( n66399 , n66398 );
not ( n66400 , n61434 );
or ( n66401 , n66399 , n66400 );
nand ( n66402 , n41656 , n28430 );
nand ( n66403 , n66401 , n66402 );
buf ( n66404 , n66403 );
not ( n66405 , n66404 );
buf ( n66406 , n64413 );
not ( n66407 , n66406 );
or ( n66408 , n66405 , n66407 );
buf ( n66409 , n64407 );
buf ( n66410 , n62582 );
nand ( n66411 , n66409 , n66410 );
buf ( n66412 , n66411 );
buf ( n66413 , n66412 );
nand ( n66414 , n66408 , n66413 );
buf ( n66415 , n66414 );
buf ( n66416 , n66415 );
not ( n66417 , n66416 );
buf ( n66418 , n66417 );
buf ( n66419 , n66418 );
xor ( n66420 , n66395 , n66419 );
and ( n66421 , n42336 , n65238 );
buf ( n66422 , n42366 );
not ( n66423 , n66422 );
buf ( n66424 , n13662 );
not ( n66425 , n66424 );
buf ( n66426 , n66425 );
buf ( n66427 , n66426 );
not ( n66428 , n66427 );
or ( n66429 , n66423 , n66428 );
buf ( n66430 , n13662 );
buf ( n66431 , n63913 );
nand ( n66432 , n66430 , n66431 );
buf ( n66433 , n66432 );
buf ( n66434 , n66433 );
nand ( n66435 , n66429 , n66434 );
buf ( n66436 , n66435 );
buf ( n66437 , n66436 );
not ( n66438 , n66437 );
buf ( n66439 , n42375 );
nor ( n66440 , n66438 , n66439 );
buf ( n66441 , n66440 );
nor ( n66442 , n66421 , n66441 );
buf ( n66443 , n66442 );
and ( n66444 , n66420 , n66443 );
and ( n66445 , n66395 , n66419 );
or ( n66446 , n66444 , n66445 );
buf ( n66447 , n66446 );
buf ( n66448 , n66447 );
nand ( n66449 , n66389 , n66448 );
buf ( n66450 , n66449 );
buf ( n66451 , n66450 );
not ( n66452 , n66451 );
xor ( n66453 , n64108 , n64111 );
xor ( n66454 , n66453 , n64115 );
xor ( n66455 , n64274 , n64383 );
xor ( n66456 , n66454 , n66455 );
buf ( n66457 , n66456 );
not ( n66458 , n66457 );
not ( n66459 , n42372 );
buf ( n66460 , n66459 );
buf ( n66461 , n29463 );
not ( n66462 , n66461 );
not ( n66463 , n24951 );
buf ( n66464 , n66463 );
not ( n66465 , n66464 );
or ( n66466 , n66462 , n66465 );
buf ( n66467 , n42366 );
buf ( n66468 , n29463 );
not ( n66469 , n66468 );
buf ( n66470 , n66469 );
buf ( n66471 , n66470 );
nand ( n66472 , n66467 , n66471 );
buf ( n66473 , n66472 );
buf ( n66474 , n66473 );
nand ( n66475 , n66466 , n66474 );
buf ( n66476 , n66475 );
buf ( n66477 , n66476 );
and ( n66478 , n66460 , n66477 );
buf ( n66479 , n66436 );
buf ( n66480 , n42333 );
not ( n66481 , n66480 );
buf ( n66482 , n66481 );
buf ( n66483 , n66482 );
and ( n66484 , n66479 , n66483 );
nor ( n66485 , n66478 , n66484 );
buf ( n66486 , n66485 );
buf ( n66487 , n66486 );
nand ( n66488 , n66458 , n66487 );
buf ( n66489 , n66488 );
buf ( n66490 , n66489 );
buf ( n66491 , n58857 );
buf ( n66492 , n58897 );
and ( n66493 , n66491 , n66492 );
buf ( n66494 , n58858 );
buf ( n66495 , n58894 );
and ( n66496 , n66494 , n66495 );
nor ( n66497 , n66493 , n66496 );
buf ( n66498 , n66497 );
buf ( n66499 , n66498 );
buf ( n66500 , n58913 );
or ( n66501 , n66499 , n66500 );
buf ( n66502 , n64251 );
buf ( n66503 , n58890 );
or ( n66504 , n66502 , n66503 );
nand ( n66505 , n66501 , n66504 );
buf ( n66506 , n66505 );
buf ( n66507 , n64219 );
buf ( n66508 , n64238 );
or ( n66509 , n66507 , n66508 );
buf ( n66510 , n64241 );
nand ( n66511 , n66509 , n66510 );
buf ( n66512 , n66511 );
xor ( n66513 , n66506 , n66512 );
buf ( n66514 , n58747 );
buf ( n66515 , n60261 );
and ( n66516 , n66514 , n66515 );
buf ( n66517 , n58841 );
buf ( n66518 , n60090 );
and ( n66519 , n66517 , n66518 );
nor ( n66520 , n66516 , n66519 );
buf ( n66521 , n66520 );
buf ( n66522 , n66521 );
buf ( n66523 , n60270 );
or ( n66524 , n66522 , n66523 );
buf ( n66525 , n64291 );
buf ( n66526 , n60100 );
or ( n66527 , n66525 , n66526 );
nand ( n66528 , n66524 , n66527 );
buf ( n66529 , n66528 );
and ( n66530 , n66513 , n66529 );
and ( n66531 , n66506 , n66512 );
or ( n66532 , n66530 , n66531 );
buf ( n66533 , n66532 );
xor ( n66534 , n64147 , n64164 );
xor ( n66535 , n66534 , n64182 );
buf ( n66536 , n66535 );
buf ( n66537 , n66536 );
xor ( n66538 , n66533 , n66537 );
buf ( n66539 , n56582 );
buf ( n66540 , n62681 );
and ( n66541 , n66539 , n66540 );
buf ( n66542 , n56585 );
buf ( n66543 , n62663 );
and ( n66544 , n66542 , n66543 );
nor ( n66545 , n66541 , n66544 );
buf ( n66546 , n66545 );
buf ( n66547 , n66546 );
buf ( n66548 , n62935 );
or ( n66549 , n66547 , n66548 );
buf ( n66550 , n64200 );
buf ( n66551 , n62676 );
or ( n66552 , n66550 , n66551 );
nand ( n66553 , n66549 , n66552 );
buf ( n66554 , n66553 );
buf ( n66555 , n66554 );
buf ( n66556 , n55113 );
buf ( n66557 , n64129 );
and ( n66558 , n66556 , n66557 );
buf ( n66559 , n56655 );
buf ( n66560 , n64133 );
and ( n66561 , n66559 , n66560 );
nor ( n66562 , n66558 , n66561 );
buf ( n66563 , n66562 );
buf ( n66564 , n66563 );
buf ( n66565 , n64141 );
or ( n66566 , n66564 , n66565 );
buf ( n66567 , n64137 );
buf ( n66568 , n63010 );
or ( n66569 , n66567 , n66568 );
nand ( n66570 , n66566 , n66569 );
buf ( n66571 , n66570 );
buf ( n66572 , n66571 );
xor ( n66573 , n66555 , n66572 );
buf ( n66574 , n64068 );
buf ( n66575 , n56652 );
and ( n66576 , n66574 , n66575 );
buf ( n66577 , n64068 );
not ( n66578 , n66577 );
buf ( n66579 , n66578 );
buf ( n66580 , n66579 );
buf ( n66581 , n55201 );
and ( n66582 , n66580 , n66581 );
nor ( n66583 , n66576 , n66582 );
buf ( n66584 , n66583 );
buf ( n66585 , n66584 );
buf ( n66586 , n56664 );
or ( n66587 , n66585 , n66586 );
buf ( n66588 , n64331 );
buf ( n66589 , n56673 );
or ( n66590 , n66588 , n66589 );
nand ( n66591 , n66587 , n66590 );
buf ( n66592 , n66591 );
buf ( n66593 , n66592 );
not ( n66594 , n54816 );
not ( n66595 , n66594 );
not ( n66596 , n55049 );
or ( n66597 , n66595 , n66596 );
not ( n66598 , n55052 );
nand ( n66599 , n66597 , n66598 );
nand ( n66600 , n54784 , n55054 );
xnor ( n66601 , n66599 , n66600 );
buf ( n66602 , n66601 );
not ( n66603 , n66602 );
buf ( n66604 , n66603 );
buf ( n66605 , n66604 );
buf ( n66606 , n56589 );
or ( n66607 , n66605 , n66606 );
buf ( n66608 , n64211 );
not ( n66609 , n66608 );
buf ( n66610 , n66609 );
buf ( n66611 , n66610 );
buf ( n66612 , n56598 );
or ( n66613 , n66611 , n66612 );
nand ( n66614 , n66607 , n66613 );
buf ( n66615 , n66614 );
buf ( n66616 , n66615 );
xor ( n66617 , n66593 , n66616 );
buf ( n66618 , n56800 );
not ( n66619 , n66618 );
buf ( n66620 , n60229 );
buf ( n66621 , n58721 );
and ( n66622 , n66620 , n66621 );
buf ( n66623 , n62652 );
buf ( n66624 , n58718 );
and ( n66625 , n66623 , n66624 );
nor ( n66626 , n66622 , n66625 );
buf ( n66627 , n66626 );
buf ( n66628 , n66627 );
not ( n66629 , n66628 );
buf ( n66630 , n66629 );
buf ( n66631 , n66630 );
not ( n66632 , n66631 );
or ( n66633 , n66619 , n66632 );
buf ( n66634 , n64349 );
buf ( n66635 , n58982 );
or ( n66636 , n66634 , n66635 );
nand ( n66637 , n66633 , n66636 );
buf ( n66638 , n66637 );
buf ( n66639 , n66638 );
and ( n66640 , n66617 , n66639 );
and ( n66641 , n66593 , n66616 );
or ( n66642 , n66640 , n66641 );
buf ( n66643 , n66642 );
buf ( n66644 , n66643 );
and ( n66645 , n66573 , n66644 );
and ( n66646 , n66555 , n66572 );
or ( n66647 , n66645 , n66646 );
buf ( n66648 , n66647 );
buf ( n66649 , n66648 );
and ( n66650 , n66538 , n66649 );
and ( n66651 , n66533 , n66537 );
or ( n66652 , n66650 , n66651 );
buf ( n66653 , n66652 );
xor ( n66654 , n64187 , n64191 );
xor ( n66655 , n66654 , n64265 );
buf ( n66656 , n66655 );
xor ( n66657 , n66653 , n66656 );
xor ( n66658 , n63974 , n63990 );
xor ( n66659 , n66658 , n64007 );
xor ( n66660 , n64280 , n64365 );
xor ( n66661 , n66659 , n66660 );
and ( n66662 , n66657 , n66661 );
and ( n66663 , n66653 , n66656 );
or ( n66664 , n66662 , n66663 );
not ( n66665 , n66664 );
not ( n66666 , n64374 );
and ( n66667 , n64379 , n66666 );
not ( n66668 , n64382 );
and ( n66669 , n64379 , n66668 );
nor ( n66670 , n66667 , n66669 );
not ( n66671 , n64370 );
not ( n66672 , n64379 );
nand ( n66673 , n66671 , n66672 , n64373 );
not ( n66674 , n64370 );
nor ( n66675 , n66674 , n64373 );
nand ( n66676 , n66672 , n66675 );
and ( n66677 , n66670 , n66673 , n66676 );
nand ( n66678 , n66665 , n66677 );
not ( n66679 , n66678 );
xor ( n66680 , n64209 , n64242 );
xor ( n66681 , n66680 , n64260 );
buf ( n66682 , n66681 );
xor ( n66683 , n64299 , n64305 );
xor ( n66684 , n66683 , n64362 );
and ( n66685 , n66682 , n66684 );
xor ( n66686 , n64323 , n64340 );
xor ( n66687 , n66686 , n64358 );
buf ( n66688 , n66687 );
and ( n66689 , n66598 , n66594 );
xor ( n66690 , n66689 , n55049 );
buf ( n66691 , n66690 );
not ( n66692 , n66691 );
buf ( n66693 , n66692 );
buf ( n66694 , n66693 );
buf ( n66695 , n56589 );
or ( n66696 , n66694 , n66695 );
buf ( n66697 , n66604 );
buf ( n66698 , n56598 );
or ( n66699 , n66697 , n66698 );
nand ( n66700 , n66696 , n66699 );
buf ( n66701 , n66700 );
buf ( n66702 , n66701 );
buf ( n66703 , n64211 );
buf ( n66704 , n56652 );
and ( n66705 , n66703 , n66704 );
buf ( n66706 , n66610 );
buf ( n66707 , n55201 );
and ( n66708 , n66706 , n66707 );
nor ( n66709 , n66705 , n66708 );
buf ( n66710 , n66709 );
buf ( n66711 , n66710 );
buf ( n66712 , n56664 );
or ( n66713 , n66711 , n66712 );
buf ( n66714 , n66584 );
buf ( n66715 , n56673 );
or ( n66716 , n66714 , n66715 );
nand ( n66717 , n66713 , n66716 );
buf ( n66718 , n66717 );
buf ( n66719 , n66718 );
and ( n66720 , n66702 , n66719 );
buf ( n66721 , n66720 );
buf ( n66722 , n66721 );
buf ( n66723 , n62782 );
buf ( n66724 , n56641 );
and ( n66725 , n66723 , n66724 );
buf ( n66726 , n62980 );
buf ( n66727 , n56631 );
and ( n66728 , n66726 , n66727 );
nor ( n66729 , n66725 , n66728 );
buf ( n66730 , n66729 );
buf ( n66731 , n66730 );
buf ( n66732 , n56626 );
or ( n66733 , n66731 , n66732 );
buf ( n66734 , n64314 );
buf ( n66735 , n56639 );
or ( n66736 , n66734 , n66735 );
nand ( n66737 , n66733 , n66736 );
buf ( n66738 , n66737 );
buf ( n66739 , n66738 );
xor ( n66740 , n66722 , n66739 );
buf ( n66741 , n55152 );
buf ( n66742 , n62999 );
buf ( n66743 , n66742 );
and ( n66744 , n66741 , n66743 );
buf ( n66745 , n55205 );
buf ( n66746 , n63000 );
and ( n66747 , n66745 , n66746 );
nor ( n66748 , n66744 , n66747 );
buf ( n66749 , n66748 );
buf ( n66750 , n66749 );
buf ( n66751 , n64230 );
or ( n66752 , n66750 , n66751 );
buf ( n66753 , n64235 );
nand ( n66754 , n66752 , n66753 );
buf ( n66755 , n66754 );
buf ( n66756 , n66755 );
and ( n66757 , n66740 , n66756 );
and ( n66758 , n66722 , n66739 );
or ( n66759 , n66757 , n66758 );
buf ( n66760 , n66759 );
xor ( n66761 , n66688 , n66760 );
buf ( n66762 , n58699 );
buf ( n66763 , n64129 );
and ( n66764 , n66762 , n66763 );
buf ( n66765 , n56594 );
buf ( n66766 , n64133 );
and ( n66767 , n66765 , n66766 );
nor ( n66768 , n66764 , n66767 );
buf ( n66769 , n66768 );
buf ( n66770 , n66769 );
buf ( n66771 , n64141 );
or ( n66772 , n66770 , n66771 );
buf ( n66773 , n66563 );
buf ( n66774 , n63010 );
or ( n66775 , n66773 , n66774 );
nand ( n66776 , n66772 , n66775 );
buf ( n66777 , n66776 );
buf ( n66778 , n66777 );
buf ( n66779 , n59009 );
buf ( n66780 , n58897 );
and ( n66781 , n66779 , n66780 );
buf ( n66782 , n60077 );
buf ( n66783 , n58894 );
and ( n66784 , n66782 , n66783 );
nor ( n66785 , n66781 , n66784 );
buf ( n66786 , n66785 );
buf ( n66787 , n66786 );
buf ( n66788 , n58913 );
or ( n66789 , n66787 , n66788 );
buf ( n66790 , n66498 );
buf ( n66791 , n58890 );
or ( n66792 , n66790 , n66791 );
nand ( n66793 , n66789 , n66792 );
buf ( n66794 , n66793 );
buf ( n66795 , n66794 );
xor ( n66796 , n66778 , n66795 );
buf ( n66797 , n60101 );
not ( n66798 , n66797 );
buf ( n66799 , n58823 );
buf ( n66800 , n60261 );
and ( n66801 , n66799 , n66800 );
buf ( n66802 , n58862 );
buf ( n66803 , n60090 );
and ( n66804 , n66802 , n66803 );
nor ( n66805 , n66801 , n66804 );
buf ( n66806 , n66805 );
buf ( n66807 , n66806 );
not ( n66808 , n66807 );
buf ( n66809 , n66808 );
buf ( n66810 , n66809 );
not ( n66811 , n66810 );
or ( n66812 , n66798 , n66811 );
buf ( n66813 , n66521 );
buf ( n66814 , n60100 );
or ( n66815 , n66813 , n66814 );
nand ( n66816 , n66812 , n66815 );
buf ( n66817 , n66816 );
buf ( n66818 , n66817 );
and ( n66819 , n66796 , n66818 );
and ( n66820 , n66778 , n66795 );
or ( n66821 , n66819 , n66820 );
buf ( n66822 , n66821 );
and ( n66823 , n66761 , n66822 );
and ( n66824 , n66688 , n66760 );
or ( n66825 , n66823 , n66824 );
xor ( n66826 , n64299 , n64305 );
xor ( n66827 , n66826 , n64362 );
and ( n66828 , n66825 , n66827 );
and ( n66829 , n66682 , n66825 );
or ( n66830 , n66685 , n66828 , n66829 );
xor ( n66831 , n66653 , n66656 );
xor ( n66832 , n66831 , n66661 );
xor ( n66833 , n66830 , n66832 );
xor ( n66834 , n66533 , n66537 );
xor ( n66835 , n66834 , n66649 );
buf ( n66836 , n66835 );
buf ( n66837 , n66836 );
xor ( n66838 , n66593 , n66616 );
xor ( n66839 , n66838 , n66639 );
buf ( n66840 , n66839 );
buf ( n66841 , n56720 );
buf ( n66842 , n62681 );
and ( n66843 , n66841 , n66842 );
buf ( n66844 , n58792 );
buf ( n66845 , n62663 );
and ( n66846 , n66844 , n66845 );
nor ( n66847 , n66843 , n66846 );
buf ( n66848 , n66847 );
buf ( n66849 , n66848 );
buf ( n66850 , n62935 );
or ( n66851 , n66849 , n66850 );
buf ( n66852 , n66546 );
buf ( n66853 , n62676 );
or ( n66854 , n66852 , n66853 );
nand ( n66855 , n66851 , n66854 );
buf ( n66856 , n66855 );
xor ( n66857 , n66840 , n66856 );
buf ( n66858 , n62643 );
buf ( n66859 , n58721 );
and ( n66860 , n66858 , n66859 );
buf ( n66861 , n62646 );
buf ( n66862 , n58718 );
and ( n66863 , n66861 , n66862 );
nor ( n66864 , n66860 , n66863 );
buf ( n66865 , n66864 );
buf ( n66866 , n66865 );
buf ( n66867 , n56799 );
or ( n66868 , n66866 , n66867 );
buf ( n66869 , n66627 );
buf ( n66870 , n58982 );
or ( n66871 , n66869 , n66870 );
nand ( n66872 , n66868 , n66871 );
buf ( n66873 , n66872 );
buf ( n66874 , n62971 );
buf ( n66875 , n56641 );
and ( n66876 , n66874 , n66875 );
buf ( n66877 , n62974 );
buf ( n66878 , n56631 );
and ( n66879 , n66877 , n66878 );
nor ( n66880 , n66876 , n66879 );
buf ( n66881 , n66880 );
buf ( n66882 , n66881 );
buf ( n66883 , n56626 );
or ( n66884 , n66882 , n66883 );
buf ( n66885 , n66730 );
buf ( n66886 , n56639 );
or ( n66887 , n66885 , n66886 );
nand ( n66888 , n66884 , n66887 );
buf ( n66889 , n66888 );
xor ( n66890 , n66873 , n66889 );
xor ( n66891 , n66702 , n66719 );
buf ( n66892 , n66891 );
and ( n66893 , n66890 , n66892 );
and ( n66894 , n66873 , n66889 );
or ( n66895 , n66893 , n66894 );
and ( n66896 , n66857 , n66895 );
and ( n66897 , n66840 , n66856 );
or ( n66898 , n66896 , n66897 );
xor ( n66899 , n66506 , n66512 );
xor ( n66900 , n66899 , n66529 );
and ( n66901 , n66898 , n66900 );
xor ( n66902 , n66555 , n66572 );
xor ( n66903 , n66902 , n66644 );
buf ( n66904 , n66903 );
xor ( n66905 , n66506 , n66512 );
xor ( n66906 , n66905 , n66529 );
and ( n66907 , n66904 , n66906 );
and ( n66908 , n66898 , n66904 );
or ( n66909 , n66901 , n66907 , n66908 );
buf ( n66910 , n66909 );
xor ( n66911 , n66837 , n66910 );
xor ( n66912 , n64299 , n64305 );
xor ( n66913 , n66912 , n64362 );
xor ( n66914 , n66682 , n66825 );
xor ( n66915 , n66913 , n66914 );
buf ( n66916 , n66915 );
and ( n66917 , n66911 , n66916 );
and ( n66918 , n66837 , n66910 );
or ( n66919 , n66917 , n66918 );
buf ( n66920 , n66919 );
and ( n66921 , n66833 , n66920 );
and ( n66922 , n66830 , n66832 );
or ( n66923 , n66921 , n66922 );
not ( n66924 , n66923 );
or ( n66925 , n66679 , n66924 );
not ( n66926 , n66677 );
nand ( n66927 , n66926 , n66664 );
nand ( n66928 , n66925 , n66927 );
buf ( n66929 , n66928 );
and ( n66930 , n66490 , n66929 );
buf ( n66931 , n66456 );
not ( n66932 , n66931 );
buf ( n66933 , n66486 );
nor ( n66934 , n66932 , n66933 );
buf ( n66935 , n66934 );
buf ( n66936 , n66935 );
nor ( n66937 , n66930 , n66936 );
buf ( n66938 , n66937 );
buf ( n66939 , n66938 );
and ( n66940 , n65268 , n42668 );
not ( n66941 , n64748 );
not ( n66942 , n61446 );
or ( n66943 , n66941 , n66942 );
buf ( n66944 , n13653 );
buf ( n66945 , n64753 );
nand ( n66946 , n66944 , n66945 );
buf ( n66947 , n66946 );
nand ( n66948 , n66943 , n66947 );
not ( n66949 , n66948 );
nor ( n66950 , n66949 , n42711 );
nor ( n66951 , n66940 , n66950 );
buf ( n66952 , n66951 );
xor ( n66953 , n66939 , n66952 );
buf ( n66954 , n42865 );
not ( n66955 , n66954 );
buf ( n66956 , n25181 );
not ( n66957 , n66956 );
or ( n66958 , n66955 , n66957 );
buf ( n66959 , n61462 );
buf ( n66960 , n42862 );
nand ( n66961 , n66959 , n66960 );
buf ( n66962 , n66961 );
buf ( n66963 , n66962 );
nand ( n66964 , n66958 , n66963 );
buf ( n66965 , n66964 );
buf ( n66966 , n66965 );
not ( n66967 , n66966 );
buf ( n66968 , n66967 );
not ( n66969 , n66968 );
not ( n66970 , n43932 );
and ( n66971 , n66969 , n66970 );
and ( n66972 , n43905 , n65247 );
nor ( n66973 , n66971 , n66972 );
buf ( n66974 , n66973 );
and ( n66975 , n66953 , n66974 );
and ( n66976 , n66939 , n66952 );
or ( n66977 , n66975 , n66976 );
buf ( n66978 , n66977 );
buf ( n66979 , n66978 );
not ( n66980 , n66979 );
buf ( n66981 , n66980 );
buf ( n66982 , n66981 );
not ( n66983 , n66982 );
or ( n66984 , n66452 , n66983 );
buf ( n66985 , n66447 );
not ( n66986 , n66985 );
buf ( n66987 , n66387 );
nand ( n66988 , n66986 , n66987 );
buf ( n66989 , n66988 );
buf ( n66990 , n66989 );
nand ( n66991 , n66984 , n66990 );
buf ( n66992 , n66991 );
buf ( n66993 , n66992 );
xor ( n66994 , n64741 , n64766 );
xnor ( n66995 , n66994 , n64789 );
buf ( n66996 , n66995 );
xor ( n66997 , n66993 , n66996 );
buf ( n66998 , n51004 );
not ( n66999 , n66998 );
buf ( n67000 , n41805 );
not ( n67001 , n67000 );
or ( n67002 , n66999 , n67001 );
buf ( n67003 , n53861 );
buf ( n67004 , n51001 );
nand ( n67005 , n67003 , n67004 );
buf ( n67006 , n67005 );
buf ( n67007 , n67006 );
nand ( n67008 , n67002 , n67007 );
buf ( n67009 , n67008 );
buf ( n67010 , n67009 );
not ( n67011 , n67010 );
buf ( n67012 , n37400 );
not ( n67013 , n67012 );
or ( n67014 , n67011 , n67013 );
buf ( n67015 , n65140 );
buf ( n67016 , n37413 );
nand ( n67017 , n67015 , n67016 );
buf ( n67018 , n67017 );
buf ( n67019 , n67018 );
nand ( n67020 , n67014 , n67019 );
buf ( n67021 , n67020 );
buf ( n67022 , n67021 );
and ( n67023 , n66997 , n67022 );
and ( n67024 , n66993 , n66996 );
or ( n67025 , n67023 , n67024 );
buf ( n67026 , n67025 );
buf ( n67027 , n67026 );
and ( n67028 , n66384 , n67027 );
and ( n67029 , n66376 , n66383 );
or ( n67030 , n67028 , n67029 );
buf ( n67031 , n67030 );
and ( n67032 , n66351 , n67031 );
and ( n67033 , n66341 , n66350 );
or ( n67034 , n67032 , n67033 );
buf ( n67035 , n65507 );
buf ( n67036 , n65437 );
xor ( n67037 , n67035 , n67036 );
buf ( n67038 , n65367 );
xor ( n67039 , n67037 , n67038 );
buf ( n67040 , n67039 );
or ( n67041 , n67034 , n67040 );
buf ( n67042 , n65081 );
not ( n67043 , n67042 );
buf ( n67044 , n65344 );
not ( n67045 , n67044 );
and ( n67046 , n67043 , n67045 );
buf ( n67047 , n65344 );
buf ( n67048 , n65081 );
and ( n67049 , n67047 , n67048 );
nor ( n67050 , n67046 , n67049 );
buf ( n67051 , n67050 );
buf ( n67052 , n67051 );
buf ( n67053 , n65059 );
and ( n67054 , n67052 , n67053 );
not ( n67055 , n67052 );
buf ( n67056 , n65352 );
and ( n67057 , n67055 , n67056 );
nor ( n67058 , n67054 , n67057 );
buf ( n67059 , n67058 );
nand ( n67060 , n67041 , n67059 );
buf ( n67061 , n67060 );
buf ( n67062 , n67040 );
buf ( n67063 , n67034 );
nand ( n67064 , n67062 , n67063 );
buf ( n67065 , n67064 );
buf ( n67066 , n67065 );
nand ( n67067 , n67061 , n67066 );
buf ( n67068 , n67067 );
not ( n67069 , n67068 );
xor ( n67070 , n65641 , n65737 );
xor ( n67071 , n67070 , n65742 );
buf ( n67072 , n67071 );
buf ( n67073 , n67072 );
not ( n67074 , n67073 );
buf ( n67075 , n67074 );
buf ( n67076 , n67075 );
xor ( n67077 , n65509 , n65361 );
buf ( n67078 , n67077 );
buf ( n67079 , n65356 );
and ( n67080 , n67078 , n67079 );
not ( n67081 , n67078 );
buf ( n67082 , n65356 );
not ( n67083 , n67082 );
buf ( n67084 , n67083 );
buf ( n67085 , n67084 );
and ( n67086 , n67081 , n67085 );
nor ( n67087 , n67080 , n67086 );
buf ( n67088 , n67087 );
buf ( n67089 , n67088 );
not ( n67090 , n67089 );
buf ( n67091 , n67090 );
buf ( n67092 , n67091 );
nand ( n67093 , n67076 , n67092 );
buf ( n67094 , n67093 );
not ( n67095 , n67094 );
or ( n67096 , n67069 , n67095 );
nand ( n67097 , n67072 , n67088 );
nand ( n67098 , n67096 , n67097 );
buf ( n67099 , n67098 );
not ( n67100 , n67099 );
not ( n67101 , n67100 );
xor ( n67102 , n65589 , n65593 );
xor ( n67103 , n67102 , n65825 );
buf ( n67104 , n67103 );
buf ( n67105 , n67104 );
not ( n67106 , n67105 );
buf ( n67107 , n67106 );
not ( n67108 , n67107 );
or ( n67109 , n67101 , n67108 );
xor ( n67110 , n65763 , n65767 );
xor ( n67111 , n67110 , n65817 );
buf ( n67112 , n67111 );
not ( n67113 , n67112 );
xor ( n67114 , n65727 , n65731 );
xor ( n67115 , n67114 , n65733 );
buf ( n67116 , n67115 );
not ( n67117 , n67116 );
xor ( n67118 , n66146 , n66151 );
xor ( n67119 , n67118 , n66170 );
buf ( n67120 , n67119 );
buf ( n67121 , n67120 );
buf ( n67122 , n56289 );
not ( n67123 , n67122 );
buf ( n67124 , n41805 );
not ( n67125 , n67124 );
or ( n67126 , n67123 , n67125 );
buf ( n67127 , n41769 );
buf ( n67128 , n52094 );
nand ( n67129 , n67127 , n67128 );
buf ( n67130 , n67129 );
buf ( n67131 , n67130 );
nand ( n67132 , n67126 , n67131 );
buf ( n67133 , n67132 );
buf ( n67134 , n67133 );
not ( n67135 , n67134 );
buf ( n67136 , n37397 );
not ( n67137 , n67136 );
or ( n67138 , n67135 , n67137 );
buf ( n67139 , n67009 );
buf ( n67140 , n37410 );
nand ( n67141 , n67139 , n67140 );
buf ( n67142 , n67141 );
buf ( n67143 , n67142 );
nand ( n67144 , n67138 , n67143 );
buf ( n67145 , n67144 );
buf ( n67146 , n67145 );
buf ( n67147 , n45730 );
not ( n67148 , n67147 );
buf ( n67149 , n67148 );
not ( n67150 , n67149 );
buf ( n67151 , n53492 );
not ( n67152 , n67151 );
buf ( n67153 , n44210 );
not ( n67154 , n67153 );
or ( n67155 , n67152 , n67154 );
buf ( n67156 , n50783 );
buf ( n67157 , n45747 );
nand ( n67158 , n67156 , n67157 );
buf ( n67159 , n67158 );
buf ( n67160 , n67159 );
nand ( n67161 , n67155 , n67160 );
buf ( n67162 , n67161 );
not ( n67163 , n67162 );
or ( n67164 , n67150 , n67163 );
not ( n67165 , n64616 );
not ( n67166 , n41763 );
or ( n67167 , n67165 , n67166 );
buf ( n67168 , n41764 );
buf ( n67169 , n45747 );
nand ( n67170 , n67168 , n67169 );
buf ( n67171 , n67170 );
nand ( n67172 , n67167 , n67171 );
nand ( n67173 , n67172 , n46225 );
nand ( n67174 , n67164 , n67173 );
buf ( n67175 , n67174 );
xor ( n67176 , n67146 , n67175 );
xor ( n67177 , n66252 , n66274 );
xor ( n67178 , n67177 , n66301 );
buf ( n67179 , n67178 );
buf ( n67180 , n67179 );
and ( n67181 , n67176 , n67180 );
and ( n67182 , n67146 , n67175 );
or ( n67183 , n67181 , n67182 );
buf ( n67184 , n67183 );
buf ( n67185 , n67184 );
xor ( n67186 , n67121 , n67185 );
buf ( n67187 , n48855 );
not ( n67188 , n67187 );
buf ( n67189 , n48808 );
not ( n67190 , n67189 );
buf ( n67191 , n47119 );
not ( n67192 , n67191 );
or ( n67193 , n67190 , n67192 );
buf ( n67194 , n39205 );
buf ( n67195 , n48818 );
nand ( n67196 , n67194 , n67195 );
buf ( n67197 , n67196 );
buf ( n67198 , n67197 );
nand ( n67199 , n67193 , n67198 );
buf ( n67200 , n67199 );
buf ( n67201 , n67200 );
not ( n67202 , n67201 );
or ( n67203 , n67188 , n67202 );
buf ( n67204 , n48808 );
not ( n67205 , n67204 );
buf ( n67206 , n44157 );
not ( n67207 , n67206 );
or ( n67208 , n67205 , n67207 );
buf ( n67209 , n37586 );
buf ( n67210 , n48821 );
nand ( n67211 , n67209 , n67210 );
buf ( n67212 , n67211 );
buf ( n67213 , n67212 );
nand ( n67214 , n67208 , n67213 );
buf ( n67215 , n67214 );
buf ( n67216 , n67215 );
buf ( n67217 , n48868 );
nand ( n67218 , n67216 , n67217 );
buf ( n67219 , n67218 );
buf ( n67220 , n67219 );
nand ( n67221 , n67203 , n67220 );
buf ( n67222 , n67221 );
buf ( n67223 , n67222 );
and ( n67224 , n67186 , n67223 );
and ( n67225 , n67121 , n67185 );
or ( n67226 , n67224 , n67225 );
buf ( n67227 , n67226 );
buf ( n67228 , n67227 );
not ( n67229 , n67228 );
buf ( n67230 , n67229 );
not ( n67231 , n67230 );
or ( n67232 , C0 , n67231 );
xor ( n67233 , n65294 , n65312 );
xor ( n67234 , n67233 , n65330 );
buf ( n67235 , n67234 );
nand ( n67236 , n67232 , n67235 );
nand ( n67237 , n67236 , C1 );
not ( n67238 , n67237 );
not ( n67239 , n67238 );
buf ( n67240 , n65199 );
not ( n67241 , n67240 );
buf ( n67242 , n65105 );
not ( n67243 , n67242 );
or ( n67244 , n67241 , n67243 );
buf ( n67245 , n65102 );
buf ( n67246 , n65202 );
nand ( n67247 , n67245 , n67246 );
buf ( n67248 , n67247 );
buf ( n67249 , n67248 );
nand ( n67250 , n67244 , n67249 );
buf ( n67251 , n67250 );
buf ( n67252 , n67251 );
buf ( n67253 , n65334 );
not ( n67254 , n67253 );
buf ( n67255 , n67254 );
buf ( n67256 , n67255 );
and ( n67257 , n67252 , n67256 );
not ( n67258 , n67252 );
buf ( n67259 , n65334 );
and ( n67260 , n67258 , n67259 );
nor ( n67261 , n67257 , n67260 );
buf ( n67262 , n67261 );
buf ( n67263 , n67262 );
buf ( n67264 , n67263 );
buf ( n67265 , n67264 );
not ( n67266 , n67265 );
and ( n67267 , n67239 , n67266 );
buf ( n67268 , n67238 );
buf ( n67269 , n67265 );
nand ( n67270 , n67268 , n67269 );
buf ( n67271 , n67270 );
not ( n67272 , n67215 );
not ( n67273 , n48855 );
or ( n67274 , n67272 , n67273 );
not ( n67275 , n65667 );
nand ( n67276 , n67275 , n48868 );
nand ( n67277 , n67274 , n67276 );
buf ( n67278 , n67277 );
not ( n67279 , n67278 );
buf ( n67280 , n67279 );
buf ( n67281 , n67280 );
not ( n67282 , n67281 );
buf ( n67283 , n37511 );
not ( n67284 , n67283 );
buf ( n67285 , n37473 );
not ( n67286 , n67285 );
buf ( n67287 , n52789 );
not ( n67288 , n67287 );
and ( n67289 , n67286 , n67288 );
buf ( n67290 , n41843 );
buf ( n67291 , n52789 );
and ( n67292 , n67290 , n67291 );
nor ( n67293 , n67289 , n67292 );
buf ( n67294 , n67293 );
buf ( n67295 , n67294 );
not ( n67296 , n67295 );
and ( n67297 , n67284 , n67296 );
buf ( n67298 , n41855 );
buf ( n67299 , n65304 );
nor ( n67300 , n67298 , n67299 );
buf ( n67301 , n67300 );
buf ( n67302 , n67301 );
nor ( n67303 , n67297 , n67302 );
buf ( n67304 , n67303 );
buf ( n67305 , n67304 );
not ( n67306 , n67305 );
buf ( n67307 , n67306 );
buf ( n67308 , n67307 );
not ( n67309 , n67308 );
buf ( n67310 , n43798 );
not ( n67311 , n67310 );
or ( n67312 , n41889 , n55841 );
nand ( n67313 , n37892 , n55841 );
nand ( n67314 , n67312 , n67313 );
buf ( n67315 , n67314 );
not ( n67316 , n67315 );
and ( n67317 , n67311 , n67316 );
buf ( n67318 , n41908 );
buf ( n67319 , n65322 );
nor ( n67320 , n67318 , n67319 );
buf ( n67321 , n67320 );
buf ( n67322 , n67321 );
nor ( n67323 , n67317 , n67322 );
buf ( n67324 , n67323 );
buf ( n67325 , n67324 );
not ( n67326 , n67325 );
buf ( n67327 , n67326 );
buf ( n67328 , n67327 );
not ( n67329 , n67328 );
or ( n67330 , n67309 , n67329 );
buf ( n67331 , n67304 );
not ( n67332 , n67331 );
buf ( n67333 , n67324 );
not ( n67334 , n67333 );
or ( n67335 , n67332 , n67334 );
buf ( n67336 , n43868 );
not ( n67337 , n67336 );
buf ( n67338 , n66215 );
not ( n67339 , n67338 );
or ( n67340 , n67337 , n67339 );
buf ( n67341 , n41605 );
not ( n67342 , n67341 );
buf ( n67343 , n50578 );
not ( n67344 , n67343 );
or ( n67345 , n67342 , n67344 );
buf ( n67346 , n47063 );
buf ( n67347 , n41604 );
nand ( n67348 , n67346 , n67347 );
buf ( n67349 , n67348 );
buf ( n67350 , n67349 );
nand ( n67351 , n67345 , n67350 );
buf ( n67352 , n67351 );
buf ( n67353 , n67352 );
not ( n67354 , n41594 );
buf ( n67355 , n67354 );
nand ( n67356 , n67353 , n67355 );
buf ( n67357 , n67356 );
buf ( n67358 , n67357 );
nand ( n67359 , n67340 , n67358 );
buf ( n67360 , n67359 );
buf ( n67361 , n67360 );
xor ( n67362 , n66387 , n66447 );
xor ( n67363 , n67362 , n66978 );
buf ( n67364 , n67363 );
xor ( n67365 , n67361 , n67364 );
buf ( n67366 , n65010 );
not ( n67367 , n67366 );
buf ( n67368 , n51250 );
not ( n67369 , n67368 );
or ( n67370 , n67367 , n67369 );
buf ( n67371 , n41822 );
buf ( n67372 , n44530 );
nand ( n67373 , n67371 , n67372 );
buf ( n67374 , n67373 );
buf ( n67375 , n67374 );
nand ( n67376 , n67370 , n67375 );
buf ( n67377 , n67376 );
not ( n67378 , n67377 );
not ( n67379 , n44517 );
or ( n67380 , n67378 , n67379 );
buf ( n67381 , n66165 );
not ( n67382 , n67381 );
buf ( n67383 , n67382 );
or ( n67384 , n67383 , n44497 );
nand ( n67385 , n67380 , n67384 );
buf ( n67386 , n67385 );
and ( n67387 , n67365 , n67386 );
and ( n67388 , n67361 , n67364 );
or ( n67389 , n67387 , n67388 );
buf ( n67390 , n67389 );
buf ( n67391 , n67390 );
nand ( n67392 , n67335 , n67391 );
buf ( n67393 , n67392 );
buf ( n67394 , n67393 );
nand ( n67395 , n67330 , n67394 );
buf ( n67396 , n67395 );
buf ( n67397 , n67396 );
not ( n67398 , n67397 );
buf ( n67399 , n67398 );
buf ( n67400 , n67399 );
not ( n67401 , n67400 );
or ( n67402 , n67282 , n67401 );
buf ( n67403 , n46907 );
not ( n67404 , n67403 );
buf ( n67405 , n46875 );
not ( n67406 , n67405 );
buf ( n67407 , n44983 );
not ( n67408 , n67407 );
or ( n67409 , n67406 , n67408 );
buf ( n67410 , n38848 );
buf ( n67411 , n46887 );
nand ( n67412 , n67410 , n67411 );
buf ( n67413 , n67412 );
buf ( n67414 , n67413 );
nand ( n67415 , n67409 , n67414 );
buf ( n67416 , n67415 );
buf ( n67417 , n67416 );
not ( n67418 , n67417 );
or ( n67419 , n67404 , n67418 );
buf ( n67420 , n66329 );
buf ( n67421 , n46912 );
nand ( n67422 , n67420 , n67421 );
buf ( n67423 , n67422 );
buf ( n67424 , n67423 );
nand ( n67425 , n67419 , n67424 );
buf ( n67426 , n67425 );
buf ( n67427 , n67426 );
not ( n67428 , n37828 );
not ( n67429 , n37472 );
or ( n67430 , n67428 , n67429 );
nand ( n67431 , n67430 , n12481 );
nand ( n67432 , n41843 , n37829 );
nand ( n67433 , n67431 , n49228 , n67432 );
buf ( n67434 , n67433 );
not ( n67435 , n67434 );
buf ( n67436 , n46619 );
not ( n67437 , n67436 );
buf ( n67438 , n50059 );
buf ( n67439 , n67438 );
buf ( n67440 , n42411 );
and ( n67441 , n67439 , n67440 );
not ( n67442 , n67439 );
buf ( n67443 , n42414 );
and ( n67444 , n67442 , n67443 );
nor ( n67445 , n67441 , n67444 );
buf ( n67446 , n67445 );
buf ( n67447 , n67446 );
not ( n67448 , n67447 );
and ( n67449 , n67437 , n67448 );
buf ( n67450 , n66138 );
not ( n67451 , n67450 );
buf ( n67452 , n38379 );
nor ( n67453 , n67451 , n67452 );
buf ( n67454 , n67453 );
buf ( n67455 , n67454 );
nor ( n67456 , n67449 , n67455 );
buf ( n67457 , n67456 );
buf ( n67458 , n67457 );
not ( n67459 , n67458 );
or ( n67460 , n67435 , n67459 );
not ( n67461 , n42625 );
buf ( n67462 , n44952 );
not ( n67463 , n67462 );
buf ( n67464 , n52670 );
not ( n67465 , n67464 );
or ( n67466 , n67463 , n67465 );
buf ( n67467 , n25159 );
buf ( n67468 , n44949 );
nand ( n67469 , n67467 , n67468 );
buf ( n67470 , n67469 );
buf ( n67471 , n67470 );
nand ( n67472 , n67466 , n67471 );
buf ( n67473 , n67472 );
buf ( n67474 , n67473 );
not ( n67475 , n67474 );
buf ( n67476 , n67475 );
not ( n67477 , n67476 );
and ( n67478 , n67461 , n67477 );
and ( n67479 , n66239 , n47872 );
nor ( n67480 , n67478 , n67479 );
buf ( n67481 , n67480 );
not ( n67482 , n67481 );
buf ( n67483 , n41596 );
not ( n67484 , n67483 );
buf ( n67485 , n41605 );
not ( n67486 , n67485 );
buf ( n67487 , n53579 );
not ( n67488 , n67487 );
or ( n67489 , n67486 , n67488 );
buf ( n67490 , n42149 );
buf ( n67491 , n41604 );
nand ( n67492 , n67490 , n67491 );
buf ( n67493 , n67492 );
buf ( n67494 , n67493 );
nand ( n67495 , n67489 , n67494 );
buf ( n67496 , n67495 );
buf ( n67497 , n67496 );
not ( n67498 , n67497 );
or ( n67499 , n67484 , n67498 );
buf ( n67500 , n67352 );
buf ( n67501 , n43868 );
nand ( n67502 , n67500 , n67501 );
buf ( n67503 , n67502 );
buf ( n67504 , n67503 );
nand ( n67505 , n67499 , n67504 );
buf ( n67506 , n67505 );
not ( n67507 , n67506 );
buf ( n67508 , n67507 );
not ( n67509 , n67508 );
or ( n67510 , n67482 , n67509 );
xor ( n67511 , n66939 , n66952 );
xor ( n67512 , n67511 , n66974 );
buf ( n67513 , n67512 );
buf ( n67514 , n67513 );
not ( n67515 , n67514 );
buf ( n67516 , n67515 );
buf ( n67517 , n67516 );
nand ( n67518 , n67510 , n67517 );
buf ( n67519 , n67518 );
buf ( n67520 , n67519 );
buf ( n67521 , n67480 );
not ( n67522 , n67521 );
buf ( n67523 , n67506 );
nand ( n67524 , n67522 , n67523 );
buf ( n67525 , n67524 );
buf ( n67526 , n67525 );
nand ( n67527 , n67520 , n67526 );
buf ( n67528 , n67527 );
buf ( n67529 , n67528 );
nand ( n67530 , n67460 , n67529 );
buf ( n67531 , n67530 );
buf ( n67532 , n67531 );
buf ( n67533 , n67457 );
not ( n67534 , n67533 );
buf ( n67535 , n67433 );
not ( n67536 , n67535 );
buf ( n67537 , n67536 );
buf ( n67538 , n67537 );
nand ( n67539 , n67534 , n67538 );
buf ( n67540 , n67539 );
buf ( n67541 , n67540 );
nand ( n67542 , n67532 , n67541 );
buf ( n67543 , n67542 );
buf ( n67544 , n67543 );
xor ( n67545 , n67427 , n67544 );
xor ( n67546 , n66200 , n66226 );
xor ( n67547 , n67546 , n66306 );
buf ( n67548 , n67547 );
buf ( n67549 , n67548 );
and ( n67550 , n67545 , n67549 );
and ( n67551 , n67427 , n67544 );
or ( n67552 , n67550 , n67551 );
buf ( n67553 , n67552 );
buf ( n67554 , n67553 );
nand ( n67555 , n67402 , n67554 );
buf ( n67556 , n67555 );
buf ( n67557 , n67556 );
buf ( n67558 , n67396 );
buf ( n67559 , n67277 );
nand ( n67560 , n67558 , n67559 );
buf ( n67561 , n67560 );
buf ( n67562 , n67561 );
nand ( n67563 , n67557 , n67562 );
buf ( n67564 , n67563 );
and ( n67565 , n67271 , n67564 );
nor ( n67566 , n67267 , n67565 );
buf ( n67567 , n67566 );
not ( n67568 , n67567 );
buf ( n67569 , n67568 );
not ( n67570 , n67569 );
or ( n67571 , n67117 , n67570 );
buf ( n67572 , n67116 );
not ( n67573 , n67572 );
buf ( n67574 , n67573 );
buf ( n67575 , n67574 );
not ( n67576 , n67575 );
buf ( n67577 , n67566 );
not ( n67578 , n67577 );
or ( n67579 , n67576 , n67578 );
buf ( n67580 , C0 );
buf ( n67581 , n65148 );
not ( n67582 , n65193 );
not ( n67583 , n65126 );
or ( n67584 , n67582 , n67583 );
or ( n67585 , n65126 , n65193 );
nand ( n67586 , n67584 , n67585 );
xor ( n67587 , n67581 , n67586 );
nand ( n67588 , n62125 , n65651 );
buf ( n67589 , n61853 );
not ( n67590 , n67589 );
buf ( n67591 , n37745 );
not ( n67592 , n67591 );
or ( n67593 , n67590 , n67592 );
buf ( n67594 , n43198 );
buf ( n67595 , n61850 );
nand ( n67596 , n67594 , n67595 );
buf ( n67597 , n67596 );
buf ( n67598 , n67597 );
nand ( n67599 , n67593 , n67598 );
buf ( n67600 , n67599 );
buf ( n67601 , n67600 );
buf ( n67602 , n51488 );
nand ( n67603 , n67601 , n67602 );
buf ( n67604 , n67603 );
nand ( n67605 , n67587 , n67588 , n67604 );
not ( n67606 , n67605 );
not ( n67607 , n46225 );
not ( n67608 , n67162 );
or ( n67609 , n67607 , n67608 );
nand ( n67610 , n65698 , n46246 );
nand ( n67611 , n67609 , n67610 );
not ( n67612 , n67611 );
xor ( n67613 , n65231 , n65278 );
buf ( n67614 , n67613 );
buf ( n67615 , n65282 );
xnor ( n67616 , n67614 , n67615 );
buf ( n67617 , n67616 );
not ( n67618 , n67617 );
not ( n67619 , n67618 );
or ( n67620 , n67612 , n67619 );
buf ( n67621 , n67611 );
not ( n67622 , n67621 );
buf ( n67623 , n67622 );
not ( n67624 , n67623 );
not ( n67625 , n67617 );
or ( n67626 , n67624 , n67625 );
xor ( n67627 , n65243 , n65260 );
xor ( n67628 , n67627 , n65274 );
buf ( n67629 , n67628 );
buf ( n67630 , n67629 );
not ( n67631 , n67630 );
buf ( n67632 , n67631 );
buf ( n67633 , n67632 );
not ( n67634 , n67633 );
not ( n67635 , n42448 );
not ( n67636 , n66187 );
or ( n67637 , n67635 , n67636 );
not ( n67638 , n47716 );
not ( n67639 , n47031 );
or ( n67640 , n67638 , n67639 );
nand ( n67641 , n47725 , n42468 );
nand ( n67642 , n67640 , n67641 );
nand ( n67643 , n47050 , n67642 );
nand ( n67644 , n67637 , n67643 );
buf ( n67645 , n67644 );
not ( n67646 , n67645 );
buf ( n67647 , n67646 );
buf ( n67648 , n67647 );
not ( n67649 , n67648 );
or ( n67650 , n67634 , n67649 );
buf ( n67651 , n42315 );
not ( n67652 , n67651 );
buf ( n67653 , n66293 );
not ( n67654 , n67653 );
or ( n67655 , n67652 , n67654 );
and ( n67656 , n28368 , n42260 );
not ( n67657 , n28368 );
and ( n67658 , n67657 , n59242 );
or ( n67659 , n67656 , n67658 );
buf ( n67660 , n67659 );
buf ( n67661 , n42252 );
nand ( n67662 , n67660 , n67661 );
buf ( n67663 , n67662 );
buf ( n67664 , n67663 );
nand ( n67665 , n67655 , n67664 );
buf ( n67666 , n67665 );
buf ( n67667 , n67666 );
not ( n67668 , n67667 );
buf ( n67669 , n67668 );
not ( n67670 , n67669 );
xor ( n67671 , n66395 , n66419 );
xor ( n67672 , n67671 , n66443 );
buf ( n67673 , n67672 );
not ( n67674 , n67673 );
or ( n67675 , n67670 , n67674 );
buf ( n67676 , n43056 );
not ( n67677 , n67676 );
buf ( n67678 , n58107 );
not ( n67679 , n67678 );
or ( n67680 , n67677 , n67679 );
buf ( n67681 , n61434 );
buf ( n67682 , n43055 );
nand ( n67683 , n67681 , n67682 );
buf ( n67684 , n67683 );
buf ( n67685 , n67684 );
nand ( n67686 , n67680 , n67685 );
buf ( n67687 , n67686 );
buf ( n67688 , n67687 );
not ( n67689 , n67688 );
buf ( n67690 , n62588 );
not ( n67691 , n67690 );
or ( n67692 , n67689 , n67691 );
buf ( n67693 , n66403 );
buf ( n67694 , n47640 );
nand ( n67695 , n67693 , n67694 );
buf ( n67696 , n67695 );
buf ( n67697 , n67696 );
nand ( n67698 , n67692 , n67697 );
buf ( n67699 , n67698 );
not ( n67700 , n67699 );
not ( n67701 , n42668 );
not ( n67702 , n66948 );
or ( n67703 , n67701 , n67702 );
not ( n67704 , n64748 );
not ( n67705 , n41733 );
or ( n67706 , n67704 , n67705 );
buf ( n67707 , n28344 );
buf ( n67708 , n64753 );
nand ( n67709 , n67707 , n67708 );
buf ( n67710 , n67709 );
nand ( n67711 , n67706 , n67710 );
buf ( n67712 , n67711 );
buf ( n67713 , n46047 );
nand ( n67714 , n67712 , n67713 );
buf ( n67715 , n67714 );
nand ( n67716 , n67703 , n67715 );
not ( n67717 , n67716 );
or ( n67718 , n67700 , n67717 );
or ( n67719 , n67699 , n67716 );
xor ( n67720 , n66928 , n66456 );
xnor ( n67721 , n67720 , n66486 );
nand ( n67722 , n67719 , n67721 );
nand ( n67723 , n67718 , n67722 );
nand ( n67724 , n67675 , n67723 );
buf ( n67725 , n67724 );
buf ( n67726 , n67673 );
not ( n67727 , n67726 );
buf ( n67728 , n67666 );
nand ( n67729 , n67727 , n67728 );
buf ( n67730 , n67729 );
buf ( n67731 , n67730 );
nand ( n67732 , n67725 , n67731 );
buf ( n67733 , n67732 );
buf ( n67734 , n67733 );
nand ( n67735 , n67650 , n67734 );
buf ( n67736 , n67735 );
buf ( n67737 , n67736 );
buf ( n67738 , n67644 );
buf ( n67739 , n67629 );
nand ( n67740 , n67738 , n67739 );
buf ( n67741 , n67740 );
buf ( n67742 , n67741 );
nand ( n67743 , n67737 , n67742 );
buf ( n67744 , n67743 );
nand ( n67745 , n67626 , n67744 );
nand ( n67746 , n67620 , n67745 );
not ( n67747 , n67746 );
or ( n67748 , n67606 , n67747 );
not ( n67749 , n67587 );
nand ( n67750 , n67588 , n67604 );
nand ( n67751 , n67749 , n67750 );
nand ( n67752 , n67748 , n67751 );
xor ( n67753 , n67580 , n67752 );
xor ( n67754 , n65488 , n65463 );
xor ( n67755 , n67754 , n65496 );
and ( n67756 , n67753 , n67755 );
or ( n67757 , n67756 , C0 );
buf ( n67758 , n67757 );
nand ( n67759 , n67579 , n67758 );
buf ( n67760 , n67759 );
nand ( n67761 , n67571 , n67760 );
not ( n67762 , n67761 );
or ( n67763 , n67113 , n67762 );
xor ( n67764 , n65814 , n65783 );
xor ( n67765 , n67764 , n65792 );
not ( n67766 , n67765 );
xor ( n67767 , n66341 , n66350 );
xor ( n67768 , n67767 , n67031 );
not ( n67769 , n67768 );
xor ( n67770 , n65672 , n65658 );
xor ( n67771 , n67770 , n65724 );
not ( n67772 , n67771 );
not ( n67773 , n65776 );
xor ( n67774 , n65771 , n67773 );
xor ( n67775 , n67774 , C0 );
nand ( n67776 , n67772 , n67775 );
not ( n67777 , n67776 );
or ( n67778 , n67769 , n67777 );
not ( n67779 , n67775 );
nand ( n67780 , n67779 , n67771 );
nand ( n67781 , n67778 , n67780 );
not ( n67782 , n67781 );
not ( n67783 , n67782 );
and ( n67784 , n67766 , n67783 );
nand ( n67785 , n67765 , n67782 );
xor ( n67786 , n66175 , n66311 );
xor ( n67787 , n67786 , n66337 );
buf ( n67788 , n67787 );
buf ( n67789 , n67788 );
buf ( n67790 , n65705 );
buf ( n67791 , n65714 );
xor ( n67792 , n67790 , n67791 );
buf ( n67793 , n65718 );
xnor ( n67794 , n67792 , n67793 );
buf ( n67795 , n67794 );
buf ( n67796 , n67795 );
xor ( n67797 , n67789 , n67796 );
xor ( n67798 , n66376 , n66383 );
xor ( n67799 , n67798 , n67027 );
buf ( n67800 , n67799 );
buf ( n67801 , n67800 );
and ( n67802 , n67797 , n67801 );
and ( n67803 , n67789 , n67796 );
or ( n67804 , n67802 , n67803 );
buf ( n67805 , n67804 );
buf ( n67806 , n67805 );
xor ( n67807 , n67746 , n67750 );
xor ( n67808 , n67807 , n67587 );
not ( n67809 , n67808 );
or ( n67810 , C0 , n67809 );
buf ( n67811 , C0 );
buf ( n67812 , n67811 );
xor ( n67813 , n67744 , n67623 );
xnor ( n67814 , n67813 , n67618 );
buf ( n67815 , n67814 );
xor ( n67816 , n67812 , n67815 );
buf ( n67817 , n51488 );
not ( n67818 , n67817 );
buf ( n67819 , n61853 );
not ( n67820 , n67819 );
buf ( n67821 , n37786 );
not ( n67822 , n67821 );
or ( n67823 , n67820 , n67822 );
buf ( n67824 , n38480 );
buf ( n67825 , n51493 );
nand ( n67826 , n67824 , n67825 );
buf ( n67827 , n67826 );
buf ( n67828 , n67827 );
nand ( n67829 , n67823 , n67828 );
buf ( n67830 , n67829 );
buf ( n67831 , n67830 );
not ( n67832 , n67831 );
or ( n67833 , n67818 , n67832 );
buf ( n67834 , n67600 );
buf ( n67835 , n52456 );
nand ( n67836 , n67834 , n67835 );
buf ( n67837 , n67836 );
buf ( n67838 , n67837 );
nand ( n67839 , n67833 , n67838 );
buf ( n67840 , n67839 );
buf ( n67841 , n67840 );
and ( n67842 , n67816 , n67841 );
or ( n67843 , n67842 , C0 );
buf ( n67844 , n67843 );
nand ( n67845 , n67810 , n67844 );
nand ( n67846 , C1 , n67845 );
buf ( n67847 , n67846 );
xor ( n67848 , n67806 , n67847 );
xor ( n67849 , n67580 , n67752 );
xor ( n67850 , n67849 , n67755 );
buf ( n67851 , n67850 );
and ( n67852 , n67848 , n67851 );
and ( n67853 , n67806 , n67847 );
or ( n67854 , n67852 , n67853 );
buf ( n67855 , n67854 );
and ( n67856 , n67785 , n67855 );
nor ( n67857 , n67784 , n67856 );
nor ( n67858 , n67112 , n67761 );
or ( n67859 , n67857 , n67858 );
nand ( n67860 , n67763 , n67859 );
buf ( n67861 , n67860 );
nand ( n67862 , n67109 , n67861 );
nand ( n67863 , n67099 , n67104 );
nand ( n67864 , n67862 , n67863 );
nand ( n67865 , n66133 , n67864 );
not ( n67866 , n67865 );
nand ( n67867 , n66006 , n65911 );
nand ( n67868 , n67866 , n67867 );
nand ( n67869 , n66095 , n66130 , n67868 );
not ( n67870 , n66093 );
nand ( n67871 , n67870 , n66087 );
not ( n67872 , n67871 );
buf ( n67873 , n66118 );
buf ( n67874 , n66126 );
nand ( n67875 , n67873 , n67874 );
buf ( n67876 , n67875 );
not ( n67877 , n67876 );
or ( n67878 , n67872 , n67877 );
nand ( n67879 , n67878 , n66130 );
buf ( n67880 , n62096 );
buf ( n67881 , n63469 );
xor ( n67882 , n67880 , n67881 );
buf ( n67883 , n62073 );
xnor ( n67884 , n67882 , n67883 );
buf ( n67885 , n67884 );
xor ( n67886 , n66106 , n66112 );
and ( n67887 , n67886 , n66116 );
and ( n67888 , n66106 , n66112 );
or ( n67889 , n67887 , n67888 );
buf ( n67890 , n67889 );
nand ( n67891 , n67885 , n67890 );
nand ( n67892 , n67869 , n67879 , n67891 );
buf ( n67893 , n67104 );
not ( n67894 , n67893 );
not ( n67895 , n67098 );
not ( n67896 , n67860 );
or ( n67897 , n67895 , n67896 );
or ( n67898 , n67860 , n67098 );
nand ( n67899 , n67897 , n67898 );
buf ( n67900 , n67899 );
not ( n67901 , n67900 );
and ( n67902 , n67894 , n67901 );
buf ( n67903 , n67104 );
buf ( n67904 , n67899 );
and ( n67905 , n67903 , n67904 );
nor ( n67906 , n67902 , n67905 );
buf ( n67907 , n67906 );
buf ( n67908 , n67068 );
not ( n67909 , n67908 );
buf ( n67910 , n67091 );
not ( n67911 , n67910 );
or ( n67912 , n67909 , n67911 );
buf ( n67913 , n67068 );
not ( n67914 , n67913 );
buf ( n67915 , n67088 );
nand ( n67916 , n67914 , n67915 );
buf ( n67917 , n67916 );
buf ( n67918 , n67917 );
nand ( n67919 , n67912 , n67918 );
buf ( n67920 , n67919 );
buf ( n67921 , n67920 );
buf ( n67922 , n67075 );
and ( n67923 , n67921 , n67922 );
not ( n67924 , n67921 );
buf ( n67925 , n67072 );
and ( n67926 , n67924 , n67925 );
nor ( n67927 , n67923 , n67926 );
buf ( n67928 , n67927 );
buf ( n67929 , n67928 );
buf ( n67930 , n67034 );
buf ( n67931 , n67040 );
xor ( n67932 , n67930 , n67931 );
buf ( n67933 , n67059 );
xnor ( n67934 , n67932 , n67933 );
buf ( n67935 , n67934 );
buf ( n67936 , n67935 );
buf ( n67937 , n67757 );
buf ( n67938 , n67116 );
xor ( n67939 , n67937 , n67938 );
buf ( n67940 , n67569 );
xnor ( n67941 , n67939 , n67940 );
buf ( n67942 , n67941 );
buf ( n67943 , n67942 );
xor ( n67944 , n67936 , n67943 );
xor ( n67945 , n67789 , n67796 );
xor ( n67946 , n67945 , n67801 );
buf ( n67947 , n67946 );
buf ( n67948 , n67947 );
xor ( n67949 , n67121 , n67185 );
xor ( n67950 , n67949 , n67223 );
buf ( n67951 , n67950 );
not ( n67952 , n67951 );
buf ( n67953 , C1 );
nand ( n67954 , n67952 , n67953 );
not ( n67955 , n67954 );
xor ( n67956 , n67361 , n67364 );
xor ( n67957 , n67956 , n67386 );
buf ( n67958 , n67957 );
buf ( n67959 , n67958 );
xor ( n67960 , n67537 , n67528 );
xnor ( n67961 , n67960 , n67457 );
buf ( n67962 , n67961 );
xor ( n67963 , n67959 , n67962 );
buf ( n67964 , n52780 );
not ( n67965 , n67964 );
buf ( n67966 , n45270 );
not ( n67967 , n67966 );
or ( n67968 , n67965 , n67967 );
buf ( n67969 , n41769 );
buf ( n67970 , n52789 );
nand ( n67971 , n67969 , n67970 );
buf ( n67972 , n67971 );
buf ( n67973 , n67972 );
nand ( n67974 , n67968 , n67973 );
buf ( n67975 , n67974 );
buf ( n67976 , n67975 );
not ( n67977 , n67976 );
buf ( n67978 , n37400 );
not ( n67979 , n67978 );
or ( n67980 , n67977 , n67979 );
buf ( n67981 , n67133 );
buf ( n67982 , n37413 );
nand ( n67983 , n67981 , n67982 );
buf ( n67984 , n67983 );
buf ( n67985 , n67984 );
nand ( n67986 , n67980 , n67985 );
buf ( n67987 , n67986 );
not ( n67988 , n67987 );
buf ( n67989 , n46390 );
not ( n67990 , n67989 );
buf ( n67991 , n47857 );
not ( n67992 , n67991 );
or ( n67993 , n67990 , n67992 );
buf ( n67994 , n50598 );
buf ( n67995 , n46393 );
nand ( n67996 , n67994 , n67995 );
buf ( n67997 , n67996 );
buf ( n67998 , n67997 );
nand ( n67999 , n67993 , n67998 );
buf ( n68000 , n67999 );
buf ( n68001 , n68000 );
not ( n68002 , n68001 );
buf ( n68003 , n64777 );
not ( n68004 , n68003 );
or ( n68005 , n68002 , n68004 );
buf ( n68006 , n66264 );
buf ( n68007 , n48975 );
nand ( n68008 , n68006 , n68007 );
buf ( n68009 , n68008 );
buf ( n68010 , n68009 );
nand ( n68011 , n68005 , n68010 );
buf ( n68012 , n68011 );
buf ( n68013 , n42847 );
not ( n68014 , n68013 );
buf ( n68015 , n25181 );
not ( n68016 , n68015 );
or ( n68017 , n68014 , n68016 );
buf ( n68018 , n52724 );
buf ( n68019 , n46691 );
nand ( n68020 , n68018 , n68019 );
buf ( n68021 , n68020 );
buf ( n68022 , n68021 );
nand ( n68023 , n68017 , n68022 );
buf ( n68024 , n68023 );
not ( n68025 , n68024 );
not ( n68026 , n53628 );
or ( n68027 , n68025 , n68026 );
buf ( n68028 , n66965 );
buf ( n68029 , n43905 );
nand ( n68030 , n68028 , n68029 );
buf ( n68031 , n68030 );
nand ( n68032 , n68027 , n68031 );
not ( n68033 , n68032 );
buf ( n68034 , n42315 );
not ( n68035 , n68034 );
buf ( n68036 , n67659 );
not ( n68037 , n68036 );
or ( n68038 , n68035 , n68037 );
xor ( n68039 , n59242 , n29754 );
buf ( n68040 , n68039 );
buf ( n68041 , n42252 );
nand ( n68042 , n68040 , n68041 );
buf ( n68043 , n68042 );
buf ( n68044 , n68043 );
nand ( n68045 , n68038 , n68044 );
buf ( n68046 , n68045 );
buf ( n68047 , n68046 );
not ( n68048 , n68047 );
buf ( n68049 , n68048 );
nand ( n68050 , n68033 , n68049 );
not ( n68051 , n68050 );
not ( n68052 , n46047 );
and ( n68053 , n13662 , n64753 );
not ( n68054 , n13662 );
and ( n68055 , n68054 , n64748 );
or ( n68056 , n68053 , n68055 );
not ( n68057 , n68056 );
or ( n68058 , n68052 , n68057 );
nand ( n68059 , n67711 , n42665 );
nand ( n68060 , n68058 , n68059 );
not ( n68061 , n66459 );
buf ( n68062 , n24951 );
not ( n68063 , n68062 );
not ( n68064 , n66398 );
or ( n68065 , n68063 , n68064 );
nand ( n68066 , n63913 , n28430 );
nand ( n68067 , n68065 , n68066 );
not ( n68068 , n68067 );
or ( n68069 , n68061 , n68068 );
nand ( n68070 , n66476 , n66482 );
nand ( n68071 , n68069 , n68070 );
or ( n68072 , n68060 , n68071 );
buf ( n68073 , n68072 );
xor ( n68074 , n66664 , n66677 );
xnor ( n68075 , n68074 , n66923 );
buf ( n68076 , n68075 );
and ( n68077 , n68073 , n68076 );
and ( n68078 , n68060 , n68071 );
buf ( n68079 , n68078 );
nor ( n68080 , n68077 , n68079 );
buf ( n68081 , n68080 );
buf ( n68082 , n68081 );
not ( n68083 , n68082 );
buf ( n68084 , n68083 );
not ( n68085 , n68084 );
or ( n68086 , n68051 , n68085 );
buf ( n68087 , n68046 );
buf ( n68088 , n68032 );
nand ( n68089 , n68087 , n68088 );
buf ( n68090 , n68089 );
nand ( n68091 , n68086 , n68090 );
xor ( n68092 , n68012 , n68091 );
buf ( n68093 , n48323 );
not ( n68094 , n68093 );
buf ( n68095 , n42471 );
not ( n68096 , n68095 );
or ( n68097 , n68094 , n68096 );
buf ( n68098 , n38979 );
buf ( n68099 , n48320 );
nand ( n68100 , n68098 , n68099 );
buf ( n68101 , n68100 );
buf ( n68102 , n68101 );
nand ( n68103 , n68097 , n68102 );
buf ( n68104 , n68103 );
buf ( n68105 , n68104 );
not ( n68106 , n68105 );
buf ( n68107 , n47050 );
not ( n68108 , n68107 );
or ( n68109 , n68106 , n68108 );
buf ( n68110 , n67642 );
buf ( n68111 , n52595 );
nand ( n68112 , n68110 , n68111 );
buf ( n68113 , n68112 );
buf ( n68114 , n68113 );
nand ( n68115 , n68109 , n68114 );
buf ( n68116 , n68115 );
buf ( n68117 , n68116 );
not ( n68118 , n68117 );
buf ( n68119 , n68118 );
xor ( n68120 , n68092 , n68119 );
nand ( n68121 , n67988 , n68120 );
not ( n68122 , n68121 );
and ( n68123 , n52724 , n44949 );
not ( n68124 , n52724 );
and ( n68125 , n68124 , n44952 );
or ( n68126 , n68123 , n68125 );
buf ( n68127 , n68126 );
not ( n68128 , n68127 );
buf ( n68129 , n53628 );
not ( n68130 , n68129 );
or ( n68131 , n68128 , n68130 );
buf ( n68132 , n43904 );
not ( n68133 , n68132 );
buf ( n68134 , n68024 );
nand ( n68135 , n68133 , n68134 );
buf ( n68136 , n68135 );
buf ( n68137 , n68136 );
nand ( n68138 , n68131 , n68137 );
buf ( n68139 , n68138 );
buf ( n68140 , n68139 );
not ( n68141 , n68140 );
buf ( n68142 , n68141 );
not ( n68143 , n68142 );
xor ( n68144 , n68075 , n68071 );
xor ( n68145 , n68144 , n68060 );
not ( n68146 , n68145 );
not ( n68147 , n68146 );
or ( n68148 , n68143 , n68147 );
not ( n68149 , n42374 );
not ( n68150 , n66463 );
not ( n68151 , n43056 );
or ( n68152 , n68150 , n68151 );
buf ( n68153 , n42366 );
buf ( n68154 , n43055 );
nand ( n68155 , n68153 , n68154 );
buf ( n68156 , n68155 );
nand ( n68157 , n68152 , n68156 );
not ( n68158 , n68157 );
or ( n68159 , n68149 , n68158 );
nand ( n68160 , n66482 , n68067 );
nand ( n68161 , n68159 , n68160 );
xor ( n68162 , n66688 , n66760 );
xor ( n68163 , n68162 , n66822 );
buf ( n68164 , n60068 );
buf ( n68165 , n58897 );
and ( n68166 , n68164 , n68165 );
buf ( n68167 , n60071 );
buf ( n68168 , n58897 );
not ( n68169 , n68168 );
buf ( n68170 , n68169 );
buf ( n68171 , n68170 );
and ( n68172 , n68167 , n68171 );
nor ( n68173 , n68166 , n68172 );
buf ( n68174 , n68173 );
buf ( n68175 , n68174 );
buf ( n68176 , n58913 );
or ( n68177 , n68175 , n68176 );
buf ( n68178 , n66786 );
buf ( n68179 , n58890 );
or ( n68180 , n68178 , n68179 );
nand ( n68181 , n68177 , n68180 );
buf ( n68182 , n68181 );
buf ( n68183 , n68182 );
buf ( n68184 , n55201 );
buf ( n68185 , n66601 );
and ( n68186 , n68184 , n68185 );
not ( n68187 , n68184 );
buf ( n68188 , n66604 );
and ( n68189 , n68187 , n68188 );
nor ( n68190 , n68186 , n68189 );
buf ( n68191 , n68190 );
buf ( n68192 , n68191 );
not ( n68193 , n68192 );
buf ( n68194 , n68193 );
buf ( n68195 , n68194 );
buf ( n68196 , n56664 );
or ( n68197 , n68195 , n68196 );
buf ( n68198 , n66710 );
buf ( n68199 , n56673 );
or ( n68200 , n68198 , n68199 );
nand ( n68201 , n68197 , n68200 );
buf ( n68202 , n68201 );
buf ( n68203 , n68202 );
not ( n68204 , n55045 );
not ( n68205 , n68204 );
not ( n68206 , n54884 );
nand ( n68207 , n68206 , n55042 );
not ( n68208 , n68207 );
or ( n68209 , n68205 , n68208 );
nand ( n68210 , n55047 , n54850 );
nand ( n68211 , n68209 , n68210 );
not ( n68212 , n68206 );
not ( n68213 , n55042 );
or ( n68214 , n68212 , n68213 );
nor ( n68215 , n55045 , n68210 );
nand ( n68216 , n68214 , n68215 );
nand ( n68217 , n68211 , n68216 );
buf ( n68218 , n68217 );
not ( n68219 , n68218 );
buf ( n68220 , n68219 );
buf ( n68221 , n68220 );
buf ( n68222 , n56589 );
or ( n68223 , n68221 , n68222 );
buf ( n68224 , n66693 );
buf ( n68225 , n56598 );
or ( n68226 , n68224 , n68225 );
nand ( n68227 , n68223 , n68226 );
buf ( n68228 , n68227 );
buf ( n68229 , n68228 );
xor ( n68230 , n68203 , n68229 );
nand ( n68231 , n68206 , n68204 );
xnor ( n68232 , n55042 , n68231 );
buf ( n68233 , n68232 );
not ( n68234 , n68233 );
buf ( n68235 , n68234 );
buf ( n68236 , n68235 );
buf ( n68237 , n55129 );
or ( n68238 , n68236 , n68237 );
buf ( n68239 , n56598 );
buf ( n68240 , n68220 );
or ( n68241 , n68239 , n68240 );
nand ( n68242 , n68238 , n68241 );
buf ( n68243 , n68242 );
buf ( n68244 , n68243 );
buf ( n68245 , n56670 );
not ( n68246 , n68245 );
buf ( n68247 , n68191 );
not ( n68248 , n68247 );
or ( n68249 , n68246 , n68248 );
buf ( n68250 , n55201 );
buf ( n68251 , n66693 );
and ( n68252 , n68250 , n68251 );
not ( n68253 , n68250 );
buf ( n68254 , n66690 );
and ( n68255 , n68253 , n68254 );
nor ( n68256 , n68252 , n68255 );
buf ( n68257 , n68256 );
buf ( n68258 , n68257 );
buf ( n68259 , n56664 );
or ( n68260 , n68258 , n68259 );
nand ( n68261 , n68249 , n68260 );
buf ( n68262 , n68261 );
buf ( n68263 , n68262 );
and ( n68264 , n68244 , n68263 );
buf ( n68265 , n68264 );
buf ( n68266 , n68265 );
and ( n68267 , n68230 , n68266 );
and ( n68268 , n68203 , n68229 );
or ( n68269 , n68267 , n68268 );
buf ( n68270 , n68269 );
buf ( n68271 , n68270 );
xor ( n68272 , n68183 , n68271 );
not ( n68273 , n63010 );
not ( n68274 , n68273 );
not ( n68275 , n66769 );
not ( n68276 , n68275 );
or ( n68277 , n68274 , n68276 );
and ( n68278 , n56585 , n64133 );
and ( n68279 , n64129 , n56582 );
nor ( n68280 , n68278 , n68279 );
not ( n68281 , n68280 );
nand ( n68282 , n68281 , n63013 );
nand ( n68283 , n68277 , n68282 );
buf ( n68284 , n68283 );
and ( n68285 , n68272 , n68284 );
and ( n68286 , n68183 , n68271 );
or ( n68287 , n68285 , n68286 );
buf ( n68288 , n68287 );
buf ( n68289 , n68288 );
xor ( n68290 , n66722 , n66739 );
xor ( n68291 , n68290 , n66756 );
buf ( n68292 , n68291 );
buf ( n68293 , n68292 );
xor ( n68294 , n68289 , n68293 );
buf ( n68295 , n58835 );
buf ( n68296 , n62681 );
and ( n68297 , n68295 , n68296 );
buf ( n68298 , n58841 );
buf ( n68299 , n62663 );
and ( n68300 , n68298 , n68299 );
nor ( n68301 , n68297 , n68300 );
buf ( n68302 , n68301 );
buf ( n68303 , n68302 );
buf ( n68304 , n62935 );
or ( n68305 , n68303 , n68304 );
buf ( n68306 , n66848 );
buf ( n68307 , n62676 );
or ( n68308 , n68306 , n68307 );
nand ( n68309 , n68305 , n68308 );
buf ( n68310 , n68309 );
buf ( n68311 , n68310 );
buf ( n68312 , n55113 );
buf ( n68313 , n66742 );
and ( n68314 , n68312 , n68313 );
buf ( n68315 , n56655 );
buf ( n68316 , n63000 );
and ( n68317 , n68315 , n68316 );
nor ( n68318 , n68314 , n68317 );
buf ( n68319 , n68318 );
buf ( n68320 , n68319 );
buf ( n68321 , n64230 );
or ( n68322 , n68320 , n68321 );
buf ( n68323 , n66749 );
buf ( n68324 , n64227 );
or ( n68325 , n68323 , n68324 );
nand ( n68326 , n68322 , n68325 );
buf ( n68327 , n68326 );
buf ( n68328 , n68327 );
xor ( n68329 , n68311 , n68328 );
buf ( n68330 , n62782 );
buf ( n68331 , n58721 );
and ( n68332 , n68330 , n68331 );
buf ( n68333 , n62980 );
buf ( n68334 , n58718 );
and ( n68335 , n68333 , n68334 );
nor ( n68336 , n68332 , n68335 );
buf ( n68337 , n68336 );
buf ( n68338 , n68337 );
buf ( n68339 , n56799 );
or ( n68340 , n68338 , n68339 );
buf ( n68341 , n66865 );
buf ( n68342 , n58982 );
or ( n68343 , n68341 , n68342 );
nand ( n68344 , n68340 , n68343 );
buf ( n68345 , n68344 );
buf ( n68346 , n68345 );
buf ( n68347 , n64068 );
buf ( n68348 , n56641 );
and ( n68349 , n68347 , n68348 );
buf ( n68350 , n66579 );
buf ( n68351 , n56631 );
and ( n68352 , n68350 , n68351 );
nor ( n68353 , n68349 , n68352 );
buf ( n68354 , n68353 );
buf ( n68355 , n68354 );
buf ( n68356 , n56626 );
or ( n68357 , n68355 , n68356 );
buf ( n68358 , n66881 );
buf ( n68359 , n56639 );
or ( n68360 , n68358 , n68359 );
nand ( n68361 , n68357 , n68360 );
buf ( n68362 , n68361 );
buf ( n68363 , n68362 );
xor ( n68364 , n68346 , n68363 );
buf ( n68365 , n58887 );
not ( n68366 , n68365 );
buf ( n68367 , n68174 );
not ( n68368 , n68367 );
buf ( n68369 , n68368 );
buf ( n68370 , n68369 );
not ( n68371 , n68370 );
or ( n68372 , n68366 , n68371 );
buf ( n68373 , n62652 );
buf ( n68374 , n68170 );
or ( n68375 , n68373 , n68374 );
buf ( n68376 , n60229 );
buf ( n68377 , n58897 );
or ( n68378 , n68376 , n68377 );
nand ( n68379 , n68375 , n68378 );
buf ( n68380 , n68379 );
buf ( n68381 , n68380 );
not ( n68382 , n68381 );
buf ( n68383 , n68382 );
buf ( n68384 , n68383 );
buf ( n68385 , n58913 );
or ( n68386 , n68384 , n68385 );
nand ( n68387 , n68372 , n68386 );
buf ( n68388 , n68387 );
buf ( n68389 , n68388 );
and ( n68390 , n68364 , n68389 );
and ( n68391 , n68346 , n68363 );
or ( n68392 , n68390 , n68391 );
buf ( n68393 , n68392 );
buf ( n68394 , n68393 );
and ( n68395 , n68329 , n68394 );
and ( n68396 , n68311 , n68328 );
or ( n68397 , n68395 , n68396 );
buf ( n68398 , n68397 );
buf ( n68399 , n68398 );
and ( n68400 , n68294 , n68399 );
and ( n68401 , n68289 , n68293 );
or ( n68402 , n68400 , n68401 );
buf ( n68403 , n68402 );
xor ( n68404 , n66506 , n66512 );
xor ( n68405 , n68404 , n66529 );
xor ( n68406 , n66898 , n66904 );
xor ( n68407 , n68405 , n68406 );
xor ( n68408 , n68403 , n68407 );
xor ( n68409 , n68163 , n68408 );
not ( n68410 , n68409 );
and ( n68411 , n60077 , n60090 );
and ( n68412 , n59009 , n60261 );
nor ( n68413 , n68411 , n68412 );
or ( n68414 , n68413 , n60270 );
and ( n68415 , n58858 , n60090 );
and ( n68416 , n58857 , n60261 );
nor ( n68417 , n68415 , n68416 );
or ( n68418 , n68417 , n60100 );
nand ( n68419 , n68414 , n68418 );
xor ( n68420 , n68203 , n68229 );
xor ( n68421 , n68420 , n68266 );
buf ( n68422 , n68421 );
xor ( n68423 , n68419 , n68422 );
not ( n68424 , n63013 );
buf ( n68425 , n56720 );
buf ( n68426 , n64129 );
and ( n68427 , n68425 , n68426 );
buf ( n68428 , n58792 );
buf ( n68429 , n64133 );
and ( n68430 , n68428 , n68429 );
nor ( n68431 , n68427 , n68430 );
buf ( n68432 , n68431 );
buf ( n68433 , n68432 );
not ( n68434 , n68433 );
buf ( n68435 , n68434 );
not ( n68436 , n68435 );
or ( n68437 , n68424 , n68436 );
or ( n68438 , n68280 , n63010 );
nand ( n68439 , n68437 , n68438 );
and ( n68440 , n68423 , n68439 );
and ( n68441 , n68419 , n68422 );
or ( n68442 , n68440 , n68441 );
buf ( n68443 , n68442 );
or ( n68444 , n68302 , n62676 );
not ( n68445 , n62935 );
and ( n68446 , n58862 , n60096 );
and ( n68447 , n58823 , n62663 );
nor ( n68448 , n68446 , n68447 );
nand ( n68449 , n68445 , n68448 );
nand ( n68450 , n68444 , n68449 );
buf ( n68451 , n68450 );
buf ( n68452 , n55249 );
buf ( n68453 , n66742 );
and ( n68454 , n68452 , n68453 );
buf ( n68455 , n56594 );
buf ( n68456 , n63000 );
and ( n68457 , n68455 , n68456 );
nor ( n68458 , n68454 , n68457 );
buf ( n68459 , n68458 );
or ( n68460 , n68459 , n64230 );
not ( n68461 , n68319 );
nand ( n68462 , n68461 , n1664 );
nand ( n68463 , n68460 , n68462 );
buf ( n68464 , n68463 );
xor ( n68465 , n68451 , n68464 );
xor ( n68466 , n68244 , n68263 );
buf ( n68467 , n68466 );
buf ( n68468 , n68467 );
buf ( n68469 , n64211 );
buf ( n68470 , n56641 );
and ( n68471 , n68469 , n68470 );
buf ( n68472 , n66610 );
buf ( n68473 , n56631 );
and ( n68474 , n68472 , n68473 );
nor ( n68475 , n68471 , n68474 );
buf ( n68476 , n68475 );
buf ( n68477 , n68476 );
buf ( n68478 , n56626 );
or ( n68479 , n68477 , n68478 );
buf ( n68480 , n68354 );
buf ( n68481 , n56639 );
or ( n68482 , n68480 , n68481 );
nand ( n68483 , n68479 , n68482 );
buf ( n68484 , n68483 );
buf ( n68485 , n68484 );
xor ( n68486 , n68468 , n68485 );
buf ( n68487 , n58887 );
not ( n68488 , n68487 );
buf ( n68489 , n68380 );
not ( n68490 , n68489 );
or ( n68491 , n68488 , n68490 );
buf ( n68492 , n62643 );
buf ( n68493 , n58897 );
and ( n68494 , n68492 , n68493 );
buf ( n68495 , n62646 );
buf ( n68496 , n58894 );
and ( n68497 , n68495 , n68496 );
nor ( n68498 , n68494 , n68497 );
buf ( n68499 , n68498 );
buf ( n68500 , n68499 );
buf ( n68501 , n58913 );
or ( n68502 , n68500 , n68501 );
nand ( n68503 , n68491 , n68502 );
buf ( n68504 , n68503 );
buf ( n68505 , n68504 );
and ( n68506 , n68486 , n68505 );
and ( n68507 , n68468 , n68485 );
or ( n68508 , n68506 , n68507 );
buf ( n68509 , n68508 );
buf ( n68510 , n68509 );
and ( n68511 , n68465 , n68510 );
and ( n68512 , n68451 , n68464 );
or ( n68513 , n68511 , n68512 );
buf ( n68514 , n68513 );
buf ( n68515 , n68514 );
xor ( n68516 , n68443 , n68515 );
xor ( n68517 , n68311 , n68328 );
xor ( n68518 , n68517 , n68394 );
buf ( n68519 , n68518 );
buf ( n68520 , n68519 );
and ( n68521 , n68516 , n68520 );
and ( n68522 , n68443 , n68515 );
or ( n68523 , n68521 , n68522 );
buf ( n68524 , n68523 );
buf ( n68525 , n68524 );
xor ( n68526 , n68289 , n68293 );
xor ( n68527 , n68526 , n68399 );
buf ( n68528 , n68527 );
buf ( n68529 , n68528 );
xor ( n68530 , n68525 , n68529 );
xor ( n68531 , n66840 , n66856 );
xor ( n68532 , n68531 , n66895 );
xor ( n68533 , n66778 , n66795 );
xor ( n68534 , n68533 , n66818 );
buf ( n68535 , n68534 );
or ( n68536 , n66806 , n60100 );
or ( n68537 , n68417 , n60270 );
nand ( n68538 , n68536 , n68537 );
xor ( n68539 , n66873 , n66889 );
xor ( n68540 , n68539 , n66892 );
and ( n68541 , n68538 , n68540 );
xor ( n68542 , n68183 , n68271 );
xor ( n68543 , n68542 , n68284 );
buf ( n68544 , n68543 );
xor ( n68545 , n66873 , n66889 );
xor ( n68546 , n68545 , n66892 );
and ( n68547 , n68544 , n68546 );
and ( n68548 , n68538 , n68544 );
or ( n68549 , n68541 , n68547 , n68548 );
xor ( n68550 , n68535 , n68549 );
xor ( n68551 , n68532 , n68550 );
buf ( n68552 , n68551 );
and ( n68553 , n68530 , n68552 );
and ( n68554 , n68525 , n68529 );
or ( n68555 , n68553 , n68554 );
buf ( n68556 , n68555 );
not ( n68557 , n68556 );
xor ( n68558 , n66840 , n66856 );
xor ( n68559 , n68558 , n66895 );
and ( n68560 , n68535 , n68559 );
xor ( n68561 , n66840 , n66856 );
xor ( n68562 , n68561 , n66895 );
and ( n68563 , n68549 , n68562 );
and ( n68564 , n68535 , n68549 );
or ( n68565 , n68560 , n68563 , n68564 );
not ( n68566 , n68565 );
nand ( n68567 , n68557 , n68566 );
not ( n68568 , n68567 );
or ( n68569 , n68410 , n68568 );
nand ( n68570 , n68556 , n68565 );
nand ( n68571 , n68569 , n68570 );
not ( n68572 , n68571 );
xor ( n68573 , n66837 , n66910 );
xor ( n68574 , n68573 , n66916 );
buf ( n68575 , n68574 );
not ( n68576 , n68575 );
xor ( n68577 , n66688 , n66760 );
xor ( n68578 , n68577 , n66822 );
and ( n68579 , n68403 , n68578 );
xor ( n68580 , n66688 , n66760 );
xor ( n68581 , n68580 , n66822 );
and ( n68582 , n68407 , n68581 );
and ( n68583 , n68403 , n68407 );
or ( n68584 , n68579 , n68582 , n68583 );
not ( n68585 , n68584 );
nand ( n68586 , n68576 , n68585 );
not ( n68587 , n68586 );
or ( n68588 , n68572 , n68587 );
nor ( n68589 , n68576 , n68585 );
not ( n68590 , n68589 );
nand ( n68591 , n68588 , n68590 );
buf ( n68592 , n68591 );
xor ( n68593 , n66830 , n66832 );
xor ( n68594 , n68593 , n66920 );
buf ( n68595 , n68594 );
xor ( n68596 , n68592 , n68595 );
buf ( n68597 , n68596 );
xor ( n68598 , n68161 , n68597 );
not ( n68599 , n68598 );
buf ( n68600 , n46047 );
buf ( n68601 , n64748 );
not ( n68602 , n68601 );
buf ( n68603 , n66470 );
not ( n68604 , n68603 );
or ( n68605 , n68602 , n68604 );
not ( n68606 , n25226 );
buf ( n68607 , n68606 );
buf ( n68608 , n29463 );
nand ( n68609 , n68607 , n68608 );
buf ( n68610 , n68609 );
buf ( n68611 , n68610 );
nand ( n68612 , n68605 , n68611 );
buf ( n68613 , n68612 );
buf ( n68614 , n68613 );
nand ( n68615 , n68600 , n68614 );
buf ( n68616 , n68615 );
nand ( n68617 , n68056 , n42665 );
nand ( n68618 , n68616 , n68617 );
not ( n68619 , n68618 );
not ( n68620 , n59928 );
buf ( n68621 , n61434 );
not ( n68622 , n68621 );
buf ( n68623 , n46691 );
not ( n68624 , n68623 );
and ( n68625 , n68622 , n68624 );
buf ( n68626 , n61442 );
buf ( n68627 , n46691 );
and ( n68628 , n68626 , n68627 );
nor ( n68629 , n68625 , n68628 );
buf ( n68630 , n68629 );
not ( n68631 , n68630 );
not ( n68632 , n68631 );
or ( n68633 , n68620 , n68632 );
buf ( n68634 , n42862 );
buf ( n68635 , n61434 );
and ( n68636 , n68634 , n68635 );
not ( n68637 , n68634 );
buf ( n68638 , n62598 );
and ( n68639 , n68637 , n68638 );
nor ( n68640 , n68636 , n68639 );
buf ( n68641 , n68640 );
or ( n68642 , n68641 , n62579 );
nand ( n68643 , n68633 , n68642 );
not ( n68644 , n68643 );
nand ( n68645 , n68619 , n68644 );
not ( n68646 , n68645 );
or ( n68647 , n68599 , n68646 );
nand ( n68648 , n68643 , n68618 );
nand ( n68649 , n68647 , n68648 );
nand ( n68650 , n68148 , n68649 );
buf ( n68651 , n68650 );
buf ( n68652 , n68146 );
not ( n68653 , n68652 );
buf ( n68654 , n68139 );
nand ( n68655 , n68653 , n68654 );
buf ( n68656 , n68655 );
buf ( n68657 , n68656 );
nand ( n68658 , n68651 , n68657 );
buf ( n68659 , n68658 );
buf ( n68660 , n68659 );
buf ( n68661 , n50060 );
not ( n68662 , n68661 );
buf ( n68663 , n38994 );
not ( n68664 , n68663 );
or ( n68665 , n68662 , n68664 );
buf ( n68666 , n42468 );
buf ( n68667 , n67438 );
nand ( n68668 , n68666 , n68667 );
buf ( n68669 , n68668 );
buf ( n68670 , n68669 );
nand ( n68671 , n68665 , n68670 );
buf ( n68672 , n68671 );
buf ( n68673 , n68672 );
not ( n68674 , n68673 );
buf ( n68675 , n47050 );
not ( n68676 , n68675 );
or ( n68677 , n68674 , n68676 );
buf ( n68678 , n68104 );
buf ( n68679 , n50104 );
nand ( n68680 , n68678 , n68679 );
buf ( n68681 , n68680 );
buf ( n68682 , n68681 );
nand ( n68683 , n68677 , n68682 );
buf ( n68684 , n68683 );
buf ( n68685 , n68684 );
xor ( n68686 , n68660 , n68685 );
buf ( n68687 , n44496 );
not ( n68688 , n68687 );
buf ( n68689 , n65010 );
not ( n68690 , n68689 );
buf ( n68691 , n41915 );
not ( n68692 , n68691 );
or ( n68693 , n68690 , n68692 );
buf ( n68694 , n59291 );
buf ( n68695 , n44530 );
nand ( n68696 , n68694 , n68695 );
buf ( n68697 , n68696 );
buf ( n68698 , n68697 );
nand ( n68699 , n68693 , n68698 );
buf ( n68700 , n68699 );
buf ( n68701 , n68700 );
not ( n68702 , n68701 );
or ( n68703 , n68688 , n68702 );
buf ( n68704 , n65010 );
not ( n68705 , n68704 );
buf ( n68706 , n41873 );
not ( n68707 , n68706 );
or ( n68708 , n68705 , n68707 );
buf ( n68709 , n50575 );
buf ( n68710 , n44530 );
nand ( n68711 , n68709 , n68710 );
buf ( n68712 , n68711 );
buf ( n68713 , n68712 );
nand ( n68714 , n68708 , n68713 );
buf ( n68715 , n68714 );
buf ( n68716 , n68715 );
buf ( n68717 , n44517 );
nand ( n68718 , n68716 , n68717 );
buf ( n68719 , n68718 );
buf ( n68720 , n68719 );
nand ( n68721 , n68703 , n68720 );
buf ( n68722 , n68721 );
buf ( n68723 , n68722 );
and ( n68724 , n68686 , n68723 );
and ( n68725 , n68660 , n68685 );
or ( n68726 , n68724 , n68725 );
buf ( n68727 , n68726 );
not ( n68728 , n68727 );
or ( n68729 , n68122 , n68728 );
buf ( n68730 , n67987 );
buf ( n68731 , n68120 );
not ( n68732 , n68731 );
buf ( n68733 , n68732 );
buf ( n68734 , n68733 );
nand ( n68735 , n68730 , n68734 );
buf ( n68736 , n68735 );
nand ( n68737 , n68729 , n68736 );
buf ( n68738 , n68737 );
and ( n68739 , n67963 , n68738 );
and ( n68740 , n67959 , n67962 );
or ( n68741 , n68739 , n68740 );
buf ( n68742 , n68741 );
not ( n68743 , n68742 );
or ( n68744 , n67955 , n68743 );
buf ( n68745 , C1 );
nand ( n68746 , n68744 , n68745 );
buf ( n68747 , n68746 );
xor ( n68748 , n67948 , n68747 );
not ( n68749 , n67227 );
and ( n68750 , n68749 , C1 );
nor ( n68751 , C0 , n68750 );
buf ( n68752 , n68751 );
buf ( n68753 , n67235 );
xor ( n68754 , n68752 , n68753 );
buf ( n68755 , n68754 );
buf ( n68756 , n68755 );
and ( n68757 , n68748 , n68756 );
and ( n68758 , n67948 , n68747 );
or ( n68759 , n68757 , n68758 );
buf ( n68760 , n68759 );
buf ( n68761 , n68760 );
not ( n68762 , n68761 );
buf ( n68763 , n68762 );
not ( n68764 , n68763 );
xor ( n68765 , n67564 , n67262 );
and ( n68766 , n68765 , n67238 );
not ( n68767 , n68765 );
and ( n68768 , n68767 , n67237 );
nor ( n68769 , n68766 , n68768 );
not ( n68770 , n68769 );
not ( n68771 , n68770 );
and ( n68772 , n68764 , n68771 );
buf ( n68773 , n68763 );
buf ( n68774 , n68770 );
nand ( n68775 , n68773 , n68774 );
buf ( n68776 , n68775 );
buf ( n68777 , n67277 );
not ( n68778 , n68777 );
buf ( n68779 , n67399 );
not ( n68780 , n68779 );
or ( n68781 , n68778 , n68780 );
buf ( n68782 , n67396 );
buf ( n68783 , n67280 );
nand ( n68784 , n68782 , n68783 );
buf ( n68785 , n68784 );
buf ( n68786 , n68785 );
nand ( n68787 , n68781 , n68786 );
buf ( n68788 , n68787 );
xnor ( n68789 , n68788 , n67553 );
buf ( n68790 , n68789 );
not ( n68791 , n68790 );
buf ( n68792 , n68791 );
buf ( n68793 , n68792 );
not ( n68794 , n68793 );
and ( n68795 , n67390 , n67304 );
not ( n68796 , n67390 );
and ( n68797 , n68796 , n67307 );
or ( n68798 , n68795 , n68797 );
xnor ( n68799 , n68798 , n67327 );
not ( n68800 , n68799 );
xor ( n68801 , n67427 , n67544 );
xor ( n68802 , n68801 , n67549 );
buf ( n68803 , n68802 );
buf ( n68804 , n68803 );
not ( n68805 , n68804 );
buf ( n68806 , n68805 );
not ( n68807 , n68806 );
and ( n68808 , n68800 , n68807 );
buf ( n68809 , n68799 );
buf ( n68810 , n68806 );
nand ( n68811 , n68809 , n68810 );
buf ( n68812 , n68811 );
not ( n68813 , n48868 );
not ( n68814 , n67200 );
or ( n68815 , n68813 , n68814 );
buf ( n68816 , n48808 );
not ( n68817 , n68816 );
buf ( n68818 , n42461 );
not ( n68819 , n68818 );
or ( n68820 , n68817 , n68819 );
buf ( n68821 , n38821 );
buf ( n68822 , n48818 );
nand ( n68823 , n68821 , n68822 );
buf ( n68824 , n68823 );
buf ( n68825 , n68824 );
nand ( n68826 , n68820 , n68825 );
buf ( n68827 , n68826 );
buf ( n68828 , n68827 );
buf ( n68829 , n48855 );
nand ( n68830 , n68828 , n68829 );
buf ( n68831 , n68830 );
nand ( n68832 , n68815 , n68831 );
not ( n68833 , n68832 );
not ( n68834 , n67507 );
not ( n68835 , n67516 );
or ( n68836 , n68834 , n68835 );
nand ( n68837 , n67513 , n67506 );
nand ( n68838 , n68836 , n68837 );
not ( n68839 , n67480 );
and ( n68840 , n68838 , n68839 );
not ( n68841 , n68838 );
and ( n68842 , n68841 , n67480 );
nor ( n68843 , n68840 , n68842 );
not ( n68844 , n50608 );
buf ( n68845 , n47716 );
not ( n68846 , n68845 );
buf ( n68847 , n47857 );
not ( n68848 , n68847 );
or ( n68849 , n68846 , n68848 );
buf ( n68850 , n24092 );
buf ( n68851 , n47713 );
nand ( n68852 , n68850 , n68851 );
buf ( n68853 , n68852 );
buf ( n68854 , n68853 );
nand ( n68855 , n68849 , n68854 );
buf ( n68856 , n68855 );
not ( n68857 , n68856 );
or ( n68858 , n68844 , n68857 );
buf ( n68859 , n68000 );
buf ( n68860 , n46633 );
nand ( n68861 , n68859 , n68860 );
buf ( n68862 , n68861 );
nand ( n68863 , n68858 , n68862 );
not ( n68864 , n68863 );
not ( n68865 , n43868 );
not ( n68866 , n67496 );
or ( n68867 , n68865 , n68866 );
and ( n68868 , n47434 , n47432 );
and ( n68869 , n41605 , n68868 );
not ( n68870 , n41605 );
and ( n68871 , n68870 , n50624 );
or ( n68872 , n68869 , n68871 );
nand ( n68873 , n68872 , n67354 );
nand ( n68874 , n68867 , n68873 );
not ( n68875 , n68874 );
or ( n68876 , n68864 , n68875 );
buf ( n68877 , n68863 );
not ( n68878 , n68877 );
buf ( n68879 , n68878 );
not ( n68880 , n68879 );
buf ( n68881 , n68874 );
not ( n68882 , n68881 );
buf ( n68883 , n68882 );
not ( n68884 , n68883 );
or ( n68885 , n68880 , n68884 );
not ( n68886 , n68084 );
not ( n68887 , n68049 );
or ( n68888 , n68886 , n68887 );
buf ( n68889 , n68046 );
buf ( n68890 , n68081 );
nand ( n68891 , n68889 , n68890 );
buf ( n68892 , n68891 );
nand ( n68893 , n68888 , n68892 );
buf ( n68894 , n68032 );
xor ( n68895 , n68893 , n68894 );
nand ( n68896 , n68885 , n68895 );
nand ( n68897 , n68876 , n68896 );
not ( n68898 , n68897 );
buf ( n68899 , n46875 );
not ( n68900 , n68899 );
buf ( n68901 , n39671 );
not ( n68902 , n68901 );
or ( n68903 , n68900 , n68902 );
buf ( n68904 , n42434 );
buf ( n68905 , n46887 );
nand ( n68906 , n68904 , n68905 );
buf ( n68907 , n68906 );
buf ( n68908 , n68907 );
nand ( n68909 , n68903 , n68908 );
buf ( n68910 , n68909 );
nand ( n68911 , n68910 , n46912 );
nand ( n68912 , n41799 , n46875 );
not ( n68913 , n68912 );
buf ( n68914 , n29290 );
buf ( n68915 , n46887 );
nand ( n68916 , n68914 , n68915 );
buf ( n68917 , n68916 );
not ( n68918 , n68917 );
or ( n68919 , n68913 , n68918 );
nand ( n68920 , n68919 , n46907 );
nand ( n68921 , n68898 , n68911 , n68920 );
and ( n68922 , n68843 , n68921 );
nand ( n68923 , n68911 , n68920 );
and ( n68924 , n68923 , n68897 );
nor ( n68925 , n68922 , n68924 );
nand ( n68926 , n68833 , n68925 );
not ( n68927 , n68926 );
not ( n68928 , n44496 );
not ( n68929 , n67377 );
or ( n68930 , n68928 , n68929 );
buf ( n68931 , n68700 );
buf ( n68932 , n44517 );
nand ( n68933 , n68931 , n68932 );
buf ( n68934 , n68933 );
nand ( n68935 , n68930 , n68934 );
not ( n68936 , n68935 );
not ( n68937 , n67669 );
not ( n68938 , n67673 );
not ( n68939 , n68938 );
or ( n68940 , n68937 , n68939 );
nand ( n68941 , n67673 , n67666 );
nand ( n68942 , n68940 , n68941 );
and ( n68943 , n68942 , n67723 );
not ( n68944 , n68942 );
not ( n68945 , n67723 );
and ( n68946 , n68944 , n68945 );
nor ( n68947 , n68943 , n68946 );
not ( n68948 , n68947 );
nand ( n68949 , n68936 , n68948 );
not ( n68950 , n68949 );
not ( n68951 , n52174 );
not ( n68952 , n67446 );
not ( n68953 , n68952 );
or ( n68954 , n68951 , n68953 );
buf ( n68955 , n51004 );
not ( n68956 , n68955 );
buf ( n68957 , n45069 );
not ( n68958 , n68957 );
or ( n68959 , n68956 , n68958 );
buf ( n68960 , n42411 );
buf ( n68961 , n51001 );
nand ( n68962 , n68960 , n68961 );
buf ( n68963 , n68962 );
buf ( n68964 , n68963 );
nand ( n68965 , n68959 , n68964 );
buf ( n68966 , n68965 );
nand ( n68967 , n68966 , n38404 );
nand ( n68968 , n68954 , n68967 );
not ( n68969 , n68968 );
or ( n68970 , n68950 , n68969 );
nand ( n68971 , n68947 , n68935 );
nand ( n68972 , n68970 , n68971 );
not ( n68973 , n68972 );
or ( n68974 , n68927 , n68973 );
not ( n68975 , n68925 );
nand ( n68976 , n68975 , n68832 );
nand ( n68977 , n68974 , n68976 );
buf ( n68978 , n68977 );
buf ( n68979 , n68978 );
buf ( n68980 , n68979 );
and ( n68981 , n68812 , n68980 );
nor ( n68982 , n68808 , n68981 );
buf ( n68983 , n68982 );
not ( n68984 , n68983 );
buf ( n68985 , n68984 );
buf ( n68986 , n68985 );
not ( n68987 , n68986 );
or ( n68988 , n68794 , n68987 );
buf ( n68989 , n68789 );
not ( n68990 , n68989 );
buf ( n68991 , n68982 );
not ( n68992 , n68991 );
or ( n68993 , n68990 , n68992 );
xor ( n68994 , n66993 , n66996 );
xor ( n68995 , n68994 , n67022 );
buf ( n68996 , n68995 );
buf ( n68997 , n68996 );
not ( n68998 , n68997 );
buf ( n68999 , n68998 );
buf ( n69000 , n68999 );
not ( n69001 , n69000 );
buf ( n69002 , n67294 );
not ( n69003 , n69002 );
buf ( n69004 , n41973 );
not ( n69005 , n69004 );
and ( n69006 , n69003 , n69005 );
buf ( n69007 , n43766 );
buf ( n69008 , n53539 );
not ( n69009 , n69008 );
buf ( n69010 , n37472 );
not ( n69011 , n69010 );
or ( n69012 , n69009 , n69011 );
buf ( n69013 , n41981 );
buf ( n69014 , n53548 );
nand ( n69015 , n69013 , n69014 );
buf ( n69016 , n69015 );
buf ( n69017 , n69016 );
nand ( n69018 , n69012 , n69017 );
buf ( n69019 , n69018 );
buf ( n69020 , n69019 );
and ( n69021 , n69007 , n69020 );
nor ( n69022 , n69006 , n69021 );
buf ( n69023 , n69022 );
not ( n69024 , n69023 );
buf ( n69025 , n12481 );
buf ( n69026 , n43813 );
and ( n69027 , n69025 , n69026 );
not ( n69028 , n69025 );
buf ( n69029 , n41890 );
and ( n69030 , n69028 , n69029 );
nor ( n69031 , n69027 , n69030 );
buf ( n69032 , n69031 );
buf ( n69033 , n69032 );
not ( n69034 , n69033 );
buf ( n69035 , n37872 );
not ( n69036 , n69035 );
or ( n69037 , n69034 , n69036 );
buf ( n69038 , n67314 );
not ( n69039 , n69038 );
buf ( n69040 , n42175 );
nand ( n69041 , n69039 , n69040 );
buf ( n69042 , n69041 );
buf ( n69043 , n69042 );
nand ( n69044 , n69037 , n69043 );
buf ( n69045 , n69044 );
buf ( n69046 , n69045 );
not ( n69047 , n69046 );
buf ( n69048 , n69047 );
not ( n69049 , n69048 );
and ( n69050 , n69024 , n69049 );
buf ( n69051 , n69023 );
buf ( n69052 , n69048 );
nand ( n69053 , n69051 , n69052 );
buf ( n69054 , n69053 );
not ( n69055 , n68012 );
nand ( n69056 , n69055 , n68119 );
not ( n69057 , n69056 );
not ( n69058 , n68091 );
or ( n69059 , n69057 , n69058 );
buf ( n69060 , n68116 );
buf ( n69061 , n68012 );
nand ( n69062 , n69060 , n69061 );
buf ( n69063 , n69062 );
nand ( n69064 , n69059 , n69063 );
and ( n69065 , n69054 , n69064 );
nor ( n69066 , n69050 , n69065 );
buf ( n69067 , n69066 );
not ( n69068 , n69067 );
or ( n69069 , n69001 , n69068 );
xor ( n69070 , n67632 , n67733 );
xnor ( n69071 , n69070 , n67647 );
buf ( n69072 , n69071 );
not ( n69073 , n69072 );
buf ( n69074 , n69073 );
buf ( n69075 , n69074 );
not ( n69076 , n69075 );
buf ( n69077 , n46912 );
not ( n69078 , n69077 );
buf ( n69079 , n67416 );
not ( n69080 , n69079 );
or ( n69081 , n69078 , n69080 );
buf ( n69082 , n68910 );
buf ( n69083 , n46907 );
nand ( n69084 , n69082 , n69083 );
buf ( n69085 , n69084 );
buf ( n69086 , n69085 );
nand ( n69087 , n69081 , n69086 );
buf ( n69088 , n69087 );
buf ( n69089 , n69088 );
not ( n69090 , n69089 );
or ( n69091 , n69076 , n69090 );
buf ( n69092 , n69088 );
not ( n69093 , n69092 );
buf ( n69094 , n69093 );
buf ( n69095 , n69094 );
not ( n69096 , n69095 );
buf ( n69097 , n69071 );
not ( n69098 , n69097 );
or ( n69099 , n69096 , n69098 );
buf ( n69100 , n46117 );
not ( n69101 , n69100 );
buf ( n69102 , n52670 );
not ( n69103 , n69102 );
or ( n69104 , n69101 , n69103 );
buf ( n69105 , n25159 );
buf ( n69106 , n46126 );
nand ( n69107 , n69105 , n69106 );
buf ( n69108 , n69107 );
buf ( n69109 , n69108 );
nand ( n69110 , n69104 , n69109 );
buf ( n69111 , n69110 );
buf ( n69112 , n69111 );
not ( n69113 , n69112 );
buf ( n69114 , n50128 );
not ( n69115 , n69114 );
or ( n69116 , n69113 , n69115 );
buf ( n69117 , n47872 );
buf ( n69118 , n67473 );
nand ( n69119 , n69117 , n69118 );
buf ( n69120 , n69119 );
buf ( n69121 , n69120 );
nand ( n69122 , n69116 , n69121 );
buf ( n69123 , n69122 );
not ( n69124 , n69123 );
buf ( n69125 , n68641 );
not ( n69126 , n69125 );
buf ( n69127 , n69126 );
buf ( n69128 , n69127 );
not ( n69129 , n69128 );
buf ( n69130 , n61454 );
not ( n69131 , n69130 );
or ( n69132 , n69129 , n69131 );
buf ( n69133 , n67687 );
buf ( n69134 , n62582 );
nand ( n69135 , n69133 , n69134 );
buf ( n69136 , n69135 );
buf ( n69137 , n69136 );
nand ( n69138 , n69132 , n69137 );
buf ( n69139 , n69138 );
or ( n69140 , n68591 , n68594 );
not ( n69141 , n69140 );
not ( n69142 , n68161 );
or ( n69143 , n69141 , n69142 );
nand ( n69144 , n68591 , n68594 );
nand ( n69145 , n69143 , n69144 );
xor ( n69146 , n69139 , n69145 );
buf ( n69147 , n42315 );
not ( n69148 , n69147 );
buf ( n69149 , n68039 );
not ( n69150 , n69149 );
or ( n69151 , n69148 , n69150 );
and ( n69152 , n13653 , n42260 );
not ( n69153 , n13653 );
and ( n69154 , n69153 , n59242 );
or ( n69155 , n69152 , n69154 );
buf ( n69156 , n69155 );
buf ( n69157 , n42252 );
nand ( n69158 , n69156 , n69157 );
buf ( n69159 , n69158 );
buf ( n69160 , n69159 );
nand ( n69161 , n69151 , n69160 );
buf ( n69162 , n69161 );
and ( n69163 , n69146 , n69162 );
and ( n69164 , n69139 , n69145 );
or ( n69165 , n69163 , n69164 );
not ( n69166 , n69165 );
or ( n69167 , n69124 , n69166 );
buf ( n69168 , n69165 );
not ( n69169 , n69168 );
buf ( n69170 , n69169 );
not ( n69171 , n69170 );
buf ( n69172 , n69123 );
not ( n69173 , n69172 );
buf ( n69174 , n69173 );
not ( n69175 , n69174 );
or ( n69176 , n69171 , n69175 );
xor ( n69177 , n67716 , n67699 );
xnor ( n69178 , n69177 , n67721 );
buf ( n69179 , n69178 );
not ( n69180 , n69179 );
buf ( n69181 , n69180 );
nand ( n69182 , n69176 , n69181 );
nand ( n69183 , n69167 , n69182 );
buf ( n69184 , n69183 );
buf ( n69185 , n46225 );
not ( n69186 , n69185 );
buf ( n69187 , n45747 );
buf ( n69188 , n44025 );
and ( n69189 , n69187 , n69188 );
not ( n69190 , n69187 );
buf ( n69191 , n28305 );
and ( n69192 , n69190 , n69191 );
nor ( n69193 , n69189 , n69192 );
buf ( n69194 , n69193 );
buf ( n69195 , n69194 );
not ( n69196 , n69195 );
or ( n69197 , n69186 , n69196 );
nand ( n69198 , n67172 , n67149 );
buf ( n69199 , n69198 );
nand ( n69200 , n69197 , n69199 );
buf ( n69201 , n69200 );
buf ( n69202 , n69201 );
xor ( n69203 , n69184 , n69202 );
buf ( n69204 , n41908 );
buf ( n69205 , n56325 );
nor ( n69206 , n69204 , n69205 );
buf ( n69207 , n69206 );
buf ( n69208 , n69207 );
and ( n69209 , n69203 , n69208 );
and ( n69210 , n69184 , n69202 );
or ( n69211 , n69209 , n69210 );
buf ( n69212 , n69211 );
buf ( n69213 , n69212 );
nand ( n69214 , n69099 , n69213 );
buf ( n69215 , n69214 );
buf ( n69216 , n69215 );
nand ( n69217 , n69091 , n69216 );
buf ( n69218 , n69217 );
buf ( n69219 , n69218 );
nand ( n69220 , n69069 , n69219 );
buf ( n69221 , n69220 );
buf ( n69222 , n69221 );
buf ( n69223 , n68999 );
not ( n69224 , n69223 );
buf ( n69225 , n69066 );
not ( n69226 , n69225 );
buf ( n69227 , n69226 );
buf ( n69228 , n69227 );
nand ( n69229 , n69224 , n69228 );
buf ( n69230 , n69229 );
buf ( n69231 , n69230 );
nand ( n69232 , n69222 , n69231 );
buf ( n69233 , n69232 );
buf ( n69234 , n69233 );
nand ( n69235 , n68993 , n69234 );
buf ( n69236 , n69235 );
buf ( n69237 , n69236 );
nand ( n69238 , n68988 , n69237 );
buf ( n69239 , n69238 );
buf ( n69240 , n69239 );
not ( n69241 , n69240 );
buf ( n69242 , n69241 );
buf ( n69243 , n69242 );
not ( n69244 , n69243 );
buf ( n69245 , n69244 );
and ( n69246 , n68776 , n69245 );
nor ( n69247 , n68772 , n69246 );
buf ( n69248 , n69247 );
and ( n69249 , n67944 , n69248 );
and ( n69250 , n67936 , n67943 );
or ( n69251 , n69249 , n69250 );
buf ( n69252 , n69251 );
buf ( n69253 , n69252 );
xor ( n69254 , n67929 , n69253 );
not ( n69255 , n67761 );
buf ( n69256 , n67112 );
not ( n69257 , n69256 );
buf ( n69258 , n69257 );
not ( n69259 , n69258 );
or ( n69260 , n69255 , n69259 );
not ( n69261 , n67761 );
nand ( n69262 , n69261 , n67112 );
nand ( n69263 , n69260 , n69262 );
xor ( n69264 , n69263 , n67857 );
buf ( n69265 , n69264 );
and ( n69266 , n69254 , n69265 );
and ( n69267 , n67929 , n69253 );
or ( n69268 , n69266 , n69267 );
buf ( n69269 , n69268 );
nand ( n69270 , n67907 , n69269 );
buf ( n69271 , n69270 );
xor ( n69272 , n67929 , n69253 );
xor ( n69273 , n69272 , n69265 );
buf ( n69274 , n69273 );
buf ( n69275 , n69274 );
not ( n69276 , n67782 );
buf ( n69277 , n67765 );
not ( n69278 , n69277 );
buf ( n69279 , n69278 );
not ( n69280 , n69279 );
or ( n69281 , n69276 , n69280 );
nand ( n69282 , n67765 , n67781 );
nand ( n69283 , n69281 , n69282 );
buf ( n69284 , n69283 );
buf ( n69285 , n67855 );
not ( n69286 , n69285 );
buf ( n69287 , n69286 );
buf ( n69288 , n69287 );
and ( n69289 , n69284 , n69288 );
not ( n69290 , n69284 );
buf ( n69291 , n67855 );
and ( n69292 , n69290 , n69291 );
nor ( n69293 , n69289 , n69292 );
buf ( n69294 , n69293 );
buf ( n69295 , n69294 );
buf ( n69296 , n68769 );
buf ( n69297 , n69239 );
and ( n69298 , n69296 , n69297 );
not ( n69299 , n69296 );
buf ( n69300 , n69242 );
and ( n69301 , n69299 , n69300 );
nor ( n69302 , n69298 , n69301 );
buf ( n69303 , n69302 );
buf ( n69304 , n69303 );
buf ( n69305 , n68760 );
and ( n69306 , n69304 , n69305 );
not ( n69307 , n69304 );
buf ( n69308 , n68763 );
and ( n69309 , n69307 , n69308 );
nor ( n69310 , n69306 , n69309 );
buf ( n69311 , n69310 );
buf ( n69312 , n69311 );
xor ( n69313 , n67806 , n67847 );
xor ( n69314 , n69313 , n67851 );
buf ( n69315 , n69314 );
not ( n69316 , n69315 );
buf ( n69317 , n69316 );
buf ( n69318 , n67771 );
buf ( n69319 , n67768 );
xor ( n69320 , n69318 , n69319 );
buf ( n69321 , n67779 );
xnor ( n69322 , n69320 , n69321 );
buf ( n69323 , n69322 );
buf ( n69324 , n69323 );
nand ( n69325 , n69317 , n69324 );
buf ( n69326 , n69325 );
buf ( n69327 , n69326 );
nand ( n69328 , n69312 , n69327 );
buf ( n69329 , n69328 );
buf ( n69330 , n69329 );
buf ( n69331 , n69316 );
buf ( n69332 , n69323 );
or ( n69333 , n69331 , n69332 );
buf ( n69334 , n69333 );
buf ( n69335 , n69334 );
and ( n69336 , n69330 , n69335 );
buf ( n69337 , n69336 );
buf ( n69338 , n69337 );
xor ( n69339 , n69295 , n69338 );
xor ( n69340 , n67936 , n67943 );
xor ( n69341 , n69340 , n69248 );
buf ( n69342 , n69341 );
buf ( n69343 , n69342 );
and ( n69344 , n69339 , n69343 );
and ( n69345 , n69295 , n69338 );
or ( n69346 , n69344 , n69345 );
buf ( n69347 , n69346 );
buf ( n69348 , n69347 );
nand ( n69349 , n69275 , n69348 );
buf ( n69350 , n69349 );
buf ( n69351 , n69350 );
xor ( n69352 , n69295 , n69338 );
xor ( n69353 , n69352 , n69343 );
buf ( n69354 , n69353 );
buf ( n69355 , n69354 );
xor ( n69356 , n69323 , n69315 );
xnor ( n69357 , n69356 , n69311 );
buf ( n69358 , n69357 );
buf ( n69359 , n69358 );
buf ( n69360 , n69359 );
buf ( n69361 , n69360 );
not ( n69362 , n67808 );
not ( n69363 , n67844 );
nand ( n69364 , n69362 , n69363 , C1 );
nand ( n69365 , n67808 , n67844 , C1 );
nand ( n69366 , n69364 , n69365 , C1 , C1 );
xor ( n69367 , n67146 , n67175 );
xor ( n69368 , n69367 , n67180 );
buf ( n69369 , n69368 );
buf ( n69370 , n69369 );
buf ( n69371 , C0 );
buf ( n69372 , n69371 );
xor ( n69373 , n69370 , n69372 );
buf ( n69374 , n55841 );
not ( n69375 , n69374 );
buf ( n69376 , n41982 );
not ( n69377 , n69376 );
or ( n69378 , n69375 , n69377 );
buf ( n69379 , n37473 );
buf ( n69380 , n55840 );
nand ( n69381 , n69379 , n69380 );
buf ( n69382 , n69381 );
buf ( n69383 , n69382 );
nand ( n69384 , n69378 , n69383 );
buf ( n69385 , n69384 );
buf ( n69386 , n69385 );
not ( n69387 , n69386 );
buf ( n69388 , n41966 );
not ( n69389 , n69388 );
or ( n69390 , n69387 , n69389 );
buf ( n69391 , n69019 );
buf ( n69392 , n44253 );
nand ( n69393 , n69391 , n69392 );
buf ( n69394 , n69393 );
buf ( n69395 , n69394 );
nand ( n69396 , n69390 , n69395 );
buf ( n69397 , n69396 );
buf ( n69398 , n69397 );
buf ( n69399 , n48855 );
not ( n69400 , n69399 );
and ( n69401 , n48808 , n44989 );
not ( n69402 , n48808 );
and ( n69403 , n69402 , n30187 );
or ( n69404 , n69401 , n69403 );
buf ( n69405 , n69404 );
not ( n69406 , n69405 );
or ( n69407 , n69400 , n69406 );
buf ( n69408 , n68827 );
buf ( n69409 , n48868 );
nand ( n69410 , n69408 , n69409 );
buf ( n69411 , n69410 );
buf ( n69412 , n69411 );
nand ( n69413 , n69407 , n69412 );
buf ( n69414 , n69413 );
buf ( n69415 , n69414 );
xor ( n69416 , n69398 , n69415 );
buf ( n69417 , n43442 );
not ( n69418 , n69417 );
buf ( n69419 , n37437 );
not ( n69420 , n69419 );
or ( n69421 , n69418 , n69420 );
buf ( n69422 , n12481 );
nand ( n69423 , n69421 , n69422 );
buf ( n69424 , n69423 );
buf ( n69425 , n69424 );
buf ( n69426 , n41843 );
buf ( n69427 , n37437 );
not ( n69428 , n69427 );
buf ( n69429 , n41779 );
nand ( n69430 , n69428 , n69429 );
buf ( n69431 , n69430 );
buf ( n69432 , n69431 );
nand ( n69433 , n69425 , n69426 , n69432 );
buf ( n69434 , n69433 );
buf ( n69435 , n69434 );
not ( n69436 , n69435 );
buf ( n69437 , n69436 );
buf ( n69438 , n69437 );
not ( n69439 , n69438 );
buf ( n69440 , n67149 );
not ( n69441 , n69440 );
buf ( n69442 , n69194 );
not ( n69443 , n69442 );
or ( n69444 , n69441 , n69443 );
not ( n69445 , n41817 );
not ( n69446 , n45747 );
and ( n69447 , n29323 , n69446 );
not ( n69448 , n29323 );
not ( n69449 , n53492 );
and ( n69450 , n69448 , n69449 );
or ( n69451 , n69447 , n69450 );
and ( n69452 , n69445 , n69451 );
not ( n69453 , n69445 );
not ( n69454 , n45747 );
and ( n69455 , n29313 , n69454 );
not ( n69456 , n29313 );
not ( n69457 , n53492 );
and ( n69458 , n69456 , n69457 );
or ( n69459 , n69455 , n69458 );
and ( n69460 , n69453 , n69459 );
or ( n69461 , n69452 , n69460 );
nand ( n69462 , n69461 , n46225 );
buf ( n69463 , n69462 );
nand ( n69464 , n69444 , n69463 );
buf ( n69465 , n69464 );
buf ( n69466 , n69465 );
not ( n69467 , n69466 );
or ( n69468 , n69439 , n69467 );
buf ( n69469 , n69434 );
not ( n69470 , n69469 );
buf ( n69471 , n69465 );
not ( n69472 , n69471 );
buf ( n69473 , n69472 );
buf ( n69474 , n69473 );
not ( n69475 , n69474 );
or ( n69476 , n69470 , n69475 );
not ( n69477 , n44496 );
not ( n69478 , n68715 );
or ( n69479 , n69477 , n69478 );
not ( n69480 , n46657 );
not ( n69481 , n65010 );
or ( n69482 , n69480 , n69481 );
or ( n69483 , n53579 , n65010 );
nand ( n69484 , n69482 , n69483 );
nand ( n69485 , n69484 , n44517 );
nand ( n69486 , n69479 , n69485 );
not ( n69487 , n43868 );
not ( n69488 , n68872 );
or ( n69489 , n69487 , n69488 );
buf ( n69490 , n41605 );
not ( n69491 , n69490 );
buf ( n69492 , n42072 );
not ( n69493 , n69492 );
or ( n69494 , n69491 , n69493 );
buf ( n69495 , n28368 );
buf ( n69496 , n41604 );
nand ( n69497 , n69495 , n69496 );
buf ( n69498 , n69497 );
buf ( n69499 , n69498 );
nand ( n69500 , n69494 , n69499 );
buf ( n69501 , n69500 );
buf ( n69502 , n69501 );
buf ( n69503 , n41596 );
nand ( n69504 , n69502 , n69503 );
buf ( n69505 , n69504 );
nand ( n69506 , n69489 , n69505 );
or ( n69507 , n69486 , n69506 );
xor ( n69508 , n69139 , n69145 );
xor ( n69509 , n69508 , n69162 );
nand ( n69510 , n69507 , n69509 );
buf ( n69511 , n69510 );
buf ( n69512 , n69486 );
buf ( n69513 , n69506 );
nand ( n69514 , n69512 , n69513 );
buf ( n69515 , n69514 );
buf ( n69516 , n69515 );
and ( n69517 , n69511 , n69516 );
buf ( n69518 , n69517 );
buf ( n69519 , n69518 );
not ( n69520 , n69519 );
buf ( n69521 , n69520 );
buf ( n69522 , n69521 );
nand ( n69523 , n69476 , n69522 );
buf ( n69524 , n69523 );
buf ( n69525 , n69524 );
nand ( n69526 , n69468 , n69525 );
buf ( n69527 , n69526 );
buf ( n69528 , n69527 );
and ( n69529 , n69416 , n69528 );
and ( n69530 , n69398 , n69415 );
or ( n69531 , n69529 , n69530 );
buf ( n69532 , n69531 );
buf ( n69533 , n69532 );
and ( n69534 , n69373 , n69533 );
or ( n69535 , n69534 , C0 );
buf ( n69536 , n69535 );
buf ( n69537 , n69536 );
not ( n69538 , n69537 );
xor ( n69539 , n67812 , n67815 );
xor ( n69540 , n69539 , n67841 );
buf ( n69541 , n69540 );
buf ( n69542 , n69541 );
buf ( n69543 , n69542 );
buf ( n69544 , n69543 );
buf ( n69545 , n69544 );
not ( n69546 , n69545 );
or ( n69547 , n69538 , n69546 );
buf ( n69548 , n69544 );
buf ( n69549 , n69536 );
or ( n69550 , n69548 , n69549 );
buf ( n69551 , n68996 );
buf ( n69552 , n69218 );
xor ( n69553 , n69551 , n69552 );
buf ( n69554 , n69227 );
xor ( n69555 , n69553 , n69554 );
buf ( n69556 , n69555 );
buf ( n69557 , n69556 );
nand ( n69558 , n69550 , n69557 );
buf ( n69559 , n69558 );
buf ( n69560 , n69559 );
nand ( n69561 , n69547 , n69560 );
buf ( n69562 , n69561 );
xor ( n69563 , n69366 , n69562 );
buf ( n69564 , n62125 );
not ( n69565 , n69564 );
buf ( n69566 , n67830 );
not ( n69567 , n69566 );
or ( n69568 , n69565 , n69567 );
not ( n69569 , n51493 );
not ( n69570 , n39489 );
or ( n69571 , n69569 , n69570 );
nand ( n69572 , n44157 , n48836 );
nand ( n69573 , n69571 , n69572 );
buf ( n69574 , n69573 );
buf ( n69575 , n51488 );
nand ( n69576 , n69574 , n69575 );
buf ( n69577 , n69576 );
buf ( n69578 , n69577 );
nand ( n69579 , n69568 , n69578 );
buf ( n69580 , n69579 );
buf ( n69581 , n69580 );
buf ( n69582 , n69064 );
buf ( n69583 , n69045 );
xor ( n69584 , n69582 , n69583 );
buf ( n69585 , n69023 );
xnor ( n69586 , n69584 , n69585 );
buf ( n69587 , n69586 );
buf ( n69588 , n69587 );
xor ( n69589 , n69581 , n69588 );
buf ( n69590 , n68863 );
not ( n69591 , n69590 );
buf ( n69592 , n68883 );
not ( n69593 , n69592 );
or ( n69594 , n69591 , n69593 );
buf ( n69595 , n68874 );
buf ( n69596 , n68879 );
nand ( n69597 , n69595 , n69596 );
buf ( n69598 , n69597 );
buf ( n69599 , n69598 );
nand ( n69600 , n69594 , n69599 );
buf ( n69601 , n69600 );
buf ( n69602 , n69601 );
buf ( n69603 , n68895 );
not ( n69604 , n69603 );
buf ( n69605 , n69604 );
buf ( n69606 , n69605 );
and ( n69607 , n69602 , n69606 );
not ( n69608 , n69602 );
buf ( n69609 , n68895 );
and ( n69610 , n69608 , n69609 );
nor ( n69611 , n69607 , n69610 );
buf ( n69612 , n69611 );
buf ( n69613 , n69612 );
not ( n69614 , n69613 );
buf ( n69615 , n69614 );
not ( n69616 , n69615 );
buf ( n69617 , n46875 );
buf ( n69618 , n41763 );
and ( n69619 , n69617 , n69618 );
not ( n69620 , n69617 );
buf ( n69621 , n41762 );
and ( n69622 , n69620 , n69621 );
nor ( n69623 , n69619 , n69622 );
buf ( n69624 , n69623 );
not ( n69625 , n69624 );
not ( n69626 , n46910 );
and ( n69627 , n69625 , n69626 );
nand ( n69628 , n68917 , n68912 );
and ( n69629 , n69628 , n46912 );
nor ( n69630 , n69627 , n69629 );
buf ( n69631 , n69630 );
not ( n69632 , n69631 );
buf ( n69633 , n69632 );
not ( n69634 , n69633 );
or ( n69635 , n69616 , n69634 );
not ( n69636 , n69630 );
not ( n69637 , n69612 );
or ( n69638 , n69636 , n69637 );
buf ( n69639 , n69170 );
not ( n69640 , n69639 );
buf ( n69641 , n69181 );
not ( n69642 , n69641 );
or ( n69643 , n69640 , n69642 );
buf ( n69644 , n69178 );
buf ( n69645 , n69165 );
nand ( n69646 , n69644 , n69645 );
buf ( n69647 , n69646 );
buf ( n69648 , n69647 );
nand ( n69649 , n69643 , n69648 );
buf ( n69650 , n69649 );
and ( n69651 , n69650 , n69174 );
not ( n69652 , n69650 );
and ( n69653 , n69652 , n69123 );
nor ( n69654 , n69651 , n69653 );
buf ( n69655 , n69654 );
not ( n69656 , n69655 );
buf ( n69657 , n69656 );
nand ( n69658 , n69638 , n69657 );
nand ( n69659 , n69635 , n69658 );
buf ( n69660 , n48323 );
not ( n69661 , n69660 );
buf ( n69662 , n55743 );
not ( n69663 , n69662 );
or ( n69664 , n69661 , n69663 );
buf ( n69665 , n50591 );
buf ( n69666 , n48320 );
nand ( n69667 , n69665 , n69666 );
buf ( n69668 , n69667 );
buf ( n69669 , n69668 );
nand ( n69670 , n69664 , n69669 );
buf ( n69671 , n69670 );
buf ( n69672 , n69671 );
not ( n69673 , n69672 );
buf ( n69674 , n52537 );
not ( n69675 , n69674 );
or ( n69676 , n69673 , n69675 );
buf ( n69677 , n68856 );
buf ( n69678 , n48975 );
nand ( n69679 , n69677 , n69678 );
buf ( n69680 , n69679 );
buf ( n69681 , n69680 );
nand ( n69682 , n69676 , n69681 );
buf ( n69683 , n69682 );
not ( n69684 , n69683 );
buf ( n69685 , n46390 );
not ( n69686 , n69685 );
buf ( n69687 , n52670 );
not ( n69688 , n69687 );
or ( n69689 , n69686 , n69688 );
buf ( n69690 , n25159 );
buf ( n69691 , n46393 );
nand ( n69692 , n69690 , n69691 );
buf ( n69693 , n69692 );
buf ( n69694 , n69693 );
nand ( n69695 , n69689 , n69694 );
buf ( n69696 , n69695 );
buf ( n69697 , n69696 );
not ( n69698 , n69697 );
buf ( n69699 , n42628 );
not ( n69700 , n69699 );
or ( n69701 , n69698 , n69700 );
buf ( n69702 , n69111 );
buf ( n69703 , n42564 );
nand ( n69704 , n69702 , n69703 );
buf ( n69705 , n69704 );
buf ( n69706 , n69705 );
nand ( n69707 , n69701 , n69706 );
buf ( n69708 , n69707 );
not ( n69709 , n69708 );
or ( n69710 , n69684 , n69709 );
buf ( n69711 , n69708 );
buf ( n69712 , n69683 );
nor ( n69713 , n69711 , n69712 );
buf ( n69714 , n69713 );
buf ( n69715 , n46117 );
not ( n69716 , n69715 );
buf ( n69717 , n52725 );
not ( n69718 , n69717 );
or ( n69719 , n69716 , n69718 );
buf ( n69720 , n25182 );
buf ( n69721 , n46126 );
nand ( n69722 , n69720 , n69721 );
buf ( n69723 , n69722 );
buf ( n69724 , n69723 );
nand ( n69725 , n69719 , n69724 );
buf ( n69726 , n69725 );
buf ( n69727 , n69726 );
not ( n69728 , n69727 );
buf ( n69729 , n43935 );
not ( n69730 , n69729 );
or ( n69731 , n69728 , n69730 );
buf ( n69732 , n68126 );
buf ( n69733 , n43905 );
nand ( n69734 , n69732 , n69733 );
buf ( n69735 , n69734 );
buf ( n69736 , n69735 );
nand ( n69737 , n69731 , n69736 );
buf ( n69738 , n69737 );
buf ( n69739 , n69738 );
buf ( n69740 , n69155 );
buf ( n69741 , n42309 );
and ( n69742 , n69740 , n69741 );
buf ( n69743 , n59242 );
not ( n69744 , n69743 );
buf ( n69745 , n60330 );
not ( n69746 , n69745 );
or ( n69747 , n69744 , n69746 );
buf ( n69748 , n60327 );
buf ( n69749 , n42260 );
nand ( n69750 , n69748 , n69749 );
buf ( n69751 , n69750 );
buf ( n69752 , n69751 );
nand ( n69753 , n69747 , n69752 );
buf ( n69754 , n69753 );
and ( n69755 , n69754 , n42246 );
buf ( n69756 , n69755 );
nor ( n69757 , n69742 , n69756 );
buf ( n69758 , n69757 );
buf ( n69759 , n69758 );
not ( n69760 , n69759 );
buf ( n69761 , n69760 );
buf ( n69762 , n69761 );
or ( n69763 , n69739 , n69762 );
and ( n69764 , n68571 , n68589 );
not ( n69765 , n68571 );
nor ( n69766 , n68575 , n68585 );
and ( n69767 , n69765 , n69766 );
nor ( n69768 , n69764 , n69767 );
and ( n69769 , n68571 , n68586 );
not ( n69770 , n68571 );
nand ( n69771 , n68575 , n68585 );
and ( n69772 , n69770 , n69771 );
or ( n69773 , n69769 , n69772 );
nand ( n69774 , n69768 , n69773 );
buf ( n69775 , n69774 );
and ( n69776 , n28430 , n62510 );
not ( n69777 , n28430 );
and ( n69778 , n69777 , n25226 );
or ( n69779 , n69776 , n69778 );
buf ( n69780 , n69779 );
not ( n69781 , n69780 );
buf ( n69782 , n46047 );
not ( n69783 , n69782 );
or ( n69784 , n69781 , n69783 );
buf ( n69785 , n68613 );
buf ( n69786 , n42665 );
nand ( n69787 , n69785 , n69786 );
buf ( n69788 , n69787 );
buf ( n69789 , n69788 );
nand ( n69790 , n69784 , n69789 );
buf ( n69791 , n69790 );
buf ( n69792 , n69791 );
xor ( n69793 , n69775 , n69792 );
buf ( n69794 , n42856 );
not ( n69795 , n69794 );
buf ( n69796 , n42366 );
not ( n69797 , n69796 );
buf ( n69798 , n69797 );
buf ( n69799 , n69798 );
not ( n69800 , n69799 );
or ( n69801 , n69795 , n69800 );
buf ( n69802 , n63913 );
not ( n69803 , n69802 );
buf ( n69804 , n69803 );
buf ( n69805 , n69804 );
buf ( n69806 , n42862 );
nand ( n69807 , n69805 , n69806 );
buf ( n69808 , n69807 );
buf ( n69809 , n69808 );
nand ( n69810 , n69801 , n69809 );
buf ( n69811 , n69810 );
buf ( n69812 , n69811 );
not ( n69813 , n69812 );
buf ( n69814 , n66459 );
not ( n69815 , n69814 );
or ( n69816 , n69813 , n69815 );
buf ( n69817 , n66482 );
buf ( n69818 , n68157 );
nand ( n69819 , n69817 , n69818 );
buf ( n69820 , n69819 );
buf ( n69821 , n69820 );
nand ( n69822 , n69816 , n69821 );
buf ( n69823 , n69822 );
buf ( n69824 , n69823 );
and ( n69825 , n69793 , n69824 );
and ( n69826 , n69775 , n69792 );
or ( n69827 , n69825 , n69826 );
buf ( n69828 , n69827 );
buf ( n69829 , n69828 );
nand ( n69830 , n69763 , n69829 );
buf ( n69831 , n69830 );
buf ( n69832 , n69831 );
buf ( n69833 , n69738 );
buf ( n69834 , n69761 );
nand ( n69835 , n69833 , n69834 );
buf ( n69836 , n69835 );
buf ( n69837 , n69836 );
and ( n69838 , n69832 , n69837 );
buf ( n69839 , n69838 );
or ( n69840 , n69714 , n69839 );
nand ( n69841 , n69710 , n69840 );
buf ( n69842 , n69841 );
buf ( n69843 , n56289 );
not ( n69844 , n69843 );
buf ( n69845 , n38412 );
not ( n69846 , n69845 );
or ( n69847 , n69844 , n69846 );
buf ( n69848 , n48984 );
buf ( n69849 , n52094 );
nand ( n69850 , n69848 , n69849 );
buf ( n69851 , n69850 );
buf ( n69852 , n69851 );
nand ( n69853 , n69847 , n69852 );
buf ( n69854 , n69853 );
buf ( n69855 , n69854 );
not ( n69856 , n69855 );
buf ( n69857 , n44042 );
not ( n69858 , n69857 );
or ( n69859 , n69856 , n69858 );
buf ( n69860 , n68966 );
buf ( n69861 , n38380 );
nand ( n69862 , n69860 , n69861 );
buf ( n69863 , n69862 );
buf ( n69864 , n69863 );
nand ( n69865 , n69859 , n69864 );
buf ( n69866 , n69865 );
buf ( n69867 , n69866 );
xor ( n69868 , n69842 , n69867 );
buf ( n69869 , n53539 );
not ( n69870 , n69869 );
buf ( n69871 , n37328 );
not ( n69872 , n69871 );
or ( n69873 , n69870 , n69872 );
buf ( n69874 , n43434 );
buf ( n69875 , n53548 );
nand ( n69876 , n69874 , n69875 );
buf ( n69877 , n69876 );
buf ( n69878 , n69877 );
nand ( n69879 , n69873 , n69878 );
buf ( n69880 , n69879 );
buf ( n69881 , n69880 );
not ( n69882 , n69881 );
buf ( n69883 , n37400 );
not ( n69884 , n69883 );
or ( n69885 , n69882 , n69884 );
buf ( n69886 , n67975 );
buf ( n69887 , n42135 );
nand ( n69888 , n69886 , n69887 );
buf ( n69889 , n69888 );
buf ( n69890 , n69889 );
nand ( n69891 , n69885 , n69890 );
buf ( n69892 , n69891 );
buf ( n69893 , n69892 );
and ( n69894 , n69868 , n69893 );
and ( n69895 , n69842 , n69867 );
or ( n69896 , n69894 , n69895 );
buf ( n69897 , n69896 );
xor ( n69898 , n69659 , n69897 );
xor ( n69899 , n69184 , n69202 );
xor ( n69900 , n69899 , n69208 );
buf ( n69901 , n69900 );
and ( n69902 , n69898 , n69901 );
and ( n69903 , n69659 , n69897 );
or ( n69904 , n69902 , n69903 );
buf ( n69905 , n69904 );
and ( n69906 , n69589 , n69905 );
and ( n69907 , n69581 , n69588 );
or ( n69908 , n69906 , n69907 );
buf ( n69909 , n69908 );
buf ( n69910 , n69909 );
xor ( n69911 , n68803 , n68977 );
xnor ( n69912 , n69911 , n68799 );
buf ( n69913 , n69912 );
xor ( n69914 , n69910 , n69913 );
xor ( n69915 , n69088 , n69071 );
xnor ( n69916 , n69915 , n69212 );
buf ( n69917 , n69916 );
not ( n69918 , n52456 );
not ( n69919 , n69573 );
or ( n69920 , n69918 , n69919 );
and ( n69921 , n39205 , n51493 );
not ( n69922 , n39205 );
and ( n69923 , n69922 , n61853 );
or ( n69924 , n69921 , n69923 );
nand ( n69925 , n69924 , n51488 );
nand ( n69926 , n69920 , n69925 );
not ( n69927 , n68968 );
and ( n69928 , n68948 , n68935 );
nand ( n69929 , n69927 , n69928 );
not ( n69930 , n68949 );
nand ( n69931 , n69930 , n68968 );
and ( n69932 , n68936 , n68947 );
nand ( n69933 , n69932 , n69927 );
nand ( n69934 , n68968 , n68947 , n68935 );
nand ( n69935 , n69929 , n69931 , n69933 , n69934 );
xor ( n69936 , n69926 , n69935 );
not ( n69937 , n68923 );
and ( n69938 , n68898 , n69937 );
not ( n69939 , n68898 );
and ( n69940 , n69939 , n68923 );
nor ( n69941 , n69938 , n69940 );
and ( n69942 , n69941 , n68843 );
not ( n69943 , n69941 );
not ( n69944 , n68843 );
and ( n69945 , n69943 , n69944 );
nor ( n69946 , n69942 , n69945 );
and ( n69947 , n69936 , n69946 );
and ( n69948 , n69926 , n69935 );
or ( n69949 , n69947 , n69948 );
buf ( n69950 , n69949 );
xor ( n69951 , n69917 , n69950 );
xor ( n69952 , n67959 , n67962 );
xor ( n69953 , n69952 , n68738 );
buf ( n69954 , n69953 );
buf ( n69955 , n69954 );
and ( n69956 , n69951 , n69955 );
and ( n69957 , n69917 , n69950 );
or ( n69958 , n69956 , n69957 );
buf ( n69959 , n69958 );
buf ( n69960 , n69959 );
and ( n69961 , n69914 , n69960 );
and ( n69962 , n69910 , n69913 );
or ( n69963 , n69961 , n69962 );
buf ( n69964 , n69963 );
and ( n69965 , n69563 , n69964 );
and ( n69966 , n69366 , n69562 );
or ( n69967 , n69965 , n69966 );
buf ( n69968 , n69967 );
buf ( n69969 , n69233 );
buf ( n69970 , n68792 );
xor ( n69971 , n69969 , n69970 );
buf ( n69972 , n68985 );
xor ( n69973 , n69971 , n69972 );
buf ( n69974 , n69973 );
buf ( n69975 , n69974 );
xor ( n69976 , n67948 , n68747 );
xor ( n69977 , n69976 , n68756 );
buf ( n69978 , n69977 );
buf ( n69979 , n69978 );
xor ( n69980 , n69975 , n69979 );
and ( n69981 , n68833 , n68972 );
not ( n69982 , n68833 );
not ( n69983 , n68972 );
and ( n69984 , n69982 , n69983 );
nor ( n69985 , n69981 , n69984 );
not ( n69986 , n68975 );
and ( n69987 , n69985 , n69986 );
not ( n69988 , n69985 );
and ( n69989 , n69988 , n68975 );
nor ( n69990 , n69987 , n69989 );
buf ( n69991 , n69990 );
not ( n69992 , n46851 );
buf ( n69993 , C0 );
buf ( n69994 , n69993 );
xor ( n69995 , n69991 , n69994 );
buf ( n69996 , n68120 );
not ( n69997 , n69996 );
buf ( n69998 , n67987 );
not ( n69999 , n69998 );
or ( n70000 , n69997 , n69999 );
buf ( n70001 , n67987 );
buf ( n70002 , n68120 );
or ( n70003 , n70001 , n70002 );
nand ( n70004 , n70000 , n70003 );
buf ( n70005 , n70004 );
xor ( n70006 , n68727 , n70005 );
nor ( n70007 , C0 , n70006 );
buf ( n70008 , n48868 );
not ( n70009 , n70008 );
buf ( n70010 , n69404 );
not ( n70011 , n70010 );
or ( n70012 , n70009 , n70011 );
and ( n70013 , n48808 , n42437 );
not ( n70014 , n48808 );
and ( n70015 , n70014 , n42428 );
or ( n70016 , n70013 , n70015 );
buf ( n70017 , n70016 );
buf ( n70018 , n48855 );
nand ( n70019 , n70017 , n70018 );
buf ( n70020 , n70019 );
buf ( n70021 , n70020 );
nand ( n70022 , n70012 , n70021 );
buf ( n70023 , n70022 );
buf ( n70024 , n70023 );
not ( n70025 , n70024 );
buf ( n70026 , n70025 );
buf ( n70027 , n70026 );
not ( n70028 , n70027 );
buf ( n70029 , n37514 );
not ( n70030 , n70029 );
buf ( n70031 , n56325 );
buf ( n70032 , n41828 );
and ( n70033 , n70031 , n70032 );
not ( n70034 , n70031 );
buf ( n70035 , n37475 );
and ( n70036 , n70034 , n70035 );
nor ( n70037 , n70033 , n70036 );
buf ( n70038 , n70037 );
buf ( n70039 , n70038 );
not ( n70040 , n70039 );
and ( n70041 , n70030 , n70040 );
not ( n70042 , n69385 );
nor ( n70043 , n70042 , n37449 );
buf ( n70044 , n70043 );
nor ( n70045 , n70041 , n70044 );
buf ( n70046 , n70045 );
buf ( n70047 , n70046 );
not ( n70048 , n70047 );
or ( n70049 , n70028 , n70048 );
buf ( n70050 , n37440 );
buf ( n70051 , n12481 );
nand ( n70052 , n70050 , n70051 );
buf ( n70053 , n70052 );
not ( n70054 , n70053 );
buf ( n70055 , n50995 );
not ( n70056 , n70055 );
buf ( n70057 , n42471 );
not ( n70058 , n70057 );
or ( n70059 , n70056 , n70058 );
buf ( n70060 , n42468 );
buf ( n70061 , n50998 );
nand ( n70062 , n70060 , n70061 );
buf ( n70063 , n70062 );
buf ( n70064 , n70063 );
nand ( n70065 , n70059 , n70064 );
buf ( n70066 , n70065 );
buf ( n70067 , n70066 );
not ( n70068 , n70067 );
buf ( n70069 , n47014 );
not ( n70070 , n70069 );
or ( n70071 , n70068 , n70070 );
buf ( n70072 , n68672 );
buf ( n70073 , n52595 );
nand ( n70074 , n70072 , n70073 );
buf ( n70075 , n70074 );
buf ( n70076 , n70075 );
nand ( n70077 , n70071 , n70076 );
buf ( n70078 , n70077 );
nor ( n70079 , n70054 , n70078 );
not ( n70080 , n68649 );
not ( n70081 , n68146 );
not ( n70082 , n68139 );
or ( n70083 , n70081 , n70082 );
nand ( n70084 , n68145 , n68142 );
nand ( n70085 , n70083 , n70084 );
not ( n70086 , n70085 );
or ( n70087 , n70080 , n70086 );
not ( n70088 , n68146 );
not ( n70089 , n68139 );
or ( n70090 , n70088 , n70089 );
nand ( n70091 , n70090 , n70084 );
or ( n70092 , n68649 , n70091 );
nand ( n70093 , n70087 , n70092 );
or ( n70094 , n70079 , n70093 );
not ( n70095 , n70053 );
nand ( n70096 , n70095 , n70078 );
nand ( n70097 , n70094 , n70096 );
buf ( n70098 , n70097 );
nand ( n70099 , n70049 , n70098 );
buf ( n70100 , n70099 );
buf ( n70101 , n70100 );
buf ( n70102 , n70046 );
not ( n70103 , n70102 );
buf ( n70104 , n70103 );
buf ( n70105 , n70104 );
buf ( n70106 , n70023 );
nand ( n70107 , n70105 , n70106 );
buf ( n70108 , n70107 );
buf ( n70109 , n70108 );
nand ( n70110 , n70101 , n70109 );
buf ( n70111 , n70110 );
not ( n70112 , n70111 );
or ( n70113 , n70007 , n70112 );
nand ( n70114 , n70113 , C1 );
buf ( n70115 , n70114 );
and ( n70116 , n69995 , n70115 );
or ( n70117 , n70116 , C0 );
buf ( n70118 , n70117 );
buf ( n70119 , n70118 );
xor ( n70120 , n67951 , n67953 );
not ( n70121 , n68742 );
xor ( n70122 , n70120 , n70121 );
buf ( n70123 , n70122 );
xor ( n70124 , n70119 , n70123 );
xor ( n70125 , n69370 , n69372 );
xor ( n70126 , n70125 , n69533 );
buf ( n70127 , n70126 );
buf ( n70128 , n70127 );
buf ( n70129 , C0 );
buf ( n70130 , n70129 );
xor ( n70131 , n69398 , n69415 );
xor ( n70132 , n70131 , n69528 );
buf ( n70133 , n70132 );
buf ( n70134 , n70133 );
xor ( n70135 , n70130 , n70134 );
xor ( n70136 , n68660 , n68685 );
xor ( n70137 , n70136 , n68723 );
buf ( n70138 , n70137 );
buf ( n70139 , n70138 );
not ( n70140 , n70139 );
buf ( n70141 , n50060 );
not ( n70142 , n70141 );
buf ( n70143 , n50599 );
not ( n70144 , n70143 );
or ( n70145 , n70142 , n70144 );
buf ( n70146 , n50591 );
buf ( n70147 , n67438 );
nand ( n70148 , n70146 , n70147 );
buf ( n70149 , n70148 );
buf ( n70150 , n70149 );
nand ( n70151 , n70145 , n70150 );
buf ( n70152 , n70151 );
buf ( n70153 , n70152 );
not ( n70154 , n70153 );
buf ( n70155 , n50608 );
not ( n70156 , n70155 );
or ( n70157 , n70154 , n70156 );
buf ( n70158 , n69671 );
buf ( n70159 , n39983 );
nand ( n70160 , n70158 , n70159 );
buf ( n70161 , n70160 );
buf ( n70162 , n70161 );
nand ( n70163 , n70157 , n70162 );
buf ( n70164 , n70163 );
buf ( n70165 , n70164 );
not ( n70166 , n70165 );
buf ( n70167 , n70166 );
buf ( n70168 , n70167 );
not ( n70169 , n70168 );
buf ( n70170 , n42408 );
not ( n70171 , n70170 );
buf ( n70172 , n37369 );
nand ( n70173 , n70171 , n70172 );
buf ( n70174 , n70173 );
and ( n70175 , n70174 , n12481 );
and ( n70176 , n46623 , n37389 );
nor ( n70177 , n70175 , n70176 );
nand ( n70178 , n42114 , n70177 );
buf ( n70179 , n70178 );
not ( n70180 , n70179 );
or ( n70181 , n70169 , n70180 );
buf ( n70182 , n44496 );
not ( n70183 , n70182 );
buf ( n70184 , n69484 );
not ( n70185 , n70184 );
or ( n70186 , n70183 , n70185 );
buf ( n70187 , n65010 );
not ( n70188 , n70187 );
buf ( n70189 , n43362 );
not ( n70190 , n70189 );
or ( n70191 , n70188 , n70190 );
buf ( n70192 , n50624 );
buf ( n70193 , n44530 );
nand ( n70194 , n70192 , n70193 );
buf ( n70195 , n70194 );
buf ( n70196 , n70195 );
nand ( n70197 , n70191 , n70196 );
buf ( n70198 , n70197 );
buf ( n70199 , n70198 );
buf ( n70200 , n44517 );
nand ( n70201 , n70199 , n70200 );
buf ( n70202 , n70201 );
buf ( n70203 , n70202 );
nand ( n70204 , n70186 , n70203 );
buf ( n70205 , n70204 );
buf ( n70206 , n70205 );
nand ( n70207 , n70181 , n70206 );
buf ( n70208 , n70207 );
buf ( n70209 , n70208 );
buf ( n70210 , n70178 );
not ( n70211 , n70210 );
buf ( n70212 , n70164 );
nand ( n70213 , n70211 , n70212 );
buf ( n70214 , n70213 );
buf ( n70215 , n70214 );
nand ( n70216 , n70209 , n70215 );
buf ( n70217 , n70216 );
buf ( n70218 , n70217 );
buf ( n70219 , n69506 );
buf ( n70220 , n69509 );
xor ( n70221 , n70219 , n70220 );
buf ( n70222 , n69486 );
xor ( n70223 , n70221 , n70222 );
buf ( n70224 , n70223 );
buf ( n70225 , n70224 );
xor ( n70226 , n70218 , n70225 );
not ( n70227 , n48855 );
and ( n70228 , n48808 , n43777 );
not ( n70229 , n48808 );
and ( n70230 , n70229 , n39653 );
or ( n70231 , n70228 , n70230 );
not ( n70232 , n70231 );
or ( n70233 , n70227 , n70232 );
buf ( n70234 , n70016 );
buf ( n70235 , n48868 );
nand ( n70236 , n70234 , n70235 );
buf ( n70237 , n70236 );
nand ( n70238 , n70233 , n70237 );
buf ( n70239 , n70238 );
and ( n70240 , n70226 , n70239 );
and ( n70241 , n70218 , n70225 );
or ( n70242 , n70240 , n70241 );
buf ( n70243 , n70242 );
buf ( n70244 , n70243 );
not ( n70245 , n70244 );
or ( n70246 , n70140 , n70245 );
buf ( n70247 , n70243 );
buf ( n70248 , n70138 );
or ( n70249 , n70247 , n70248 );
xor ( n70250 , n68566 , n68556 );
xnor ( n70251 , n70250 , n68409 );
not ( n70252 , n70251 );
buf ( n70253 , n43056 );
not ( n70254 , n70253 );
buf ( n70255 , n68606 );
not ( n70256 , n70255 );
or ( n70257 , n70254 , n70256 );
buf ( n70258 , n25226 );
buf ( n70259 , n44125 );
nand ( n70260 , n70258 , n70259 );
buf ( n70261 , n70260 );
buf ( n70262 , n70261 );
nand ( n70263 , n70257 , n70262 );
buf ( n70264 , n70263 );
not ( n70265 , n70264 );
buf ( n70266 , n42710 );
not ( n70267 , n70266 );
buf ( n70268 , n70267 );
not ( n70269 , n70268 );
or ( n70270 , n70265 , n70269 );
buf ( n70271 , n69779 );
buf ( n70272 , n42665 );
nand ( n70273 , n70271 , n70272 );
buf ( n70274 , n70273 );
nand ( n70275 , n70270 , n70274 );
not ( n70276 , n70275 );
or ( n70277 , n70252 , n70276 );
not ( n70278 , n70251 );
not ( n70279 , n70278 );
not ( n70280 , n70275 );
not ( n70281 , n70280 );
or ( n70282 , n70279 , n70281 );
xor ( n70283 , n68525 , n68529 );
xor ( n70284 , n70283 , n68552 );
buf ( n70285 , n70284 );
xor ( n70286 , n66873 , n66889 );
xor ( n70287 , n70286 , n66892 );
xor ( n70288 , n68538 , n68544 );
xor ( n70289 , n70287 , n70288 );
buf ( n70290 , n62971 );
buf ( n70291 , n58721 );
and ( n70292 , n70290 , n70291 );
buf ( n70293 , n62974 );
buf ( n70294 , n58718 );
and ( n70295 , n70293 , n70294 );
nor ( n70296 , n70292 , n70295 );
buf ( n70297 , n70296 );
buf ( n70298 , n70297 );
buf ( n70299 , n56799 );
or ( n70300 , n70298 , n70299 );
buf ( n70301 , n68337 );
buf ( n70302 , n58982 );
or ( n70303 , n70301 , n70302 );
nand ( n70304 , n70300 , n70303 );
buf ( n70305 , n70304 );
buf ( n70306 , n70305 );
buf ( n70307 , n68220 );
buf ( n70308 , n55198 );
or ( n70309 , n70307 , n70308 );
buf ( n70310 , n68217 );
buf ( n70311 , n55195 );
or ( n70312 , n70310 , n70311 );
nand ( n70313 , n70309 , n70312 );
buf ( n70314 , n70313 );
buf ( n70315 , n70314 );
not ( n70316 , n70315 );
buf ( n70317 , n70316 );
buf ( n70318 , n70317 );
buf ( n70319 , n56664 );
or ( n70320 , n70318 , n70319 );
buf ( n70321 , n68257 );
buf ( n70322 , n56673 );
or ( n70323 , n70321 , n70322 );
nand ( n70324 , n70320 , n70323 );
buf ( n70325 , n70324 );
buf ( n70326 , n70325 );
nand ( n70327 , n54904 , n55040 );
not ( n70328 , n54926 );
not ( n70329 , n55035 );
or ( n70330 , n70328 , n70329 );
not ( n70331 , n55038 );
nand ( n70332 , n70330 , n70331 );
xnor ( n70333 , n70327 , n70332 );
buf ( n70334 , n70333 );
not ( n70335 , n70334 );
buf ( n70336 , n70335 );
buf ( n70337 , n70336 );
buf ( n70338 , n55129 );
or ( n70339 , n70337 , n70338 );
buf ( n70340 , n68235 );
buf ( n70341 , n56598 );
or ( n70342 , n70340 , n70341 );
nand ( n70343 , n70339 , n70342 );
buf ( n70344 , n70343 );
buf ( n70345 , n70344 );
xor ( n70346 , n70326 , n70345 );
and ( n70347 , n70331 , n54926 );
xor ( n70348 , n70347 , n55035 );
buf ( n70349 , n70348 );
not ( n70350 , n70349 );
buf ( n70351 , n70350 );
buf ( n70352 , n70351 );
buf ( n70353 , n56589 );
or ( n70354 , n70352 , n70353 );
buf ( n70355 , n70336 );
buf ( n70356 , n56598 );
or ( n70357 , n70355 , n70356 );
nand ( n70358 , n70354 , n70357 );
buf ( n70359 , n70358 );
buf ( n70360 , n70359 );
buf ( n70361 , n56670 );
not ( n70362 , n70361 );
buf ( n70363 , n70314 );
not ( n70364 , n70363 );
or ( n70365 , n70362 , n70364 );
buf ( n70366 , n55195 );
buf ( n70367 , n68232 );
and ( n70368 , n70366 , n70367 );
not ( n70369 , n70366 );
buf ( n70370 , n68235 );
and ( n70371 , n70369 , n70370 );
nor ( n70372 , n70368 , n70371 );
buf ( n70373 , n70372 );
buf ( n70374 , n70373 );
buf ( n70375 , n56664 );
or ( n70376 , n70374 , n70375 );
nand ( n70377 , n70365 , n70376 );
buf ( n70378 , n70377 );
buf ( n70379 , n70378 );
and ( n70380 , n70360 , n70379 );
buf ( n70381 , n70380 );
buf ( n70382 , n70381 );
and ( n70383 , n70346 , n70382 );
and ( n70384 , n70326 , n70345 );
or ( n70385 , n70383 , n70384 );
buf ( n70386 , n70385 );
buf ( n70387 , n70386 );
xor ( n70388 , n70306 , n70387 );
buf ( n70389 , n60068 );
buf ( n70390 , n60261 );
and ( n70391 , n70389 , n70390 );
buf ( n70392 , n60071 );
buf ( n70393 , n60090 );
and ( n70394 , n70392 , n70393 );
nor ( n70395 , n70391 , n70394 );
buf ( n70396 , n70395 );
or ( n70397 , n70396 , n60270 );
or ( n70398 , n68413 , n60100 );
nand ( n70399 , n70397 , n70398 );
buf ( n70400 , n70399 );
and ( n70401 , n70388 , n70400 );
and ( n70402 , n70306 , n70387 );
or ( n70403 , n70401 , n70402 );
buf ( n70404 , n70403 );
buf ( n70405 , n70404 );
xor ( n70406 , n68346 , n68363 );
xor ( n70407 , n70406 , n68389 );
buf ( n70408 , n70407 );
buf ( n70409 , n70408 );
xor ( n70410 , n70405 , n70409 );
xor ( n70411 , n68419 , n68422 );
xor ( n70412 , n70411 , n68439 );
buf ( n70413 , n70412 );
and ( n70414 , n70410 , n70413 );
and ( n70415 , n70405 , n70409 );
or ( n70416 , n70414 , n70415 );
buf ( n70417 , n70416 );
xor ( n70418 , n70289 , n70417 );
xor ( n70419 , n68443 , n68515 );
xor ( n70420 , n70419 , n68520 );
buf ( n70421 , n70420 );
and ( n70422 , n70418 , n70421 );
and ( n70423 , n70289 , n70417 );
or ( n70424 , n70422 , n70423 );
or ( n70425 , n70285 , n70424 );
not ( n70426 , n70425 );
xor ( n70427 , n68468 , n68485 );
xor ( n70428 , n70427 , n68505 );
buf ( n70429 , n70428 );
not ( n70430 , n62691 );
not ( n70431 , n68448 );
or ( n70432 , n70430 , n70431 );
buf ( n70433 , n58857 );
buf ( n70434 , n62681 );
and ( n70435 , n70433 , n70434 );
buf ( n70436 , n58858 );
buf ( n70437 , n62663 );
and ( n70438 , n70436 , n70437 );
nor ( n70439 , n70435 , n70438 );
buf ( n70440 , n70439 );
not ( n70441 , n70440 );
nand ( n70442 , n70441 , n62679 );
nand ( n70443 , n70432 , n70442 );
xor ( n70444 , n70429 , n70443 );
buf ( n70445 , n60229 );
buf ( n70446 , n60261 );
and ( n70447 , n70445 , n70446 );
buf ( n70448 , n62652 );
buf ( n70449 , n60090 );
and ( n70450 , n70448 , n70449 );
nor ( n70451 , n70447 , n70450 );
buf ( n70452 , n70451 );
buf ( n70453 , n70452 );
buf ( n70454 , n60270 );
or ( n70455 , n70453 , n70454 );
buf ( n70456 , n70396 );
buf ( n70457 , n60100 );
or ( n70458 , n70456 , n70457 );
nand ( n70459 , n70455 , n70458 );
buf ( n70460 , n70459 );
buf ( n70461 , n70460 );
buf ( n70462 , n62782 );
buf ( n70463 , n58897 );
and ( n70464 , n70462 , n70463 );
buf ( n70465 , n62980 );
buf ( n70466 , n68170 );
and ( n70467 , n70465 , n70466 );
nor ( n70468 , n70464 , n70467 );
buf ( n70469 , n70468 );
buf ( n70470 , n70469 );
buf ( n70471 , n58913 );
or ( n70472 , n70470 , n70471 );
buf ( n70473 , n68499 );
buf ( n70474 , n58890 );
or ( n70475 , n70473 , n70474 );
nand ( n70476 , n70472 , n70475 );
buf ( n70477 , n70476 );
buf ( n70478 , n70477 );
xor ( n70479 , n70461 , n70478 );
xor ( n70480 , n70360 , n70379 );
buf ( n70481 , n70480 );
buf ( n70482 , n70481 );
buf ( n70483 , n66690 );
buf ( n70484 , n56641 );
and ( n70485 , n70483 , n70484 );
buf ( n70486 , n66693 );
buf ( n70487 , n56631 );
and ( n70488 , n70486 , n70487 );
nor ( n70489 , n70485 , n70488 );
buf ( n70490 , n70489 );
buf ( n70491 , n70490 );
buf ( n70492 , n56626 );
or ( n70493 , n70491 , n70492 );
buf ( n70494 , n66601 );
buf ( n70495 , n56641 );
and ( n70496 , n70494 , n70495 );
buf ( n70497 , n66604 );
buf ( n70498 , n56631 );
and ( n70499 , n70497 , n70498 );
nor ( n70500 , n70496 , n70499 );
buf ( n70501 , n70500 );
buf ( n70502 , n70501 );
buf ( n70503 , n56639 );
or ( n70504 , n70502 , n70503 );
nand ( n70505 , n70493 , n70504 );
buf ( n70506 , n70505 );
buf ( n70507 , n70506 );
xor ( n70508 , n70482 , n70507 );
buf ( n70509 , n70333 );
buf ( n70510 , n55195 );
and ( n70511 , n70509 , n70510 );
buf ( n70512 , n70336 );
buf ( n70513 , n55198 );
and ( n70514 , n70512 , n70513 );
nor ( n70515 , n70511 , n70514 );
buf ( n70516 , n70515 );
buf ( n70517 , n70516 );
buf ( n70518 , n56664 );
or ( n70519 , n70517 , n70518 );
buf ( n70520 , n70373 );
buf ( n70521 , n56673 );
or ( n70522 , n70520 , n70521 );
nand ( n70523 , n70519 , n70522 );
buf ( n70524 , n70523 );
buf ( n70525 , n70524 );
and ( n70526 , n55034 , n54952 );
xor ( n70527 , n70526 , n55030 );
buf ( n70528 , n70527 );
not ( n70529 , n70528 );
buf ( n70530 , n70529 );
buf ( n70531 , n70530 );
buf ( n70532 , n56589 );
or ( n70533 , n70531 , n70532 );
buf ( n70534 , n70351 );
buf ( n70535 , n56598 );
or ( n70536 , n70534 , n70535 );
nand ( n70537 , n70533 , n70536 );
buf ( n70538 , n70537 );
buf ( n70539 , n70538 );
xor ( n70540 , n70525 , n70539 );
buf ( n70541 , n56629 );
not ( n70542 , n70541 );
buf ( n70543 , n68217 );
buf ( n70544 , n56641 );
and ( n70545 , n70543 , n70544 );
buf ( n70546 , n68220 );
buf ( n70547 , n56631 );
and ( n70548 , n70546 , n70547 );
nor ( n70549 , n70545 , n70548 );
buf ( n70550 , n70549 );
buf ( n70551 , n70550 );
not ( n70552 , n70551 );
buf ( n70553 , n70552 );
buf ( n70554 , n70553 );
not ( n70555 , n70554 );
or ( n70556 , n70542 , n70555 );
buf ( n70557 , n70490 );
buf ( n70558 , n56639 );
or ( n70559 , n70557 , n70558 );
nand ( n70560 , n70556 , n70559 );
buf ( n70561 , n70560 );
buf ( n70562 , n70561 );
and ( n70563 , n70540 , n70562 );
and ( n70564 , n70525 , n70539 );
or ( n70565 , n70563 , n70564 );
buf ( n70566 , n70565 );
buf ( n70567 , n70566 );
and ( n70568 , n70508 , n70567 );
and ( n70569 , n70482 , n70507 );
or ( n70570 , n70568 , n70569 );
buf ( n70571 , n70570 );
buf ( n70572 , n70571 );
and ( n70573 , n70479 , n70572 );
and ( n70574 , n70461 , n70478 );
or ( n70575 , n70573 , n70574 );
buf ( n70576 , n70575 );
and ( n70577 , n70444 , n70576 );
and ( n70578 , n70429 , n70443 );
or ( n70579 , n70577 , n70578 );
buf ( n70580 , n70579 );
buf ( n70581 , n56582 );
buf ( n70582 , n66742 );
and ( n70583 , n70581 , n70582 );
buf ( n70584 , n56585 );
buf ( n70585 , n63000 );
and ( n70586 , n70584 , n70585 );
nor ( n70587 , n70583 , n70586 );
buf ( n70588 , n70587 );
buf ( n70589 , n70588 );
buf ( n70590 , n64230 );
or ( n70591 , n70589 , n70590 );
buf ( n70592 , n68459 );
buf ( n70593 , n64227 );
or ( n70594 , n70592 , n70593 );
nand ( n70595 , n70591 , n70594 );
buf ( n70596 , n70595 );
buf ( n70597 , n70596 );
buf ( n70598 , n64068 );
buf ( n70599 , n58721 );
and ( n70600 , n70598 , n70599 );
buf ( n70601 , n66579 );
buf ( n70602 , n58718 );
and ( n70603 , n70601 , n70602 );
nor ( n70604 , n70600 , n70603 );
buf ( n70605 , n70604 );
buf ( n70606 , n70605 );
buf ( n70607 , n56799 );
or ( n70608 , n70606 , n70607 );
buf ( n70609 , n70297 );
buf ( n70610 , n58982 );
or ( n70611 , n70609 , n70610 );
nand ( n70612 , n70608 , n70611 );
buf ( n70613 , n70612 );
buf ( n70614 , n70613 );
buf ( n70615 , n70501 );
buf ( n70616 , n56626 );
or ( n70617 , n70615 , n70616 );
buf ( n70618 , n68476 );
buf ( n70619 , n56639 );
or ( n70620 , n70618 , n70619 );
nand ( n70621 , n70617 , n70620 );
buf ( n70622 , n70621 );
buf ( n70623 , n70622 );
xor ( n70624 , n70614 , n70623 );
xor ( n70625 , n70326 , n70345 );
xor ( n70626 , n70625 , n70382 );
buf ( n70627 , n70626 );
buf ( n70628 , n70627 );
and ( n70629 , n70624 , n70628 );
and ( n70630 , n70614 , n70623 );
or ( n70631 , n70629 , n70630 );
buf ( n70632 , n70631 );
buf ( n70633 , n70632 );
xor ( n70634 , n70597 , n70633 );
buf ( n70635 , n63013 );
not ( n70636 , n70635 );
buf ( n70637 , n58747 );
buf ( n70638 , n64129 );
and ( n70639 , n70637 , n70638 );
buf ( n70640 , n58841 );
buf ( n70641 , n64133 );
and ( n70642 , n70640 , n70641 );
nor ( n70643 , n70639 , n70642 );
buf ( n70644 , n70643 );
buf ( n70645 , n70644 );
not ( n70646 , n70645 );
buf ( n70647 , n70646 );
buf ( n70648 , n70647 );
not ( n70649 , n70648 );
or ( n70650 , n70636 , n70649 );
buf ( n70651 , n68432 );
buf ( n70652 , n63010 );
or ( n70653 , n70651 , n70652 );
nand ( n70654 , n70650 , n70653 );
buf ( n70655 , n70654 );
buf ( n70656 , n70655 );
and ( n70657 , n70634 , n70656 );
and ( n70658 , n70597 , n70633 );
or ( n70659 , n70657 , n70658 );
buf ( n70660 , n70659 );
buf ( n70661 , n70660 );
xor ( n70662 , n70580 , n70661 );
xor ( n70663 , n68451 , n68464 );
xor ( n70664 , n70663 , n68510 );
buf ( n70665 , n70664 );
buf ( n70666 , n70665 );
and ( n70667 , n70662 , n70666 );
and ( n70668 , n70580 , n70661 );
or ( n70669 , n70667 , n70668 );
buf ( n70670 , n70669 );
xor ( n70671 , n70289 , n70417 );
xor ( n70672 , n70671 , n70421 );
and ( n70673 , n70670 , n70672 );
or ( n70674 , n70588 , n64227 );
not ( n70675 , n64230 );
and ( n70676 , n58792 , n62999 );
and ( n70677 , n56720 , n63000 );
nor ( n70678 , n70676 , n70677 );
nand ( n70679 , n70675 , n70678 );
nand ( n70680 , n70674 , n70679 );
buf ( n70681 , n70680 );
buf ( n70682 , n59009 );
buf ( n70683 , n62681 );
and ( n70684 , n70682 , n70683 );
buf ( n70685 , n60077 );
buf ( n70686 , n62663 );
and ( n70687 , n70685 , n70686 );
nor ( n70688 , n70684 , n70687 );
buf ( n70689 , n70688 );
buf ( n70690 , n70689 );
buf ( n70691 , n62935 );
or ( n70692 , n70690 , n70691 );
buf ( n70693 , n70440 );
buf ( n70694 , n62676 );
or ( n70695 , n70693 , n70694 );
nand ( n70696 , n70692 , n70695 );
buf ( n70697 , n70696 );
buf ( n70698 , n70697 );
xor ( n70699 , n70681 , n70698 );
xor ( n70700 , n70614 , n70623 );
xor ( n70701 , n70700 , n70628 );
buf ( n70702 , n70701 );
buf ( n70703 , n70702 );
and ( n70704 , n70699 , n70703 );
and ( n70705 , n70681 , n70698 );
or ( n70706 , n70704 , n70705 );
buf ( n70707 , n70706 );
buf ( n70708 , n70707 );
xor ( n70709 , n70306 , n70387 );
xor ( n70710 , n70709 , n70400 );
buf ( n70711 , n70710 );
buf ( n70712 , n70711 );
xor ( n70713 , n70708 , n70712 );
xor ( n70714 , n70597 , n70633 );
xor ( n70715 , n70714 , n70656 );
buf ( n70716 , n70715 );
buf ( n70717 , n70716 );
and ( n70718 , n70713 , n70717 );
and ( n70719 , n70708 , n70712 );
or ( n70720 , n70718 , n70719 );
buf ( n70721 , n70720 );
xor ( n70722 , n70405 , n70409 );
xor ( n70723 , n70722 , n70413 );
buf ( n70724 , n70723 );
xor ( n70725 , n70721 , n70724 );
xor ( n70726 , n70580 , n70661 );
xor ( n70727 , n70726 , n70666 );
buf ( n70728 , n70727 );
and ( n70729 , n70725 , n70728 );
and ( n70730 , n70721 , n70724 );
or ( n70731 , n70729 , n70730 );
xor ( n70732 , n70289 , n70417 );
xor ( n70733 , n70732 , n70421 );
and ( n70734 , n70731 , n70733 );
and ( n70735 , n70670 , n70731 );
or ( n70736 , n70673 , n70734 , n70735 );
not ( n70737 , n70736 );
or ( n70738 , n70426 , n70737 );
nand ( n70739 , n70285 , n70424 );
nand ( n70740 , n70738 , n70739 );
nand ( n70741 , n70282 , n70740 );
nand ( n70742 , n70277 , n70741 );
buf ( n70743 , n70742 );
buf ( n70744 , n42309 );
not ( n70745 , n70744 );
buf ( n70746 , n69754 );
not ( n70747 , n70746 );
or ( n70748 , n70745 , n70747 );
and ( n70749 , n13662 , n42260 );
not ( n70750 , n13662 );
and ( n70751 , n70750 , n59242 );
or ( n70752 , n70749 , n70751 );
buf ( n70753 , n70752 );
buf ( n70754 , n42246 );
nand ( n70755 , n70753 , n70754 );
buf ( n70756 , n70755 );
buf ( n70757 , n70756 );
nand ( n70758 , n70748 , n70757 );
buf ( n70759 , n70758 );
buf ( n70760 , n70759 );
xor ( n70761 , n70743 , n70760 );
not ( n70762 , n44952 );
not ( n70763 , n41657 );
or ( n70764 , n70762 , n70763 );
buf ( n70765 , n61442 );
buf ( n70766 , n44949 );
nand ( n70767 , n70765 , n70766 );
buf ( n70768 , n70767 );
nand ( n70769 , n70764 , n70768 );
not ( n70770 , n70769 );
not ( n70771 , n61454 );
or ( n70772 , n70770 , n70771 );
buf ( n70773 , n68630 );
not ( n70774 , n70773 );
buf ( n70775 , n48671 );
nand ( n70776 , n70774 , n70775 );
buf ( n70777 , n70776 );
nand ( n70778 , n70772 , n70777 );
buf ( n70779 , n70778 );
and ( n70780 , n70761 , n70779 );
and ( n70781 , n70743 , n70760 );
or ( n70782 , n70780 , n70781 );
buf ( n70783 , n70782 );
buf ( n70784 , n70783 );
buf ( n70785 , n43868 );
not ( n70786 , n70785 );
buf ( n70787 , n69501 );
not ( n70788 , n70787 );
or ( n70789 , n70786 , n70788 );
and ( n70790 , n29754 , n41604 );
not ( n70791 , n29754 );
and ( n70792 , n70791 , n41605 );
or ( n70793 , n70790 , n70792 );
buf ( n70794 , n70793 );
buf ( n70795 , n41596 );
nand ( n70796 , n70794 , n70795 );
buf ( n70797 , n70796 );
buf ( n70798 , n70797 );
nand ( n70799 , n70789 , n70798 );
buf ( n70800 , n70799 );
buf ( n70801 , n70800 );
xor ( n70802 , n70784 , n70801 );
xor ( n70803 , n69775 , n69792 );
xor ( n70804 , n70803 , n69824 );
buf ( n70805 , n70804 );
buf ( n70806 , n70805 );
buf ( n70807 , n43868 );
not ( n70808 , n70807 );
buf ( n70809 , n70793 );
not ( n70810 , n70809 );
or ( n70811 , n70808 , n70810 );
buf ( n70812 , n41605 );
not ( n70813 , n70812 );
buf ( n70814 , n63906 );
not ( n70815 , n70814 );
or ( n70816 , n70813 , n70815 );
buf ( n70817 , n13653 );
buf ( n70818 , n41604 );
nand ( n70819 , n70817 , n70818 );
buf ( n70820 , n70819 );
buf ( n70821 , n70820 );
nand ( n70822 , n70816 , n70821 );
buf ( n70823 , n70822 );
buf ( n70824 , n70823 );
buf ( n70825 , n41596 );
nand ( n70826 , n70824 , n70825 );
buf ( n70827 , n70826 );
buf ( n70828 , n70827 );
nand ( n70829 , n70811 , n70828 );
buf ( n70830 , n70829 );
buf ( n70831 , n70830 );
xor ( n70832 , n70806 , n70831 );
not ( n70833 , n70278 );
not ( n70834 , n70740 );
or ( n70835 , n70833 , n70834 );
or ( n70836 , n70740 , n70278 );
nand ( n70837 , n70835 , n70836 );
and ( n70838 , n70275 , n70837 );
not ( n70839 , n70275 );
buf ( n70840 , n70837 );
not ( n70841 , n70840 );
buf ( n70842 , n70841 );
and ( n70843 , n70839 , n70842 );
nor ( n70844 , n70838 , n70843 );
buf ( n70845 , n70844 );
buf ( n70846 , n42309 );
not ( n70847 , n70846 );
buf ( n70848 , n70752 );
not ( n70849 , n70848 );
or ( n70850 , n70847 , n70849 );
buf ( n70851 , n59242 );
not ( n70852 , n70851 );
buf ( n70853 , n29463 );
not ( n70854 , n70853 );
buf ( n70855 , n70854 );
buf ( n70856 , n70855 );
not ( n70857 , n70856 );
or ( n70858 , n70852 , n70857 );
buf ( n70859 , n29463 );
buf ( n70860 , n42260 );
nand ( n70861 , n70859 , n70860 );
buf ( n70862 , n70861 );
buf ( n70863 , n70862 );
nand ( n70864 , n70858 , n70863 );
buf ( n70865 , n70864 );
buf ( n70866 , n70865 );
buf ( n70867 , n42246 );
nand ( n70868 , n70866 , n70867 );
buf ( n70869 , n70868 );
buf ( n70870 , n70869 );
nand ( n70871 , n70850 , n70870 );
buf ( n70872 , n70871 );
buf ( n70873 , n70872 );
xor ( n70874 , n70845 , n70873 );
buf ( n70875 , n42847 );
not ( n70876 , n70875 );
buf ( n70877 , n69798 );
not ( n70878 , n70877 );
or ( n70879 , n70876 , n70878 );
buf ( n70880 , n46691 );
buf ( n70881 , n69804 );
nand ( n70882 , n70880 , n70881 );
buf ( n70883 , n70882 );
buf ( n70884 , n70883 );
nand ( n70885 , n70879 , n70884 );
buf ( n70886 , n70885 );
buf ( n70887 , n70886 );
not ( n70888 , n70887 );
buf ( n70889 , n66459 );
not ( n70890 , n70889 );
or ( n70891 , n70888 , n70890 );
buf ( n70892 , n69811 );
buf ( n70893 , n66482 );
nand ( n70894 , n70892 , n70893 );
buf ( n70895 , n70894 );
buf ( n70896 , n70895 );
nand ( n70897 , n70891 , n70896 );
buf ( n70898 , n70897 );
buf ( n70899 , n70898 );
and ( n70900 , n70874 , n70899 );
and ( n70901 , n70845 , n70873 );
or ( n70902 , n70900 , n70901 );
buf ( n70903 , n70902 );
buf ( n70904 , n70903 );
and ( n70905 , n70832 , n70904 );
and ( n70906 , n70806 , n70831 );
or ( n70907 , n70905 , n70906 );
buf ( n70908 , n70907 );
buf ( n70909 , n70908 );
and ( n70910 , n70802 , n70909 );
and ( n70911 , n70784 , n70801 );
or ( n70912 , n70910 , n70911 );
buf ( n70913 , n70912 );
buf ( n70914 , n70913 );
buf ( n70915 , n46225 );
not ( n70916 , n70915 );
buf ( n70917 , n64616 );
not ( n70918 , n70917 );
buf ( n70919 , n41915 );
not ( n70920 , n70919 );
or ( n70921 , n70918 , n70920 );
buf ( n70922 , n41912 );
buf ( n70923 , n45747 );
nand ( n70924 , n70922 , n70923 );
buf ( n70925 , n70924 );
buf ( n70926 , n70925 );
nand ( n70927 , n70921 , n70926 );
buf ( n70928 , n70927 );
buf ( n70929 , n70928 );
not ( n70930 , n70929 );
or ( n70931 , n70916 , n70930 );
buf ( n70932 , n69461 );
buf ( n70933 , n67149 );
nand ( n70934 , n70932 , n70933 );
buf ( n70935 , n70934 );
buf ( n70936 , n70935 );
nand ( n70937 , n70931 , n70936 );
buf ( n70938 , n70937 );
buf ( n70939 , n70938 );
xor ( n70940 , n70914 , n70939 );
not ( n70941 , n38404 );
buf ( n70942 , n42411 );
not ( n70943 , n70942 );
buf ( n70944 , n52789 );
not ( n70945 , n70944 );
and ( n70946 , n70943 , n70945 );
buf ( n70947 , n48984 );
buf ( n70948 , n52789 );
and ( n70949 , n70947 , n70948 );
nor ( n70950 , n70946 , n70949 );
buf ( n70951 , n70950 );
buf ( n70952 , n70951 );
not ( n70953 , n70952 );
buf ( n70954 , n70953 );
not ( n70955 , n70954 );
or ( n70956 , n70941 , n70955 );
buf ( n70957 , n69854 );
buf ( n70958 , n38380 );
nand ( n70959 , n70957 , n70958 );
buf ( n70960 , n70959 );
nand ( n70961 , n70956 , n70960 );
buf ( n70962 , n70961 );
and ( n70963 , n70940 , n70962 );
and ( n70964 , n70914 , n70939 );
or ( n70965 , n70963 , n70964 );
buf ( n70966 , n70965 );
buf ( n70967 , n70966 );
nand ( n70968 , n70249 , n70967 );
buf ( n70969 , n70968 );
buf ( n70970 , n70969 );
nand ( n70971 , n70246 , n70970 );
buf ( n70972 , n70971 );
buf ( n70973 , n70972 );
and ( n70974 , n70135 , n70973 );
or ( n70975 , n70974 , C0 );
buf ( n70976 , n70975 );
buf ( n70977 , n70976 );
xor ( n70978 , n70128 , n70977 );
xor ( n70979 , n69581 , n69588 );
xor ( n70980 , n70979 , n69905 );
buf ( n70981 , n70980 );
buf ( n70982 , n70981 );
and ( n70983 , n70978 , n70982 );
and ( n70984 , n70128 , n70977 );
or ( n70985 , n70983 , n70984 );
buf ( n70986 , n70985 );
buf ( n70987 , n70986 );
and ( n70988 , n70124 , n70987 );
and ( n70989 , n70119 , n70123 );
or ( n70990 , n70988 , n70989 );
buf ( n70991 , n70990 );
buf ( n70992 , n70991 );
and ( n70993 , n69980 , n70992 );
and ( n70994 , n69975 , n69979 );
or ( n70995 , n70993 , n70994 );
buf ( n70996 , n70995 );
buf ( n70997 , n70996 );
or ( n70998 , n69968 , n70997 );
buf ( n70999 , n70998 );
buf ( n71000 , n70999 );
and ( n71001 , n69361 , n71000 );
buf ( n71002 , n69967 );
buf ( n71003 , n70996 );
and ( n71004 , n71002 , n71003 );
buf ( n71005 , n71004 );
buf ( n71006 , n71005 );
nor ( n71007 , n71001 , n71006 );
buf ( n71008 , n71007 );
buf ( n71009 , n71008 );
nand ( n71010 , n69355 , n71009 );
buf ( n71011 , n71010 );
buf ( n71012 , n71011 );
and ( n71013 , n69271 , n69351 , n71012 );
buf ( n71014 , n71013 );
not ( n71015 , n71014 );
buf ( n71016 , n67149 );
not ( n71017 , n71016 );
buf ( n71018 , n53492 );
not ( n71019 , n71018 );
buf ( n71020 , n42072 );
not ( n71021 , n71020 );
or ( n71022 , n71019 , n71021 );
buf ( n71023 , n28368 );
buf ( n71024 , n45747 );
nand ( n71025 , n71023 , n71024 );
buf ( n71026 , n71025 );
buf ( n71027 , n71026 );
nand ( n71028 , n71022 , n71027 );
buf ( n71029 , n71028 );
buf ( n71030 , n71029 );
not ( n71031 , n71030 );
or ( n71032 , n71017 , n71031 );
buf ( n71033 , n53492 );
not ( n71034 , n71033 );
buf ( n71035 , n56545 );
not ( n71036 , n71035 );
or ( n71037 , n71034 , n71036 );
buf ( n71038 , n42049 );
buf ( n71039 , n45747 );
nand ( n71040 , n71038 , n71039 );
buf ( n71041 , n71040 );
buf ( n71042 , n71041 );
nand ( n71043 , n71037 , n71042 );
buf ( n71044 , n71043 );
buf ( n71045 , n71044 );
buf ( n71046 , n45742 );
not ( n71047 , n71046 );
buf ( n71048 , n71047 );
buf ( n71049 , n71048 );
nand ( n71050 , n71045 , n71049 );
buf ( n71051 , n71050 );
buf ( n71052 , n71051 );
nand ( n71053 , n71032 , n71052 );
buf ( n71054 , n71053 );
buf ( n71055 , n71054 );
buf ( n71056 , n38979 );
buf ( n71057 , n50599 );
not ( n71058 , n71057 );
buf ( n71059 , n38969 );
not ( n71060 , n71059 );
or ( n71061 , n71058 , n71060 );
buf ( n71062 , n12481 );
nand ( n71063 , n71061 , n71062 );
buf ( n71064 , n71063 );
buf ( n71065 , n71064 );
buf ( n71066 , n38969 );
not ( n71067 , n71066 );
buf ( n71068 , n24092 );
nand ( n71069 , n71067 , n71068 );
buf ( n71070 , n71069 );
buf ( n71071 , n71070 );
and ( n71072 , n71056 , n71065 , n71071 );
buf ( n71073 , n71072 );
buf ( n71074 , n71073 );
xor ( n71075 , n71055 , n71074 );
buf ( n71076 , n48320 );
not ( n71077 , n71076 );
buf ( n71078 , n71077 );
buf ( n71079 , n71078 );
not ( n71080 , n71079 );
buf ( n71081 , n58107 );
not ( n71082 , n71081 );
or ( n71083 , n71080 , n71082 );
buf ( n71084 , n61442 );
buf ( n71085 , n48320 );
nand ( n71086 , n71084 , n71085 );
buf ( n71087 , n71086 );
buf ( n71088 , n71087 );
nand ( n71089 , n71083 , n71088 );
buf ( n71090 , n71089 );
buf ( n71091 , n71090 );
not ( n71092 , n71091 );
buf ( n71093 , n59928 );
not ( n71094 , n71093 );
or ( n71095 , n71092 , n71094 );
buf ( n71096 , n47716 );
not ( n71097 , n71096 );
buf ( n71098 , n62598 );
not ( n71099 , n71098 );
or ( n71100 , n71097 , n71099 );
buf ( n71101 , n61434 );
buf ( n71102 , n47725 );
nand ( n71103 , n71101 , n71102 );
buf ( n71104 , n71103 );
buf ( n71105 , n71104 );
nand ( n71106 , n71100 , n71105 );
buf ( n71107 , n71106 );
buf ( n71108 , n71107 );
buf ( n71109 , n62582 );
nand ( n71110 , n71108 , n71109 );
buf ( n71111 , n71110 );
buf ( n71112 , n71111 );
nand ( n71113 , n71095 , n71112 );
buf ( n71114 , n71113 );
buf ( n71115 , n71114 );
buf ( n71116 , n42856 );
not ( n71117 , n71116 );
buf ( n71118 , n42260 );
not ( n71119 , n71118 );
or ( n71120 , n71117 , n71119 );
buf ( n71121 , n25303 );
not ( n71122 , n71121 );
buf ( n71123 , n71122 );
buf ( n71124 , n71123 );
buf ( n71125 , n42859 );
nand ( n71126 , n71124 , n71125 );
buf ( n71127 , n71126 );
buf ( n71128 , n71127 );
nand ( n71129 , n71120 , n71128 );
buf ( n71130 , n71129 );
buf ( n71131 , n71130 );
buf ( n71132 , n42309 );
nand ( n71133 , n71131 , n71132 );
buf ( n71134 , n71133 );
not ( n71135 , n71134 );
buf ( n71136 , n42847 );
buf ( n71137 , n25306 );
and ( n71138 , n71136 , n71137 );
not ( n71139 , n71136 );
buf ( n71140 , n25303 );
and ( n71141 , n71139 , n71140 );
nor ( n71142 , n71138 , n71141 );
buf ( n71143 , n71142 );
not ( n71144 , n71143 );
nor ( n71145 , n71144 , n42243 );
nor ( n71146 , n71135 , n71145 );
buf ( n71147 , n58823 );
buf ( n71148 , n66742 );
and ( n71149 , n71147 , n71148 );
buf ( n71150 , n58862 );
buf ( n71151 , n63000 );
and ( n71152 , n71150 , n71151 );
nor ( n71153 , n71149 , n71152 );
buf ( n71154 , n71153 );
buf ( n71155 , n71154 );
buf ( n71156 , n64230 );
or ( n71157 , n71155 , n71156 );
buf ( n71158 , n58835 );
buf ( n71159 , n66742 );
and ( n71160 , n71158 , n71159 );
buf ( n71161 , n58841 );
buf ( n71162 , n63000 );
and ( n71163 , n71161 , n71162 );
nor ( n71164 , n71160 , n71163 );
buf ( n71165 , n71164 );
buf ( n71166 , n71165 );
buf ( n71167 , n64227 );
or ( n71168 , n71166 , n71167 );
nand ( n71169 , n71157 , n71168 );
buf ( n71170 , n71169 );
buf ( n71171 , n71170 );
buf ( n71172 , n64211 );
buf ( n71173 , n58897 );
and ( n71174 , n71172 , n71173 );
buf ( n71175 , n66610 );
buf ( n71176 , n58894 );
and ( n71177 , n71175 , n71176 );
nor ( n71178 , n71174 , n71177 );
buf ( n71179 , n71178 );
buf ( n71180 , n71179 );
buf ( n71181 , n58913 );
or ( n71182 , n71180 , n71181 );
buf ( n71183 , n64068 );
buf ( n71184 , n58897 );
and ( n71185 , n71183 , n71184 );
buf ( n71186 , n66579 );
buf ( n71187 , n68170 );
and ( n71188 , n71186 , n71187 );
nor ( n71189 , n71185 , n71188 );
buf ( n71190 , n71189 );
buf ( n71191 , n71190 );
buf ( n71192 , n58890 );
or ( n71193 , n71191 , n71192 );
nand ( n71194 , n71182 , n71193 );
buf ( n71195 , n71194 );
buf ( n71196 , n71195 );
buf ( n71197 , n70527 );
buf ( n71198 , n55195 );
and ( n71199 , n71197 , n71198 );
buf ( n71200 , n70530 );
buf ( n71201 , n55198 );
and ( n71202 , n71200 , n71201 );
nor ( n71203 , n71199 , n71202 );
buf ( n71204 , n71203 );
buf ( n71205 , n71204 );
buf ( n71206 , n56664 );
or ( n71207 , n71205 , n71206 );
buf ( n71208 , n70348 );
buf ( n71209 , n55195 );
and ( n71210 , n71208 , n71209 );
buf ( n71211 , n70351 );
buf ( n71212 , n55201 );
and ( n71213 , n71211 , n71212 );
nor ( n71214 , n71210 , n71213 );
buf ( n71215 , n71214 );
buf ( n71216 , n71215 );
buf ( n71217 , n56673 );
or ( n71218 , n71216 , n71217 );
nand ( n71219 , n71207 , n71218 );
buf ( n71220 , n71219 );
buf ( n71221 , n71220 );
buf ( n71222 , n55129 );
not ( n71223 , n54986 );
nor ( n71224 , n71223 , n55025 );
xor ( n71225 , n55022 , n71224 );
buf ( n71226 , n71225 );
not ( n71227 , n71226 );
buf ( n71228 , n71227 );
buf ( n71229 , n71228 );
or ( n71230 , n71222 , n71229 );
xor ( n71231 , n54966 , n54968 );
xor ( n71232 , n71231 , n55027 );
buf ( n71233 , n71232 );
not ( n71234 , n71233 );
buf ( n71235 , n71234 );
buf ( n71236 , n71235 );
buf ( n71237 , n56598 );
or ( n71238 , n71236 , n71237 );
nand ( n71239 , n71230 , n71238 );
buf ( n71240 , n71239 );
buf ( n71241 , n71240 );
xor ( n71242 , n71221 , n71241 );
buf ( n71243 , n56611 );
not ( n71244 , n71243 );
buf ( n71245 , n68232 );
buf ( n71246 , n56641 );
and ( n71247 , n71245 , n71246 );
buf ( n71248 , n68235 );
buf ( n71249 , n56631 );
and ( n71250 , n71248 , n71249 );
nor ( n71251 , n71247 , n71250 );
buf ( n71252 , n71251 );
buf ( n71253 , n71252 );
not ( n71254 , n71253 );
buf ( n71255 , n71254 );
buf ( n71256 , n71255 );
not ( n71257 , n71256 );
or ( n71258 , n71244 , n71257 );
buf ( n71259 , n70333 );
buf ( n71260 , n56641 );
and ( n71261 , n71259 , n71260 );
buf ( n71262 , n70336 );
buf ( n71263 , n56631 );
and ( n71264 , n71262 , n71263 );
nor ( n71265 , n71261 , n71264 );
buf ( n71266 , n71265 );
buf ( n71267 , n71266 );
buf ( n71268 , n56626 );
or ( n71269 , n71267 , n71268 );
nand ( n71270 , n71258 , n71269 );
buf ( n71271 , n71270 );
buf ( n71272 , n71271 );
and ( n71273 , n71242 , n71272 );
and ( n71274 , n71221 , n71241 );
or ( n71275 , n71273 , n71274 );
buf ( n71276 , n71275 );
buf ( n71277 , n71276 );
xor ( n71278 , n71196 , n71277 );
buf ( n71279 , n68217 );
buf ( n71280 , n58721 );
and ( n71281 , n71279 , n71280 );
buf ( n71282 , n68220 );
buf ( n71283 , n58718 );
and ( n71284 , n71282 , n71283 );
nor ( n71285 , n71281 , n71284 );
buf ( n71286 , n71285 );
buf ( n71287 , n71286 );
buf ( n71288 , n56799 );
or ( n71289 , n71287 , n71288 );
buf ( n71290 , n66690 );
buf ( n71291 , n58721 );
and ( n71292 , n71290 , n71291 );
buf ( n71293 , n66693 );
buf ( n71294 , n58718 );
and ( n71295 , n71293 , n71294 );
nor ( n71296 , n71292 , n71295 );
buf ( n71297 , n71296 );
buf ( n71298 , n71297 );
buf ( n71299 , n58982 );
or ( n71300 , n71298 , n71299 );
nand ( n71301 , n71289 , n71300 );
buf ( n71302 , n71301 );
buf ( n71303 , n71302 );
buf ( n71304 , n55129 );
not ( n71305 , n55019 );
nand ( n71306 , n71305 , n55021 );
xor ( n71307 , n71306 , n55015 );
buf ( n71308 , n71307 );
not ( n71309 , n71308 );
buf ( n71310 , n71309 );
buf ( n71311 , n71310 );
or ( n71312 , n71304 , n71311 );
buf ( n71313 , n56598 );
buf ( n71314 , n71228 );
or ( n71315 , n71313 , n71314 );
nand ( n71316 , n71312 , n71315 );
buf ( n71317 , n71316 );
buf ( n71318 , n71317 );
buf ( n71319 , n56670 );
not ( n71320 , n71319 );
buf ( n71321 , n71204 );
not ( n71322 , n71321 );
buf ( n71323 , n71322 );
buf ( n71324 , n71323 );
not ( n71325 , n71324 );
or ( n71326 , n71320 , n71325 );
buf ( n71327 , n55195 );
buf ( n71328 , n71232 );
and ( n71329 , n71327 , n71328 );
not ( n71330 , n71327 );
buf ( n71331 , n71235 );
and ( n71332 , n71330 , n71331 );
nor ( n71333 , n71329 , n71332 );
buf ( n71334 , n71333 );
buf ( n71335 , n71334 );
buf ( n71336 , n56664 );
or ( n71337 , n71335 , n71336 );
nand ( n71338 , n71326 , n71337 );
buf ( n71339 , n71338 );
buf ( n71340 , n71339 );
and ( n71341 , n71318 , n71340 );
buf ( n71342 , n71341 );
buf ( n71343 , n71342 );
xor ( n71344 , n71303 , n71343 );
xor ( n71345 , n71221 , n71241 );
xor ( n71346 , n71345 , n71272 );
buf ( n71347 , n71346 );
buf ( n71348 , n71347 );
and ( n71349 , n71344 , n71348 );
and ( n71350 , n71303 , n71343 );
or ( n71351 , n71349 , n71350 );
buf ( n71352 , n71351 );
buf ( n71353 , n71352 );
and ( n71354 , n71278 , n71353 );
and ( n71355 , n71196 , n71277 );
or ( n71356 , n71354 , n71355 );
buf ( n71357 , n71356 );
buf ( n71358 , n71357 );
xor ( n71359 , n71171 , n71358 );
buf ( n71360 , n62643 );
buf ( n71361 , n62681 );
and ( n71362 , n71360 , n71361 );
buf ( n71363 , n62646 );
buf ( n71364 , n62663 );
and ( n71365 , n71363 , n71364 );
nor ( n71366 , n71362 , n71365 );
buf ( n71367 , n71366 );
buf ( n71368 , n71367 );
buf ( n71369 , n62935 );
or ( n71370 , n71368 , n71369 );
buf ( n71371 , n60229 );
buf ( n71372 , n62681 );
and ( n71373 , n71371 , n71372 );
buf ( n71374 , n62652 );
buf ( n71375 , n62663 );
and ( n71376 , n71374 , n71375 );
nor ( n71377 , n71373 , n71376 );
buf ( n71378 , n71377 );
buf ( n71379 , n71378 );
buf ( n71380 , n62676 );
or ( n71381 , n71379 , n71380 );
nand ( n71382 , n71370 , n71381 );
buf ( n71383 , n71382 );
buf ( n71384 , n71383 );
buf ( n71385 , n62971 );
buf ( n71386 , n60261 );
and ( n71387 , n71385 , n71386 );
buf ( n71388 , n62974 );
buf ( n71389 , n60090 );
and ( n71390 , n71388 , n71389 );
nor ( n71391 , n71387 , n71390 );
buf ( n71392 , n71391 );
buf ( n71393 , n71392 );
buf ( n71394 , n60270 );
or ( n71395 , n71393 , n71394 );
buf ( n71396 , n62782 );
buf ( n71397 , n60261 );
and ( n71398 , n71396 , n71397 );
buf ( n71399 , n62980 );
buf ( n71400 , n60090 );
and ( n71401 , n71399 , n71400 );
nor ( n71402 , n71398 , n71401 );
buf ( n71403 , n71402 );
buf ( n71404 , n71403 );
buf ( n71405 , n60100 );
or ( n71406 , n71404 , n71405 );
nand ( n71407 , n71395 , n71406 );
buf ( n71408 , n71407 );
buf ( n71409 , n71408 );
xor ( n71410 , n71384 , n71409 );
buf ( n71411 , n55129 );
buf ( n71412 , n71235 );
or ( n71413 , n71411 , n71412 );
buf ( n71414 , n70530 );
buf ( n71415 , n56598 );
or ( n71416 , n71414 , n71415 );
nand ( n71417 , n71413 , n71416 );
buf ( n71418 , n71417 );
buf ( n71419 , n71418 );
buf ( n71420 , n71215 );
buf ( n71421 , n56664 );
or ( n71422 , n71420 , n71421 );
buf ( n71423 , n70516 );
buf ( n71424 , n56673 );
or ( n71425 , n71423 , n71424 );
nand ( n71426 , n71422 , n71425 );
buf ( n71427 , n71426 );
buf ( n71428 , n71427 );
xor ( n71429 , n71419 , n71428 );
buf ( n71430 , n71429 );
buf ( n71431 , n71430 );
buf ( n71432 , n71252 );
buf ( n71433 , n56626 );
or ( n71434 , n71432 , n71433 );
buf ( n71435 , n70550 );
buf ( n71436 , n56639 );
or ( n71437 , n71435 , n71436 );
nand ( n71438 , n71434 , n71437 );
buf ( n71439 , n71438 );
buf ( n71440 , n71439 );
xor ( n71441 , n71431 , n71440 );
buf ( n71442 , n71297 );
buf ( n71443 , n56799 );
or ( n71444 , n71442 , n71443 );
buf ( n71445 , n66601 );
buf ( n71446 , n58721 );
and ( n71447 , n71445 , n71446 );
buf ( n71448 , n66604 );
buf ( n71449 , n58718 );
and ( n71450 , n71448 , n71449 );
nor ( n71451 , n71447 , n71450 );
buf ( n71452 , n71451 );
buf ( n71453 , n71452 );
buf ( n71454 , n58982 );
or ( n71455 , n71453 , n71454 );
nand ( n71456 , n71444 , n71455 );
buf ( n71457 , n71456 );
buf ( n71458 , n71457 );
xor ( n71459 , n71441 , n71458 );
buf ( n71460 , n71459 );
buf ( n71461 , n71460 );
and ( n71462 , n71410 , n71461 );
and ( n71463 , n71384 , n71409 );
or ( n71464 , n71462 , n71463 );
buf ( n71465 , n71464 );
buf ( n71466 , n71465 );
and ( n71467 , n71359 , n71466 );
and ( n71468 , n71171 , n71358 );
or ( n71469 , n71467 , n71468 );
buf ( n71470 , n71469 );
buf ( n71471 , n58857 );
buf ( n71472 , n64129 );
and ( n71473 , n71471 , n71472 );
buf ( n71474 , n58858 );
buf ( n71475 , n64133 );
and ( n71476 , n71474 , n71475 );
nor ( n71477 , n71473 , n71476 );
buf ( n71478 , n71477 );
buf ( n71479 , n71478 );
buf ( n71480 , n64141 );
or ( n71481 , n71479 , n71480 );
buf ( n71482 , n58823 );
buf ( n71483 , n64129 );
and ( n71484 , n71482 , n71483 );
buf ( n71485 , n58862 );
buf ( n71486 , n64133 );
and ( n71487 , n71485 , n71486 );
nor ( n71488 , n71484 , n71487 );
buf ( n71489 , n71488 );
buf ( n71490 , n71489 );
buf ( n71491 , n63010 );
or ( n71492 , n71490 , n71491 );
nand ( n71493 , n71481 , n71492 );
buf ( n71494 , n71493 );
or ( n71495 , n71165 , n64230 );
not ( n71496 , n64227 );
nand ( n71497 , n71496 , n70678 );
nand ( n71498 , n71495 , n71497 );
xor ( n71499 , n71494 , n71498 );
xor ( n71500 , n71431 , n71440 );
and ( n71501 , n71500 , n71458 );
and ( n71502 , n71431 , n71440 );
or ( n71503 , n71501 , n71502 );
buf ( n71504 , n71503 );
buf ( n71505 , n71504 );
buf ( n71506 , n71190 );
buf ( n71507 , n58913 );
or ( n71508 , n71506 , n71507 );
buf ( n71509 , n62971 );
buf ( n71510 , n58897 );
and ( n71511 , n71509 , n71510 );
buf ( n71512 , n62974 );
buf ( n71513 , n68170 );
and ( n71514 , n71512 , n71513 );
nor ( n71515 , n71511 , n71514 );
buf ( n71516 , n71515 );
buf ( n71517 , n71516 );
buf ( n71518 , n58890 );
or ( n71519 , n71517 , n71518 );
nand ( n71520 , n71508 , n71519 );
buf ( n71521 , n71520 );
buf ( n71522 , n71521 );
xor ( n71523 , n71505 , n71522 );
buf ( n71524 , n71378 );
buf ( n71525 , n62935 );
or ( n71526 , n71524 , n71525 );
buf ( n71527 , n60068 );
buf ( n71528 , n62681 );
and ( n71529 , n71527 , n71528 );
buf ( n71530 , n60071 );
buf ( n71531 , n62663 );
and ( n71532 , n71530 , n71531 );
nor ( n71533 , n71529 , n71532 );
buf ( n71534 , n71533 );
buf ( n71535 , n71534 );
buf ( n71536 , n62676 );
or ( n71537 , n71535 , n71536 );
nand ( n71538 , n71526 , n71537 );
buf ( n71539 , n71538 );
buf ( n71540 , n71539 );
and ( n71541 , n71523 , n71540 );
and ( n71542 , n71505 , n71522 );
or ( n71543 , n71541 , n71542 );
buf ( n71544 , n71543 );
xor ( n71545 , n71499 , n71544 );
and ( n71546 , n71470 , n71545 );
buf ( n71547 , n71452 );
buf ( n71548 , n56799 );
or ( n71549 , n71547 , n71548 );
buf ( n71550 , n64211 );
buf ( n71551 , n58721 );
and ( n71552 , n71550 , n71551 );
buf ( n71553 , n66610 );
buf ( n71554 , n58718 );
and ( n71555 , n71553 , n71554 );
nor ( n71556 , n71552 , n71555 );
buf ( n71557 , n71556 );
buf ( n71558 , n71557 );
buf ( n71559 , n58982 );
or ( n71560 , n71558 , n71559 );
nand ( n71561 , n71549 , n71560 );
buf ( n71562 , n71561 );
buf ( n71563 , n71562 );
and ( n71564 , n71419 , n71428 );
buf ( n71565 , n71564 );
buf ( n71566 , n71565 );
xor ( n71567 , n71563 , n71566 );
xor ( n71568 , n70525 , n70539 );
xor ( n71569 , n71568 , n70562 );
buf ( n71570 , n71569 );
buf ( n71571 , n71570 );
xor ( n71572 , n71567 , n71571 );
buf ( n71573 , n71572 );
buf ( n71574 , n71403 );
buf ( n71575 , n60270 );
or ( n71576 , n71574 , n71575 );
buf ( n71577 , n62643 );
buf ( n71578 , n60261 );
and ( n71579 , n71577 , n71578 );
buf ( n71580 , n62646 );
buf ( n71581 , n60090 );
and ( n71582 , n71580 , n71581 );
nor ( n71583 , n71579 , n71582 );
buf ( n71584 , n71583 );
buf ( n71585 , n71584 );
buf ( n71586 , n60100 );
or ( n71587 , n71585 , n71586 );
nand ( n71588 , n71576 , n71587 );
buf ( n71589 , n71588 );
xor ( n71590 , n71573 , n71589 );
buf ( n71591 , n59009 );
buf ( n71592 , n64129 );
and ( n71593 , n71591 , n71592 );
buf ( n71594 , n60077 );
buf ( n71595 , n64133 );
and ( n71596 , n71594 , n71595 );
nor ( n71597 , n71593 , n71596 );
buf ( n71598 , n71597 );
buf ( n71599 , n71598 );
buf ( n71600 , n64141 );
or ( n71601 , n71599 , n71600 );
buf ( n71602 , n71478 );
buf ( n71603 , n63010 );
or ( n71604 , n71602 , n71603 );
nand ( n71605 , n71601 , n71604 );
buf ( n71606 , n71605 );
and ( n71607 , n71590 , n71606 );
and ( n71608 , n71573 , n71589 );
or ( n71609 , n71607 , n71608 );
buf ( n71610 , n71609 );
buf ( n71611 , n71516 );
buf ( n71612 , n58913 );
or ( n71613 , n71611 , n71612 );
buf ( n71614 , n70469 );
buf ( n71615 , n58890 );
or ( n71616 , n71614 , n71615 );
nand ( n71617 , n71613 , n71616 );
buf ( n71618 , n71617 );
buf ( n71619 , n71618 );
buf ( n71620 , n71557 );
buf ( n71621 , n56799 );
or ( n71622 , n71620 , n71621 );
buf ( n71623 , n70605 );
buf ( n71624 , n58982 );
or ( n71625 , n71623 , n71624 );
nand ( n71626 , n71622 , n71625 );
buf ( n71627 , n71626 );
buf ( n71628 , n71627 );
xor ( n71629 , n71619 , n71628 );
buf ( n71630 , n71584 );
buf ( n71631 , n60270 );
or ( n71632 , n71630 , n71631 );
buf ( n71633 , n70452 );
buf ( n71634 , n60100 );
or ( n71635 , n71633 , n71634 );
nand ( n71636 , n71632 , n71635 );
buf ( n71637 , n71636 );
buf ( n71638 , n71637 );
xor ( n71639 , n71629 , n71638 );
buf ( n71640 , n71639 );
buf ( n71641 , n71640 );
xor ( n71642 , n71610 , n71641 );
xor ( n71643 , n70482 , n70507 );
xor ( n71644 , n71643 , n70567 );
buf ( n71645 , n71644 );
buf ( n71646 , n71645 );
xor ( n71647 , n71563 , n71566 );
and ( n71648 , n71647 , n71571 );
and ( n71649 , n71563 , n71566 );
or ( n71650 , n71648 , n71649 );
buf ( n71651 , n71650 );
buf ( n71652 , n71651 );
xor ( n71653 , n71646 , n71652 );
buf ( n71654 , n71534 );
buf ( n71655 , n62935 );
or ( n71656 , n71654 , n71655 );
buf ( n71657 , n70689 );
buf ( n71658 , n62676 );
or ( n71659 , n71657 , n71658 );
nand ( n71660 , n71656 , n71659 );
buf ( n71661 , n71660 );
buf ( n71662 , n71661 );
xor ( n71663 , n71653 , n71662 );
buf ( n71664 , n71663 );
buf ( n71665 , n71664 );
xor ( n71666 , n71642 , n71665 );
buf ( n71667 , n71666 );
xor ( n71668 , n71494 , n71498 );
xor ( n71669 , n71668 , n71544 );
and ( n71670 , n71667 , n71669 );
and ( n71671 , n71470 , n71667 );
or ( n71672 , n71546 , n71670 , n71671 );
not ( n71673 , n71672 );
xor ( n71674 , n71610 , n71641 );
and ( n71675 , n71674 , n71665 );
and ( n71676 , n71610 , n71641 );
or ( n71677 , n71675 , n71676 );
buf ( n71678 , n71677 );
buf ( n71679 , n71678 );
xor ( n71680 , n71619 , n71628 );
and ( n71681 , n71680 , n71638 );
and ( n71682 , n71619 , n71628 );
or ( n71683 , n71681 , n71682 );
buf ( n71684 , n71683 );
buf ( n71685 , n71684 );
buf ( n71686 , n71489 );
buf ( n71687 , n64141 );
or ( n71688 , n71686 , n71687 );
buf ( n71689 , n70644 );
buf ( n71690 , n63010 );
or ( n71691 , n71689 , n71690 );
nand ( n71692 , n71688 , n71691 );
buf ( n71693 , n71692 );
buf ( n71694 , n71693 );
xor ( n71695 , n71685 , n71694 );
xor ( n71696 , n70461 , n70478 );
xor ( n71697 , n71696 , n70572 );
buf ( n71698 , n71697 );
buf ( n71699 , n71698 );
xor ( n71700 , n71695 , n71699 );
buf ( n71701 , n71700 );
buf ( n71702 , n71701 );
xor ( n71703 , n71679 , n71702 );
xor ( n71704 , n71494 , n71498 );
and ( n71705 , n71704 , n71544 );
and ( n71706 , n71494 , n71498 );
or ( n71707 , n71705 , n71706 );
buf ( n71708 , n71707 );
xor ( n71709 , n71646 , n71652 );
and ( n71710 , n71709 , n71662 );
and ( n71711 , n71646 , n71652 );
or ( n71712 , n71710 , n71711 );
buf ( n71713 , n71712 );
buf ( n71714 , n71713 );
xor ( n71715 , n71708 , n71714 );
xor ( n71716 , n70681 , n70698 );
xor ( n71717 , n71716 , n70703 );
buf ( n71718 , n71717 );
buf ( n71719 , n71718 );
xor ( n71720 , n71715 , n71719 );
buf ( n71721 , n71720 );
buf ( n71722 , n71721 );
xor ( n71723 , n71703 , n71722 );
buf ( n71724 , n71723 );
not ( n71725 , n71724 );
or ( n71726 , n71673 , n71725 );
not ( n71727 , n71672 );
not ( n71728 , n71724 );
and ( n71729 , n71727 , n71728 );
not ( n71730 , n71729 );
xor ( n71731 , n71494 , n71498 );
xor ( n71732 , n71731 , n71544 );
xor ( n71733 , n71470 , n71667 );
xor ( n71734 , n71732 , n71733 );
buf ( n71735 , n71734 );
xor ( n71736 , n71505 , n71522 );
xor ( n71737 , n71736 , n71540 );
buf ( n71738 , n71737 );
xor ( n71739 , n71573 , n71589 );
xor ( n71740 , n71739 , n71606 );
and ( n71741 , n71738 , n71740 );
buf ( n71742 , n60068 );
buf ( n71743 , n64129 );
and ( n71744 , n71742 , n71743 );
buf ( n71745 , n60071 );
buf ( n71746 , n64133 );
and ( n71747 , n71745 , n71746 );
nor ( n71748 , n71744 , n71747 );
buf ( n71749 , n71748 );
buf ( n71750 , n71749 );
buf ( n71751 , n64141 );
or ( n71752 , n71750 , n71751 );
buf ( n71753 , n71598 );
buf ( n71754 , n63010 );
or ( n71755 , n71753 , n71754 );
nand ( n71756 , n71752 , n71755 );
buf ( n71757 , n71756 );
buf ( n71758 , n71757 );
buf ( n71759 , n70348 );
buf ( n71760 , n56641 );
and ( n71761 , n71759 , n71760 );
buf ( n71762 , n70351 );
buf ( n71763 , n56631 );
and ( n71764 , n71762 , n71763 );
nor ( n71765 , n71761 , n71764 );
buf ( n71766 , n71765 );
buf ( n71767 , n71766 );
buf ( n71768 , n56626 );
or ( n71769 , n71767 , n71768 );
buf ( n71770 , n71266 );
buf ( n71771 , n56639 );
or ( n71772 , n71770 , n71771 );
nand ( n71773 , n71769 , n71772 );
buf ( n71774 , n71773 );
buf ( n71775 , n71774 );
buf ( n71776 , n56664 );
buf ( n71777 , n71225 );
buf ( n71778 , n55195 );
and ( n71779 , n71777 , n71778 );
buf ( n71780 , n71228 );
buf ( n71781 , n55184 );
and ( n71782 , n71780 , n71781 );
nor ( n71783 , n71779 , n71782 );
buf ( n71784 , n71783 );
buf ( n71785 , n71784 );
or ( n71786 , n71776 , n71785 );
buf ( n71787 , n71334 );
buf ( n71788 , n56673 );
or ( n71789 , n71787 , n71788 );
nand ( n71790 , n71786 , n71789 );
buf ( n71791 , n71790 );
buf ( n71792 , n55129 );
not ( n71793 , n55013 );
nor ( n71794 , n71793 , n55004 );
not ( n71795 , n71794 );
not ( n71796 , n54991 );
nor ( n71797 , n71796 , n55011 );
not ( n71798 , n71797 );
or ( n71799 , n71795 , n71798 );
or ( n71800 , n71797 , n71794 );
nand ( n71801 , n71799 , n71800 );
buf ( n71802 , n71801 );
not ( n71803 , n71802 );
buf ( n71804 , n71803 );
buf ( n71805 , n71804 );
or ( n71806 , n71792 , n71805 );
buf ( n71807 , n55125 );
buf ( n71808 , n71310 );
or ( n71809 , n71807 , n71808 );
nand ( n71810 , n71806 , n71809 );
buf ( n71811 , n71810 );
xor ( n71812 , n71791 , n71811 );
buf ( n71813 , n55129 );
not ( n71814 , n55011 );
or ( n71815 , n55008 , n621 );
nand ( n71816 , n71815 , n55009 , n55010 );
nand ( n71817 , n71814 , n71816 );
xnor ( n71818 , n71817 , n54990 );
buf ( n71819 , n71818 );
not ( n71820 , n71819 );
buf ( n71821 , n71820 );
buf ( n71822 , n71821 );
or ( n71823 , n71813 , n71822 );
buf ( n71824 , n55125 );
buf ( n71825 , n71804 );
or ( n71826 , n71824 , n71825 );
nand ( n71827 , n71823 , n71826 );
buf ( n71828 , n71827 );
buf ( n71829 , n71828 );
buf ( n71830 , n56664 );
buf ( n71831 , n55195 );
buf ( n71832 , n71307 );
and ( n71833 , n71831 , n71832 );
buf ( n71834 , n55184 );
buf ( n71835 , n71310 );
and ( n71836 , n71834 , n71835 );
nor ( n71837 , n71833 , n71836 );
buf ( n71838 , n71837 );
buf ( n71839 , n71838 );
or ( n71840 , n71830 , n71839 );
buf ( n71841 , n71784 );
buf ( n71842 , n55166 );
or ( n71843 , n71841 , n71842 );
nand ( n71844 , n71840 , n71843 );
buf ( n71845 , n71844 );
buf ( n71846 , n71845 );
and ( n71847 , n71829 , n71846 );
buf ( n71848 , n71847 );
and ( n71849 , n71812 , n71848 );
and ( n71850 , n71791 , n71811 );
or ( n71851 , n71849 , n71850 );
buf ( n71852 , n71851 );
xor ( n71853 , n71775 , n71852 );
xor ( n71854 , n71318 , n71340 );
buf ( n71855 , n71854 );
buf ( n71856 , n71855 );
and ( n71857 , n71853 , n71856 );
and ( n71858 , n71775 , n71852 );
or ( n71859 , n71857 , n71858 );
buf ( n71860 , n71859 );
buf ( n71861 , n66601 );
buf ( n71862 , n58897 );
and ( n71863 , n71861 , n71862 );
buf ( n71864 , n66604 );
buf ( n71865 , n68170 );
and ( n71866 , n71864 , n71865 );
nor ( n71867 , n71863 , n71866 );
buf ( n71868 , n71867 );
buf ( n71869 , n71868 );
buf ( n71870 , n58913 );
or ( n71871 , n71869 , n71870 );
buf ( n71872 , n71179 );
buf ( n71873 , n58890 );
or ( n71874 , n71872 , n71873 );
nand ( n71875 , n71871 , n71874 );
buf ( n71876 , n71875 );
xor ( n71877 , n71860 , n71876 );
buf ( n71878 , n64068 );
buf ( n71879 , n60261 );
and ( n71880 , n71878 , n71879 );
buf ( n71881 , n66579 );
buf ( n71882 , n60090 );
and ( n71883 , n71881 , n71882 );
nor ( n71884 , n71880 , n71883 );
buf ( n71885 , n71884 );
buf ( n71886 , n71885 );
buf ( n71887 , n60270 );
or ( n71888 , n71886 , n71887 );
buf ( n71889 , n71392 );
buf ( n71890 , n60100 );
or ( n71891 , n71889 , n71890 );
nand ( n71892 , n71888 , n71891 );
buf ( n71893 , n71892 );
and ( n71894 , n71877 , n71893 );
and ( n71895 , n71860 , n71876 );
or ( n71896 , n71894 , n71895 );
buf ( n71897 , n71896 );
xor ( n71898 , n71758 , n71897 );
xor ( n71899 , n71196 , n71277 );
xor ( n71900 , n71899 , n71353 );
buf ( n71901 , n71900 );
buf ( n71902 , n71901 );
and ( n71903 , n71898 , n71902 );
and ( n71904 , n71758 , n71897 );
or ( n71905 , n71903 , n71904 );
buf ( n71906 , n71905 );
xor ( n71907 , n71573 , n71589 );
xor ( n71908 , n71907 , n71606 );
and ( n71909 , n71906 , n71908 );
and ( n71910 , n71738 , n71906 );
or ( n71911 , n71741 , n71909 , n71910 );
buf ( n71912 , n71911 );
xor ( n71913 , n71735 , n71912 );
buf ( n71914 , n60229 );
buf ( n71915 , n64129 );
and ( n71916 , n71914 , n71915 );
buf ( n71917 , n62652 );
buf ( n71918 , n64133 );
and ( n71919 , n71917 , n71918 );
nor ( n71920 , n71916 , n71919 );
buf ( n71921 , n71920 );
buf ( n71922 , n71921 );
buf ( n71923 , n64141 );
or ( n71924 , n71922 , n71923 );
buf ( n71925 , n71749 );
buf ( n71926 , n63010 );
or ( n71927 , n71925 , n71926 );
nand ( n71928 , n71924 , n71927 );
buf ( n71929 , n71928 );
buf ( n71930 , n71929 );
xor ( n71931 , n71303 , n71343 );
xor ( n71932 , n71931 , n71348 );
buf ( n71933 , n71932 );
buf ( n71934 , n71933 );
xor ( n71935 , n71930 , n71934 );
buf ( n71936 , n66690 );
buf ( n71937 , n58897 );
and ( n71938 , n71936 , n71937 );
buf ( n71939 , n66693 );
buf ( n71940 , n68170 );
and ( n71941 , n71939 , n71940 );
nor ( n71942 , n71938 , n71941 );
buf ( n71943 , n71942 );
buf ( n71944 , n71943 );
buf ( n71945 , n58913 );
or ( n71946 , n71944 , n71945 );
buf ( n71947 , n71868 );
buf ( n71948 , n58890 );
or ( n71949 , n71947 , n71948 );
nand ( n71950 , n71946 , n71949 );
buf ( n71951 , n71950 );
buf ( n71952 , n71951 );
buf ( n71953 , n68235 );
buf ( n71954 , n58718 );
or ( n71955 , n71953 , n71954 );
buf ( n71956 , n68232 );
buf ( n71957 , n56777 );
or ( n71958 , n71956 , n71957 );
nand ( n71959 , n71955 , n71958 );
buf ( n71960 , n71959 );
buf ( n71961 , n71960 );
not ( n71962 , n71961 );
buf ( n71963 , n71962 );
buf ( n71964 , n71963 );
buf ( n71965 , n56799 );
or ( n71966 , n71964 , n71965 );
buf ( n71967 , n71286 );
buf ( n71968 , n58982 );
or ( n71969 , n71967 , n71968 );
nand ( n71970 , n71966 , n71969 );
buf ( n71971 , n71970 );
buf ( n71972 , n71971 );
xor ( n71973 , n71952 , n71972 );
buf ( n71974 , n70527 );
buf ( n71975 , n56641 );
and ( n71976 , n71974 , n71975 );
buf ( n71977 , n70530 );
buf ( n71978 , n56631 );
and ( n71979 , n71977 , n71978 );
nor ( n71980 , n71976 , n71979 );
buf ( n71981 , n71980 );
buf ( n71982 , n71981 );
buf ( n71983 , n56626 );
or ( n71984 , n71982 , n71983 );
buf ( n71985 , n71766 );
buf ( n71986 , n56639 );
or ( n71987 , n71985 , n71986 );
nand ( n71988 , n71984 , n71987 );
buf ( n71989 , n71988 );
xor ( n71990 , n71791 , n71811 );
xor ( n71991 , n71990 , n71848 );
and ( n71992 , n71989 , n71991 );
buf ( n71993 , n56811 );
not ( n71994 , n71993 );
buf ( n71995 , n71960 );
not ( n71996 , n71995 );
or ( n71997 , n71994 , n71996 );
buf ( n71998 , n70333 );
buf ( n71999 , n56777 );
and ( n72000 , n71998 , n71999 );
buf ( n72001 , n70336 );
buf ( n72002 , n58718 );
and ( n72003 , n72001 , n72002 );
nor ( n72004 , n72000 , n72003 );
buf ( n72005 , n72004 );
buf ( n72006 , n72005 );
buf ( n72007 , n56799 );
or ( n72008 , n72006 , n72007 );
nand ( n72009 , n71997 , n72008 );
buf ( n72010 , n72009 );
xor ( n72011 , n71791 , n71811 );
xor ( n72012 , n72011 , n71848 );
and ( n72013 , n72010 , n72012 );
and ( n72014 , n71989 , n72010 );
or ( n72015 , n71992 , n72013 , n72014 );
buf ( n72016 , n72015 );
and ( n72017 , n71973 , n72016 );
and ( n72018 , n71952 , n71972 );
or ( n72019 , n72017 , n72018 );
buf ( n72020 , n72019 );
buf ( n72021 , n72020 );
and ( n72022 , n71935 , n72021 );
and ( n72023 , n71930 , n71934 );
or ( n72024 , n72022 , n72023 );
buf ( n72025 , n72024 );
buf ( n72026 , n72025 );
buf ( n72027 , n58857 );
buf ( n72028 , n66742 );
and ( n72029 , n72027 , n72028 );
buf ( n72030 , n58858 );
buf ( n72031 , n63000 );
and ( n72032 , n72030 , n72031 );
nor ( n72033 , n72029 , n72032 );
buf ( n72034 , n72033 );
buf ( n72035 , n72034 );
buf ( n72036 , n64230 );
or ( n72037 , n72035 , n72036 );
buf ( n72038 , n71154 );
buf ( n72039 , n64227 );
or ( n72040 , n72038 , n72039 );
nand ( n72041 , n72037 , n72040 );
buf ( n72042 , n72041 );
buf ( n72043 , n72042 );
xor ( n72044 , n72026 , n72043 );
xor ( n72045 , n71384 , n71409 );
xor ( n72046 , n72045 , n71461 );
buf ( n72047 , n72046 );
buf ( n72048 , n72047 );
and ( n72049 , n72044 , n72048 );
and ( n72050 , n72026 , n72043 );
or ( n72051 , n72049 , n72050 );
buf ( n72052 , n72051 );
xor ( n72053 , n71171 , n71358 );
xor ( n72054 , n72053 , n71466 );
buf ( n72055 , n72054 );
xor ( n72056 , n72052 , n72055 );
xor ( n72057 , n71573 , n71589 );
xor ( n72058 , n72057 , n71606 );
xor ( n72059 , n71738 , n71906 );
xor ( n72060 , n72058 , n72059 );
and ( n72061 , n72056 , n72060 );
and ( n72062 , n72052 , n72055 );
or ( n72063 , n72061 , n72062 );
buf ( n72064 , n72063 );
and ( n72065 , n71913 , n72064 );
and ( n72066 , n71735 , n71912 );
or ( n72067 , n72065 , n72066 );
buf ( n72068 , n72067 );
nand ( n72069 , n71730 , n72068 );
nand ( n72070 , n71726 , n72069 );
xor ( n72071 , n71679 , n71702 );
and ( n72072 , n72071 , n71722 );
and ( n72073 , n71679 , n71702 );
or ( n72074 , n72072 , n72073 );
buf ( n72075 , n72074 );
xor ( n72076 , n70429 , n70443 );
xor ( n72077 , n72076 , n70576 );
xor ( n72078 , n71685 , n71694 );
and ( n72079 , n72078 , n71699 );
and ( n72080 , n71685 , n71694 );
or ( n72081 , n72079 , n72080 );
buf ( n72082 , n72081 );
xor ( n72083 , n70708 , n70712 );
xor ( n72084 , n72083 , n70717 );
buf ( n72085 , n72084 );
xor ( n72086 , n72082 , n72085 );
xor ( n72087 , n72077 , n72086 );
xor ( n72088 , n71708 , n71714 );
and ( n72089 , n72088 , n71719 );
and ( n72090 , n71708 , n71714 );
or ( n72091 , n72089 , n72090 );
buf ( n72092 , n72091 );
or ( n72093 , n72087 , n72092 );
not ( n72094 , n72093 );
and ( n72095 , n72075 , n72094 );
nand ( n72096 , n72087 , n72092 );
not ( n72097 , n72096 );
and ( n72098 , n72097 , n72075 );
nor ( n72099 , n72095 , n72098 );
not ( n72100 , n72087 );
not ( n72101 , n72075 );
nand ( n72102 , n72100 , n72101 , n72092 );
not ( n72103 , n72092 );
nand ( n72104 , n72103 , n72101 , n72087 );
and ( n72105 , n72099 , n72102 , n72104 );
and ( n72106 , n72070 , n72105 );
not ( n72107 , n72070 );
not ( n72108 , n72105 );
and ( n72109 , n72107 , n72108 );
nor ( n72110 , n72106 , n72109 );
and ( n72111 , n71146 , n72110 );
not ( n72112 , n71146 );
not ( n72113 , n72110 );
and ( n72114 , n72112 , n72113 );
nor ( n72115 , n72111 , n72114 );
buf ( n72116 , n72115 );
buf ( n72117 , n44496 );
not ( n72118 , n72117 );
buf ( n72119 , n44533 );
not ( n72120 , n72119 );
buf ( n72121 , n66426 );
not ( n72122 , n72121 );
or ( n72123 , n72120 , n72122 );
buf ( n72124 , n13662 );
buf ( n72125 , n44530 );
nand ( n72126 , n72124 , n72125 );
buf ( n72127 , n72126 );
buf ( n72128 , n72127 );
nand ( n72129 , n72123 , n72128 );
buf ( n72130 , n72129 );
buf ( n72131 , n72130 );
not ( n72132 , n72131 );
or ( n72133 , n72118 , n72132 );
buf ( n72134 , n44533 );
not ( n72135 , n72134 );
buf ( n72136 , n63633 );
not ( n72137 , n72136 );
or ( n72138 , n72135 , n72137 );
buf ( n72139 , n29463 );
buf ( n72140 , n44530 );
nand ( n72141 , n72139 , n72140 );
buf ( n72142 , n72141 );
buf ( n72143 , n72142 );
nand ( n72144 , n72138 , n72143 );
buf ( n72145 , n72144 );
buf ( n72146 , n72145 );
buf ( n72147 , n44517 );
nand ( n72148 , n72146 , n72147 );
buf ( n72149 , n72148 );
buf ( n72150 , n72149 );
nand ( n72151 , n72133 , n72150 );
buf ( n72152 , n72151 );
buf ( n72153 , n72152 );
xor ( n72154 , n72116 , n72153 );
and ( n72155 , n47716 , n42366 );
not ( n72156 , n47716 );
and ( n72157 , n72156 , n63913 );
nor ( n72158 , n72155 , n72157 );
not ( n72159 , n72158 );
not ( n72160 , n42374 );
or ( n72161 , n72159 , n72160 );
or ( n72162 , n42342 , n46393 );
or ( n72163 , n46390 , n24951 );
nand ( n72164 , n72162 , n72163 );
or ( n72165 , n42333 , n72164 );
nand ( n72166 , n72161 , n72165 );
buf ( n72167 , n72166 );
and ( n72168 , n72154 , n72167 );
and ( n72169 , n72116 , n72153 );
or ( n72170 , n72168 , n72169 );
buf ( n72171 , n72170 );
buf ( n72172 , n72171 );
xor ( n72173 , n71115 , n72172 );
buf ( n72174 , n67149 );
not ( n72175 , n72174 );
buf ( n72176 , n71044 );
not ( n72177 , n72176 );
or ( n72178 , n72175 , n72177 );
buf ( n72179 , n45746 );
not ( n72180 , n72179 );
buf ( n72181 , n63906 );
not ( n72182 , n72181 );
or ( n72183 , n72180 , n72182 );
buf ( n72184 , n13653 );
buf ( n72185 , n45747 );
nand ( n72186 , n72184 , n72185 );
buf ( n72187 , n72186 );
buf ( n72188 , n72187 );
nand ( n72189 , n72183 , n72188 );
buf ( n72190 , n72189 );
buf ( n72191 , n72190 );
buf ( n72192 , n71048 );
nand ( n72193 , n72191 , n72192 );
buf ( n72194 , n72193 );
buf ( n72195 , n72194 );
nand ( n72196 , n72178 , n72195 );
buf ( n72197 , n72196 );
buf ( n72198 , n72197 );
and ( n72199 , n72173 , n72198 );
and ( n72200 , n71115 , n72172 );
or ( n72201 , n72199 , n72200 );
buf ( n72202 , n72201 );
buf ( n72203 , n72202 );
xor ( n72204 , n71075 , n72203 );
buf ( n72205 , n72204 );
buf ( n72206 , n72205 );
xor ( n72207 , n71727 , n71728 );
xor ( n72208 , n72207 , n72068 );
buf ( n72209 , n41574 );
not ( n72210 , n72209 );
buf ( n72211 , n41605 );
not ( n72212 , n72211 );
not ( n72213 , n43056 );
buf ( n72214 , n72213 );
not ( n72215 , n72214 );
or ( n72216 , n72212 , n72215 );
buf ( n72217 , n43056 );
buf ( n72218 , n41604 );
nand ( n72219 , n72217 , n72218 );
buf ( n72220 , n72219 );
buf ( n72221 , n72220 );
nand ( n72222 , n72216 , n72221 );
buf ( n72223 , n72222 );
buf ( n72224 , n72223 );
not ( n72225 , n72224 );
or ( n72226 , n72210 , n72225 );
buf ( n72227 , n41596 );
buf ( n72228 , n42228 );
not ( n72229 , n72228 );
buf ( n72230 , n42859 );
not ( n72231 , n72230 );
or ( n72232 , n72229 , n72231 );
buf ( n72233 , n42856 );
not ( n72234 , n72233 );
buf ( n72235 , n72234 );
buf ( n72236 , n72235 );
not ( n72237 , n72236 );
buf ( n72238 , n42228 );
not ( n72239 , n72238 );
buf ( n72240 , n72239 );
buf ( n72241 , n72240 );
nand ( n72242 , n72237 , n72241 );
buf ( n72243 , n72242 );
buf ( n72244 , n72243 );
nand ( n72245 , n72232 , n72244 );
buf ( n72246 , n72245 );
buf ( n72247 , n72246 );
nand ( n72248 , n72227 , n72247 );
buf ( n72249 , n72248 );
buf ( n72250 , n72249 );
nand ( n72251 , n72226 , n72250 );
buf ( n72252 , n72251 );
xor ( n72253 , n72208 , n72252 );
buf ( n72254 , n44949 );
buf ( n72255 , n25303 );
and ( n72256 , n72254 , n72255 );
not ( n72257 , n72254 );
buf ( n72258 , n71123 );
and ( n72259 , n72257 , n72258 );
nor ( n72260 , n72256 , n72259 );
buf ( n72261 , n72260 );
buf ( n72262 , n72261 );
not ( n72263 , n72262 );
buf ( n72264 , n42246 );
not ( n72265 , n72264 );
or ( n72266 , n72263 , n72265 );
buf ( n72267 , n71143 );
buf ( n72268 , n42309 );
nand ( n72269 , n72267 , n72268 );
buf ( n72270 , n72269 );
buf ( n72271 , n72270 );
nand ( n72272 , n72266 , n72271 );
buf ( n72273 , n72272 );
xor ( n72274 , n72253 , n72273 );
not ( n72275 , n72274 );
not ( n72276 , n72275 );
not ( n72277 , n66459 );
buf ( n72278 , n71078 );
not ( n72279 , n72278 );
buf ( n72280 , n42342 );
not ( n72281 , n72280 );
or ( n72282 , n72279 , n72281 );
buf ( n72283 , n65236 );
buf ( n72284 , n48320 );
nand ( n72285 , n72283 , n72284 );
buf ( n72286 , n72285 );
buf ( n72287 , n72286 );
nand ( n72288 , n72282 , n72287 );
buf ( n72289 , n72288 );
not ( n72290 , n72289 );
or ( n72291 , n72277 , n72290 );
buf ( n72292 , n72158 );
buf ( n72293 , n66482 );
nand ( n72294 , n72292 , n72293 );
buf ( n72295 , n72294 );
nand ( n72296 , n72291 , n72295 );
not ( n72297 , n72296 );
not ( n72298 , n72297 );
and ( n72299 , n72276 , n72298 );
not ( n72300 , n72296 );
nand ( n72301 , n72300 , n72275 );
buf ( n72302 , n46114 );
not ( n72303 , n72302 );
buf ( n72304 , n25303 );
not ( n72305 , n72304 );
or ( n72306 , n72303 , n72305 );
buf ( n72307 , n25306 );
buf ( n72308 , n46114 );
not ( n72309 , n72308 );
buf ( n72310 , n72309 );
buf ( n72311 , n72310 );
nand ( n72312 , n72307 , n72311 );
buf ( n72313 , n72312 );
buf ( n72314 , n72313 );
nand ( n72315 , n72306 , n72314 );
buf ( n72316 , n72315 );
buf ( n72317 , n72316 );
not ( n72318 , n72317 );
buf ( n72319 , n42246 );
not ( n72320 , n72319 );
or ( n72321 , n72318 , n72320 );
buf ( n72322 , n72261 );
buf ( n72323 , n42309 );
nand ( n72324 , n72322 , n72323 );
buf ( n72325 , n72324 );
buf ( n72326 , n72325 );
nand ( n72327 , n72321 , n72326 );
buf ( n72328 , n72327 );
buf ( n72329 , n72328 );
xor ( n72330 , n71758 , n71897 );
xor ( n72331 , n72330 , n71902 );
buf ( n72332 , n72331 );
buf ( n72333 , n62782 );
buf ( n72334 , n62681 );
and ( n72335 , n72333 , n72334 );
buf ( n72336 , n62980 );
buf ( n72337 , n62663 );
and ( n72338 , n72336 , n72337 );
nor ( n72339 , n72335 , n72338 );
buf ( n72340 , n72339 );
buf ( n72341 , n72340 );
buf ( n72342 , n62935 );
or ( n72343 , n72341 , n72342 );
buf ( n72344 , n71367 );
buf ( n72345 , n62676 );
or ( n72346 , n72344 , n72345 );
nand ( n72347 , n72343 , n72346 );
buf ( n72348 , n72347 );
xor ( n72349 , n71860 , n71876 );
xor ( n72350 , n72349 , n71893 );
and ( n72351 , n72348 , n72350 );
buf ( n72352 , n59009 );
buf ( n72353 , n66742 );
and ( n72354 , n72352 , n72353 );
buf ( n72355 , n60077 );
buf ( n72356 , n63000 );
and ( n72357 , n72355 , n72356 );
nor ( n72358 , n72354 , n72357 );
buf ( n72359 , n72358 );
buf ( n72360 , n72359 );
buf ( n72361 , n64230 );
or ( n72362 , n72360 , n72361 );
buf ( n72363 , n72034 );
buf ( n72364 , n64227 );
or ( n72365 , n72363 , n72364 );
nand ( n72366 , n72362 , n72365 );
buf ( n72367 , n72366 );
xor ( n72368 , n71860 , n71876 );
xor ( n72369 , n72368 , n71893 );
and ( n72370 , n72367 , n72369 );
and ( n72371 , n72348 , n72367 );
or ( n72372 , n72351 , n72370 , n72371 );
xor ( n72373 , n72332 , n72372 );
xor ( n72374 , n72026 , n72043 );
xor ( n72375 , n72374 , n72048 );
buf ( n72376 , n72375 );
and ( n72377 , n72373 , n72376 );
and ( n72378 , n72332 , n72372 );
or ( n72379 , n72377 , n72378 );
xor ( n72380 , n72052 , n72055 );
xor ( n72381 , n72380 , n72060 );
and ( n72382 , n72379 , n72381 );
buf ( n72383 , n68217 );
buf ( n72384 , n58897 );
and ( n72385 , n72383 , n72384 );
buf ( n72386 , n68220 );
buf ( n72387 , n58894 );
and ( n72388 , n72386 , n72387 );
nor ( n72389 , n72385 , n72388 );
buf ( n72390 , n72389 );
buf ( n72391 , n72390 );
buf ( n72392 , n58913 );
or ( n72393 , n72391 , n72392 );
buf ( n72394 , n71943 );
buf ( n72395 , n58890 );
or ( n72396 , n72394 , n72395 );
nand ( n72397 , n72393 , n72396 );
buf ( n72398 , n72397 );
buf ( n72399 , n72398 );
buf ( n72400 , n71235 );
buf ( n72401 , n56631 );
or ( n72402 , n72400 , n72401 );
buf ( n72403 , n71232 );
buf ( n72404 , n16469 );
or ( n72405 , n72403 , n72404 );
nand ( n72406 , n72402 , n72405 );
buf ( n72407 , n72406 );
buf ( n72408 , n72407 );
not ( n72409 , n72408 );
buf ( n72410 , n72409 );
buf ( n72411 , n72410 );
buf ( n72412 , n56626 );
or ( n72413 , n72411 , n72412 );
buf ( n72414 , n71981 );
buf ( n72415 , n56639 );
or ( n72416 , n72414 , n72415 );
nand ( n72417 , n72413 , n72416 );
buf ( n72418 , n72417 );
buf ( n72419 , n72418 );
xor ( n72420 , n71829 , n71846 );
buf ( n72421 , n72420 );
buf ( n72422 , n72421 );
xor ( n72423 , n72419 , n72422 );
buf ( n72424 , n56664 );
buf ( n72425 , n55184 );
not ( n72426 , n72425 );
buf ( n72427 , n72426 );
buf ( n72428 , n72427 );
buf ( n72429 , n71801 );
and ( n72430 , n72428 , n72429 );
buf ( n72431 , n55184 );
buf ( n72432 , n71804 );
and ( n72433 , n72431 , n72432 );
nor ( n72434 , n72430 , n72433 );
buf ( n72435 , n72434 );
buf ( n72436 , n72435 );
or ( n72437 , n72424 , n72436 );
buf ( n72438 , n71838 );
buf ( n72439 , n55166 );
or ( n72440 , n72438 , n72439 );
nand ( n72441 , n72437 , n72440 );
buf ( n72442 , n72441 );
buf ( n72443 , n72442 );
buf ( n72444 , n55129 );
xor ( n72445 , n54989 , n54988 );
buf ( n72446 , n72445 );
not ( n72447 , n72446 );
buf ( n72448 , n72447 );
buf ( n72449 , n72448 );
or ( n72450 , n72444 , n72449 );
buf ( n72451 , n55125 );
buf ( n72452 , n71821 );
or ( n72453 , n72451 , n72452 );
nand ( n72454 , n72450 , n72453 );
buf ( n72455 , n72454 );
buf ( n72456 , n72455 );
xor ( n72457 , n72443 , n72456 );
buf ( n72458 , n56611 );
not ( n72459 , n72458 );
buf ( n72460 , n72407 );
not ( n72461 , n72460 );
or ( n72462 , n72459 , n72461 );
buf ( n72463 , n56626 );
buf ( n72464 , n71225 );
buf ( n72465 , n16469 );
and ( n72466 , n72464 , n72465 );
buf ( n72467 , n71228 );
buf ( n72468 , n16472 );
and ( n72469 , n72467 , n72468 );
nor ( n72470 , n72466 , n72469 );
buf ( n72471 , n72470 );
buf ( n72472 , n72471 );
or ( n72473 , n72463 , n72472 );
nand ( n72474 , n72462 , n72473 );
buf ( n72475 , n72474 );
buf ( n72476 , n72475 );
and ( n72477 , n72457 , n72476 );
and ( n72478 , n72443 , n72456 );
or ( n72479 , n72477 , n72478 );
buf ( n72480 , n72479 );
buf ( n72481 , n72480 );
and ( n72482 , n72423 , n72481 );
and ( n72483 , n72419 , n72422 );
or ( n72484 , n72482 , n72483 );
buf ( n72485 , n72484 );
buf ( n72486 , n72485 );
xor ( n72487 , n72399 , n72486 );
buf ( n72488 , n60104 );
not ( n72489 , n72488 );
buf ( n72490 , n64211 );
buf ( n72491 , n60261 );
and ( n72492 , n72490 , n72491 );
buf ( n72493 , n66610 );
buf ( n72494 , n60090 );
and ( n72495 , n72493 , n72494 );
nor ( n72496 , n72492 , n72495 );
buf ( n72497 , n72496 );
buf ( n72498 , n72497 );
not ( n72499 , n72498 );
buf ( n72500 , n72499 );
buf ( n72501 , n72500 );
not ( n72502 , n72501 );
or ( n72503 , n72489 , n72502 );
buf ( n72504 , n66601 );
buf ( n72505 , n60261 );
and ( n72506 , n72504 , n72505 );
buf ( n72507 , n66604 );
buf ( n72508 , n60090 );
and ( n72509 , n72507 , n72508 );
nor ( n72510 , n72506 , n72509 );
buf ( n72511 , n72510 );
buf ( n72512 , n72511 );
buf ( n72513 , n60270 );
or ( n72514 , n72512 , n72513 );
nand ( n72515 , n72503 , n72514 );
buf ( n72516 , n72515 );
buf ( n72517 , n72516 );
and ( n72518 , n72487 , n72517 );
and ( n72519 , n72399 , n72486 );
or ( n72520 , n72518 , n72519 );
buf ( n72521 , n72520 );
buf ( n72522 , n72521 );
buf ( n72523 , n62971 );
buf ( n72524 , n62681 );
and ( n72525 , n72523 , n72524 );
buf ( n72526 , n62974 );
buf ( n72527 , n62663 );
and ( n72528 , n72526 , n72527 );
nor ( n72529 , n72525 , n72528 );
buf ( n72530 , n72529 );
buf ( n72531 , n72530 );
buf ( n72532 , n62935 );
or ( n72533 , n72531 , n72532 );
buf ( n72534 , n72340 );
buf ( n72535 , n62676 );
or ( n72536 , n72534 , n72535 );
nand ( n72537 , n72533 , n72536 );
buf ( n72538 , n72537 );
buf ( n72539 , n72538 );
xor ( n72540 , n72522 , n72539 );
xor ( n72541 , n71952 , n71972 );
xor ( n72542 , n72541 , n72016 );
buf ( n72543 , n72542 );
buf ( n72544 , n72543 );
and ( n72545 , n72540 , n72544 );
and ( n72546 , n72522 , n72539 );
or ( n72547 , n72545 , n72546 );
buf ( n72548 , n72547 );
buf ( n72549 , n72548 );
buf ( n72550 , n72497 );
buf ( n72551 , n60270 );
or ( n72552 , n72550 , n72551 );
buf ( n72553 , n71885 );
buf ( n72554 , n60100 );
or ( n72555 , n72553 , n72554 );
nand ( n72556 , n72552 , n72555 );
buf ( n72557 , n72556 );
buf ( n72558 , n72557 );
xor ( n72559 , n71775 , n71852 );
xor ( n72560 , n72559 , n71856 );
buf ( n72561 , n72560 );
buf ( n72562 , n72561 );
xor ( n72563 , n72558 , n72562 );
buf ( n72564 , n63013 );
not ( n72565 , n72564 );
buf ( n72566 , n62643 );
buf ( n72567 , n64129 );
and ( n72568 , n72566 , n72567 );
buf ( n72569 , n62646 );
buf ( n72570 , n64133 );
and ( n72571 , n72569 , n72570 );
nor ( n72572 , n72568 , n72571 );
buf ( n72573 , n72572 );
buf ( n72574 , n72573 );
not ( n72575 , n72574 );
buf ( n72576 , n72575 );
buf ( n72577 , n72576 );
not ( n72578 , n72577 );
or ( n72579 , n72565 , n72578 );
buf ( n72580 , n71921 );
buf ( n72581 , n63010 );
or ( n72582 , n72580 , n72581 );
nand ( n72583 , n72579 , n72582 );
buf ( n72584 , n72583 );
buf ( n72585 , n72584 );
and ( n72586 , n72563 , n72585 );
and ( n72587 , n72558 , n72562 );
or ( n72588 , n72586 , n72587 );
buf ( n72589 , n72588 );
buf ( n72590 , n72589 );
xor ( n72591 , n72549 , n72590 );
xor ( n72592 , n71930 , n71934 );
xor ( n72593 , n72592 , n72021 );
buf ( n72594 , n72593 );
buf ( n72595 , n72594 );
and ( n72596 , n72591 , n72595 );
and ( n72597 , n72549 , n72590 );
or ( n72598 , n72596 , n72597 );
buf ( n72599 , n72598 );
xor ( n72600 , n72332 , n72372 );
xor ( n72601 , n72600 , n72376 );
and ( n72602 , n72599 , n72601 );
xor ( n72603 , n71860 , n71876 );
xor ( n72604 , n72603 , n71893 );
xor ( n72605 , n72348 , n72367 );
xor ( n72606 , n72604 , n72605 );
buf ( n72607 , n68232 );
buf ( n72608 , n58897 );
and ( n72609 , n72607 , n72608 );
buf ( n72610 , n68235 );
buf ( n72611 , n58894 );
and ( n72612 , n72610 , n72611 );
nor ( n72613 , n72609 , n72612 );
buf ( n72614 , n72613 );
buf ( n72615 , n72614 );
buf ( n72616 , n58913 );
or ( n72617 , n72615 , n72616 );
buf ( n72618 , n72390 );
buf ( n72619 , n58890 );
or ( n72620 , n72618 , n72619 );
nand ( n72621 , n72617 , n72620 );
buf ( n72622 , n72621 );
buf ( n72623 , n72622 );
buf ( n72624 , n70348 );
buf ( n72625 , n56777 );
and ( n72626 , n72624 , n72625 );
buf ( n72627 , n70351 );
buf ( n72628 , n56804 );
and ( n72629 , n72627 , n72628 );
nor ( n72630 , n72626 , n72629 );
buf ( n72631 , n72630 );
buf ( n72632 , n72631 );
buf ( n72633 , n56799 );
or ( n72634 , n72632 , n72633 );
buf ( n72635 , n72005 );
buf ( n72636 , n58982 );
or ( n72637 , n72635 , n72636 );
nand ( n72638 , n72634 , n72637 );
buf ( n72639 , n72638 );
buf ( n72640 , n72639 );
xor ( n72641 , n72623 , n72640 );
xor ( n72642 , n72419 , n72422 );
xor ( n72643 , n72642 , n72481 );
buf ( n72644 , n72643 );
buf ( n72645 , n72644 );
and ( n72646 , n72641 , n72645 );
and ( n72647 , n72623 , n72640 );
or ( n72648 , n72646 , n72647 );
buf ( n72649 , n72648 );
xor ( n72650 , n71791 , n71811 );
xor ( n72651 , n72650 , n71848 );
xor ( n72652 , n71989 , n72010 );
xor ( n72653 , n72651 , n72652 );
xor ( n72654 , n72649 , n72653 );
buf ( n72655 , n62679 );
not ( n72656 , n72655 );
buf ( n72657 , n64068 );
buf ( n72658 , n62681 );
and ( n72659 , n72657 , n72658 );
buf ( n72660 , n66579 );
buf ( n72661 , n62663 );
and ( n72662 , n72660 , n72661 );
nor ( n72663 , n72659 , n72662 );
buf ( n72664 , n72663 );
buf ( n72665 , n72664 );
not ( n72666 , n72665 );
buf ( n72667 , n72666 );
buf ( n72668 , n72667 );
not ( n72669 , n72668 );
or ( n72670 , n72656 , n72669 );
buf ( n72671 , n72530 );
buf ( n72672 , n62676 );
or ( n72673 , n72671 , n72672 );
nand ( n72674 , n72670 , n72673 );
buf ( n72675 , n72674 );
and ( n72676 , n72654 , n72675 );
and ( n72677 , n72649 , n72653 );
or ( n72678 , n72676 , n72677 );
buf ( n72679 , n72678 );
buf ( n72680 , n60068 );
buf ( n72681 , n66742 );
and ( n72682 , n72680 , n72681 );
buf ( n72683 , n60071 );
buf ( n72684 , n63000 );
and ( n72685 , n72683 , n72684 );
nor ( n72686 , n72682 , n72685 );
buf ( n72687 , n72686 );
buf ( n72688 , n72687 );
buf ( n72689 , n64230 );
or ( n72690 , n72688 , n72689 );
buf ( n72691 , n72359 );
buf ( n72692 , n64227 );
or ( n72693 , n72691 , n72692 );
nand ( n72694 , n72690 , n72693 );
buf ( n72695 , n72694 );
buf ( n72696 , n72695 );
xor ( n72697 , n72679 , n72696 );
xor ( n72698 , n72558 , n72562 );
xor ( n72699 , n72698 , n72585 );
buf ( n72700 , n72699 );
buf ( n72701 , n72700 );
and ( n72702 , n72697 , n72701 );
and ( n72703 , n72679 , n72696 );
or ( n72704 , n72702 , n72703 );
buf ( n72705 , n72704 );
xor ( n72706 , n72606 , n72705 );
xor ( n72707 , n72549 , n72590 );
xor ( n72708 , n72707 , n72595 );
buf ( n72709 , n72708 );
and ( n72710 , n72706 , n72709 );
and ( n72711 , n72606 , n72705 );
or ( n72712 , n72710 , n72711 );
xor ( n72713 , n72332 , n72372 );
xor ( n72714 , n72713 , n72376 );
and ( n72715 , n72712 , n72714 );
and ( n72716 , n72599 , n72712 );
or ( n72717 , n72602 , n72715 , n72716 );
xor ( n72718 , n72052 , n72055 );
xor ( n72719 , n72718 , n72060 );
and ( n72720 , n72717 , n72719 );
and ( n72721 , n72379 , n72717 );
or ( n72722 , n72382 , n72720 , n72721 );
buf ( n72723 , n72722 );
xor ( n72724 , n71735 , n71912 );
xor ( n72725 , n72724 , n72064 );
buf ( n72726 , n72725 );
buf ( n72727 , n72726 );
xor ( n72728 , n72723 , n72727 );
and ( n72729 , n42844 , n72240 );
not ( n72730 , n42844 );
and ( n72731 , n72730 , n42228 );
or ( n72732 , n72729 , n72731 );
buf ( n72733 , n72732 );
not ( n72734 , n72733 );
buf ( n72735 , n41596 );
not ( n72736 , n72735 );
or ( n72737 , n72734 , n72736 );
buf ( n72738 , n72246 );
buf ( n72739 , n41574 );
nand ( n72740 , n72738 , n72739 );
buf ( n72741 , n72740 );
buf ( n72742 , n72741 );
nand ( n72743 , n72737 , n72742 );
buf ( n72744 , n72743 );
buf ( n72745 , n72744 );
xor ( n72746 , n72728 , n72745 );
buf ( n72747 , n72746 );
buf ( n72748 , n72747 );
xor ( n72749 , n72329 , n72748 );
buf ( n72750 , n44496 );
not ( n72751 , n72750 );
buf ( n72752 , n44524 );
not ( n72753 , n72752 );
buf ( n72754 , n28430 );
not ( n72755 , n72754 );
buf ( n72756 , n72755 );
buf ( n72757 , n72756 );
not ( n72758 , n72757 );
or ( n72759 , n72753 , n72758 );
buf ( n72760 , n66398 );
not ( n72761 , n72760 );
buf ( n72762 , n44527 );
nand ( n72763 , n72761 , n72762 );
buf ( n72764 , n72763 );
buf ( n72765 , n72764 );
nand ( n72766 , n72759 , n72765 );
buf ( n72767 , n72766 );
buf ( n72768 , n72767 );
not ( n72769 , n72768 );
or ( n72770 , n72751 , n72769 );
buf ( n72771 , n44524 );
not ( n72772 , n72771 );
buf ( n72773 , n43055 );
not ( n72774 , n72773 );
or ( n72775 , n72772 , n72774 );
not ( n72776 , n43055 );
buf ( n72777 , n72776 );
buf ( n72778 , n44527 );
nand ( n72779 , n72777 , n72778 );
buf ( n72780 , n72779 );
buf ( n72781 , n72780 );
nand ( n72782 , n72775 , n72781 );
buf ( n72783 , n72782 );
buf ( n72784 , n72783 );
buf ( n72785 , n44517 );
nand ( n72786 , n72784 , n72785 );
buf ( n72787 , n72786 );
buf ( n72788 , n72787 );
nand ( n72789 , n72770 , n72788 );
buf ( n72790 , n72789 );
buf ( n72791 , n72790 );
and ( n72792 , n72749 , n72791 );
and ( n72793 , n72329 , n72748 );
or ( n72794 , n72792 , n72793 );
buf ( n72795 , n72794 );
buf ( n72796 , n72795 );
and ( n72797 , n72301 , n72796 );
nor ( n72798 , n72299 , n72797 );
buf ( n72799 , n72798 );
not ( n72800 , n72799 );
buf ( n72801 , n72800 );
buf ( n72802 , n72801 );
not ( n72803 , n72802 );
buf ( n72804 , n67149 );
not ( n72805 , n72804 );
buf ( n72806 , n72190 );
not ( n72807 , n72806 );
or ( n72808 , n72805 , n72807 );
buf ( n72809 , n45746 );
not ( n72810 , n72809 );
buf ( n72811 , n41733 );
not ( n72812 , n72811 );
or ( n72813 , n72810 , n72812 );
buf ( n72814 , n60327 );
buf ( n72815 , n45747 );
nand ( n72816 , n72814 , n72815 );
buf ( n72817 , n72816 );
buf ( n72818 , n72817 );
nand ( n72819 , n72813 , n72818 );
buf ( n72820 , n72819 );
buf ( n72821 , n72820 );
buf ( n72822 , n71048 );
nand ( n72823 , n72821 , n72822 );
buf ( n72824 , n72823 );
buf ( n72825 , n72824 );
nand ( n72826 , n72808 , n72825 );
buf ( n72827 , n72826 );
buf ( n72828 , n72827 );
not ( n72829 , n72828 );
or ( n72830 , n72803 , n72829 );
buf ( n72831 , n72827 );
buf ( n72832 , n72801 );
or ( n72833 , n72831 , n72832 );
xor ( n72834 , n72116 , n72153 );
xor ( n72835 , n72834 , n72167 );
buf ( n72836 , n72835 );
buf ( n72837 , n72836 );
nand ( n72838 , n72833 , n72837 );
buf ( n72839 , n72838 );
buf ( n72840 , n72839 );
nand ( n72841 , n72830 , n72840 );
buf ( n72842 , n72841 );
buf ( n72843 , n72842 );
buf ( n72844 , n52780 );
buf ( n72845 , n52673 );
and ( n72846 , n72844 , n72845 );
not ( n72847 , n72844 );
buf ( n72848 , n51804 );
and ( n72849 , n72847 , n72848 );
or ( n72850 , n72846 , n72849 );
buf ( n72851 , n72850 );
buf ( n72852 , n72851 );
not ( n72853 , n72852 );
buf ( n72854 , n72853 );
buf ( n72855 , n72854 );
not ( n72856 , n72855 );
buf ( n72857 , n42628 );
not ( n72858 , n72857 );
or ( n72859 , n72856 , n72858 );
buf ( n72860 , n56289 );
not ( n72861 , n72860 );
buf ( n72862 , n51804 );
not ( n72863 , n72862 );
or ( n72864 , n72861 , n72863 );
buf ( n72865 , n25159 );
buf ( n72866 , n52094 );
nand ( n72867 , n72865 , n72866 );
buf ( n72868 , n72867 );
buf ( n72869 , n72868 );
nand ( n72870 , n72864 , n72869 );
buf ( n72871 , n72870 );
buf ( n72872 , n72871 );
buf ( n72873 , n47872 );
nand ( n72874 , n72872 , n72873 );
buf ( n72875 , n72874 );
buf ( n72876 , n72875 );
nand ( n72877 , n72859 , n72876 );
buf ( n72878 , n72877 );
buf ( n72879 , n72878 );
xor ( n72880 , n72843 , n72879 );
buf ( n72881 , n48868 );
not ( n72882 , n72881 );
buf ( n72883 , n48808 );
not ( n72884 , n72883 );
buf ( n72885 , n41879 );
not ( n72886 , n72885 );
or ( n72887 , n72884 , n72886 );
buf ( n72888 , n50583 );
buf ( n72889 , n48808 );
not ( n72890 , n72889 );
buf ( n72891 , n72890 );
buf ( n72892 , n72891 );
nand ( n72893 , n72888 , n72892 );
buf ( n72894 , n72893 );
buf ( n72895 , n72894 );
nand ( n72896 , n72887 , n72895 );
buf ( n72897 , n72896 );
buf ( n72898 , n72897 );
not ( n72899 , n72898 );
or ( n72900 , n72882 , n72899 );
buf ( n72901 , n48808 );
not ( n72902 , n72901 );
buf ( n72903 , n47836 );
not ( n72904 , n72903 );
or ( n72905 , n72902 , n72904 );
buf ( n72906 , n42152 );
buf ( n72907 , n72891 );
nand ( n72908 , n72906 , n72907 );
buf ( n72909 , n72908 );
buf ( n72910 , n72909 );
nand ( n72911 , n72905 , n72910 );
buf ( n72912 , n72911 );
buf ( n72913 , n72912 );
buf ( n72914 , n48855 );
nand ( n72915 , n72913 , n72914 );
buf ( n72916 , n72915 );
buf ( n72917 , n72916 );
nand ( n72918 , n72900 , n72917 );
buf ( n72919 , n72918 );
buf ( n72920 , n72919 );
and ( n72921 , n72880 , n72920 );
and ( n72922 , n72843 , n72879 );
or ( n72923 , n72921 , n72922 );
buf ( n72924 , n72923 );
buf ( n72925 , n72924 );
xor ( n72926 , n72206 , n72925 );
buf ( n72927 , n62125 );
not ( n72928 , n72927 );
buf ( n72929 , n43806 );
not ( n72930 , n72929 );
not ( n72931 , n48836 );
buf ( n72932 , n72931 );
not ( n72933 , n72932 );
and ( n72934 , n72930 , n72933 );
buf ( n72935 , n43806 );
buf ( n72936 , n72931 );
and ( n72937 , n72935 , n72936 );
nor ( n72938 , n72934 , n72937 );
buf ( n72939 , n72938 );
buf ( n72940 , n72939 );
not ( n72941 , n72940 );
buf ( n72942 , n72941 );
buf ( n72943 , n72942 );
not ( n72944 , n72943 );
or ( n72945 , n72928 , n72944 );
and ( n72946 , n48836 , n41951 );
not ( n72947 , n48836 );
and ( n72948 , n72947 , n41823 );
or ( n72949 , n72946 , n72948 );
buf ( n72950 , n72949 );
buf ( n72951 , n51488 );
nand ( n72952 , n72950 , n72951 );
buf ( n72953 , n72952 );
buf ( n72954 , n72953 );
nand ( n72955 , n72945 , n72954 );
buf ( n72956 , n72955 );
buf ( n72957 , n72956 );
xor ( n72958 , n72926 , n72957 );
buf ( n72959 , n72958 );
buf ( n72960 , n72959 );
xor ( n72961 , n71115 , n72172 );
xor ( n72962 , n72961 , n72198 );
buf ( n72963 , n72962 );
buf ( n72964 , n72963 );
buf ( n72965 , n55841 );
not ( n72966 , n72965 );
buf ( n72967 , n47857 );
not ( n72968 , n72967 );
or ( n72969 , n72966 , n72968 );
buf ( n72970 , n50591 );
buf ( n72971 , n58361 );
nand ( n72972 , n72970 , n72971 );
buf ( n72973 , n72972 );
buf ( n72974 , n72973 );
nand ( n72975 , n72969 , n72974 );
buf ( n72976 , n72975 );
buf ( n72977 , n72976 );
not ( n72978 , n72977 );
buf ( n72979 , n52537 );
not ( n72980 , n72979 );
or ( n72981 , n72978 , n72980 );
buf ( n72982 , n53548 );
buf ( n72983 , n55743 );
and ( n72984 , n72982 , n72983 );
not ( n72985 , n72982 );
buf ( n72986 , n50598 );
and ( n72987 , n72985 , n72986 );
nor ( n72988 , n72984 , n72987 );
buf ( n72989 , n72988 );
buf ( n72990 , n72989 );
buf ( n72991 , n48705 );
nand ( n72992 , n72990 , n72991 );
buf ( n72993 , n72992 );
buf ( n72994 , n72993 );
nand ( n72995 , n72981 , n72994 );
buf ( n72996 , n72995 );
buf ( n72997 , n72996 );
xor ( n72998 , n72964 , n72997 );
buf ( n72999 , n41574 );
not ( n73000 , n72999 );
and ( n73001 , n41605 , n70855 );
not ( n73002 , n41605 );
and ( n73003 , n73002 , n29463 );
or ( n73004 , n73001 , n73003 );
buf ( n73005 , n73004 );
not ( n73006 , n73005 );
or ( n73007 , n73000 , n73006 );
buf ( n73008 , n41605 );
not ( n73009 , n73008 );
buf ( n73010 , n72756 );
not ( n73011 , n73010 );
or ( n73012 , n73009 , n73011 );
nand ( n73013 , n28430 , n41604 );
buf ( n73014 , n73013 );
nand ( n73015 , n73012 , n73014 );
buf ( n73016 , n73015 );
buf ( n73017 , n73016 );
buf ( n73018 , n41596 );
nand ( n73019 , n73017 , n73018 );
buf ( n73020 , n73019 );
buf ( n73021 , n73020 );
nand ( n73022 , n73007 , n73021 );
buf ( n73023 , n73022 );
buf ( n73024 , n73023 );
not ( n73025 , n72108 );
not ( n73026 , n71146 );
not ( n73027 , n73026 );
or ( n73028 , n73025 , n73027 );
not ( n73029 , n71145 );
nand ( n73030 , n73029 , n71134 , n72105 );
nand ( n73031 , n73030 , n72070 );
nand ( n73032 , n73028 , n73031 );
buf ( n73033 , n73032 );
xor ( n73034 , n73024 , n73033 );
buf ( n73035 , n66459 );
not ( n73036 , n73035 );
buf ( n73037 , n73036 );
buf ( n73038 , n73037 );
buf ( n73039 , n72164 );
or ( n73040 , n73038 , n73039 );
buf ( n73041 , n46117 );
buf ( n73042 , n63913 );
xnor ( n73043 , n73041 , n73042 );
buf ( n73044 , n73043 );
buf ( n73045 , n73044 );
not ( n73046 , n73045 );
buf ( n73047 , n73046 );
buf ( n73048 , n73047 );
buf ( n73049 , n42333 );
or ( n73050 , n73048 , n73049 );
nand ( n73051 , n73040 , n73050 );
buf ( n73052 , n73051 );
buf ( n73053 , n73052 );
xor ( n73054 , n73034 , n73053 );
buf ( n73055 , n73054 );
buf ( n73056 , n73055 );
buf ( n73057 , n50995 );
not ( n73058 , n73057 );
buf ( n73059 , n57599 );
not ( n73060 , n73059 );
or ( n73061 , n73058 , n73060 );
buf ( n73062 , n42560 );
buf ( n73063 , n50998 );
nand ( n73064 , n73062 , n73063 );
buf ( n73065 , n73064 );
buf ( n73066 , n73065 );
nand ( n73067 , n73061 , n73066 );
buf ( n73068 , n73067 );
buf ( n73069 , n73068 );
not ( n73070 , n73069 );
buf ( n73071 , n43938 );
not ( n73072 , n73071 );
or ( n73073 , n73070 , n73072 );
buf ( n73074 , n50060 );
not ( n73075 , n73074 );
buf ( n73076 , n52725 );
not ( n73077 , n73076 );
or ( n73078 , n73075 , n73077 );
buf ( n73079 , n58185 );
buf ( n73080 , n67438 );
nand ( n73081 , n73079 , n73080 );
buf ( n73082 , n73081 );
buf ( n73083 , n73082 );
nand ( n73084 , n73078 , n73083 );
buf ( n73085 , n73084 );
buf ( n73086 , n73085 );
buf ( n73087 , n43905 );
nand ( n73088 , n73086 , n73087 );
buf ( n73089 , n73088 );
buf ( n73090 , n73089 );
nand ( n73091 , n73073 , n73090 );
buf ( n73092 , n73091 );
buf ( n73093 , n73092 );
xor ( n73094 , n73056 , n73093 );
xor ( n73095 , n72723 , n72727 );
and ( n73096 , n73095 , n72745 );
and ( n73097 , n72723 , n72727 );
or ( n73098 , n73096 , n73097 );
buf ( n73099 , n73098 );
buf ( n73100 , n73099 );
buf ( n73101 , n46390 );
not ( n73102 , n73101 );
buf ( n73103 , n62510 );
not ( n73104 , n73103 );
or ( n73105 , n73102 , n73104 );
buf ( n73106 , n64748 );
buf ( n73107 , n46387 );
nand ( n73108 , n73106 , n73107 );
buf ( n73109 , n73108 );
buf ( n73110 , n73109 );
nand ( n73111 , n73105 , n73110 );
buf ( n73112 , n73111 );
buf ( n73113 , n73112 );
not ( n73114 , n73113 );
buf ( n73115 , n46047 );
not ( n73116 , n73115 );
or ( n73117 , n73114 , n73116 );
and ( n73118 , n46117 , n68606 );
not ( n73119 , n46117 );
and ( n73120 , n73119 , n64748 );
or ( n73121 , n73118 , n73120 );
buf ( n73122 , n73121 );
buf ( n73123 , n42665 );
nand ( n73124 , n73122 , n73123 );
buf ( n73125 , n73124 );
buf ( n73126 , n73125 );
nand ( n73127 , n73117 , n73126 );
buf ( n73128 , n73127 );
buf ( n73129 , n73128 );
xor ( n73130 , n73100 , n73129 );
buf ( n73131 , n44496 );
not ( n73132 , n73131 );
buf ( n73133 , n72145 );
not ( n73134 , n73133 );
or ( n73135 , n73132 , n73134 );
buf ( n73136 , n72767 );
buf ( n73137 , n44517 );
nand ( n73138 , n73136 , n73137 );
buf ( n73139 , n73138 );
buf ( n73140 , n73139 );
nand ( n73141 , n73135 , n73140 );
buf ( n73142 , n73141 );
buf ( n73143 , n73142 );
and ( n73144 , n73130 , n73143 );
and ( n73145 , n73100 , n73129 );
or ( n73146 , n73144 , n73145 );
buf ( n73147 , n73146 );
buf ( n73148 , n73147 );
buf ( n73149 , n41574 );
not ( n73150 , n73149 );
buf ( n73151 , n73016 );
not ( n73152 , n73151 );
or ( n73153 , n73150 , n73152 );
buf ( n73154 , n72223 );
buf ( n73155 , n41596 );
nand ( n73156 , n73154 , n73155 );
buf ( n73157 , n73156 );
buf ( n73158 , n73157 );
nand ( n73159 , n73153 , n73158 );
buf ( n73160 , n73159 );
buf ( n73161 , n73121 );
not ( n73162 , n73161 );
not ( n73163 , n42708 );
buf ( n73164 , n73163 );
not ( n73165 , n73164 );
or ( n73166 , n73162 , n73165 );
buf ( n73167 , n44952 );
not ( n73168 , n73167 );
buf ( n73169 , n62510 );
not ( n73170 , n73169 );
or ( n73171 , n73168 , n73170 );
buf ( n73172 , n25226 );
buf ( n73173 , n44949 );
nand ( n73174 , n73172 , n73173 );
buf ( n73175 , n73174 );
buf ( n73176 , n73175 );
nand ( n73177 , n73171 , n73176 );
buf ( n73178 , n73177 );
buf ( n73179 , n73178 );
buf ( n73180 , n42665 );
nand ( n73181 , n73179 , n73180 );
buf ( n73182 , n73181 );
buf ( n73183 , n73182 );
nand ( n73184 , n73166 , n73183 );
buf ( n73185 , n73184 );
xor ( n73186 , n73160 , n73185 );
xor ( n73187 , n72208 , n72252 );
and ( n73188 , n73187 , n72273 );
and ( n73189 , n72208 , n72252 );
or ( n73190 , n73188 , n73189 );
xor ( n73191 , n73186 , n73190 );
buf ( n73192 , n73191 );
xor ( n73193 , n73148 , n73192 );
buf ( n73194 , n50060 );
not ( n73195 , n73194 );
buf ( n73196 , n41657 );
not ( n73197 , n73196 );
or ( n73198 , n73195 , n73197 );
buf ( n73199 , n61442 );
buf ( n73200 , n67438 );
nand ( n73201 , n73199 , n73200 );
buf ( n73202 , n73201 );
buf ( n73203 , n73202 );
nand ( n73204 , n73198 , n73203 );
buf ( n73205 , n73204 );
buf ( n73206 , n73205 );
not ( n73207 , n73206 );
buf ( n73208 , n59928 );
not ( n73209 , n73208 );
or ( n73210 , n73207 , n73209 );
buf ( n73211 , n71090 );
buf ( n73212 , n62582 );
nand ( n73213 , n73211 , n73212 );
buf ( n73214 , n73213 );
buf ( n73215 , n73214 );
nand ( n73216 , n73210 , n73215 );
buf ( n73217 , n73216 );
buf ( n73218 , n73217 );
and ( n73219 , n73193 , n73218 );
and ( n73220 , n73148 , n73192 );
or ( n73221 , n73219 , n73220 );
buf ( n73222 , n73221 );
buf ( n73223 , n73222 );
xor ( n73224 , n73094 , n73223 );
buf ( n73225 , n73224 );
buf ( n73226 , n73225 );
and ( n73227 , n72998 , n73226 );
and ( n73228 , n72964 , n72997 );
or ( n73229 , n73227 , n73228 );
buf ( n73230 , n73229 );
buf ( n73231 , n73230 );
buf ( n73232 , n72871 );
not ( n73233 , n73232 );
buf ( n73234 , n42628 );
not ( n73235 , n73234 );
or ( n73236 , n73233 , n73235 );
buf ( n73237 , n50995 );
not ( n73238 , n73237 );
buf ( n73239 , n46356 );
not ( n73240 , n73239 );
or ( n73241 , n73238 , n73240 );
buf ( n73242 , n25159 );
buf ( n73243 , n50998 );
nand ( n73244 , n73242 , n73243 );
buf ( n73245 , n73244 );
buf ( n73246 , n73245 );
nand ( n73247 , n73241 , n73246 );
buf ( n73248 , n73247 );
buf ( n73249 , n73248 );
buf ( n73250 , n42564 );
nand ( n73251 , n73249 , n73250 );
buf ( n73252 , n73251 );
buf ( n73253 , n73252 );
nand ( n73254 , n73236 , n73253 );
buf ( n73255 , n73254 );
not ( n73256 , n73255 );
buf ( n73257 , n46912 );
not ( n73258 , n73257 );
buf ( n73259 , n46875 );
not ( n73260 , n73259 );
buf ( n73261 , n28411 );
not ( n73262 , n73261 );
buf ( n73263 , n73262 );
buf ( n73264 , n73263 );
not ( n73265 , n73264 );
or ( n73266 , n73260 , n73265 );
buf ( n73267 , n46660 );
buf ( n73268 , n46887 );
nand ( n73269 , n73267 , n73268 );
buf ( n73270 , n73269 );
buf ( n73271 , n73270 );
nand ( n73272 , n73266 , n73271 );
buf ( n73273 , n73272 );
buf ( n73274 , n73273 );
not ( n73275 , n73274 );
or ( n73276 , n73258 , n73275 );
buf ( n73277 , n46887 );
buf ( n73278 , n47436 );
and ( n73279 , n73277 , n73278 );
not ( n73280 , n73277 );
buf ( n73281 , n50624 );
and ( n73282 , n73280 , n73281 );
or ( n73283 , n73279 , n73282 );
buf ( n73284 , n73283 );
buf ( n73285 , n73284 );
not ( n73286 , n73285 );
buf ( n73287 , n46907 );
nand ( n73288 , n73286 , n73287 );
buf ( n73289 , n73288 );
buf ( n73290 , n73289 );
nand ( n73291 , n73276 , n73290 );
buf ( n73292 , n73291 );
not ( n73293 , n73292 );
xor ( n73294 , n73256 , n73293 );
not ( n73295 , n48975 );
and ( n73296 , n50599 , n52780 );
not ( n73297 , n50599 );
and ( n73298 , n73297 , n52789 );
or ( n73299 , n73296 , n73298 );
not ( n73300 , n73299 );
or ( n73301 , n73295 , n73300 );
nand ( n73302 , n72989 , n50608 );
nand ( n73303 , n73301 , n73302 );
xor ( n73304 , n73294 , n73303 );
buf ( n73305 , n73304 );
xor ( n73306 , n73231 , n73305 );
buf ( n73307 , C0 );
buf ( n73308 , n73307 );
xor ( n73309 , n73306 , n73308 );
buf ( n73310 , n73309 );
buf ( n73311 , n73310 );
xor ( n73312 , n72960 , n73311 );
buf ( n73313 , n46887 );
not ( n73314 , n73313 );
buf ( n73315 , n56548 );
not ( n73316 , n73315 );
or ( n73317 , n73314 , n73316 );
buf ( n73318 , n29754 );
not ( n73319 , n73318 );
buf ( n73320 , n46875 );
nand ( n73321 , n73319 , n73320 );
buf ( n73322 , n73321 );
buf ( n73323 , n73322 );
nand ( n73324 , n73317 , n73323 );
buf ( n73325 , n73324 );
and ( n73326 , n73325 , n46912 );
and ( n73327 , n63906 , n46875 );
not ( n73328 , n63906 );
and ( n73329 , n73328 , n46887 );
or ( n73330 , n73327 , n73329 );
and ( n73331 , n73330 , n46907 );
nor ( n73332 , n73326 , n73331 );
buf ( n73333 , n73332 );
not ( n73334 , n73333 );
buf ( n73335 , n48705 );
buf ( n73336 , n12481 );
nand ( n73337 , n73335 , n73336 );
buf ( n73338 , n73337 );
buf ( n73339 , n73338 );
not ( n73340 , n73339 );
or ( n73341 , n73334 , n73340 );
and ( n73342 , n52780 , n52725 );
not ( n73343 , n52780 );
and ( n73344 , n73343 , n54068 );
or ( n73345 , n73342 , n73344 );
buf ( n73346 , n73345 );
not ( n73347 , n73346 );
buf ( n73348 , n43935 );
not ( n73349 , n73348 );
or ( n73350 , n73347 , n73349 );
and ( n73351 , n56289 , n25181 );
not ( n73352 , n56289 );
and ( n73353 , n73352 , n42560 );
or ( n73354 , n73351 , n73353 );
buf ( n73355 , n73354 );
buf ( n73356 , n43905 );
nand ( n73357 , n73355 , n73356 );
buf ( n73358 , n73357 );
buf ( n73359 , n73358 );
nand ( n73360 , n73350 , n73359 );
buf ( n73361 , n73360 );
buf ( n73362 , n73361 );
nand ( n73363 , n73341 , n73362 );
buf ( n73364 , n73363 );
buf ( n73365 , n73364 );
buf ( n73366 , n73332 );
not ( n73367 , n73366 );
buf ( n73368 , n73338 );
not ( n73369 , n73368 );
buf ( n73370 , n73369 );
buf ( n73371 , n73370 );
nand ( n73372 , n73367 , n73371 );
buf ( n73373 , n73372 );
buf ( n73374 , n73373 );
nand ( n73375 , n73365 , n73374 );
buf ( n73376 , n73375 );
buf ( n73377 , n73376 );
and ( n73378 , n72827 , n72798 );
not ( n73379 , n72827 );
and ( n73380 , n73379 , n72801 );
or ( n73381 , n73378 , n73380 );
xor ( n73382 , n73381 , n72836 );
buf ( n73383 , n73382 );
xor ( n73384 , n73377 , n73383 );
and ( n73385 , n25226 , n48320 );
not ( n73386 , n25226 );
and ( n73387 , n73386 , n71078 );
or ( n73388 , n73385 , n73387 );
buf ( n73389 , n73388 );
not ( n73390 , n73389 );
buf ( n73391 , n70268 );
not ( n73392 , n73391 );
or ( n73393 , n73390 , n73392 );
buf ( n73394 , n47716 );
not ( n73395 , n73394 );
buf ( n73396 , n42324 );
not ( n73397 , n73396 );
or ( n73398 , n73395 , n73397 );
buf ( n73399 , n42325 );
buf ( n73400 , n47725 );
nand ( n73401 , n73399 , n73400 );
buf ( n73402 , n73401 );
buf ( n73403 , n73402 );
nand ( n73404 , n73398 , n73403 );
buf ( n73405 , n73404 );
buf ( n73406 , n73405 );
buf ( n73407 , n42665 );
nand ( n73408 , n73406 , n73407 );
buf ( n73409 , n73408 );
buf ( n73410 , n73409 );
nand ( n73411 , n73393 , n73410 );
buf ( n73412 , n73411 );
buf ( n73413 , n73412 );
xor ( n73414 , n72052 , n72055 );
xor ( n73415 , n73414 , n72060 );
xor ( n73416 , n72379 , n72717 );
xor ( n73417 , n73415 , n73416 );
buf ( n73418 , n73417 );
and ( n73419 , n44946 , n42228 );
not ( n73420 , n44946 );
and ( n73421 , n73420 , n41586 );
nor ( n73422 , n73419 , n73421 );
buf ( n73423 , n73422 );
not ( n73424 , n73423 );
buf ( n73425 , n73424 );
buf ( n73426 , n73425 );
not ( n73427 , n73426 );
buf ( n73428 , n41596 );
not ( n73429 , n73428 );
or ( n73430 , n73427 , n73429 );
buf ( n73431 , n72732 );
buf ( n73432 , n41574 );
nand ( n73433 , n73431 , n73432 );
buf ( n73434 , n73433 );
buf ( n73435 , n73434 );
nand ( n73436 , n73430 , n73435 );
buf ( n73437 , n73436 );
buf ( n73438 , n73437 );
xor ( n73439 , n73418 , n73438 );
buf ( n73440 , n44496 );
not ( n73441 , n73440 );
buf ( n73442 , n72783 );
not ( n73443 , n73442 );
or ( n73444 , n73441 , n73443 );
buf ( n73445 , n44524 );
not ( n73446 , n73445 );
buf ( n73447 , n72235 );
not ( n73448 , n73447 );
or ( n73449 , n73446 , n73448 );
buf ( n73450 , n42856 );
buf ( n73451 , n44527 );
nand ( n73452 , n73450 , n73451 );
buf ( n73453 , n73452 );
buf ( n73454 , n73453 );
nand ( n73455 , n73449 , n73454 );
buf ( n73456 , n73455 );
buf ( n73457 , n73456 );
buf ( n73458 , n44517 );
nand ( n73459 , n73457 , n73458 );
buf ( n73460 , n73459 );
buf ( n73461 , n73460 );
nand ( n73462 , n73444 , n73461 );
buf ( n73463 , n73462 );
buf ( n73464 , n73463 );
xor ( n73465 , n73439 , n73464 );
buf ( n73466 , n73465 );
buf ( n73467 , n73466 );
xor ( n73468 , n73413 , n73467 );
buf ( n73469 , n67149 );
not ( n73470 , n73469 );
and ( n73471 , n45746 , n70855 );
not ( n73472 , n45746 );
and ( n73473 , n73472 , n29463 );
or ( n73474 , n73471 , n73473 );
buf ( n73475 , n73474 );
not ( n73476 , n73475 );
or ( n73477 , n73470 , n73476 );
and ( n73478 , n45746 , n66398 );
not ( n73479 , n45746 );
and ( n73480 , n73479 , n28430 );
or ( n73481 , n73478 , n73480 );
buf ( n73482 , n73481 );
buf ( n73483 , n71048 );
nand ( n73484 , n73482 , n73483 );
buf ( n73485 , n73484 );
buf ( n73486 , n73485 );
nand ( n73487 , n73477 , n73486 );
buf ( n73488 , n73487 );
buf ( n73489 , n73488 );
and ( n73490 , n73468 , n73489 );
and ( n73491 , n73413 , n73467 );
or ( n73492 , n73490 , n73491 );
buf ( n73493 , n73492 );
buf ( n73494 , n73493 );
buf ( n73495 , n56289 );
not ( n73496 , n73495 );
buf ( n73497 , n58107 );
not ( n73498 , n73497 );
or ( n73499 , n73496 , n73498 );
buf ( n73500 , n61434 );
buf ( n73501 , n52094 );
nand ( n73502 , n73500 , n73501 );
buf ( n73503 , n73502 );
buf ( n73504 , n73503 );
nand ( n73505 , n73499 , n73504 );
buf ( n73506 , n73505 );
buf ( n73507 , n73506 );
not ( n73508 , n73507 );
buf ( n73509 , n62588 );
not ( n73510 , n73509 );
or ( n73511 , n73508 , n73510 );
buf ( n73512 , n50995 );
not ( n73513 , n73512 );
buf ( n73514 , n58107 );
not ( n73515 , n73514 );
or ( n73516 , n73513 , n73515 );
buf ( n73517 , n61434 );
buf ( n73518 , n50998 );
nand ( n73519 , n73517 , n73518 );
buf ( n73520 , n73519 );
buf ( n73521 , n73520 );
nand ( n73522 , n73516 , n73521 );
buf ( n73523 , n73522 );
buf ( n73524 , n73523 );
buf ( n73525 , n62582 );
nand ( n73526 , n73524 , n73525 );
buf ( n73527 , n73526 );
buf ( n73528 , n73527 );
nand ( n73529 , n73511 , n73528 );
buf ( n73530 , n73529 );
buf ( n73531 , n73530 );
xor ( n73532 , n73494 , n73531 );
xor ( n73533 , n73418 , n73438 );
and ( n73534 , n73533 , n73464 );
and ( n73535 , n73418 , n73438 );
or ( n73536 , n73534 , n73535 );
buf ( n73537 , n73536 );
buf ( n73538 , n73537 );
buf ( n73539 , n73405 );
not ( n73540 , n73539 );
buf ( n73541 , n73163 );
not ( n73542 , n73541 );
or ( n73543 , n73540 , n73542 );
buf ( n73544 , n73112 );
buf ( n73545 , n42665 );
nand ( n73546 , n73544 , n73545 );
buf ( n73547 , n73546 );
buf ( n73548 , n73547 );
nand ( n73549 , n73543 , n73548 );
buf ( n73550 , n73549 );
buf ( n73551 , n73550 );
xor ( n73552 , n73538 , n73551 );
xor ( n73553 , n72329 , n72748 );
xor ( n73554 , n73553 , n72791 );
buf ( n73555 , n73554 );
buf ( n73556 , n73555 );
xor ( n73557 , n73552 , n73556 );
buf ( n73558 , n73557 );
buf ( n73559 , n73558 );
and ( n73560 , n73532 , n73559 );
and ( n73561 , n73494 , n73531 );
or ( n73562 , n73560 , n73561 );
buf ( n73563 , n73562 );
buf ( n73564 , n73563 );
buf ( n73565 , n48865 );
not ( n73566 , n73565 );
buf ( n73567 , n48808 );
not ( n73568 , n73567 );
buf ( n73569 , n47436 );
not ( n73570 , n73569 );
or ( n73571 , n73568 , n73570 );
buf ( n73572 , n50624 );
buf ( n73573 , n72891 );
nand ( n73574 , n73572 , n73573 );
buf ( n73575 , n73574 );
buf ( n73576 , n73575 );
nand ( n73577 , n73571 , n73576 );
buf ( n73578 , n73577 );
buf ( n73579 , n73578 );
not ( n73580 , n73579 );
or ( n73581 , n73566 , n73580 );
buf ( n73582 , n48808 );
not ( n73583 , n73582 );
buf ( n73584 , n42072 );
not ( n73585 , n73584 );
or ( n73586 , n73583 , n73585 );
buf ( n73587 , n56342 );
not ( n73588 , n73587 );
buf ( n73589 , n72891 );
nand ( n73590 , n73588 , n73589 );
buf ( n73591 , n73590 );
buf ( n73592 , n73591 );
nand ( n73593 , n73586 , n73592 );
buf ( n73594 , n73593 );
buf ( n73595 , n73594 );
buf ( n73596 , n48852 );
nand ( n73597 , n73595 , n73596 );
buf ( n73598 , n73597 );
buf ( n73599 , n73598 );
nand ( n73600 , n73581 , n73599 );
buf ( n73601 , n73600 );
buf ( n73602 , n73601 );
xor ( n73603 , n73564 , n73602 );
xor ( n73604 , n73100 , n73129 );
xor ( n73605 , n73604 , n73143 );
buf ( n73606 , n73605 );
buf ( n73607 , n73606 );
buf ( n73608 , n73523 );
not ( n73609 , n73608 );
buf ( n73610 , n61454 );
not ( n73611 , n73610 );
or ( n73612 , n73609 , n73611 );
buf ( n73613 , n73205 );
buf ( n73614 , n48671 );
nand ( n73615 , n73613 , n73614 );
buf ( n73616 , n73615 );
buf ( n73617 , n73616 );
nand ( n73618 , n73612 , n73617 );
buf ( n73619 , n73618 );
buf ( n73620 , n73619 );
xor ( n73621 , n73607 , n73620 );
buf ( n73622 , n67149 );
not ( n73623 , n73622 );
buf ( n73624 , n72820 );
not ( n73625 , n73624 );
or ( n73626 , n73623 , n73625 );
buf ( n73627 , n66426 );
not ( n73628 , n73627 );
buf ( n73629 , n45747 );
nand ( n73630 , n73628 , n73629 );
buf ( n73631 , n73630 );
not ( n73632 , n73631 );
nand ( n73633 , n66426 , n45746 );
not ( n73634 , n73633 );
or ( n73635 , n73632 , n73634 );
nand ( n73636 , n73635 , n71048 );
buf ( n73637 , n73636 );
nand ( n73638 , n73626 , n73637 );
buf ( n73639 , n73638 );
buf ( n73640 , n73639 );
xor ( n73641 , n73621 , n73640 );
buf ( n73642 , n73641 );
buf ( n73643 , n73642 );
and ( n73644 , n73603 , n73643 );
and ( n73645 , n73564 , n73602 );
or ( n73646 , n73644 , n73645 );
buf ( n73647 , n73646 );
buf ( n73648 , n73647 );
and ( n73649 , n73384 , n73648 );
and ( n73650 , n73377 , n73383 );
or ( n73651 , n73649 , n73650 );
buf ( n73652 , n73651 );
buf ( n73653 , n73652 );
not ( n73654 , n73653 );
buf ( n73655 , n46912 );
not ( n73656 , n73655 );
not ( n73657 , n46875 );
not ( n73658 , n42072 );
or ( n73659 , n73657 , n73658 );
buf ( n73660 , n28368 );
buf ( n73661 , n46887 );
nand ( n73662 , n73660 , n73661 );
buf ( n73663 , n73662 );
nand ( n73664 , n73659 , n73663 );
buf ( n73665 , n73664 );
not ( n73666 , n73665 );
or ( n73667 , n73656 , n73666 );
buf ( n73668 , n73325 );
buf ( n73669 , n46907 );
nand ( n73670 , n73668 , n73669 );
buf ( n73671 , n73670 );
buf ( n73672 , n73671 );
nand ( n73673 , n73667 , n73672 );
buf ( n73674 , n73673 );
buf ( n73675 , n73674 );
not ( n73676 , n73675 );
buf ( n73677 , n39994 );
not ( n73678 , n73677 );
buf ( n73679 , n51804 );
not ( n73680 , n73679 );
or ( n73681 , n73678 , n73680 );
buf ( n73682 , n12481 );
nand ( n73683 , n73681 , n73682 );
buf ( n73684 , n73683 );
buf ( n73685 , n73684 );
buf ( n73686 , n24092 );
buf ( n73687 , n25159 );
buf ( n73688 , n25098 );
nand ( n73689 , n73687 , n73688 );
buf ( n73690 , n73689 );
buf ( n73691 , n73690 );
nand ( n73692 , n73685 , n73686 , n73691 );
buf ( n73693 , n73692 );
buf ( n73694 , n73693 );
nand ( n73695 , n73676 , n73694 );
buf ( n73696 , n73695 );
not ( n73697 , n73696 );
buf ( n73698 , n73354 );
not ( n73699 , n73698 );
buf ( n73700 , n43938 );
not ( n73701 , n73700 );
or ( n73702 , n73699 , n73701 );
buf ( n73703 , n73068 );
buf ( n73704 , n43905 );
nand ( n73705 , n73703 , n73704 );
buf ( n73706 , n73705 );
buf ( n73707 , n73706 );
nand ( n73708 , n73702 , n73707 );
buf ( n73709 , n73708 );
not ( n73710 , n73709 );
or ( n73711 , n73697 , n73710 );
buf ( n73712 , n73693 );
not ( n73713 , n73712 );
buf ( n73714 , n73674 );
nand ( n73715 , n73713 , n73714 );
buf ( n73716 , n73715 );
nand ( n73717 , n73711 , n73716 );
buf ( n73718 , n73717 );
xor ( n73719 , n70721 , n70724 );
xor ( n73720 , n73719 , n70728 );
xor ( n73721 , n70429 , n70443 );
xor ( n73722 , n73721 , n70576 );
and ( n73723 , n72082 , n73722 );
xor ( n73724 , n70429 , n70443 );
xor ( n73725 , n73724 , n70576 );
and ( n73726 , n72085 , n73725 );
and ( n73727 , n72082 , n72085 );
or ( n73728 , n73723 , n73726 , n73727 );
not ( n73729 , n72075 );
not ( n73730 , n72093 );
or ( n73731 , n73729 , n73730 );
nand ( n73732 , n73731 , n72096 );
xor ( n73733 , n73728 , n73732 );
xor ( n73734 , n73720 , n73733 );
buf ( n73735 , n73734 );
buf ( n73736 , n71130 );
not ( n73737 , n73736 );
buf ( n73738 , n42246 );
not ( n73739 , n73738 );
or ( n73740 , n73737 , n73739 );
buf ( n73741 , n25290 );
buf ( n73742 , n72776 );
and ( n73743 , n73741 , n73742 );
not ( n73744 , n73741 );
buf ( n73745 , n43055 );
and ( n73746 , n73744 , n73745 );
nor ( n73747 , n73743 , n73746 );
buf ( n73748 , n73747 );
buf ( n73749 , n73748 );
buf ( n73750 , n42309 );
nand ( n73751 , n73749 , n73750 );
buf ( n73752 , n73751 );
buf ( n73753 , n73752 );
nand ( n73754 , n73740 , n73753 );
buf ( n73755 , n73754 );
buf ( n73756 , n73755 );
xor ( n73757 , n73735 , n73756 );
buf ( n73758 , n73178 );
not ( n73759 , n73758 );
buf ( n73760 , n70268 );
not ( n73761 , n73760 );
or ( n73762 , n73759 , n73761 );
buf ( n73763 , n42847 );
not ( n73764 , n73763 );
buf ( n73765 , n68606 );
not ( n73766 , n73765 );
or ( n73767 , n73764 , n73766 );
buf ( n73768 , n25226 );
buf ( n73769 , n46691 );
nand ( n73770 , n73768 , n73769 );
buf ( n73771 , n73770 );
buf ( n73772 , n73771 );
nand ( n73773 , n73767 , n73772 );
buf ( n73774 , n73773 );
buf ( n73775 , n73774 );
buf ( n73776 , n42665 );
nand ( n73777 , n73775 , n73776 );
buf ( n73778 , n73777 );
buf ( n73779 , n73778 );
nand ( n73780 , n73762 , n73779 );
buf ( n73781 , n73780 );
buf ( n73782 , n73781 );
xor ( n73783 , n73757 , n73782 );
buf ( n73784 , n73783 );
buf ( n73785 , n73784 );
not ( n73786 , n73185 );
not ( n73787 , n73160 );
nand ( n73788 , n73786 , n73787 );
not ( n73789 , n73788 );
not ( n73790 , n73190 );
or ( n73791 , n73789 , n73790 );
not ( n73792 , n73787 );
nand ( n73793 , n73792 , n73185 );
nand ( n73794 , n73791 , n73793 );
buf ( n73795 , n73794 );
xor ( n73796 , n73785 , n73795 );
buf ( n73797 , n44496 );
not ( n73798 , n73797 );
buf ( n73799 , n65010 );
not ( n73800 , n73799 );
buf ( n73801 , n60330 );
not ( n73802 , n73801 );
or ( n73803 , n73800 , n73802 );
buf ( n73804 , n41736 );
buf ( n73805 , n44530 );
nand ( n73806 , n73804 , n73805 );
buf ( n73807 , n73806 );
buf ( n73808 , n73807 );
nand ( n73809 , n73803 , n73808 );
buf ( n73810 , n73809 );
buf ( n73811 , n73810 );
not ( n73812 , n73811 );
or ( n73813 , n73798 , n73812 );
buf ( n73814 , n72130 );
buf ( n73815 , n44517 );
nand ( n73816 , n73814 , n73815 );
buf ( n73817 , n73816 );
buf ( n73818 , n73817 );
nand ( n73819 , n73813 , n73818 );
buf ( n73820 , n73819 );
buf ( n73821 , n73820 );
xor ( n73822 , n73796 , n73821 );
buf ( n73823 , n73822 );
buf ( n73824 , n73823 );
buf ( n73825 , n38973 );
buf ( n73826 , n56325 );
nor ( n73827 , n73825 , n73826 );
buf ( n73828 , n73827 );
buf ( n73829 , n73828 );
xor ( n73830 , n73824 , n73829 );
buf ( n73831 , n46907 );
not ( n73832 , n73831 );
buf ( n73833 , n73664 );
not ( n73834 , n73833 );
or ( n73835 , n73832 , n73834 );
buf ( n73836 , n73284 );
buf ( n73837 , n46915 );
or ( n73838 , n73836 , n73837 );
nand ( n73839 , n73835 , n73838 );
buf ( n73840 , n73839 );
buf ( n73841 , n73840 );
xor ( n73842 , n73830 , n73841 );
buf ( n73843 , n73842 );
buf ( n73844 , n73843 );
xor ( n73845 , n73718 , n73844 );
buf ( n73846 , n51488 );
not ( n73847 , n73846 );
buf ( n73848 , n48836 );
buf ( n73849 , n44179 );
and ( n73850 , n73848 , n73849 );
not ( n73851 , n73848 );
buf ( n73852 , n41915 );
and ( n73853 , n73851 , n73852 );
nor ( n73854 , n73850 , n73853 );
buf ( n73855 , n73854 );
buf ( n73856 , n73855 );
not ( n73857 , n73856 );
or ( n73858 , n73847 , n73857 );
buf ( n73859 , n72949 );
buf ( n73860 , n62125 );
nand ( n73861 , n73859 , n73860 );
buf ( n73862 , n73861 );
buf ( n73863 , n73862 );
nand ( n73864 , n73858 , n73863 );
buf ( n73865 , n73864 );
buf ( n73866 , n73865 );
xor ( n73867 , n73845 , n73866 );
buf ( n73868 , n73867 );
buf ( n73869 , n73868 );
not ( n73870 , n73869 );
or ( n73871 , n73654 , n73870 );
buf ( n73872 , n73652 );
buf ( n73873 , n73868 );
or ( n73874 , n73872 , n73873 );
nand ( n73875 , n73696 , n73716 );
xor ( n73876 , n73875 , n73709 );
buf ( n73877 , n73876 );
not ( n73878 , n73877 );
buf ( n73879 , n62125 );
not ( n73880 , n73879 );
buf ( n73881 , n73855 );
not ( n73882 , n73881 );
or ( n73883 , n73880 , n73882 );
buf ( n73884 , n72931 );
buf ( n73885 , n50578 );
and ( n73886 , n73884 , n73885 );
not ( n73887 , n73884 );
buf ( n73888 , n41876 );
and ( n73889 , n73887 , n73888 );
nor ( n73890 , n73886 , n73889 );
buf ( n73891 , n73890 );
buf ( n73892 , n73891 );
buf ( n73893 , n51488 );
nand ( n73894 , n73892 , n73893 );
buf ( n73895 , n73894 );
buf ( n73896 , n73895 );
nand ( n73897 , n73883 , n73896 );
buf ( n73898 , n73897 );
buf ( n73899 , n73898 );
not ( n73900 , n73899 );
buf ( n73901 , n73900 );
buf ( n73902 , n73901 );
not ( n73903 , n73902 );
or ( n73904 , n73878 , n73903 );
xor ( n73905 , n73607 , n73620 );
and ( n73906 , n73905 , n73640 );
and ( n73907 , n73607 , n73620 );
or ( n73908 , n73906 , n73907 );
buf ( n73909 , n73908 );
buf ( n73910 , n73909 );
xor ( n73911 , n73148 , n73192 );
xor ( n73912 , n73911 , n73218 );
buf ( n73913 , n73912 );
buf ( n73914 , n73913 );
xor ( n73915 , n73910 , n73914 );
xor ( n73916 , n73538 , n73551 );
and ( n73917 , n73916 , n73556 );
and ( n73918 , n73538 , n73551 );
or ( n73919 , n73917 , n73918 );
buf ( n73920 , n73919 );
and ( n73921 , n72275 , n72795 );
not ( n73922 , n72275 );
not ( n73923 , n72795 );
and ( n73924 , n73922 , n73923 );
nor ( n73925 , n73921 , n73924 );
and ( n73926 , n73925 , n72297 );
not ( n73927 , n73925 );
and ( n73928 , n73927 , n72296 );
nor ( n73929 , n73926 , n73928 );
xor ( n73930 , n73920 , n73929 );
buf ( n73931 , n46390 );
not ( n73932 , n73931 );
buf ( n73933 , n25293 );
not ( n73934 , n73933 );
or ( n73935 , n73932 , n73934 );
buf ( n73936 , n25290 );
buf ( n73937 , n46387 );
nand ( n73938 , n73936 , n73937 );
buf ( n73939 , n73938 );
buf ( n73940 , n73939 );
nand ( n73941 , n73935 , n73940 );
buf ( n73942 , n73941 );
not ( n73943 , n73942 );
not ( n73944 , n42246 );
or ( n73945 , n73943 , n73944 );
buf ( n73946 , n72316 );
buf ( n73947 , n42309 );
nand ( n73948 , n73946 , n73947 );
buf ( n73949 , n73948 );
nand ( n73950 , n73945 , n73949 );
not ( n73951 , n73950 );
xor ( n73952 , n72332 , n72372 );
xor ( n73953 , n73952 , n72376 );
xor ( n73954 , n72599 , n72712 );
xor ( n73955 , n73953 , n73954 );
buf ( n73956 , n73955 );
xor ( n73957 , n72522 , n72539 );
xor ( n73958 , n73957 , n72544 );
buf ( n73959 , n73958 );
buf ( n73960 , n73959 );
buf ( n73961 , n62782 );
buf ( n73962 , n64129 );
and ( n73963 , n73961 , n73962 );
buf ( n73964 , n62980 );
buf ( n73965 , n64133 );
and ( n73966 , n73964 , n73965 );
nor ( n73967 , n73963 , n73966 );
buf ( n73968 , n73967 );
buf ( n73969 , n73968 );
buf ( n73970 , n64141 );
or ( n73971 , n73969 , n73970 );
buf ( n73972 , n72573 );
buf ( n73973 , n63010 );
or ( n73974 , n73972 , n73973 );
nand ( n73975 , n73971 , n73974 );
buf ( n73976 , n73975 );
buf ( n73977 , n73976 );
xor ( n73978 , n72399 , n72486 );
xor ( n73979 , n73978 , n72517 );
buf ( n73980 , n73979 );
buf ( n73981 , n73980 );
xor ( n73982 , n73977 , n73981 );
buf ( n73983 , n1664 );
not ( n73984 , n73983 );
buf ( n73985 , n72687 );
not ( n73986 , n73985 );
buf ( n73987 , n73986 );
buf ( n73988 , n73987 );
not ( n73989 , n73988 );
or ( n73990 , n73984 , n73989 );
buf ( n73991 , n60229 );
buf ( n73992 , n66742 );
and ( n73993 , n73991 , n73992 );
buf ( n73994 , n62652 );
buf ( n73995 , n63000 );
and ( n73996 , n73994 , n73995 );
nor ( n73997 , n73993 , n73996 );
buf ( n73998 , n73997 );
buf ( n73999 , n73998 );
buf ( n74000 , n64230 );
or ( n74001 , n73999 , n74000 );
nand ( n74002 , n73990 , n74001 );
buf ( n74003 , n74002 );
buf ( n74004 , n74003 );
and ( n74005 , n73982 , n74004 );
and ( n74006 , n73977 , n73981 );
or ( n74007 , n74005 , n74006 );
buf ( n74008 , n74007 );
buf ( n74009 , n74008 );
xor ( n74010 , n73960 , n74009 );
buf ( n74011 , n66690 );
buf ( n74012 , n60261 );
and ( n74013 , n74011 , n74012 );
buf ( n74014 , n66693 );
buf ( n74015 , n60090 );
and ( n74016 , n74014 , n74015 );
nor ( n74017 , n74013 , n74016 );
buf ( n74018 , n74017 );
buf ( n74019 , n74018 );
buf ( n74020 , n60270 );
or ( n74021 , n74019 , n74020 );
buf ( n74022 , n72511 );
buf ( n74023 , n60100 );
or ( n74024 , n74022 , n74023 );
nand ( n74025 , n74021 , n74024 );
buf ( n74026 , n74025 );
buf ( n74027 , n74026 );
buf ( n74028 , n70527 );
buf ( n74029 , n56777 );
and ( n74030 , n74028 , n74029 );
buf ( n74031 , n70530 );
buf ( n74032 , n56804 );
and ( n74033 , n74031 , n74032 );
nor ( n74034 , n74030 , n74033 );
buf ( n74035 , n74034 );
buf ( n74036 , n74035 );
buf ( n74037 , n56799 );
or ( n74038 , n74036 , n74037 );
buf ( n74039 , n72631 );
buf ( n74040 , n58982 );
or ( n74041 , n74039 , n74040 );
nand ( n74042 , n74038 , n74041 );
buf ( n74043 , n74042 );
buf ( n74044 , n74043 );
buf ( n74045 , n56664 );
buf ( n74046 , n55195 );
buf ( n74047 , n71818 );
and ( n74048 , n74046 , n74047 );
buf ( n74049 , n55184 );
buf ( n74050 , n71821 );
and ( n74051 , n74049 , n74050 );
nor ( n74052 , n74048 , n74051 );
buf ( n74053 , n74052 );
buf ( n74054 , n74053 );
or ( n74055 , n74045 , n74054 );
buf ( n74056 , n72435 );
buf ( n74057 , n56673 );
or ( n74058 , n74056 , n74057 );
nand ( n74059 , n74055 , n74058 );
buf ( n74060 , n74059 );
buf ( n74061 , n74060 );
buf ( n74062 , n16469 );
buf ( n74063 , n71307 );
and ( n74064 , n74062 , n74063 );
buf ( n74065 , n56631 );
buf ( n74066 , n71310 );
and ( n74067 , n74065 , n74066 );
nor ( n74068 , n74064 , n74067 );
buf ( n74069 , n74068 );
buf ( n74070 , n74069 );
not ( n74071 , n74070 );
buf ( n74072 , n74071 );
buf ( n74073 , n74072 );
not ( n74074 , n74073 );
buf ( n74075 , n56629 );
not ( n74076 , n74075 );
or ( n74077 , n74074 , n74076 );
buf ( n74078 , n72471 );
buf ( n74079 , n56639 );
or ( n74080 , n74078 , n74079 );
nand ( n74081 , n74077 , n74080 );
buf ( n74082 , n74081 );
buf ( n74083 , n74082 );
and ( n74084 , n74061 , n74083 );
buf ( n74085 , n74084 );
buf ( n74086 , n74085 );
xor ( n74087 , n74044 , n74086 );
xor ( n74088 , n72443 , n72456 );
xor ( n74089 , n74088 , n72476 );
buf ( n74090 , n74089 );
buf ( n74091 , n74090 );
and ( n74092 , n74087 , n74091 );
and ( n74093 , n74044 , n74086 );
or ( n74094 , n74092 , n74093 );
buf ( n74095 , n74094 );
buf ( n74096 , n74095 );
xor ( n74097 , n74027 , n74096 );
buf ( n74098 , n71232 );
buf ( n74099 , n56777 );
and ( n74100 , n74098 , n74099 );
buf ( n74101 , n71235 );
buf ( n74102 , n56804 );
and ( n74103 , n74101 , n74102 );
nor ( n74104 , n74100 , n74103 );
buf ( n74105 , n74104 );
buf ( n74106 , n74105 );
buf ( n74107 , n56799 );
or ( n74108 , n74106 , n74107 );
buf ( n74109 , n74035 );
buf ( n74110 , n58982 );
or ( n74111 , n74109 , n74110 );
nand ( n74112 , n74108 , n74111 );
buf ( n74113 , n74112 );
buf ( n74114 , n55129 );
and ( n74115 , n54989 , n622 );
buf ( n74116 , n74115 );
not ( n74117 , n74116 );
buf ( n74118 , n74117 );
buf ( n74119 , n74118 );
or ( n74120 , n74114 , n74119 );
buf ( n74121 , n56598 );
buf ( n74122 , n72448 );
or ( n74123 , n74121 , n74122 );
nand ( n74124 , n74120 , n74123 );
buf ( n74125 , n74124 );
xor ( n74126 , n74113 , n74125 );
xor ( n74127 , n74061 , n74083 );
buf ( n74128 , n74127 );
and ( n74129 , n74126 , n74128 );
and ( n74130 , n74113 , n74125 );
or ( n74131 , n74129 , n74130 );
buf ( n74132 , n70333 );
buf ( n74133 , n58897 );
and ( n74134 , n74132 , n74133 );
buf ( n74135 , n70336 );
buf ( n74136 , n58894 );
and ( n74137 , n74135 , n74136 );
nor ( n74138 , n74134 , n74137 );
buf ( n74139 , n74138 );
buf ( n74140 , n74139 );
buf ( n74141 , n58913 );
or ( n74142 , n74140 , n74141 );
buf ( n74143 , n72614 );
buf ( n74144 , n58890 );
or ( n74145 , n74143 , n74144 );
nand ( n74146 , n74142 , n74145 );
buf ( n74147 , n74146 );
xor ( n74148 , n74131 , n74147 );
buf ( n74149 , n60101 );
not ( n74150 , n74149 );
buf ( n74151 , n68220 );
buf ( n74152 , n58880 );
or ( n74153 , n74151 , n74152 );
buf ( n74154 , n68217 );
buf ( n74155 , n15265 );
or ( n74156 , n74154 , n74155 );
nand ( n74157 , n74153 , n74156 );
buf ( n74158 , n74157 );
buf ( n74159 , n74158 );
not ( n74160 , n74159 );
or ( n74161 , n74150 , n74160 );
buf ( n74162 , n74018 );
buf ( n74163 , n60100 );
or ( n74164 , n74162 , n74163 );
nand ( n74165 , n74161 , n74164 );
buf ( n74166 , n74165 );
and ( n74167 , n74148 , n74166 );
and ( n74168 , n74131 , n74147 );
or ( n74169 , n74167 , n74168 );
buf ( n74170 , n74169 );
and ( n74171 , n74097 , n74170 );
and ( n74172 , n74027 , n74096 );
or ( n74173 , n74171 , n74172 );
buf ( n74174 , n74173 );
xor ( n74175 , n72649 , n72653 );
xor ( n74176 , n74175 , n72675 );
and ( n74177 , n74174 , n74176 );
xor ( n74178 , n72623 , n72640 );
xor ( n74179 , n74178 , n72645 );
buf ( n74180 , n74179 );
buf ( n74181 , n74180 );
buf ( n74182 , n64211 );
buf ( n74183 , n62681 );
and ( n74184 , n74182 , n74183 );
buf ( n74185 , n66610 );
buf ( n74186 , n62663 );
and ( n74187 , n74185 , n74186 );
nor ( n74188 , n74184 , n74187 );
buf ( n74189 , n74188 );
buf ( n74190 , n74189 );
buf ( n74191 , n62935 );
or ( n74192 , n74190 , n74191 );
buf ( n74193 , n72664 );
buf ( n74194 , n62676 );
or ( n74195 , n74193 , n74194 );
nand ( n74196 , n74192 , n74195 );
buf ( n74197 , n74196 );
buf ( n74198 , n74197 );
xor ( n74199 , n74181 , n74198 );
buf ( n74200 , n1664 );
not ( n74201 , n74200 );
buf ( n74202 , n73998 );
not ( n74203 , n74202 );
buf ( n74204 , n74203 );
buf ( n74205 , n74204 );
not ( n74206 , n74205 );
or ( n74207 , n74201 , n74206 );
buf ( n74208 , n62643 );
buf ( n74209 , n66742 );
and ( n74210 , n74208 , n74209 );
buf ( n74211 , n62646 );
buf ( n74212 , n63000 );
and ( n74213 , n74211 , n74212 );
nor ( n74214 , n74210 , n74213 );
buf ( n74215 , n74214 );
buf ( n74216 , n74215 );
buf ( n74217 , n64230 );
or ( n74218 , n74216 , n74217 );
nand ( n74219 , n74207 , n74218 );
buf ( n74220 , n74219 );
buf ( n74221 , n74220 );
and ( n74222 , n74199 , n74221 );
and ( n74223 , n74181 , n74198 );
or ( n74224 , n74222 , n74223 );
buf ( n74225 , n74224 );
xor ( n74226 , n72649 , n72653 );
xor ( n74227 , n74226 , n72675 );
and ( n74228 , n74225 , n74227 );
and ( n74229 , n74174 , n74225 );
or ( n74230 , n74177 , n74228 , n74229 );
buf ( n74231 , n74230 );
and ( n74232 , n74010 , n74231 );
and ( n74233 , n73960 , n74009 );
or ( n74234 , n74232 , n74233 );
buf ( n74235 , n74234 );
xor ( n74236 , n72606 , n72705 );
xor ( n74237 , n74236 , n72709 );
and ( n74238 , n74235 , n74237 );
xor ( n74239 , n73977 , n73981 );
xor ( n74240 , n74239 , n74004 );
buf ( n74241 , n74240 );
buf ( n74242 , n62971 );
buf ( n74243 , n64129 );
and ( n74244 , n74242 , n74243 );
buf ( n74245 , n62974 );
buf ( n74246 , n64133 );
and ( n74247 , n74245 , n74246 );
nor ( n74248 , n74244 , n74247 );
buf ( n74249 , n74248 );
buf ( n74250 , n74249 );
buf ( n74251 , n64141 );
or ( n74252 , n74250 , n74251 );
buf ( n74253 , n73968 );
buf ( n74254 , n63010 );
or ( n74255 , n74253 , n74254 );
nand ( n74256 , n74252 , n74255 );
buf ( n74257 , n74256 );
buf ( n74258 , n74257 );
buf ( n74259 , n66601 );
buf ( n74260 , n62681 );
and ( n74261 , n74259 , n74260 );
buf ( n74262 , n66604 );
buf ( n74263 , n62663 );
and ( n74264 , n74262 , n74263 );
nor ( n74265 , n74261 , n74264 );
buf ( n74266 , n74265 );
buf ( n74267 , n74266 );
buf ( n74268 , n62935 );
or ( n74269 , n74267 , n74268 );
buf ( n74270 , n74189 );
buf ( n74271 , n62676 );
or ( n74272 , n74270 , n74271 );
nand ( n74273 , n74269 , n74272 );
buf ( n74274 , n74273 );
buf ( n74275 , n74274 );
xor ( n74276 , n74044 , n74086 );
xor ( n74277 , n74276 , n74091 );
buf ( n74278 , n74277 );
buf ( n74279 , n74278 );
xor ( n74280 , n74275 , n74279 );
buf ( n74281 , n70348 );
buf ( n74282 , n58897 );
and ( n74283 , n74281 , n74282 );
buf ( n74284 , n70351 );
buf ( n74285 , n58894 );
and ( n74286 , n74284 , n74285 );
nor ( n74287 , n74283 , n74286 );
buf ( n74288 , n74287 );
buf ( n74289 , n74288 );
buf ( n74290 , n58913 );
or ( n74291 , n74289 , n74290 );
buf ( n74292 , n74139 );
buf ( n74293 , n58890 );
or ( n74294 , n74292 , n74293 );
nand ( n74295 , n74291 , n74294 );
buf ( n74296 , n74295 );
buf ( n74297 , n74296 );
buf ( n74298 , n56664 );
buf ( n74299 , n55195 );
buf ( n74300 , n72445 );
and ( n74301 , n74299 , n74300 );
buf ( n74302 , n55184 );
buf ( n74303 , n72448 );
and ( n74304 , n74302 , n74303 );
nor ( n74305 , n74301 , n74304 );
buf ( n74306 , n74305 );
buf ( n74307 , n74306 );
or ( n74308 , n74298 , n74307 );
buf ( n74309 , n74053 );
buf ( n74310 , n55166 );
or ( n74311 , n74309 , n74310 );
nand ( n74312 , n74308 , n74311 );
buf ( n74313 , n74312 );
buf ( n74314 , n74313 );
buf ( n74315 , n55125 );
buf ( n74316 , n74118 );
nor ( n74317 , n74315 , n74316 );
buf ( n74318 , n74317 );
buf ( n74319 , n74318 );
xor ( n74320 , n74314 , n74319 );
buf ( n74321 , n56626 );
buf ( n74322 , n56641 );
buf ( n74323 , n71801 );
and ( n74324 , n74322 , n74323 );
buf ( n74325 , n16472 );
buf ( n74326 , n71804 );
and ( n74327 , n74325 , n74326 );
nor ( n74328 , n74324 , n74327 );
buf ( n74329 , n74328 );
buf ( n74330 , n74329 );
or ( n74331 , n74321 , n74330 );
buf ( n74332 , n74069 );
buf ( n74333 , n56639 );
or ( n74334 , n74332 , n74333 );
nand ( n74335 , n74331 , n74334 );
buf ( n74336 , n74335 );
buf ( n74337 , n74336 );
and ( n74338 , n74320 , n74337 );
and ( n74339 , n74314 , n74319 );
or ( n74340 , n74338 , n74339 );
buf ( n74341 , n74340 );
buf ( n74342 , n74341 );
xor ( n74343 , n74297 , n74342 );
buf ( n74344 , n60104 );
not ( n74345 , n74344 );
buf ( n74346 , n74158 );
not ( n74347 , n74346 );
or ( n74348 , n74345 , n74347 );
buf ( n74349 , n68232 );
buf ( n74350 , n60261 );
and ( n74351 , n74349 , n74350 );
buf ( n74352 , n68235 );
buf ( n74353 , n58880 );
and ( n74354 , n74352 , n74353 );
nor ( n74355 , n74351 , n74354 );
buf ( n74356 , n74355 );
buf ( n74357 , n74356 );
buf ( n74358 , n60270 );
or ( n74359 , n74357 , n74358 );
nand ( n74360 , n74348 , n74359 );
buf ( n74361 , n74360 );
buf ( n74362 , n74361 );
and ( n74363 , n74343 , n74362 );
and ( n74364 , n74297 , n74342 );
or ( n74365 , n74363 , n74364 );
buf ( n74366 , n74365 );
buf ( n74367 , n74366 );
and ( n74368 , n74280 , n74367 );
and ( n74369 , n74275 , n74279 );
or ( n74370 , n74368 , n74369 );
buf ( n74371 , n74370 );
buf ( n74372 , n74371 );
xor ( n74373 , n74258 , n74372 );
xor ( n74374 , n74027 , n74096 );
xor ( n74375 , n74374 , n74170 );
buf ( n74376 , n74375 );
buf ( n74377 , n74376 );
and ( n74378 , n74373 , n74377 );
and ( n74379 , n74258 , n74372 );
or ( n74380 , n74378 , n74379 );
buf ( n74381 , n74380 );
xor ( n74382 , n74241 , n74381 );
xor ( n74383 , n72649 , n72653 );
xor ( n74384 , n74383 , n72675 );
xor ( n74385 , n74174 , n74225 );
xor ( n74386 , n74384 , n74385 );
and ( n74387 , n74382 , n74386 );
and ( n74388 , n74241 , n74381 );
or ( n74389 , n74387 , n74388 );
buf ( n74390 , n74389 );
xor ( n74391 , n72679 , n72696 );
xor ( n74392 , n74391 , n72701 );
buf ( n74393 , n74392 );
buf ( n74394 , n74393 );
xor ( n74395 , n74390 , n74394 );
xor ( n74396 , n73960 , n74009 );
xor ( n74397 , n74396 , n74231 );
buf ( n74398 , n74397 );
buf ( n74399 , n74398 );
and ( n74400 , n74395 , n74399 );
and ( n74401 , n74390 , n74394 );
or ( n74402 , n74400 , n74401 );
buf ( n74403 , n74402 );
xor ( n74404 , n72606 , n72705 );
xor ( n74405 , n74404 , n72709 );
and ( n74406 , n74403 , n74405 );
and ( n74407 , n74235 , n74403 );
or ( n74408 , n74238 , n74406 , n74407 );
buf ( n74409 , n74408 );
xor ( n74410 , n73956 , n74409 );
buf ( n74411 , n41595 );
buf ( n74412 , n25977 );
not ( n74413 , n74412 );
buf ( n74414 , n74413 );
buf ( n74415 , n74414 );
not ( n74416 , n74415 );
buf ( n74417 , n74416 );
buf ( n74418 , n74417 );
not ( n74419 , n74418 );
buf ( n74420 , n41586 );
not ( n74421 , n74420 );
or ( n74422 , n74419 , n74421 );
buf ( n74423 , n41586 );
not ( n74424 , n74423 );
buf ( n74425 , n74424 );
buf ( n74426 , n74425 );
buf ( n74427 , n72310 );
nand ( n74428 , n74426 , n74427 );
buf ( n74429 , n74428 );
buf ( n74430 , n74429 );
nand ( n74431 , n74422 , n74430 );
buf ( n74432 , n74431 );
buf ( n74433 , n74432 );
not ( n74434 , n74433 );
buf ( n74435 , n74434 );
buf ( n74436 , n74435 );
or ( n74437 , n74411 , n74436 );
buf ( n74438 , n73422 );
buf ( n74439 , n41577 );
or ( n74440 , n74438 , n74439 );
nand ( n74441 , n74437 , n74440 );
buf ( n74442 , n74441 );
buf ( n74443 , n74442 );
and ( n74444 , n74410 , n74443 );
and ( n74445 , n73956 , n74409 );
or ( n74446 , n74444 , n74445 );
buf ( n74447 , n74446 );
not ( n74448 , n74447 );
nand ( n74449 , n73951 , n74448 );
not ( n74450 , n74449 );
buf ( n74451 , n44496 );
not ( n74452 , n74451 );
buf ( n74453 , n73456 );
not ( n74454 , n74453 );
or ( n74455 , n74452 , n74454 );
buf ( n74456 , n41570 );
not ( n74457 , n74456 );
buf ( n74458 , n26033 );
not ( n74459 , n74458 );
buf ( n74460 , n74459 );
buf ( n74461 , n74460 );
not ( n74462 , n74461 );
or ( n74463 , n74457 , n74462 );
buf ( n74464 , n42844 );
buf ( n74465 , n25382 );
nand ( n74466 , n74464 , n74465 );
buf ( n74467 , n74466 );
buf ( n74468 , n74467 );
nand ( n74469 , n74463 , n74468 );
buf ( n74470 , n74469 );
buf ( n74471 , n74470 );
buf ( n74472 , n44517 );
nand ( n74473 , n74471 , n74472 );
buf ( n74474 , n74473 );
buf ( n74475 , n74474 );
nand ( n74476 , n74455 , n74475 );
buf ( n74477 , n74476 );
buf ( n74478 , n74477 );
not ( n74479 , n74478 );
buf ( n74480 , n44496 );
not ( n74481 , n74480 );
buf ( n74482 , n74470 );
not ( n74483 , n74482 );
or ( n74484 , n74481 , n74483 );
nand ( n74485 , n44503 , n24835 );
not ( n74486 , n74485 );
nor ( n74487 , n74486 , n44514 );
buf ( n74488 , n74487 );
buf ( n74489 , n74488 );
buf ( n74490 , n41570 );
not ( n74491 , n74490 );
buf ( n74492 , n74491 );
buf ( n74493 , n74492 );
not ( n74494 , n74493 );
buf ( n74495 , n25997 );
not ( n74496 , n74495 );
or ( n74497 , n74494 , n74496 );
buf ( n74498 , n25997 );
buf ( n74499 , n74498 );
buf ( n74500 , n74499 );
buf ( n74501 , n74500 );
not ( n74502 , n74501 );
buf ( n74503 , n74502 );
buf ( n74504 , n74503 );
buf ( n74505 , n25385 );
nand ( n74506 , n74504 , n74505 );
buf ( n74507 , n74506 );
buf ( n74508 , n74507 );
nand ( n74509 , n74497 , n74508 );
buf ( n74510 , n74509 );
buf ( n74511 , n74510 );
nand ( n74512 , n74489 , n74511 );
buf ( n74513 , n74512 );
buf ( n74514 , n74513 );
nand ( n74515 , n74484 , n74514 );
buf ( n74516 , n74515 );
not ( n74517 , n74516 );
not ( n74518 , n74517 );
xor ( n74519 , n72606 , n72705 );
xor ( n74520 , n74519 , n72709 );
xor ( n74521 , n74235 , n74403 );
xor ( n74522 , n74520 , n74521 );
not ( n74523 , n74522 );
not ( n74524 , n74523 );
or ( n74525 , n74518 , n74524 );
buf ( n74526 , n46390 );
not ( n74527 , n74526 );
buf ( n74528 , n25336 );
not ( n74529 , n74528 );
buf ( n74530 , n74529 );
buf ( n74531 , n74530 );
not ( n74532 , n74531 );
or ( n74533 , n74527 , n74532 );
buf ( n74534 , n74425 );
buf ( n74535 , n46387 );
nand ( n74536 , n74534 , n74535 );
buf ( n74537 , n74536 );
buf ( n74538 , n74537 );
nand ( n74539 , n74533 , n74538 );
buf ( n74540 , n74539 );
not ( n74541 , n74540 );
not ( n74542 , n67354 );
or ( n74543 , n74541 , n74542 );
buf ( n74544 , n74432 );
buf ( n74545 , n41574 );
nand ( n74546 , n74544 , n74545 );
buf ( n74547 , n74546 );
nand ( n74548 , n74543 , n74547 );
nand ( n74549 , n74525 , n74548 );
not ( n74550 , n74523 );
nand ( n74551 , n74550 , n74516 );
nand ( n74552 , n74549 , n74551 );
buf ( n74553 , n74552 );
not ( n74554 , n74553 );
or ( n74555 , n74479 , n74554 );
buf ( n74556 , n74552 );
buf ( n74557 , n74477 );
or ( n74558 , n74556 , n74557 );
xor ( n74559 , n73956 , n74409 );
xor ( n74560 , n74559 , n74443 );
buf ( n74561 , n74560 );
buf ( n74562 , n74561 );
nand ( n74563 , n74558 , n74562 );
buf ( n74564 , n74563 );
buf ( n74565 , n74564 );
nand ( n74566 , n74555 , n74565 );
buf ( n74567 , n74566 );
not ( n74568 , n74567 );
or ( n74569 , n74450 , n74568 );
nand ( n74570 , n73950 , n74447 );
nand ( n74571 , n74569 , n74570 );
buf ( n74572 , n74571 );
not ( n74573 , n67149 );
nand ( n74574 , n73631 , n73633 );
not ( n74575 , n74574 );
or ( n74576 , n74573 , n74575 );
buf ( n74577 , n73474 );
buf ( n74578 , n71048 );
nand ( n74579 , n74577 , n74578 );
buf ( n74580 , n74579 );
nand ( n74581 , n74576 , n74580 );
buf ( n74582 , n74581 );
xor ( n74583 , n74572 , n74582 );
buf ( n74584 , n50060 );
not ( n74585 , n74584 );
buf ( n74586 , n42342 );
not ( n74587 , n74586 );
or ( n74588 , n74585 , n74587 );
buf ( n74589 , n42366 );
buf ( n74590 , n67438 );
nand ( n74591 , n74589 , n74590 );
buf ( n74592 , n74591 );
buf ( n74593 , n74592 );
nand ( n74594 , n74588 , n74593 );
buf ( n74595 , n74594 );
buf ( n74596 , n74595 );
not ( n74597 , n74596 );
buf ( n74598 , n66459 );
not ( n74599 , n74598 );
or ( n74600 , n74597 , n74599 );
buf ( n74601 , n72289 );
buf ( n74602 , n66482 );
nand ( n74603 , n74601 , n74602 );
buf ( n74604 , n74603 );
buf ( n74605 , n74604 );
nand ( n74606 , n74600 , n74605 );
buf ( n74607 , n74606 );
buf ( n74608 , n74607 );
and ( n74609 , n74583 , n74608 );
and ( n74610 , n74572 , n74582 );
or ( n74611 , n74609 , n74610 );
buf ( n74612 , n74611 );
and ( n74613 , n73930 , n74612 );
and ( n74614 , n73920 , n73929 );
or ( n74615 , n74613 , n74614 );
buf ( n74616 , n74615 );
xor ( n74617 , n73915 , n74616 );
buf ( n74618 , n74617 );
buf ( n74619 , n74618 );
nand ( n74620 , n73904 , n74619 );
buf ( n74621 , n74620 );
buf ( n74622 , n74621 );
buf ( n74623 , n73876 );
not ( n74624 , n74623 );
buf ( n74625 , n73898 );
nand ( n74626 , n74624 , n74625 );
buf ( n74627 , n74626 );
buf ( n74628 , n74627 );
nand ( n74629 , n74622 , n74628 );
buf ( n74630 , n74629 );
buf ( n74631 , n74630 );
nand ( n74632 , n73874 , n74631 );
buf ( n74633 , n74632 );
buf ( n74634 , n74633 );
nand ( n74635 , n73871 , n74634 );
buf ( n74636 , n74635 );
buf ( n74637 , n74636 );
xor ( n74638 , n73312 , n74637 );
buf ( n74639 , n74638 );
buf ( n74640 , n74639 );
not ( n74641 , n74640 );
buf ( n74642 , n74641 );
buf ( n74643 , n74642 );
not ( n74644 , n74643 );
xor ( n74645 , n73024 , n73033 );
and ( n74646 , n74645 , n73053 );
and ( n74647 , n73024 , n73033 );
or ( n74648 , n74646 , n74647 );
buf ( n74649 , n74648 );
buf ( n74650 , n74649 );
buf ( n74651 , n42710 );
buf ( n74652 , n74651 );
buf ( n74653 , n73774 );
not ( n74654 , n74653 );
buf ( n74655 , n74654 );
buf ( n74656 , n74655 );
or ( n74657 , n74652 , n74656 );
buf ( n74658 , n42856 );
not ( n74659 , n74658 );
buf ( n74660 , n25227 );
not ( n74661 , n74660 );
or ( n74662 , n74659 , n74661 );
buf ( n74663 , n25226 );
buf ( n74664 , n42859 );
nand ( n74665 , n74663 , n74664 );
buf ( n74666 , n74665 );
buf ( n74667 , n74666 );
nand ( n74668 , n74662 , n74667 );
buf ( n74669 , n74668 );
buf ( n74670 , n74669 );
not ( n74671 , n74670 );
buf ( n74672 , n74671 );
buf ( n74673 , n74672 );
buf ( n74674 , n42664 );
buf ( n74675 , n74674 );
or ( n74676 , n74673 , n74675 );
nand ( n74677 , n74657 , n74676 );
buf ( n74678 , n74677 );
buf ( n74679 , n74678 );
xor ( n74680 , n70289 , n70417 );
xor ( n74681 , n74680 , n70421 );
xor ( n74682 , n70670 , n70731 );
xor ( n74683 , n74681 , n74682 );
buf ( n74684 , n74683 );
xor ( n74685 , n70721 , n70724 );
xor ( n74686 , n74685 , n70728 );
and ( n74687 , n73728 , n74686 );
xor ( n74688 , n70721 , n70724 );
xor ( n74689 , n74688 , n70728 );
and ( n74690 , n73732 , n74689 );
and ( n74691 , n73728 , n73732 );
or ( n74692 , n74687 , n74690 , n74691 );
buf ( n74693 , n74692 );
xor ( n74694 , n74684 , n74693 );
buf ( n74695 , n42309 );
not ( n74696 , n74695 );
buf ( n74697 , n25306 );
not ( n74698 , n74697 );
buf ( n74699 , n66398 );
not ( n74700 , n74699 );
or ( n74701 , n74698 , n74700 );
buf ( n74702 , n71123 );
not ( n74703 , n74702 );
buf ( n74704 , n28430 );
nand ( n74705 , n74703 , n74704 );
buf ( n74706 , n74705 );
buf ( n74707 , n74706 );
nand ( n74708 , n74701 , n74707 );
buf ( n74709 , n74708 );
buf ( n74710 , n74709 );
not ( n74711 , n74710 );
or ( n74712 , n74696 , n74711 );
buf ( n74713 , n42246 );
buf ( n74714 , n73748 );
nand ( n74715 , n74713 , n74714 );
buf ( n74716 , n74715 );
buf ( n74717 , n74716 );
nand ( n74718 , n74712 , n74717 );
buf ( n74719 , n74718 );
buf ( n74720 , n74719 );
xor ( n74721 , n74694 , n74720 );
buf ( n74722 , n74721 );
buf ( n74723 , n74722 );
xor ( n74724 , n74679 , n74723 );
buf ( n74725 , n73044 );
not ( n74726 , n74725 );
buf ( n74727 , n66459 );
not ( n74728 , n74727 );
or ( n74729 , n74726 , n74728 );
buf ( n74730 , n44952 );
not ( n74731 , n74730 );
buf ( n74732 , n66463 );
not ( n74733 , n74732 );
or ( n74734 , n74731 , n74733 );
buf ( n74735 , n69804 );
buf ( n74736 , n44949 );
nand ( n74737 , n74735 , n74736 );
buf ( n74738 , n74737 );
buf ( n74739 , n74738 );
nand ( n74740 , n74734 , n74739 );
buf ( n74741 , n74740 );
buf ( n74742 , n74741 );
buf ( n74743 , n66482 );
nand ( n74744 , n74742 , n74743 );
buf ( n74745 , n74744 );
buf ( n74746 , n74745 );
nand ( n74747 , n74729 , n74746 );
buf ( n74748 , n74747 );
buf ( n74749 , n74748 );
xor ( n74750 , n74724 , n74749 );
buf ( n74751 , n74750 );
buf ( n74752 , n74751 );
xor ( n74753 , n74650 , n74752 );
not ( n74754 , n73810 );
not ( n74755 , n44517 );
or ( n74756 , n74754 , n74755 );
buf ( n74757 , n65010 );
not ( n74758 , n74757 );
buf ( n74759 , n63906 );
not ( n74760 , n74759 );
or ( n74761 , n74758 , n74760 );
buf ( n74762 , n13653 );
buf ( n74763 , n44530 );
nand ( n74764 , n74762 , n74763 );
buf ( n74765 , n74764 );
buf ( n74766 , n74765 );
nand ( n74767 , n74761 , n74766 );
buf ( n74768 , n74767 );
buf ( n74769 , n74768 );
not ( n74770 , n74769 );
buf ( n74771 , n74770 );
or ( n74772 , n74771 , n44497 );
nand ( n74773 , n74756 , n74772 );
buf ( n74774 , n74773 );
xor ( n74775 , n74753 , n74774 );
buf ( n74776 , n74775 );
buf ( n74777 , n74776 );
xor ( n74778 , n73056 , n73093 );
and ( n74779 , n74778 , n73223 );
and ( n74780 , n73056 , n73093 );
or ( n74781 , n74779 , n74780 );
buf ( n74782 , n74781 );
buf ( n74783 , n74782 );
xor ( n74784 , n74777 , n74783 );
buf ( n74785 , n73085 );
not ( n74786 , n74785 );
buf ( n74787 , n53628 );
not ( n74788 , n74787 );
or ( n74789 , n74786 , n74788 );
buf ( n74790 , n48323 );
not ( n74791 , n74790 );
buf ( n74792 , n42556 );
not ( n74793 , n74792 );
or ( n74794 , n74791 , n74793 );
buf ( n74795 , n61462 );
buf ( n74796 , n48320 );
nand ( n74797 , n74795 , n74796 );
buf ( n74798 , n74797 );
buf ( n74799 , n74798 );
nand ( n74800 , n74794 , n74799 );
buf ( n74801 , n74800 );
buf ( n74802 , n74801 );
buf ( n74803 , n43905 );
nand ( n74804 , n74802 , n74803 );
buf ( n74805 , n74804 );
buf ( n74806 , n74805 );
nand ( n74807 , n74789 , n74806 );
buf ( n74808 , n74807 );
buf ( n74809 , n74808 );
not ( n74810 , n74809 );
buf ( n74811 , n74810 );
xor ( n74812 , n73785 , n73795 );
and ( n74813 , n74812 , n73821 );
and ( n74814 , n73785 , n73795 );
or ( n74815 , n74813 , n74814 );
buf ( n74816 , n74815 );
xor ( n74817 , n74811 , n74816 );
buf ( n74818 , n71107 );
not ( n74819 , n74818 );
buf ( n74820 , n62588 );
not ( n74821 , n74820 );
or ( n74822 , n74819 , n74821 );
buf ( n74823 , n46390 );
not ( n74824 , n74823 );
buf ( n74825 , n62598 );
not ( n74826 , n74825 );
or ( n74827 , n74824 , n74826 );
buf ( n74828 , n61434 );
buf ( n74829 , n46393 );
nand ( n74830 , n74828 , n74829 );
buf ( n74831 , n74830 );
buf ( n74832 , n74831 );
nand ( n74833 , n74827 , n74832 );
buf ( n74834 , n74833 );
buf ( n74835 , n74834 );
buf ( n74836 , n62582 );
nand ( n74837 , n74835 , n74836 );
buf ( n74838 , n74837 );
buf ( n74839 , n74838 );
nand ( n74840 , n74822 , n74839 );
buf ( n74841 , n74840 );
not ( n74842 , n73004 );
not ( n74843 , n41596 );
or ( n74844 , n74842 , n74843 );
buf ( n74845 , n13662 );
buf ( n74846 , n41605 );
xnor ( n74847 , n74845 , n74846 );
buf ( n74848 , n74847 );
or ( n74849 , n74848 , n41577 );
nand ( n74850 , n74844 , n74849 );
buf ( n74851 , n74850 );
not ( n74852 , n74851 );
xor ( n74853 , n73735 , n73756 );
and ( n74854 , n74853 , n73782 );
and ( n74855 , n73735 , n73756 );
or ( n74856 , n74854 , n74855 );
buf ( n74857 , n74856 );
buf ( n74858 , n74857 );
not ( n74859 , n74858 );
buf ( n74860 , n74859 );
buf ( n74861 , n74860 );
not ( n74862 , n74861 );
and ( n74863 , n74852 , n74862 );
buf ( n74864 , n74850 );
buf ( n74865 , n74860 );
and ( n74866 , n74864 , n74865 );
nor ( n74867 , n74863 , n74866 );
buf ( n74868 , n74867 );
xor ( n74869 , n74841 , n74868 );
xor ( n74870 , n74817 , n74869 );
buf ( n74871 , n74870 );
xor ( n74872 , n74784 , n74871 );
buf ( n74873 , n74872 );
xor ( n74874 , n73718 , n73844 );
and ( n74875 , n74874 , n73866 );
and ( n74876 , n73718 , n73844 );
or ( n74877 , n74875 , n74876 );
buf ( n74878 , n74877 );
xor ( n74879 , n74873 , n74878 );
buf ( n74880 , n74879 );
xor ( n74881 , n73824 , n73829 );
and ( n74882 , n74881 , n73841 );
and ( n74883 , n73824 , n73829 );
or ( n74884 , n74882 , n74883 );
buf ( n74885 , n74884 );
buf ( n74886 , n48868 );
not ( n74887 , n74886 );
buf ( n74888 , n48808 );
not ( n74889 , n74888 );
buf ( n74890 , n42195 );
not ( n74891 , n74890 );
or ( n74892 , n74889 , n74891 );
buf ( n74893 , n29360 );
buf ( n74894 , n72891 );
nand ( n74895 , n74893 , n74894 );
buf ( n74896 , n74895 );
buf ( n74897 , n74896 );
nand ( n74898 , n74892 , n74897 );
buf ( n74899 , n74898 );
buf ( n74900 , n74899 );
not ( n74901 , n74900 );
or ( n74902 , n74887 , n74901 );
buf ( n74903 , n72897 );
buf ( n74904 , n48855 );
nand ( n74905 , n74903 , n74904 );
buf ( n74906 , n74905 );
buf ( n74907 , n74906 );
nand ( n74908 , n74902 , n74907 );
buf ( n74909 , n74908 );
buf ( n74910 , n74909 );
not ( n74911 , n74910 );
buf ( n74912 , n74911 );
and ( n74913 , n74885 , n74912 );
not ( n74914 , n74885 );
and ( n74915 , n74914 , n74909 );
or ( n74916 , n74913 , n74915 );
buf ( n74917 , n74916 );
buf ( n74918 , n12481 );
buf ( n74919 , n42468 );
and ( n74920 , n74918 , n74919 );
not ( n74921 , n74918 );
buf ( n74922 , n38994 );
and ( n74923 , n74921 , n74922 );
nor ( n74924 , n74920 , n74923 );
buf ( n74925 , n74924 );
buf ( n74926 , n74925 );
not ( n74927 , n74926 );
buf ( n74928 , n45059 );
not ( n74929 , n74928 );
or ( n74930 , n74927 , n74929 );
buf ( n74931 , n55841 );
not ( n74932 , n74931 );
buf ( n74933 , n42471 );
not ( n74934 , n74933 );
or ( n74935 , n74932 , n74934 );
buf ( n74936 , n38979 );
buf ( n74937 , n55840 );
nand ( n74938 , n74936 , n74937 );
buf ( n74939 , n74938 );
buf ( n74940 , n74939 );
nand ( n74941 , n74935 , n74940 );
buf ( n74942 , n74941 );
buf ( n74943 , n74942 );
buf ( n74944 , n50104 );
nand ( n74945 , n74943 , n74944 );
buf ( n74946 , n74945 );
buf ( n74947 , n74946 );
nand ( n74948 , n74930 , n74947 );
buf ( n74949 , n74948 );
buf ( n74950 , n74949 );
not ( n74951 , n74950 );
buf ( n74952 , n74951 );
buf ( n74953 , n74952 );
and ( n74954 , n74917 , n74953 );
not ( n74955 , n74917 );
buf ( n74956 , n74949 );
and ( n74957 , n74955 , n74956 );
nor ( n74958 , n74954 , n74957 );
buf ( n74959 , n74958 );
buf ( n74960 , n74959 );
not ( n74961 , n74960 );
buf ( n74962 , n74961 );
buf ( n74963 , n74962 );
and ( n74964 , n74880 , n74963 );
not ( n74965 , n74880 );
buf ( n74966 , n74959 );
and ( n74967 , n74965 , n74966 );
nor ( n74968 , n74964 , n74967 );
buf ( n74969 , n74968 );
buf ( n74970 , n74969 );
not ( n74971 , n74970 );
buf ( n74972 , n74971 );
buf ( n74973 , n74972 );
not ( n74974 , n74973 );
buf ( n74975 , n39671 );
not ( n74976 , n74975 );
buf ( n74977 , n74976 );
xor ( n74978 , n73910 , n73914 );
and ( n74979 , n74978 , n74616 );
and ( n74980 , n73910 , n73914 );
or ( n74981 , n74979 , n74980 );
buf ( n74982 , n74981 );
buf ( n74983 , n74982 );
buf ( n74984 , n42628 );
not ( n74985 , n74984 );
buf ( n74986 , n74985 );
buf ( n74987 , n74986 );
buf ( n74988 , n53548 );
buf ( n74989 , n25159 );
and ( n74990 , n74988 , n74989 );
not ( n74991 , n74988 );
buf ( n74992 , n46356 );
and ( n74993 , n74991 , n74992 );
nor ( n74994 , n74990 , n74993 );
buf ( n74995 , n74994 );
buf ( n74996 , n74995 );
or ( n74997 , n74987 , n74996 );
buf ( n74998 , n72851 );
buf ( n74999 , n42563 );
or ( n75000 , n74998 , n74999 );
nand ( n75001 , n74997 , n75000 );
buf ( n75002 , n75001 );
buf ( n75003 , n75002 );
buf ( n75004 , n46073 );
buf ( n75005 , n12481 );
or ( n75006 , n75004 , n75005 );
buf ( n75007 , n24092 );
buf ( n75008 , n56325 );
or ( n75009 , n75007 , n75008 );
nand ( n75010 , n75006 , n75009 );
buf ( n75011 , n75010 );
buf ( n75012 , n75011 );
not ( n75013 , n75012 );
buf ( n75014 , n39999 );
not ( n75015 , n75014 );
or ( n75016 , n75013 , n75015 );
buf ( n75017 , n72976 );
buf ( n75018 , n46633 );
nand ( n75019 , n75017 , n75018 );
buf ( n75020 , n75019 );
buf ( n75021 , n75020 );
nand ( n75022 , n75016 , n75021 );
buf ( n75023 , n75022 );
buf ( n75024 , n75023 );
xor ( n75025 , n75003 , n75024 );
buf ( n75026 , n72912 );
not ( n75027 , n75026 );
buf ( n75028 , n75027 );
buf ( n75029 , n75028 );
buf ( n75030 , n48871 );
or ( n75031 , n75029 , n75030 );
buf ( n75032 , n73578 );
buf ( n75033 , n48852 );
nand ( n75034 , n75032 , n75033 );
buf ( n75035 , n75034 );
buf ( n75036 , n75035 );
nand ( n75037 , n75031 , n75036 );
buf ( n75038 , n75037 );
buf ( n75039 , n75038 );
and ( n75040 , n75025 , n75039 );
and ( n75041 , n75003 , n75024 );
or ( n75042 , n75040 , n75041 );
buf ( n75043 , n75042 );
buf ( n75044 , n75043 );
not ( n75045 , n43806 );
buf ( n75046 , C0 );
buf ( n75047 , n75046 );
and ( n75048 , n74983 , n75044 );
or ( n75049 , C0 , n75048 );
buf ( n75050 , n75049 );
buf ( n75051 , n75050 );
buf ( n75052 , C1 );
buf ( n75053 , n75052 );
nand ( n75054 , n75051 , n75053 );
buf ( n75055 , n75054 );
buf ( n75056 , n75055 );
nand ( n75057 , C1 , n75056 );
buf ( n75058 , n75057 );
buf ( n75059 , n75058 );
buf ( n75060 , C0 );
buf ( n75061 , n75060 );
xor ( n75062 , n72843 , n72879 );
xor ( n75063 , n75062 , n72920 );
buf ( n75064 , n75063 );
buf ( n75065 , n75064 );
or ( n75066 , n75061 , n75065 );
xor ( n75067 , n72964 , n72997 );
xor ( n75068 , n75067 , n73226 );
buf ( n75069 , n75068 );
buf ( n75070 , n75069 );
nand ( n75071 , n75066 , n75070 );
buf ( n75072 , n75071 );
buf ( n75073 , n75072 );
buf ( n75074 , C1 );
buf ( n75075 , n75074 );
and ( n75076 , n75073 , n75075 );
buf ( n75077 , n75076 );
buf ( n75078 , n75077 );
and ( n75079 , n75059 , n75078 );
not ( n75080 , n75059 );
buf ( n75081 , n75077 );
not ( n75082 , n75081 );
buf ( n75083 , n75082 );
buf ( n75084 , n75083 );
and ( n75085 , n75080 , n75084 );
nor ( n75086 , n75079 , n75085 );
buf ( n75087 , n75086 );
buf ( n75088 , n75087 );
not ( n75089 , n75088 );
buf ( n75090 , n75089 );
buf ( n75091 , n75090 );
not ( n75092 , n75091 );
or ( n75093 , n74974 , n75092 );
buf ( n75094 , n75087 );
buf ( n75095 , n74969 );
nand ( n75096 , n75094 , n75095 );
buf ( n75097 , n75096 );
buf ( n75098 , n75097 );
nand ( n75099 , n75093 , n75098 );
buf ( n75100 , n75099 );
buf ( n75101 , n75100 );
xor ( n75102 , n74983 , n75044 );
xor ( n75103 , n75102 , n75047 );
buf ( n75104 , n75103 );
buf ( n75105 , n75104 );
xor ( n75106 , n75003 , n75024 );
xor ( n75107 , n75106 , n75039 );
buf ( n75108 , n75107 );
buf ( n75109 , n75108 );
buf ( n75110 , C0 );
buf ( n75111 , n75110 );
xor ( n75112 , n75109 , n75111 );
xor ( n75113 , n73377 , n73383 );
xor ( n75114 , n75113 , n73648 );
buf ( n75115 , n75114 );
buf ( n75116 , n75115 );
and ( n75117 , n75112 , n75116 );
or ( n75118 , n75117 , C0 );
buf ( n75119 , n75118 );
buf ( n75120 , n75119 );
xor ( n75121 , n75105 , n75120 );
xor ( n75122 , n73920 , n73929 );
xor ( n75123 , n75122 , n74612 );
buf ( n75124 , n75123 );
not ( n75125 , n46912 );
not ( n75126 , n73330 );
or ( n75127 , n75125 , n75126 );
buf ( n75128 , n46875 );
not ( n75129 , n75128 );
buf ( n75130 , n41733 );
not ( n75131 , n75130 );
or ( n75132 , n75129 , n75131 );
buf ( n75133 , n60327 );
buf ( n75134 , n46887 );
nand ( n75135 , n75133 , n75134 );
buf ( n75136 , n75135 );
buf ( n75137 , n75136 );
nand ( n75138 , n75132 , n75137 );
buf ( n75139 , n75138 );
buf ( n75140 , n75139 );
buf ( n75141 , n46907 );
nand ( n75142 , n75140 , n75141 );
buf ( n75143 , n75142 );
nand ( n75144 , n75127 , n75143 );
buf ( n75145 , n47725 );
not ( n75146 , n75145 );
buf ( n75147 , n25290 );
not ( n75148 , n75147 );
or ( n75149 , n75146 , n75148 );
buf ( n75150 , n42257 );
not ( n75151 , n75150 );
buf ( n75152 , n75151 );
buf ( n75153 , n75152 );
not ( n75154 , n75153 );
buf ( n75155 , n47716 );
nand ( n75156 , n75154 , n75155 );
buf ( n75157 , n75156 );
buf ( n75158 , n75157 );
nand ( n75159 , n75149 , n75158 );
buf ( n75160 , n75159 );
buf ( n75161 , n75160 );
not ( n75162 , n75161 );
buf ( n75163 , n42246 );
not ( n75164 , n75163 );
or ( n75165 , n75162 , n75164 );
buf ( n75166 , n73942 );
buf ( n75167 , n42309 );
nand ( n75168 , n75166 , n75167 );
buf ( n75169 , n75168 );
buf ( n75170 , n75169 );
nand ( n75171 , n75165 , n75170 );
buf ( n75172 , n75171 );
buf ( n75173 , n75172 );
buf ( n75174 , n67149 );
not ( n75175 , n75174 );
buf ( n75176 , n73481 );
not ( n75177 , n75176 );
or ( n75178 , n75175 , n75177 );
buf ( n75179 , n45746 );
buf ( n75180 , n43056 );
and ( n75181 , n75179 , n75180 );
not ( n75182 , n75179 );
buf ( n75183 , n43055 );
and ( n75184 , n75182 , n75183 );
or ( n75185 , n75181 , n75184 );
buf ( n75186 , n75185 );
buf ( n75187 , n75186 );
not ( n75188 , n75187 );
buf ( n75189 , n71048 );
nand ( n75190 , n75188 , n75189 );
buf ( n75191 , n75190 );
buf ( n75192 , n75191 );
nand ( n75193 , n75178 , n75192 );
buf ( n75194 , n75193 );
buf ( n75195 , n75194 );
xor ( n75196 , n75173 , n75195 );
buf ( n75197 , n50060 );
not ( n75198 , n75197 );
buf ( n75199 , n42324 );
not ( n75200 , n75199 );
or ( n75201 , n75198 , n75200 );
buf ( n75202 , n25226 );
buf ( n75203 , n67438 );
nand ( n75204 , n75202 , n75203 );
buf ( n75205 , n75204 );
buf ( n75206 , n75205 );
nand ( n75207 , n75201 , n75206 );
buf ( n75208 , n75207 );
buf ( n75209 , n75208 );
not ( n75210 , n75209 );
buf ( n75211 , n73163 );
not ( n75212 , n75211 );
or ( n75213 , n75210 , n75212 );
buf ( n75214 , n73388 );
buf ( n75215 , n42665 );
nand ( n75216 , n75214 , n75215 );
buf ( n75217 , n75216 );
buf ( n75218 , n75217 );
nand ( n75219 , n75213 , n75218 );
buf ( n75220 , n75219 );
buf ( n75221 , n75220 );
and ( n75222 , n75196 , n75221 );
and ( n75223 , n75173 , n75195 );
or ( n75224 , n75222 , n75223 );
buf ( n75225 , n75224 );
not ( n75226 , n75225 );
and ( n75227 , n73951 , n74448 );
not ( n75228 , n73951 );
and ( n75229 , n75228 , n74447 );
nor ( n75230 , n75227 , n75229 );
xor ( n75231 , n74567 , n75230 );
not ( n75232 , n75231 );
or ( n75233 , n75226 , n75232 );
or ( n75234 , n75225 , n75231 );
buf ( n75235 , n50995 );
not ( n75236 , n75235 );
buf ( n75237 , n69798 );
not ( n75238 , n75237 );
or ( n75239 , n75236 , n75238 );
buf ( n75240 , n68062 );
buf ( n75241 , n50998 );
nand ( n75242 , n75240 , n75241 );
buf ( n75243 , n75242 );
buf ( n75244 , n75243 );
nand ( n75245 , n75239 , n75244 );
buf ( n75246 , n75245 );
buf ( n75247 , n75246 );
not ( n75248 , n75247 );
buf ( n75249 , n66459 );
not ( n75250 , n75249 );
or ( n75251 , n75248 , n75250 );
buf ( n75252 , n74595 );
buf ( n75253 , n66482 );
nand ( n75254 , n75252 , n75253 );
buf ( n75255 , n75254 );
buf ( n75256 , n75255 );
nand ( n75257 , n75251 , n75256 );
buf ( n75258 , n75257 );
nand ( n75259 , n75234 , n75258 );
nand ( n75260 , n75233 , n75259 );
xor ( n75261 , n75144 , n75260 );
buf ( n75262 , n54068 );
buf ( n75263 , n75262 );
buf ( n75264 , n42613 );
not ( n75265 , n75264 );
buf ( n75266 , n75265 );
buf ( n75267 , n75266 );
nand ( n75268 , n75263 , n75267 );
buf ( n75269 , n75268 );
buf ( n75270 , n75266 );
buf ( n75271 , n52724 );
or ( n75272 , n75270 , n75271 );
buf ( n75273 , n12481 );
nand ( n75274 , n75272 , n75273 );
buf ( n75275 , n75274 );
and ( n75276 , n75269 , n75275 , n25159 );
and ( n75277 , n75261 , n75276 );
and ( n75278 , n75144 , n75260 );
or ( n75279 , n75277 , n75278 );
buf ( n75280 , n75279 );
xor ( n75281 , n75124 , n75280 );
buf ( n75282 , n51488 );
not ( n75283 , n75282 );
buf ( n75284 , n48836 );
not ( n75285 , n75284 );
buf ( n75286 , n50091 );
not ( n75287 , n75286 );
or ( n75288 , n75285 , n75287 );
buf ( n75289 , n42149 );
buf ( n75290 , n72931 );
nand ( n75291 , n75289 , n75290 );
buf ( n75292 , n75291 );
buf ( n75293 , n75292 );
nand ( n75294 , n75288 , n75293 );
buf ( n75295 , n75294 );
buf ( n75296 , n75295 );
not ( n75297 , n75296 );
or ( n75298 , n75283 , n75297 );
buf ( n75299 , n73891 );
buf ( n75300 , n62125 );
nand ( n75301 , n75299 , n75300 );
buf ( n75302 , n75301 );
buf ( n75303 , n75302 );
nand ( n75304 , n75298 , n75303 );
buf ( n75305 , n75304 );
buf ( n75306 , n75305 );
and ( n75307 , n75281 , n75306 );
and ( n75308 , n75124 , n75280 );
or ( n75309 , n75307 , n75308 );
buf ( n75310 , n75309 );
buf ( n75311 , n75310 );
buf ( n75312 , n55841 );
buf ( n75313 , n42578 );
and ( n75314 , n75312 , n75313 );
not ( n75315 , n75312 );
buf ( n75316 , n46356 );
and ( n75317 , n75315 , n75316 );
nor ( n75318 , n75314 , n75317 );
buf ( n75319 , n75318 );
buf ( n75320 , n75319 );
not ( n75321 , n75320 );
buf ( n75322 , n50128 );
not ( n75323 , n75322 );
or ( n75324 , n75321 , n75323 );
buf ( n75325 , n74995 );
not ( n75326 , n75325 );
buf ( n75327 , n42566 );
nand ( n75328 , n75326 , n75327 );
buf ( n75329 , n75328 );
buf ( n75330 , n75329 );
nand ( n75331 , n75324 , n75330 );
buf ( n75332 , n75331 );
buf ( n75333 , n75332 );
buf ( n75334 , n53539 );
not ( n75335 , n75334 );
buf ( n75336 , n25181 );
not ( n75337 , n75336 );
or ( n75338 , n75335 , n75337 );
buf ( n75339 , n54068 );
buf ( n75340 , n53548 );
nand ( n75341 , n75339 , n75340 );
buf ( n75342 , n75341 );
buf ( n75343 , n75342 );
nand ( n75344 , n75338 , n75343 );
buf ( n75345 , n75344 );
buf ( n75346 , n75345 );
not ( n75347 , n75346 );
buf ( n75348 , n43938 );
not ( n75349 , n75348 );
or ( n75350 , n75347 , n75349 );
buf ( n75351 , n73345 );
buf ( n75352 , n43905 );
nand ( n75353 , n75351 , n75352 );
buf ( n75354 , n75353 );
buf ( n75355 , n75354 );
nand ( n75356 , n75350 , n75355 );
buf ( n75357 , n75356 );
buf ( n75358 , n75357 );
xor ( n75359 , n74572 , n74582 );
xor ( n75360 , n75359 , n74608 );
buf ( n75361 , n75360 );
buf ( n75362 , n75361 );
xor ( n75363 , n75358 , n75362 );
buf ( n75364 , n48868 );
not ( n75365 , n75364 );
buf ( n75366 , n73594 );
not ( n75367 , n75366 );
or ( n75368 , n75365 , n75367 );
buf ( n75369 , n48808 );
not ( n75370 , n75369 );
buf ( n75371 , n56545 );
not ( n75372 , n75371 );
or ( n75373 , n75370 , n75372 );
buf ( n75374 , n29754 );
buf ( n75375 , n48808 );
not ( n75376 , n75375 );
buf ( n75377 , n75376 );
buf ( n75378 , n75377 );
nand ( n75379 , n75374 , n75378 );
buf ( n75380 , n75379 );
buf ( n75381 , n75380 );
nand ( n75382 , n75373 , n75381 );
buf ( n75383 , n75382 );
buf ( n75384 , n75383 );
buf ( n75385 , n48852 );
nand ( n75386 , n75384 , n75385 );
buf ( n75387 , n75386 );
buf ( n75388 , n75387 );
nand ( n75389 , n75368 , n75388 );
buf ( n75390 , n75389 );
buf ( n75391 , n75390 );
and ( n75392 , n75363 , n75391 );
and ( n75393 , n75358 , n75362 );
or ( n75394 , n75392 , n75393 );
buf ( n75395 , n75394 );
buf ( n75396 , n75395 );
xor ( n75397 , n75333 , n75396 );
buf ( n75398 , n73332 );
not ( n75399 , n75398 );
buf ( n75400 , n73361 );
not ( n75401 , n75400 );
or ( n75402 , n75399 , n75401 );
buf ( n75403 , n73361 );
buf ( n75404 , n73332 );
or ( n75405 , n75403 , n75404 );
nand ( n75406 , n75402 , n75405 );
buf ( n75407 , n75406 );
buf ( n75408 , n75407 );
buf ( n75409 , n73370 );
and ( n75410 , n75408 , n75409 );
not ( n75411 , n75408 );
buf ( n75412 , n73338 );
and ( n75413 , n75411 , n75412 );
nor ( n75414 , n75410 , n75413 );
buf ( n75415 , n75414 );
buf ( n75416 , n75415 );
and ( n75417 , n75397 , n75416 );
and ( n75418 , n75333 , n75396 );
or ( n75419 , n75417 , n75418 );
buf ( n75420 , n75419 );
buf ( n75421 , n75420 );
buf ( n75422 , C0 );
buf ( n75423 , n75422 );
and ( n75424 , n75311 , n75421 );
or ( n75425 , C0 , n75424 );
buf ( n75426 , n75425 );
buf ( n75427 , n75426 );
and ( n75428 , n75121 , n75427 );
and ( n75429 , n75105 , n75120 );
or ( n75430 , n75428 , n75429 );
buf ( n75431 , n75430 );
buf ( n75432 , n75431 );
not ( n75433 , n75432 );
buf ( n75434 , n75433 );
buf ( n75435 , n75434 );
and ( n75436 , n75101 , n75435 );
not ( n75437 , n75101 );
buf ( n75438 , n75431 );
and ( n75439 , n75437 , n75438 );
nor ( n75440 , n75436 , n75439 );
buf ( n75441 , n75440 );
buf ( n75442 , n75441 );
not ( n75443 , n75442 );
or ( n75444 , n74644 , n75443 );
xor ( n75445 , n75069 , n75060 );
xnor ( n75446 , n75445 , n75064 );
buf ( n75447 , n75446 );
not ( n75448 , n75447 );
buf ( n75449 , n73652 );
buf ( n75450 , n74630 );
xor ( n75451 , n75449 , n75450 );
buf ( n75452 , n73868 );
xnor ( n75453 , n75451 , n75452 );
buf ( n75454 , n75453 );
buf ( n75455 , n75454 );
not ( n75456 , n75455 );
or ( n75457 , n75448 , n75456 );
buf ( n75458 , n46912 );
not ( n75459 , n75458 );
buf ( n75460 , n75139 );
not ( n75461 , n75460 );
or ( n75462 , n75459 , n75461 );
buf ( n75463 , n46875 );
not ( n75464 , n75463 );
buf ( n75465 , n66426 );
not ( n75466 , n75465 );
or ( n75467 , n75464 , n75466 );
buf ( n75468 , n13662 );
buf ( n75469 , n46887 );
nand ( n75470 , n75468 , n75469 );
buf ( n75471 , n75470 );
buf ( n75472 , n75471 );
nand ( n75473 , n75467 , n75472 );
buf ( n75474 , n75473 );
buf ( n75475 , n75474 );
buf ( n75476 , n46907 );
nand ( n75477 , n75475 , n75476 );
buf ( n75478 , n75477 );
buf ( n75479 , n75478 );
nand ( n75480 , n75462 , n75479 );
buf ( n75481 , n75480 );
buf ( n75482 , n75481 );
not ( n75483 , n75482 );
buf ( n75484 , n52780 );
buf ( n75485 , n41657 );
and ( n75486 , n75484 , n75485 );
not ( n75487 , n75484 );
buf ( n75488 , n61442 );
and ( n75489 , n75487 , n75488 );
nor ( n75490 , n75486 , n75489 );
buf ( n75491 , n75490 );
buf ( n75492 , n75491 );
not ( n75493 , n75492 );
buf ( n75494 , n75493 );
buf ( n75495 , n75494 );
not ( n75496 , n75495 );
buf ( n75497 , n61454 );
not ( n75498 , n75497 );
or ( n75499 , n75496 , n75498 );
buf ( n75500 , n73506 );
buf ( n75501 , n62582 );
nand ( n75502 , n75500 , n75501 );
buf ( n75503 , n75502 );
buf ( n75504 , n75503 );
nand ( n75505 , n75499 , n75504 );
buf ( n75506 , n75505 );
buf ( n75507 , n75506 );
not ( n75508 , n75507 );
or ( n75509 , n75483 , n75508 );
buf ( n75510 , n75506 );
buf ( n75511 , n75481 );
or ( n75512 , n75510 , n75511 );
xor ( n75513 , n73413 , n73467 );
xor ( n75514 , n75513 , n73489 );
buf ( n75515 , n75514 );
buf ( n75516 , n75515 );
nand ( n75517 , n75512 , n75516 );
buf ( n75518 , n75517 );
buf ( n75519 , n75518 );
nand ( n75520 , n75509 , n75519 );
buf ( n75521 , n75520 );
buf ( n75522 , n75521 );
xor ( n75523 , n73494 , n73531 );
xor ( n75524 , n75523 , n73559 );
buf ( n75525 , n75524 );
buf ( n75526 , n75525 );
xor ( n75527 , n75522 , n75526 );
buf ( n75528 , n56289 );
not ( n75529 , n75528 );
buf ( n75530 , n66463 );
not ( n75531 , n75530 );
or ( n75532 , n75529 , n75531 );
buf ( n75533 , n42366 );
buf ( n75534 , n52094 );
nand ( n75535 , n75533 , n75534 );
buf ( n75536 , n75535 );
buf ( n75537 , n75536 );
nand ( n75538 , n75532 , n75537 );
buf ( n75539 , n75538 );
buf ( n75540 , n75539 );
not ( n75541 , n75540 );
buf ( n75542 , n66459 );
not ( n75543 , n75542 );
or ( n75544 , n75541 , n75543 );
buf ( n75545 , n75246 );
buf ( n75546 , n66482 );
nand ( n75547 , n75545 , n75546 );
buf ( n75548 , n75547 );
buf ( n75549 , n75548 );
nand ( n75550 , n75544 , n75549 );
buf ( n75551 , n75550 );
buf ( n75552 , n75551 );
buf ( n75553 , n46912 );
not ( n75554 , n75553 );
buf ( n75555 , n75474 );
not ( n75556 , n75555 );
or ( n75557 , n75554 , n75556 );
buf ( n75558 , n46875 );
not ( n75559 , n75558 );
buf ( n75560 , n66470 );
not ( n75561 , n75560 );
or ( n75562 , n75559 , n75561 );
buf ( n75563 , n29463 );
buf ( n75564 , n46887 );
nand ( n75565 , n75563 , n75564 );
buf ( n75566 , n75565 );
buf ( n75567 , n75566 );
nand ( n75568 , n75562 , n75567 );
buf ( n75569 , n75568 );
buf ( n75570 , n75569 );
buf ( n75571 , n46907 );
nand ( n75572 , n75570 , n75571 );
buf ( n75573 , n75572 );
buf ( n75574 , n75573 );
nand ( n75575 , n75557 , n75574 );
buf ( n75576 , n75575 );
buf ( n75577 , n75576 );
xor ( n75578 , n75552 , n75577 );
xor ( n75579 , n75173 , n75195 );
xor ( n75580 , n75579 , n75221 );
buf ( n75581 , n75580 );
buf ( n75582 , n75581 );
and ( n75583 , n75578 , n75582 );
and ( n75584 , n75552 , n75577 );
or ( n75585 , n75583 , n75584 );
buf ( n75586 , n75585 );
buf ( n75587 , n75586 );
not ( n75588 , n75587 );
buf ( n75589 , n75588 );
not ( n75590 , n75589 );
buf ( n75591 , n48865 );
not ( n75592 , n75591 );
buf ( n75593 , n75383 );
not ( n75594 , n75593 );
or ( n75595 , n75592 , n75594 );
buf ( n75596 , n48808 );
not ( n75597 , n75596 );
buf ( n75598 , n63906 );
not ( n75599 , n75598 );
or ( n75600 , n75597 , n75599 );
buf ( n75601 , n13653 );
buf ( n75602 , n75377 );
nand ( n75603 , n75601 , n75602 );
buf ( n75604 , n75603 );
buf ( n75605 , n75604 );
nand ( n75606 , n75600 , n75605 );
buf ( n75607 , n75606 );
buf ( n75608 , n75607 );
buf ( n75609 , n48852 );
nand ( n75610 , n75608 , n75609 );
buf ( n75611 , n75610 );
buf ( n75612 , n75611 );
nand ( n75613 , n75595 , n75612 );
buf ( n75614 , n75613 );
nor ( n75615 , n75590 , n75614 );
buf ( n75616 , n48320 );
not ( n75617 , n75616 );
buf ( n75618 , n71123 );
not ( n75619 , n75618 );
or ( n75620 , n75617 , n75619 );
buf ( n75621 , n25290 );
not ( n75622 , n75621 );
buf ( n75623 , n71078 );
nand ( n75624 , n75622 , n75623 );
buf ( n75625 , n75624 );
buf ( n75626 , n75625 );
nand ( n75627 , n75620 , n75626 );
buf ( n75628 , n75627 );
buf ( n75629 , n75628 );
not ( n75630 , n75629 );
buf ( n75631 , n42246 );
not ( n75632 , n75631 );
or ( n75633 , n75630 , n75632 );
buf ( n75634 , n75160 );
buf ( n75635 , n42309 );
nand ( n75636 , n75634 , n75635 );
buf ( n75637 , n75636 );
buf ( n75638 , n75637 );
nand ( n75639 , n75633 , n75638 );
buf ( n75640 , n75639 );
buf ( n75641 , n75640 );
not ( n75642 , n75641 );
buf ( n75643 , n75642 );
buf ( n75644 , n75643 );
not ( n75645 , n75644 );
and ( n75646 , n50995 , n68606 );
not ( n75647 , n50995 );
and ( n75648 , n75647 , n42325 );
or ( n75649 , n75646 , n75648 );
buf ( n75650 , n75649 );
not ( n75651 , n75650 );
buf ( n75652 , n73163 );
not ( n75653 , n75652 );
or ( n75654 , n75651 , n75653 );
buf ( n75655 , n75208 );
buf ( n75656 , n42665 );
nand ( n75657 , n75655 , n75656 );
buf ( n75658 , n75657 );
buf ( n75659 , n75658 );
nand ( n75660 , n75654 , n75659 );
buf ( n75661 , n75660 );
buf ( n75662 , n75661 );
not ( n75663 , n75662 );
buf ( n75664 , n75663 );
buf ( n75665 , n75664 );
not ( n75666 , n75665 );
or ( n75667 , n75645 , n75666 );
xor ( n75668 , n74522 , n74548 );
xnor ( n75669 , n75668 , n74516 );
buf ( n75670 , n75669 );
not ( n75671 , n75670 );
buf ( n75672 , n75671 );
buf ( n75673 , n75672 );
nand ( n75674 , n75667 , n75673 );
buf ( n75675 , n75674 );
buf ( n75676 , n75675 );
buf ( n75677 , n75661 );
buf ( n75678 , n75640 );
nand ( n75679 , n75677 , n75678 );
buf ( n75680 , n75679 );
buf ( n75681 , n75680 );
nand ( n75682 , n75676 , n75681 );
buf ( n75683 , n75682 );
buf ( n75684 , n75683 );
not ( n75685 , n75684 );
buf ( n75686 , n75685 );
not ( n75687 , n75686 );
buf ( n75688 , n74477 );
buf ( n75689 , n74552 );
xor ( n75690 , n75688 , n75689 );
buf ( n75691 , n74561 );
xnor ( n75692 , n75690 , n75691 );
buf ( n75693 , n75692 );
not ( n75694 , n75693 );
and ( n75695 , n75687 , n75694 );
buf ( n75696 , n75686 );
buf ( n75697 , n75693 );
nand ( n75698 , n75696 , n75697 );
buf ( n75699 , n75698 );
xor ( n75700 , n74390 , n74394 );
xor ( n75701 , n75700 , n74399 );
buf ( n75702 , n75701 );
buf ( n75703 , n46114 );
not ( n75704 , n75703 );
buf ( n75705 , n74492 );
not ( n75706 , n75705 );
or ( n75707 , n75704 , n75706 );
buf ( n75708 , n25385 );
buf ( n75709 , n74414 );
nand ( n75710 , n75708 , n75709 );
buf ( n75711 , n75710 );
buf ( n75712 , n75711 );
nand ( n75713 , n75707 , n75712 );
buf ( n75714 , n75713 );
not ( n75715 , n75714 );
not ( n75716 , n74488 );
or ( n75717 , n75715 , n75716 );
buf ( n75718 , n74510 );
buf ( n75719 , n44496 );
nand ( n75720 , n75718 , n75719 );
buf ( n75721 , n75720 );
nand ( n75722 , n75717 , n75721 );
or ( n75723 , n75702 , n75722 );
xor ( n75724 , n74181 , n74198 );
xor ( n75725 , n75724 , n74221 );
buf ( n75726 , n75725 );
buf ( n75727 , n64068 );
buf ( n75728 , n64129 );
and ( n75729 , n75727 , n75728 );
buf ( n75730 , n66579 );
buf ( n75731 , n64133 );
and ( n75732 , n75730 , n75731 );
nor ( n75733 , n75729 , n75732 );
buf ( n75734 , n75733 );
buf ( n75735 , n75734 );
buf ( n75736 , n64141 );
or ( n75737 , n75735 , n75736 );
buf ( n75738 , n74249 );
buf ( n75739 , n63010 );
or ( n75740 , n75738 , n75739 );
nand ( n75741 , n75737 , n75740 );
buf ( n75742 , n75741 );
xor ( n75743 , n74131 , n74147 );
xor ( n75744 , n75743 , n74166 );
and ( n75745 , n75742 , n75744 );
buf ( n75746 , n1664 );
not ( n75747 , n75746 );
buf ( n75748 , n74215 );
not ( n75749 , n75748 );
buf ( n75750 , n75749 );
buf ( n75751 , n75750 );
not ( n75752 , n75751 );
or ( n75753 , n75747 , n75752 );
buf ( n75754 , n62782 );
buf ( n75755 , n66742 );
and ( n75756 , n75754 , n75755 );
buf ( n75757 , n62980 );
buf ( n75758 , n63000 );
and ( n75759 , n75757 , n75758 );
nor ( n75760 , n75756 , n75759 );
buf ( n75761 , n75760 );
buf ( n75762 , n75761 );
buf ( n75763 , n64230 );
or ( n75764 , n75762 , n75763 );
nand ( n75765 , n75753 , n75764 );
buf ( n75766 , n75765 );
xor ( n75767 , n74131 , n74147 );
xor ( n75768 , n75767 , n74166 );
and ( n75769 , n75766 , n75768 );
and ( n75770 , n75742 , n75766 );
or ( n75771 , n75745 , n75769 , n75770 );
xor ( n75772 , n75726 , n75771 );
xor ( n75773 , n74297 , n74342 );
xor ( n75774 , n75773 , n74362 );
buf ( n75775 , n75774 );
buf ( n75776 , n66690 );
buf ( n75777 , n62681 );
and ( n75778 , n75776 , n75777 );
buf ( n75779 , n66693 );
buf ( n75780 , n62663 );
and ( n75781 , n75779 , n75780 );
nor ( n75782 , n75778 , n75781 );
buf ( n75783 , n75782 );
buf ( n75784 , n75783 );
buf ( n75785 , n62935 );
or ( n75786 , n75784 , n75785 );
buf ( n75787 , n74266 );
buf ( n75788 , n62676 );
or ( n75789 , n75787 , n75788 );
nand ( n75790 , n75786 , n75789 );
buf ( n75791 , n75790 );
xor ( n75792 , n75775 , n75791 );
buf ( n75793 , n63013 );
not ( n75794 , n75793 );
buf ( n75795 , n64211 );
buf ( n75796 , n64129 );
and ( n75797 , n75795 , n75796 );
buf ( n75798 , n66610 );
buf ( n75799 , n64133 );
and ( n75800 , n75798 , n75799 );
nor ( n75801 , n75797 , n75800 );
buf ( n75802 , n75801 );
buf ( n75803 , n75802 );
not ( n75804 , n75803 );
buf ( n75805 , n75804 );
buf ( n75806 , n75805 );
not ( n75807 , n75806 );
or ( n75808 , n75794 , n75807 );
buf ( n75809 , n75734 );
buf ( n75810 , n63010 );
or ( n75811 , n75809 , n75810 );
nand ( n75812 , n75808 , n75811 );
buf ( n75813 , n75812 );
and ( n75814 , n75792 , n75813 );
and ( n75815 , n75775 , n75791 );
or ( n75816 , n75814 , n75815 );
buf ( n75817 , n75816 );
buf ( n75818 , n55129 );
buf ( n75819 , n623 );
not ( n75820 , n75819 );
buf ( n75821 , n75820 );
buf ( n75822 , n75821 );
nor ( n75823 , n75818 , n75822 );
buf ( n75824 , n75823 );
buf ( n75825 , n75824 );
buf ( n75826 , n56777 );
buf ( n75827 , n71307 );
and ( n75828 , n75826 , n75827 );
buf ( n75829 , n56804 );
buf ( n75830 , n71310 );
and ( n75831 , n75829 , n75830 );
nor ( n75832 , n75828 , n75831 );
buf ( n75833 , n75832 );
buf ( n75834 , n75833 );
buf ( n75835 , n56799 );
or ( n75836 , n75834 , n75835 );
buf ( n75837 , n71225 );
buf ( n75838 , n56777 );
and ( n75839 , n75837 , n75838 );
buf ( n75840 , n71228 );
buf ( n75841 , n56804 );
and ( n75842 , n75840 , n75841 );
nor ( n75843 , n75839 , n75842 );
buf ( n75844 , n75843 );
buf ( n75845 , n75844 );
buf ( n75846 , n58982 );
or ( n75847 , n75845 , n75846 );
nand ( n75848 , n75836 , n75847 );
buf ( n75849 , n75848 );
buf ( n75850 , n75849 );
and ( n75851 , n75825 , n75850 );
buf ( n75852 , n75851 );
buf ( n75853 , n75852 );
buf ( n75854 , n56799 );
buf ( n75855 , n75844 );
or ( n75856 , n75854 , n75855 );
buf ( n75857 , n74105 );
buf ( n75858 , n58982 );
or ( n75859 , n75857 , n75858 );
nand ( n75860 , n75856 , n75859 );
buf ( n75861 , n75860 );
buf ( n75862 , n75861 );
xor ( n75863 , n75853 , n75862 );
buf ( n75864 , n58887 );
not ( n75865 , n75864 );
buf ( n75866 , n74288 );
not ( n75867 , n75866 );
buf ( n75868 , n75867 );
buf ( n75869 , n75868 );
not ( n75870 , n75869 );
or ( n75871 , n75865 , n75870 );
buf ( n75872 , n70527 );
buf ( n75873 , n58897 );
and ( n75874 , n75872 , n75873 );
buf ( n75875 , n70530 );
buf ( n75876 , n58894 );
and ( n75877 , n75875 , n75876 );
nor ( n75878 , n75874 , n75877 );
buf ( n75879 , n75878 );
buf ( n75880 , n75879 );
buf ( n75881 , n58913 );
or ( n75882 , n75880 , n75881 );
nand ( n75883 , n75871 , n75882 );
buf ( n75884 , n75883 );
buf ( n75885 , n75884 );
and ( n75886 , n75863 , n75885 );
and ( n75887 , n75853 , n75862 );
or ( n75888 , n75886 , n75887 );
buf ( n75889 , n75888 );
xor ( n75890 , n74113 , n74125 );
xor ( n75891 , n75890 , n74128 );
and ( n75892 , n75889 , n75891 );
buf ( n75893 , n56626 );
buf ( n75894 , n16469 );
buf ( n75895 , n71818 );
and ( n75896 , n75894 , n75895 );
buf ( n75897 , n56631 );
buf ( n75898 , n71821 );
and ( n75899 , n75897 , n75898 );
nor ( n75900 , n75896 , n75899 );
buf ( n75901 , n75900 );
buf ( n75902 , n75901 );
or ( n75903 , n75893 , n75902 );
buf ( n75904 , n74329 );
buf ( n75905 , n56614 );
or ( n75906 , n75904 , n75905 );
nand ( n75907 , n75903 , n75906 );
buf ( n75908 , n75907 );
buf ( n75909 , n75908 );
buf ( n75910 , n56664 );
buf ( n75911 , n72427 );
buf ( n75912 , n74115 );
and ( n75913 , n75911 , n75912 );
buf ( n75914 , n55184 );
buf ( n75915 , n74118 );
and ( n75916 , n75914 , n75915 );
nor ( n75917 , n75913 , n75916 );
buf ( n75918 , n75917 );
buf ( n75919 , n75918 );
or ( n75920 , n75910 , n75919 );
buf ( n75921 , n74306 );
buf ( n75922 , n56673 );
or ( n75923 , n75921 , n75922 );
nand ( n75924 , n75920 , n75923 );
buf ( n75925 , n75924 );
buf ( n75926 , n75925 );
xor ( n75927 , n75909 , n75926 );
buf ( n75928 , n55156 );
buf ( n75929 , n623 );
and ( n75930 , n75928 , n75929 );
buf ( n75931 , n75930 );
buf ( n75932 , n75931 );
buf ( n75933 , n56799 );
buf ( n75934 , n56777 );
buf ( n75935 , n71801 );
and ( n75936 , n75934 , n75935 );
buf ( n75937 , n56804 );
buf ( n75938 , n71804 );
and ( n75939 , n75937 , n75938 );
nor ( n75940 , n75936 , n75939 );
buf ( n75941 , n75940 );
buf ( n75942 , n75941 );
or ( n75943 , n75933 , n75942 );
buf ( n75944 , n75833 );
buf ( n75945 , n56796 );
or ( n75946 , n75944 , n75945 );
nand ( n75947 , n75943 , n75946 );
buf ( n75948 , n75947 );
buf ( n75949 , n75948 );
and ( n75950 , n75932 , n75949 );
buf ( n75951 , n75950 );
buf ( n75952 , n75951 );
and ( n75953 , n75927 , n75952 );
and ( n75954 , n75909 , n75926 );
or ( n75955 , n75953 , n75954 );
buf ( n75956 , n75955 );
xor ( n75957 , n74314 , n74319 );
xor ( n75958 , n75957 , n74337 );
buf ( n75959 , n75958 );
xor ( n75960 , n75956 , n75959 );
buf ( n75961 , n60104 );
not ( n75962 , n75961 );
buf ( n75963 , n74356 );
not ( n75964 , n75963 );
buf ( n75965 , n75964 );
buf ( n75966 , n75965 );
not ( n75967 , n75966 );
or ( n75968 , n75962 , n75967 );
buf ( n75969 , n70333 );
buf ( n75970 , n60261 );
and ( n75971 , n75969 , n75970 );
buf ( n75972 , n70336 );
buf ( n75973 , n58880 );
and ( n75974 , n75972 , n75973 );
nor ( n75975 , n75971 , n75974 );
buf ( n75976 , n75975 );
buf ( n75977 , n75976 );
buf ( n75978 , n60270 );
or ( n75979 , n75977 , n75978 );
nand ( n75980 , n75968 , n75979 );
buf ( n75981 , n75980 );
and ( n75982 , n75960 , n75981 );
and ( n75983 , n75956 , n75959 );
or ( n75984 , n75982 , n75983 );
xor ( n75985 , n74113 , n74125 );
xor ( n75986 , n75985 , n74128 );
and ( n75987 , n75984 , n75986 );
and ( n75988 , n75889 , n75984 );
or ( n75989 , n75892 , n75987 , n75988 );
buf ( n75990 , n75989 );
xor ( n75991 , n75817 , n75990 );
xor ( n75992 , n74275 , n74279 );
xor ( n75993 , n75992 , n74367 );
buf ( n75994 , n75993 );
buf ( n75995 , n75994 );
and ( n75996 , n75991 , n75995 );
and ( n75997 , n75817 , n75990 );
or ( n75998 , n75996 , n75997 );
buf ( n75999 , n75998 );
and ( n76000 , n75772 , n75999 );
and ( n76001 , n75726 , n75771 );
or ( n76002 , n76000 , n76001 );
xor ( n76003 , n74241 , n74381 );
xor ( n76004 , n76003 , n74386 );
and ( n76005 , n76002 , n76004 );
xor ( n76006 , n74258 , n74372 );
xor ( n76007 , n76006 , n74377 );
buf ( n76008 , n76007 );
xor ( n76009 , n75726 , n75771 );
xor ( n76010 , n76009 , n75999 );
and ( n76011 , n76008 , n76010 );
xor ( n76012 , n74131 , n74147 );
xor ( n76013 , n76012 , n74166 );
xor ( n76014 , n75742 , n75766 );
xor ( n76015 , n76013 , n76014 );
buf ( n76016 , n62971 );
buf ( n76017 , n66742 );
and ( n76018 , n76016 , n76017 );
buf ( n76019 , n62974 );
buf ( n76020 , n63000 );
and ( n76021 , n76019 , n76020 );
nor ( n76022 , n76018 , n76021 );
buf ( n76023 , n76022 );
buf ( n76024 , n76023 );
buf ( n76025 , n64230 );
or ( n76026 , n76024 , n76025 );
buf ( n76027 , n75761 );
buf ( n76028 , n64227 );
or ( n76029 , n76027 , n76028 );
nand ( n76030 , n76026 , n76029 );
buf ( n76031 , n76030 );
buf ( n76032 , n76031 );
xor ( n76033 , n75853 , n75862 );
xor ( n76034 , n76033 , n75885 );
buf ( n76035 , n76034 );
buf ( n76036 , n76035 );
buf ( n76037 , n56786 );
buf ( n76038 , n71232 );
and ( n76039 , n76037 , n76038 );
not ( n76040 , n76037 );
buf ( n76041 , n71235 );
and ( n76042 , n76040 , n76041 );
nor ( n76043 , n76039 , n76042 );
buf ( n76044 , n76043 );
buf ( n76045 , n76044 );
not ( n76046 , n76045 );
buf ( n76047 , n76046 );
buf ( n76048 , n76047 );
buf ( n76049 , n58913 );
or ( n76050 , n76048 , n76049 );
buf ( n76051 , n75879 );
buf ( n76052 , n58884 );
or ( n76053 , n76051 , n76052 );
nand ( n76054 , n76050 , n76053 );
buf ( n76055 , n76054 );
buf ( n76056 , n76055 );
xor ( n76057 , n75825 , n75850 );
buf ( n76058 , n76057 );
buf ( n76059 , n76058 );
xor ( n76060 , n76056 , n76059 );
buf ( n76061 , n75918 );
buf ( n76062 , n55166 );
or ( n76063 , n76061 , n76062 );
buf ( n76064 , n55187 );
nand ( n76065 , n76063 , n76064 );
buf ( n76066 , n76065 );
buf ( n76067 , n76066 );
buf ( n76068 , n56626 );
buf ( n76069 , n56641 );
buf ( n76070 , n72445 );
and ( n76071 , n76069 , n76070 );
buf ( n76072 , n56631 );
buf ( n76073 , n72448 );
and ( n76074 , n76072 , n76073 );
nor ( n76075 , n76071 , n76074 );
buf ( n76076 , n76075 );
buf ( n76077 , n76076 );
or ( n76078 , n76068 , n76077 );
buf ( n76079 , n75901 );
buf ( n76080 , n56614 );
or ( n76081 , n76079 , n76080 );
nand ( n76082 , n76078 , n76081 );
buf ( n76083 , n76082 );
buf ( n76084 , n76083 );
xor ( n76085 , n76067 , n76084 );
buf ( n76086 , n58887 );
not ( n76087 , n76086 );
buf ( n76088 , n76044 );
not ( n76089 , n76088 );
or ( n76090 , n76087 , n76089 );
buf ( n76091 , n58913 );
buf ( n76092 , n56789 );
buf ( n76093 , n71225 );
and ( n76094 , n76092 , n76093 );
buf ( n76095 , n71228 );
buf ( n76096 , n56786 );
and ( n76097 , n76095 , n76096 );
nor ( n76098 , n76094 , n76097 );
buf ( n76099 , n76098 );
buf ( n76100 , n76099 );
or ( n76101 , n76091 , n76100 );
nand ( n76102 , n76090 , n76101 );
buf ( n76103 , n76102 );
buf ( n76104 , n76103 );
and ( n76105 , n76085 , n76104 );
and ( n76106 , n76067 , n76084 );
or ( n76107 , n76105 , n76106 );
buf ( n76108 , n76107 );
buf ( n76109 , n76108 );
and ( n76110 , n76060 , n76109 );
and ( n76111 , n76056 , n76059 );
or ( n76112 , n76110 , n76111 );
buf ( n76113 , n76112 );
buf ( n76114 , n76113 );
xor ( n76115 , n76036 , n76114 );
buf ( n76116 , n62679 );
not ( n76117 , n76116 );
buf ( n76118 , n68220 );
buf ( n76119 , n62663 );
or ( n76120 , n76118 , n76119 );
buf ( n76121 , n68217 );
buf ( n76122 , n62681 );
or ( n76123 , n76121 , n76122 );
nand ( n76124 , n76120 , n76123 );
buf ( n76125 , n76124 );
buf ( n76126 , n76125 );
not ( n76127 , n76126 );
or ( n76128 , n76117 , n76127 );
buf ( n76129 , n75783 );
buf ( n76130 , n62676 );
or ( n76131 , n76129 , n76130 );
nand ( n76132 , n76128 , n76131 );
buf ( n76133 , n76132 );
buf ( n76134 , n76133 );
and ( n76135 , n76115 , n76134 );
and ( n76136 , n76036 , n76114 );
or ( n76137 , n76135 , n76136 );
buf ( n76138 , n76137 );
buf ( n76139 , n76138 );
xor ( n76140 , n76032 , n76139 );
xor ( n76141 , n74113 , n74125 );
xor ( n76142 , n76141 , n74128 );
xor ( n76143 , n75889 , n75984 );
xor ( n76144 , n76142 , n76143 );
buf ( n76145 , n76144 );
and ( n76146 , n76140 , n76145 );
and ( n76147 , n76032 , n76139 );
or ( n76148 , n76146 , n76147 );
buf ( n76149 , n76148 );
xor ( n76150 , n76015 , n76149 );
xor ( n76151 , n75817 , n75990 );
xor ( n76152 , n76151 , n75995 );
buf ( n76153 , n76152 );
and ( n76154 , n76150 , n76153 );
and ( n76155 , n76015 , n76149 );
or ( n76156 , n76154 , n76155 );
xor ( n76157 , n75726 , n75771 );
xor ( n76158 , n76157 , n75999 );
and ( n76159 , n76156 , n76158 );
and ( n76160 , n76008 , n76156 );
or ( n76161 , n76011 , n76159 , n76160 );
xor ( n76162 , n74241 , n74381 );
xor ( n76163 , n76162 , n74386 );
and ( n76164 , n76161 , n76163 );
and ( n76165 , n76002 , n76161 );
or ( n76166 , n76005 , n76164 , n76165 );
nand ( n76167 , n75723 , n76166 );
nand ( n76168 , n75722 , n75702 );
nand ( n76169 , n76167 , n76168 );
buf ( n76170 , n76169 );
buf ( n76171 , n45746 );
not ( n76172 , n76171 );
buf ( n76173 , n72235 );
not ( n76174 , n76173 );
or ( n76175 , n76172 , n76174 );
buf ( n76176 , n42856 );
buf ( n76177 , n45746 );
not ( n76178 , n76177 );
buf ( n76179 , n76178 );
buf ( n76180 , n76179 );
nand ( n76181 , n76176 , n76180 );
buf ( n76182 , n76181 );
buf ( n76183 , n76182 );
nand ( n76184 , n76175 , n76183 );
buf ( n76185 , n76184 );
not ( n76186 , n76185 );
not ( n76187 , n71048 );
or ( n76188 , n76186 , n76187 );
or ( n76189 , n75186 , n45730 );
nand ( n76190 , n76188 , n76189 );
buf ( n76191 , n76190 );
xor ( n76192 , n76170 , n76191 );
buf ( n76193 , n47716 );
not ( n76194 , n76193 );
buf ( n76195 , n72240 );
not ( n76196 , n76195 );
or ( n76197 , n76194 , n76196 );
buf ( n76198 , n42228 );
buf ( n76199 , n47725 );
nand ( n76200 , n76198 , n76199 );
buf ( n76201 , n76200 );
buf ( n76202 , n76201 );
nand ( n76203 , n76197 , n76202 );
buf ( n76204 , n76203 );
buf ( n76205 , n76204 );
not ( n76206 , n76205 );
buf ( n76207 , n67354 );
not ( n76208 , n76207 );
or ( n76209 , n76206 , n76208 );
buf ( n76210 , n74540 );
buf ( n76211 , n41574 );
nand ( n76212 , n76210 , n76211 );
buf ( n76213 , n76212 );
buf ( n76214 , n76213 );
nand ( n76215 , n76209 , n76214 );
buf ( n76216 , n76215 );
buf ( n76217 , n76216 );
not ( n76218 , n75722 );
buf ( n76219 , n76166 );
buf ( n76220 , n75702 );
xnor ( n76221 , n76219 , n76220 );
buf ( n76222 , n76221 );
not ( n76223 , n76222 );
or ( n76224 , n76218 , n76223 );
or ( n76225 , n75722 , n76222 );
nand ( n76226 , n76224 , n76225 );
buf ( n76227 , n76226 );
xor ( n76228 , n76217 , n76227 );
buf ( n76229 , n67149 );
not ( n76230 , n76229 );
buf ( n76231 , n76185 );
not ( n76232 , n76231 );
or ( n76233 , n76230 , n76232 );
buf ( n76234 , n45746 );
not ( n76235 , n76234 );
buf ( n76236 , n74460 );
not ( n76237 , n76236 );
or ( n76238 , n76235 , n76237 );
buf ( n76239 , n42844 );
buf ( n76240 , n76179 );
nand ( n76241 , n76239 , n76240 );
buf ( n76242 , n76241 );
buf ( n76243 , n76242 );
nand ( n76244 , n76238 , n76243 );
buf ( n76245 , n76244 );
buf ( n76246 , n76245 );
buf ( n76247 , n71048 );
nand ( n76248 , n76246 , n76247 );
buf ( n76249 , n76248 );
buf ( n76250 , n76249 );
nand ( n76251 , n76233 , n76250 );
buf ( n76252 , n76251 );
buf ( n76253 , n76252 );
and ( n76254 , n76228 , n76253 );
and ( n76255 , n76217 , n76227 );
or ( n76256 , n76254 , n76255 );
buf ( n76257 , n76256 );
buf ( n76258 , n76257 );
and ( n76259 , n76192 , n76258 );
and ( n76260 , n76170 , n76191 );
or ( n76261 , n76259 , n76260 );
buf ( n76262 , n76261 );
and ( n76263 , n75699 , n76262 );
nor ( n76264 , n75695 , n76263 );
or ( n76265 , n75615 , n76264 );
nand ( n76266 , n75614 , n75586 );
nand ( n76267 , n76265 , n76266 );
buf ( n76268 , n76267 );
and ( n76269 , n75527 , n76268 );
and ( n76270 , n75522 , n75526 );
or ( n76271 , n76269 , n76270 );
buf ( n76272 , n76271 );
xor ( n76273 , n76272 , C0 );
xor ( n76274 , n73564 , n73602 );
xor ( n76275 , n76274 , n73643 );
buf ( n76276 , n76275 );
and ( n76277 , n76273 , n76276 );
or ( n76278 , n76277 , C0 );
buf ( n76279 , n76278 );
buf ( n76280 , C0 );
buf ( n76281 , n76280 );
buf ( n76282 , n62125 );
not ( n76283 , n76282 );
buf ( n76284 , n75295 );
not ( n76285 , n76284 );
or ( n76286 , n76283 , n76285 );
buf ( n76287 , n48836 );
buf ( n76288 , n47439 );
and ( n76289 , n76287 , n76288 );
not ( n76290 , n76287 );
buf ( n76291 , n47436 );
and ( n76292 , n76290 , n76291 );
nor ( n76293 , n76289 , n76292 );
buf ( n76294 , n76293 );
buf ( n76295 , n76294 );
buf ( n76296 , n51488 );
nand ( n76297 , n76295 , n76296 );
buf ( n76298 , n76297 );
buf ( n76299 , n76298 );
nand ( n76300 , n76286 , n76299 );
buf ( n76301 , n76300 );
buf ( n76302 , n76301 );
xor ( n76303 , n75144 , n75260 );
xor ( n76304 , n76303 , n75276 );
buf ( n76305 , n76304 );
xor ( n76306 , n76302 , n76305 );
buf ( n76307 , n42564 );
buf ( n76308 , n12481 );
nand ( n76309 , n76307 , n76308 );
buf ( n76310 , n76309 );
buf ( n76311 , n76310 );
not ( n76312 , n76311 );
buf ( n76313 , n55841 );
not ( n76314 , n76313 );
buf ( n76315 , n57599 );
not ( n76316 , n76315 );
or ( n76317 , n76314 , n76316 );
buf ( n76318 , n42560 );
buf ( n76319 , n58361 );
nand ( n76320 , n76318 , n76319 );
buf ( n76321 , n76320 );
buf ( n76322 , n76321 );
nand ( n76323 , n76317 , n76322 );
buf ( n76324 , n76323 );
buf ( n76325 , n76324 );
not ( n76326 , n76325 );
buf ( n76327 , n53628 );
not ( n76328 , n76327 );
or ( n76329 , n76326 , n76328 );
buf ( n76330 , n75345 );
buf ( n76331 , n53649 );
nand ( n76332 , n76330 , n76331 );
buf ( n76333 , n76332 );
buf ( n76334 , n76333 );
nand ( n76335 , n76329 , n76334 );
buf ( n76336 , n76335 );
buf ( n76337 , n76336 );
not ( n76338 , n76337 );
buf ( n76339 , n76338 );
buf ( n76340 , n76339 );
not ( n76341 , n76340 );
or ( n76342 , n76312 , n76341 );
xor ( n76343 , n75225 , n75231 );
xor ( n76344 , n76343 , n75258 );
buf ( n76345 , n76344 );
nand ( n76346 , n76342 , n76345 );
buf ( n76347 , n76346 );
buf ( n76348 , n76347 );
buf ( n76349 , n76310 );
not ( n76350 , n76349 );
buf ( n76351 , n76336 );
nand ( n76352 , n76350 , n76351 );
buf ( n76353 , n76352 );
buf ( n76354 , n76353 );
nand ( n76355 , n76348 , n76354 );
buf ( n76356 , n76355 );
buf ( n76357 , n76356 );
and ( n76358 , n76306 , n76357 );
and ( n76359 , n76302 , n76305 );
or ( n76360 , n76358 , n76359 );
buf ( n76361 , n76360 );
buf ( n76362 , n76361 );
xor ( n76363 , n76281 , n76362 );
xor ( n76364 , n75124 , n75280 );
xor ( n76365 , n76364 , n75306 );
buf ( n76366 , n76365 );
buf ( n76367 , n76366 );
and ( n76368 , n76363 , n76367 );
or ( n76369 , n76368 , C0 );
buf ( n76370 , n76369 );
buf ( n76371 , n76370 );
xor ( n76372 , n76279 , n76371 );
xor ( n76373 , n73876 , n74618 );
xor ( n76374 , n76373 , n73901 );
buf ( n76375 , n76374 );
and ( n76376 , n76372 , n76375 );
and ( n76377 , n76279 , n76371 );
or ( n76378 , n76376 , n76377 );
buf ( n76379 , n76378 );
buf ( n76380 , n76379 );
nand ( n76381 , n75457 , n76380 );
buf ( n76382 , n76381 );
buf ( n76383 , n76382 );
not ( n76384 , n76383 );
buf ( n76385 , n75446 );
not ( n76386 , n76385 );
buf ( n76387 , n76386 );
buf ( n76388 , n76387 );
buf ( n76389 , n75454 );
not ( n76390 , n76389 );
buf ( n76391 , n76390 );
buf ( n76392 , n76391 );
and ( n76393 , n76388 , n76392 );
buf ( n76394 , n76393 );
buf ( n76395 , n76394 );
nor ( n76396 , n76384 , n76395 );
buf ( n76397 , n76396 );
buf ( n76398 , n76397 );
not ( n76399 , n76398 );
buf ( n76400 , n76399 );
buf ( n76401 , n76400 );
nand ( n76402 , n75444 , n76401 );
buf ( n76403 , n76402 );
buf ( n76404 , n76403 );
buf ( n76405 , n75441 );
not ( n76406 , n76405 );
buf ( n76407 , n74639 );
nand ( n76408 , n76406 , n76407 );
buf ( n76409 , n76408 );
buf ( n76410 , n76409 );
nand ( n76411 , n76404 , n76410 );
buf ( n76412 , n76411 );
buf ( n76413 , n76412 );
buf ( n76414 , n67149 );
not ( n76415 , n76414 );
buf ( n76416 , n53492 );
not ( n76417 , n76416 );
buf ( n76418 , n47436 );
not ( n76419 , n76418 );
or ( n76420 , n76417 , n76419 );
buf ( n76421 , n50624 );
buf ( n76422 , n45747 );
nand ( n76423 , n76421 , n76422 );
buf ( n76424 , n76423 );
buf ( n76425 , n76424 );
nand ( n76426 , n76420 , n76425 );
buf ( n76427 , n76426 );
buf ( n76428 , n76427 );
not ( n76429 , n76428 );
or ( n76430 , n76415 , n76429 );
buf ( n76431 , n71029 );
buf ( n76432 , n71048 );
nand ( n76433 , n76431 , n76432 );
buf ( n76434 , n76433 );
buf ( n76435 , n76434 );
nand ( n76436 , n76430 , n76435 );
buf ( n76437 , n76436 );
buf ( n76438 , n76437 );
buf ( n76439 , n73248 );
not ( n76440 , n76439 );
buf ( n76441 , n42628 );
not ( n76442 , n76441 );
or ( n76443 , n76440 , n76442 );
buf ( n76444 , n50060 );
not ( n76445 , n76444 );
buf ( n76446 , n51804 );
not ( n76447 , n76446 );
or ( n76448 , n76445 , n76447 );
buf ( n76449 , n25159 );
buf ( n76450 , n67438 );
nand ( n76451 , n76449 , n76450 );
buf ( n76452 , n76451 );
buf ( n76453 , n76452 );
nand ( n76454 , n76448 , n76453 );
buf ( n76455 , n76454 );
buf ( n76456 , n76455 );
buf ( n76457 , n47872 );
nand ( n76458 , n76456 , n76457 );
buf ( n76459 , n76458 );
buf ( n76460 , n76459 );
nand ( n76461 , n76443 , n76460 );
buf ( n76462 , n76461 );
buf ( n76463 , n76462 );
xor ( n76464 , n76438 , n76463 );
buf ( n76465 , n73299 );
not ( n76466 , n76465 );
buf ( n76467 , n39999 );
not ( n76468 , n76467 );
or ( n76469 , n76466 , n76468 );
and ( n76470 , n52092 , n24092 );
not ( n76471 , n52092 );
and ( n76472 , n76471 , n50599 );
nor ( n76473 , n76470 , n76472 );
nand ( n76474 , n76473 , n48705 );
buf ( n76475 , n76474 );
nand ( n76476 , n76469 , n76475 );
buf ( n76477 , n76476 );
buf ( n76478 , n76477 );
xor ( n76479 , n76464 , n76478 );
buf ( n76480 , n76479 );
buf ( n76481 , n76480 );
buf ( n76482 , C0 );
buf ( n76483 , n76482 );
xor ( n76484 , n76481 , n76483 );
buf ( n76485 , n74949 );
not ( n76486 , n76485 );
buf ( n76487 , n74909 );
not ( n76488 , n76487 );
or ( n76489 , n76486 , n76488 );
buf ( n76490 , n74952 );
not ( n76491 , n76490 );
buf ( n76492 , n74912 );
not ( n76493 , n76492 );
or ( n76494 , n76491 , n76493 );
buf ( n76495 , n74885 );
nand ( n76496 , n76494 , n76495 );
buf ( n76497 , n76496 );
buf ( n76498 , n76497 );
nand ( n76499 , n76489 , n76498 );
buf ( n76500 , n76499 );
buf ( n76501 , n76500 );
xor ( n76502 , n76484 , n76501 );
buf ( n76503 , n76502 );
buf ( n76504 , n76503 );
buf ( n76505 , n74873 );
not ( n76506 , n76505 );
buf ( n76507 , n74959 );
nand ( n76508 , n76506 , n76507 );
buf ( n76509 , n76508 );
buf ( n76510 , n76509 );
buf ( n76511 , n74878 );
and ( n76512 , n76510 , n76511 );
buf ( n76513 , n74873 );
not ( n76514 , n76513 );
buf ( n76515 , n74959 );
nor ( n76516 , n76514 , n76515 );
buf ( n76517 , n76516 );
buf ( n76518 , n76517 );
nor ( n76519 , n76512 , n76518 );
buf ( n76520 , n76519 );
buf ( n76521 , n76520 );
not ( n76522 , n76521 );
buf ( n76523 , n76522 );
buf ( n76524 , n76523 );
xor ( n76525 , n76504 , n76524 );
buf ( n76526 , n74801 );
not ( n76527 , n76526 );
buf ( n76528 , n53628 );
not ( n76529 , n76528 );
or ( n76530 , n76527 , n76529 );
buf ( n76531 , n47716 );
not ( n76532 , n76531 );
buf ( n76533 , n52725 );
not ( n76534 , n76533 );
or ( n76535 , n76532 , n76534 );
buf ( n76536 , n61462 );
buf ( n76537 , n47713 );
nand ( n76538 , n76536 , n76537 );
buf ( n76539 , n76538 );
buf ( n76540 , n76539 );
nand ( n76541 , n76535 , n76540 );
buf ( n76542 , n76541 );
buf ( n76543 , n76542 );
buf ( n76544 , n43905 );
nand ( n76545 , n76543 , n76544 );
buf ( n76546 , n76545 );
buf ( n76547 , n76546 );
nand ( n76548 , n76530 , n76547 );
buf ( n76549 , n76548 );
buf ( n76550 , n44496 );
not ( n76551 , n76550 );
and ( n76552 , n29754 , n44530 );
not ( n76553 , n29754 );
and ( n76554 , n76553 , n65010 );
or ( n76555 , n76552 , n76554 );
buf ( n76556 , n76555 );
not ( n76557 , n76556 );
or ( n76558 , n76551 , n76557 );
buf ( n76559 , n74768 );
buf ( n76560 , n44517 );
nand ( n76561 , n76559 , n76560 );
buf ( n76562 , n76561 );
buf ( n76563 , n76562 );
nand ( n76564 , n76558 , n76563 );
buf ( n76565 , n76564 );
xor ( n76566 , n76549 , n76565 );
xor ( n76567 , n74684 , n74693 );
and ( n76568 , n76567 , n74720 );
and ( n76569 , n74684 , n74693 );
or ( n76570 , n76568 , n76569 );
buf ( n76571 , n76570 );
buf ( n76572 , n76571 );
buf ( n76573 , n74741 );
not ( n76574 , n76573 );
buf ( n76575 , n66459 );
not ( n76576 , n76575 );
or ( n76577 , n76574 , n76576 );
buf ( n76578 , n70886 );
buf ( n76579 , n66482 );
nand ( n76580 , n76578 , n76579 );
buf ( n76581 , n76580 );
buf ( n76582 , n76581 );
nand ( n76583 , n76577 , n76582 );
buf ( n76584 , n76583 );
buf ( n76585 , n76584 );
xor ( n76586 , n76572 , n76585 );
not ( n76587 , n70425 );
and ( n76588 , n70736 , n76587 );
not ( n76589 , n70739 );
and ( n76590 , n70736 , n76589 );
nor ( n76591 , n76588 , n76590 );
not ( n76592 , n70285 );
not ( n76593 , n70736 );
nand ( n76594 , n76592 , n76593 , n70424 );
not ( n76595 , n70424 );
nand ( n76596 , n76595 , n76593 , n70285 );
nand ( n76597 , n76591 , n76594 , n76596 );
buf ( n76598 , n74669 );
not ( n76599 , n76598 );
buf ( n76600 , n70268 );
not ( n76601 , n76600 );
or ( n76602 , n76599 , n76601 );
buf ( n76603 , n70264 );
buf ( n76604 , n42665 );
nand ( n76605 , n76603 , n76604 );
buf ( n76606 , n76605 );
buf ( n76607 , n76606 );
nand ( n76608 , n76602 , n76607 );
buf ( n76609 , n76608 );
xor ( n76610 , n76597 , n76609 );
buf ( n76611 , n42309 );
not ( n76612 , n76611 );
buf ( n76613 , n70865 );
not ( n76614 , n76613 );
or ( n76615 , n76612 , n76614 );
buf ( n76616 , n74709 );
buf ( n76617 , n42246 );
nand ( n76618 , n76616 , n76617 );
buf ( n76619 , n76618 );
buf ( n76620 , n76619 );
nand ( n76621 , n76615 , n76620 );
buf ( n76622 , n76621 );
xor ( n76623 , n76610 , n76622 );
buf ( n76624 , n76623 );
xnor ( n76625 , n76586 , n76624 );
buf ( n76626 , n76625 );
xnor ( n76627 , n76566 , n76626 );
buf ( n76628 , n76627 );
buf ( n76629 , n48855 );
not ( n76630 , n76629 );
buf ( n76631 , n74899 );
not ( n76632 , n76631 );
or ( n76633 , n76630 , n76632 );
buf ( n76634 , n48808 );
not ( n76635 , n76634 );
buf ( n76636 , n51250 );
not ( n76637 , n76636 );
or ( n76638 , n76635 , n76637 );
buf ( n76639 , n41822 );
buf ( n76640 , n72891 );
nand ( n76641 , n76639 , n76640 );
buf ( n76642 , n76641 );
buf ( n76643 , n76642 );
nand ( n76644 , n76638 , n76643 );
buf ( n76645 , n76644 );
buf ( n76646 , n76645 );
buf ( n76647 , n48868 );
nand ( n76648 , n76646 , n76647 );
buf ( n76649 , n76648 );
buf ( n76650 , n76649 );
nand ( n76651 , n76633 , n76650 );
buf ( n76652 , n76651 );
buf ( n76653 , n76652 );
xor ( n76654 , n76628 , n76653 );
xor ( n76655 , n71055 , n71074 );
and ( n76656 , n76655 , n72203 );
and ( n76657 , n71055 , n71074 );
or ( n76658 , n76656 , n76657 );
buf ( n76659 , n76658 );
buf ( n76660 , n76659 );
xor ( n76661 , n76654 , n76660 );
buf ( n76662 , n76661 );
buf ( n76663 , n76662 );
buf ( n76664 , C0 );
xor ( n76665 , n76663 , n76664 );
xor ( n76666 , n72206 , n72925 );
and ( n76667 , n76666 , n72957 );
and ( n76668 , n72206 , n72925 );
or ( n76669 , n76667 , n76668 );
buf ( n76670 , n76669 );
buf ( n76671 , n76670 );
xor ( n76672 , n76665 , n76671 );
buf ( n76673 , n76672 );
buf ( n76674 , n76673 );
xor ( n76675 , n76525 , n76674 );
buf ( n76676 , n76675 );
buf ( n76677 , n76676 );
buf ( n76678 , n74969 );
not ( n76679 , n76678 );
buf ( n76680 , n75090 );
not ( n76681 , n76680 );
or ( n76682 , n76679 , n76681 );
buf ( n76683 , n74972 );
not ( n76684 , n76683 );
buf ( n76685 , n75087 );
not ( n76686 , n76685 );
or ( n76687 , n76684 , n76686 );
buf ( n76688 , n75431 );
nand ( n76689 , n76687 , n76688 );
buf ( n76690 , n76689 );
buf ( n76691 , n76690 );
nand ( n76692 , n76682 , n76691 );
buf ( n76693 , n76692 );
buf ( n76694 , n76693 );
xor ( n76695 , n76677 , n76694 );
buf ( n76696 , n75077 );
not ( n76697 , n76696 );
or ( n76698 , C0 , n76697 );
buf ( n76699 , n75050 );
nand ( n76700 , n76698 , n76699 );
buf ( n76701 , n76700 );
buf ( n76702 , n76701 );
nand ( n76703 , C1 , n76702 );
buf ( n76704 , n76703 );
buf ( n76705 , n76704 );
xor ( n76706 , n72960 , n73311 );
and ( n76707 , n76706 , n74637 );
and ( n76708 , n72960 , n73311 );
or ( n76709 , n76707 , n76708 );
buf ( n76710 , n76709 );
buf ( n76711 , n76710 );
xor ( n76712 , n76705 , n76711 );
buf ( n76713 , n74942 );
not ( n76714 , n76713 );
buf ( n76715 , n47050 );
not ( n76716 , n76715 );
or ( n76717 , n76714 , n76716 );
buf ( n76718 , n53539 );
not ( n76719 , n76718 );
buf ( n76720 , n42471 );
not ( n76721 , n76720 );
or ( n76722 , n76719 , n76721 );
buf ( n76723 , n38979 );
buf ( n76724 , n53548 );
nand ( n76725 , n76723 , n76724 );
buf ( n76726 , n76725 );
buf ( n76727 , n76726 );
nand ( n76728 , n76722 , n76727 );
buf ( n76729 , n76728 );
buf ( n76730 , n76729 );
buf ( n76731 , n42448 );
nand ( n76732 , n76730 , n76731 );
buf ( n76733 , n76732 );
buf ( n76734 , n76733 );
nand ( n76735 , n76717 , n76734 );
buf ( n76736 , n76735 );
buf ( n76737 , n76736 );
buf ( n76738 , n74841 );
buf ( n76739 , n74850 );
or ( n76740 , n76738 , n76739 );
buf ( n76741 , n74857 );
nand ( n76742 , n76740 , n76741 );
buf ( n76743 , n76742 );
buf ( n76744 , n76743 );
buf ( n76745 , n74841 );
buf ( n76746 , n74850 );
nand ( n76747 , n76745 , n76746 );
buf ( n76748 , n76747 );
buf ( n76749 , n76748 );
nand ( n76750 , n76744 , n76749 );
buf ( n76751 , n76750 );
buf ( n76752 , n76751 );
buf ( n76753 , n43868 );
not ( n76754 , n76753 );
buf ( n76755 , n41605 );
not ( n76756 , n76755 );
buf ( n76757 , n60330 );
not ( n76758 , n76757 );
or ( n76759 , n76756 , n76758 );
buf ( n76760 , n60327 );
buf ( n76761 , n41604 );
nand ( n76762 , n76760 , n76761 );
buf ( n76763 , n76762 );
buf ( n76764 , n76763 );
nand ( n76765 , n76759 , n76764 );
buf ( n76766 , n76765 );
buf ( n76767 , n76766 );
not ( n76768 , n76767 );
or ( n76769 , n76754 , n76768 );
buf ( n76770 , n74848 );
not ( n76771 , n76770 );
buf ( n76772 , n41596 );
nand ( n76773 , n76771 , n76772 );
buf ( n76774 , n76773 );
buf ( n76775 , n76774 );
nand ( n76776 , n76769 , n76775 );
buf ( n76777 , n76776 );
buf ( n76778 , n76777 );
buf ( n76779 , n74834 );
not ( n76780 , n76779 );
buf ( n76781 , n61454 );
not ( n76782 , n76781 );
or ( n76783 , n76780 , n76782 );
buf ( n76784 , n46117 );
buf ( n76785 , n61442 );
and ( n76786 , n76784 , n76785 );
not ( n76787 , n76784 );
buf ( n76788 , n41657 );
and ( n76789 , n76787 , n76788 );
nor ( n76790 , n76786 , n76789 );
buf ( n76791 , n76790 );
buf ( n76792 , n76791 );
buf ( n76793 , n62582 );
nand ( n76794 , n76792 , n76793 );
buf ( n76795 , n76794 );
buf ( n76796 , n76795 );
nand ( n76797 , n76783 , n76796 );
buf ( n76798 , n76797 );
buf ( n76799 , n76798 );
xor ( n76800 , n76778 , n76799 );
xor ( n76801 , n74679 , n74723 );
and ( n76802 , n76801 , n74749 );
and ( n76803 , n74679 , n74723 );
or ( n76804 , n76802 , n76803 );
buf ( n76805 , n76804 );
buf ( n76806 , n76805 );
xor ( n76807 , n76800 , n76806 );
buf ( n76808 , n76807 );
buf ( n76809 , n76808 );
xor ( n76810 , n76752 , n76809 );
xor ( n76811 , n74650 , n74752 );
and ( n76812 , n76811 , n74774 );
and ( n76813 , n74650 , n74752 );
or ( n76814 , n76812 , n76813 );
buf ( n76815 , n76814 );
buf ( n76816 , n76815 );
xor ( n76817 , n76810 , n76816 );
buf ( n76818 , n76817 );
buf ( n76819 , n76818 );
xor ( n76820 , n76737 , n76819 );
buf ( n76821 , n72939 );
buf ( n76822 , n51489 );
or ( n76823 , n76821 , n76822 );
buf ( n76824 , n72931 );
buf ( n76825 , n41782 );
and ( n76826 , n76824 , n76825 );
not ( n76827 , n76824 );
buf ( n76828 , n41763 );
and ( n76829 , n76827 , n76828 );
nor ( n76830 , n76826 , n76829 );
buf ( n76831 , n76830 );
buf ( n76832 , n76831 );
buf ( n76833 , n51473 );
or ( n76834 , n76832 , n76833 );
nand ( n76835 , n76823 , n76834 );
buf ( n76836 , n76835 );
buf ( n76837 , n76836 );
xor ( n76838 , n76820 , n76837 );
buf ( n76839 , n76838 );
buf ( n76840 , n76839 );
and ( n76841 , n73231 , n73305 );
or ( n76842 , C0 , n76841 );
buf ( n76843 , n76842 );
buf ( n76844 , n76843 );
xor ( n76845 , n76840 , n76844 );
not ( n76846 , n73256 );
not ( n76847 , n73293 );
or ( n76848 , n76846 , n76847 );
nand ( n76849 , n76848 , n73303 );
not ( n76850 , n73293 );
nand ( n76851 , n76850 , n73255 );
nand ( n76852 , n76849 , n76851 );
buf ( n76853 , n76852 );
not ( n76854 , n76853 );
buf ( n76855 , n76854 );
and ( n76856 , n12481 , n46606 );
not ( n76857 , n74811 );
not ( n76858 , n74869 );
and ( n76859 , n76857 , n76858 );
buf ( n76860 , n74811 );
buf ( n76861 , n74869 );
nand ( n76862 , n76860 , n76861 );
buf ( n76863 , n76862 );
and ( n76864 , n76863 , n74816 );
nor ( n76865 , n76859 , n76864 );
xor ( n76866 , n76856 , n76865 );
buf ( n76867 , n73273 );
buf ( n76868 , n46907 );
and ( n76869 , n76867 , n76868 );
buf ( n76870 , n46875 );
not ( n76871 , n76870 );
buf ( n76872 , n41873 );
not ( n76873 , n76872 );
or ( n76874 , n76871 , n76873 );
buf ( n76875 , n50575 );
buf ( n76876 , n46887 );
nand ( n76877 , n76875 , n76876 );
buf ( n76878 , n76877 );
buf ( n76879 , n76878 );
nand ( n76880 , n76874 , n76879 );
buf ( n76881 , n76880 );
buf ( n76882 , n76881 );
buf ( n76883 , n46912 );
and ( n76884 , n76882 , n76883 );
nor ( n76885 , n76869 , n76884 );
buf ( n76886 , n76885 );
buf ( n76887 , n76886 );
xnor ( n76888 , n76866 , n76887 );
xor ( n76889 , n76855 , n76888 );
xor ( n76890 , n74777 , n74783 );
and ( n76891 , n76890 , n74871 );
and ( n76892 , n74777 , n74783 );
or ( n76893 , n76891 , n76892 );
buf ( n76894 , n76893 );
xor ( n76895 , n76889 , n76894 );
buf ( n76896 , n76895 );
xor ( n76897 , n76845 , n76896 );
buf ( n76898 , n76897 );
buf ( n76899 , n76898 );
xor ( n76900 , n76712 , n76899 );
buf ( n76901 , n76900 );
buf ( n76902 , n76901 );
xor ( n76903 , n76695 , n76902 );
buf ( n76904 , n76903 );
buf ( n76905 , n76904 );
xor ( n76906 , n76413 , n76905 );
buf ( n76907 , n56325 );
buf ( n76908 , n46356 );
and ( n76909 , n76907 , n76908 );
not ( n76910 , n76907 );
buf ( n76911 , n25160 );
and ( n76912 , n76910 , n76911 );
nor ( n76913 , n76909 , n76912 );
buf ( n76914 , n76913 );
buf ( n76915 , n76914 );
not ( n76916 , n76915 );
buf ( n76917 , n42628 );
not ( n76918 , n76917 );
or ( n76919 , n76916 , n76918 );
buf ( n76920 , n75319 );
buf ( n76921 , n42566 );
nand ( n76922 , n76920 , n76921 );
buf ( n76923 , n76922 );
buf ( n76924 , n76923 );
nand ( n76925 , n76919 , n76924 );
buf ( n76926 , n76925 );
buf ( n76927 , n76926 );
buf ( n76928 , C0 );
buf ( n76929 , n76928 );
xor ( n76930 , n76927 , n76929 );
xor ( n76931 , n75358 , n75362 );
xor ( n76932 , n76931 , n75391 );
buf ( n76933 , n76932 );
buf ( n76934 , n76933 );
and ( n76935 , n76930 , n76934 );
or ( n76936 , n76935 , C0 );
buf ( n76937 , n76936 );
buf ( n76938 , n76937 );
xor ( n76939 , n75333 , n75396 );
xor ( n76940 , n76939 , n75416 );
buf ( n76941 , n76940 );
buf ( n76942 , n76941 );
and ( n76943 , n76938 , n76942 );
not ( n76944 , n76938 );
buf ( n76945 , n76941 );
not ( n76946 , n76945 );
buf ( n76947 , n76946 );
buf ( n76948 , n76947 );
and ( n76949 , n76944 , n76948 );
nor ( n76950 , n76943 , n76949 );
buf ( n76951 , n76950 );
buf ( n76952 , n76951 );
buf ( n76953 , n60545 );
not ( n76954 , n76953 );
buf ( n76955 , n76294 );
not ( n76956 , n76955 );
or ( n76957 , n76954 , n76956 );
and ( n76958 , n48836 , n48169 );
not ( n76959 , n48836 );
and ( n76960 , n76959 , n28368 );
or ( n76961 , n76958 , n76960 );
buf ( n76962 , n76961 );
buf ( n76963 , n51488 );
nand ( n76964 , n76962 , n76963 );
buf ( n76965 , n76964 );
buf ( n76966 , n76965 );
nand ( n76967 , n76957 , n76966 );
buf ( n76968 , n76967 );
not ( n76969 , n76968 );
xor ( n76970 , n75481 , n75515 );
xor ( n76971 , n76970 , n75506 );
not ( n76972 , n76971 );
or ( n76973 , n76969 , n76972 );
buf ( n76974 , n76971 );
buf ( n76975 , n76968 );
or ( n76976 , n76974 , n76975 );
buf ( n76977 , n48356 );
buf ( n76978 , n41698 );
not ( n76979 , n76978 );
buf ( n76980 , n43895 );
nand ( n76981 , n76979 , n76980 );
buf ( n76982 , n76981 );
buf ( n76983 , n76982 );
buf ( n76984 , n12481 );
and ( n76985 , n76983 , n76984 );
buf ( n76986 , n61442 );
buf ( n76987 , n25028 );
and ( n76988 , n76986 , n76987 );
nor ( n76989 , n76985 , n76988 );
buf ( n76990 , n76989 );
buf ( n76991 , n76990 );
nand ( n76992 , n76977 , n76991 );
buf ( n76993 , n76992 );
buf ( n76994 , n76993 );
not ( n76995 , n76994 );
buf ( n76996 , n64410 );
buf ( n76997 , n76996 );
not ( n76998 , n76997 );
buf ( n76999 , n53548 );
buf ( n77000 , n61434 );
and ( n77001 , n76999 , n77000 );
not ( n77002 , n76999 );
buf ( n77003 , n58107 );
and ( n77004 , n77002 , n77003 );
nor ( n77005 , n77001 , n77004 );
buf ( n77006 , n77005 );
buf ( n77007 , n77006 );
not ( n77008 , n77007 );
and ( n77009 , n76998 , n77008 );
buf ( n77010 , n75491 );
buf ( n77011 , n41644 );
nor ( n77012 , n77010 , n77011 );
buf ( n77013 , n77012 );
buf ( n77014 , n77013 );
nor ( n77015 , n77009 , n77014 );
buf ( n77016 , n77015 );
buf ( n77017 , n77016 );
not ( n77018 , n77017 );
or ( n77019 , n76995 , n77018 );
buf ( n77020 , n46912 );
not ( n77021 , n77020 );
buf ( n77022 , n75569 );
not ( n77023 , n77022 );
or ( n77024 , n77021 , n77023 );
and ( n77025 , n28430 , n46887 );
not ( n77026 , n28430 );
and ( n77027 , n77026 , n46875 );
or ( n77028 , n77025 , n77027 );
buf ( n77029 , n77028 );
buf ( n77030 , n46907 );
nand ( n77031 , n77029 , n77030 );
buf ( n77032 , n77031 );
buf ( n77033 , n77032 );
nand ( n77034 , n77024 , n77033 );
buf ( n77035 , n77034 );
buf ( n77036 , n77035 );
xor ( n77037 , n76170 , n76191 );
xor ( n77038 , n77037 , n76258 );
buf ( n77039 , n77038 );
buf ( n77040 , n77039 );
xor ( n77041 , n77036 , n77040 );
xor ( n77042 , n74241 , n74381 );
xor ( n77043 , n77042 , n74386 );
xor ( n77044 , n76002 , n76161 );
xor ( n77045 , n77043 , n77044 );
buf ( n77046 , n77045 );
buf ( n77047 , n46390 );
not ( n77048 , n77047 );
buf ( n77049 , n44527 );
not ( n77050 , n77049 );
or ( n77051 , n77048 , n77050 );
buf ( n77052 , n41570 );
buf ( n77053 , n46387 );
nand ( n77054 , n77052 , n77053 );
buf ( n77055 , n77054 );
buf ( n77056 , n77055 );
nand ( n77057 , n77051 , n77056 );
buf ( n77058 , n77057 );
buf ( n77059 , n77058 );
not ( n77060 , n77059 );
buf ( n77061 , n74488 );
not ( n77062 , n77061 );
or ( n77063 , n77060 , n77062 );
buf ( n77064 , n75714 );
buf ( n77065 , n44496 );
nand ( n77066 , n77064 , n77065 );
buf ( n77067 , n77066 );
buf ( n77068 , n77067 );
nand ( n77069 , n77063 , n77068 );
buf ( n77070 , n77069 );
buf ( n77071 , n77070 );
xor ( n77072 , n77046 , n77071 );
buf ( n77073 , n71078 );
not ( n77074 , n77073 );
buf ( n77075 , n42228 );
not ( n77076 , n77075 );
buf ( n77077 , n77076 );
buf ( n77078 , n77077 );
not ( n77079 , n77078 );
or ( n77080 , n77074 , n77079 );
buf ( n77081 , n74530 );
not ( n77082 , n77081 );
buf ( n77083 , n48320 );
nand ( n77084 , n77082 , n77083 );
buf ( n77085 , n77084 );
buf ( n77086 , n77085 );
nand ( n77087 , n77080 , n77086 );
buf ( n77088 , n77087 );
buf ( n77089 , n77088 );
not ( n77090 , n77089 );
buf ( n77091 , n67354 );
not ( n77092 , n77091 );
or ( n77093 , n77090 , n77092 );
buf ( n77094 , n76204 );
buf ( n77095 , n41574 );
nand ( n77096 , n77094 , n77095 );
buf ( n77097 , n77096 );
buf ( n77098 , n77097 );
nand ( n77099 , n77093 , n77098 );
buf ( n77100 , n77099 );
buf ( n77101 , n77100 );
and ( n77102 , n77072 , n77101 );
and ( n77103 , n77046 , n77071 );
or ( n77104 , n77102 , n77103 );
buf ( n77105 , n77104 );
buf ( n77106 , n77105 );
and ( n77107 , n50060 , n42257 );
not ( n77108 , n50060 );
and ( n77109 , n77108 , n25290 );
or ( n77110 , n77107 , n77109 );
buf ( n77111 , n77110 );
not ( n77112 , n77111 );
buf ( n77113 , n42246 );
not ( n77114 , n77113 );
or ( n77115 , n77112 , n77114 );
buf ( n77116 , n75628 );
buf ( n77117 , n42309 );
nand ( n77118 , n77116 , n77117 );
buf ( n77119 , n77118 );
buf ( n77120 , n77119 );
nand ( n77121 , n77115 , n77120 );
buf ( n77122 , n77121 );
buf ( n77123 , n77122 );
xor ( n77124 , n77106 , n77123 );
buf ( n77125 , n46912 );
not ( n77126 , n77125 );
buf ( n77127 , n77028 );
not ( n77128 , n77127 );
or ( n77129 , n77126 , n77128 );
buf ( n77130 , n46875 );
not ( n77131 , n77130 );
buf ( n77132 , n72213 );
not ( n77133 , n77132 );
or ( n77134 , n77131 , n77133 );
buf ( n77135 , n72776 );
buf ( n77136 , n46887 );
nand ( n77137 , n77135 , n77136 );
buf ( n77138 , n77137 );
buf ( n77139 , n77138 );
nand ( n77140 , n77134 , n77139 );
buf ( n77141 , n77140 );
buf ( n77142 , n77141 );
buf ( n77143 , n46907 );
nand ( n77144 , n77142 , n77143 );
buf ( n77145 , n77144 );
buf ( n77146 , n77145 );
nand ( n77147 , n77129 , n77146 );
buf ( n77148 , n77147 );
buf ( n77149 , n77148 );
and ( n77150 , n77124 , n77149 );
and ( n77151 , n77106 , n77123 );
or ( n77152 , n77150 , n77151 );
buf ( n77153 , n77152 );
buf ( n77154 , n77153 );
and ( n77155 , n77041 , n77154 );
and ( n77156 , n77036 , n77040 );
or ( n77157 , n77155 , n77156 );
buf ( n77158 , n77157 );
buf ( n77159 , n77158 );
nand ( n77160 , n77019 , n77159 );
buf ( n77161 , n77160 );
buf ( n77162 , n77161 );
buf ( n77163 , n76993 );
not ( n77164 , n77163 );
buf ( n77165 , n77164 );
buf ( n77166 , n77165 );
buf ( n77167 , n77016 );
not ( n77168 , n77167 );
buf ( n77169 , n77168 );
buf ( n77170 , n77169 );
nand ( n77171 , n77166 , n77170 );
buf ( n77172 , n77171 );
buf ( n77173 , n77172 );
nand ( n77174 , n77162 , n77173 );
buf ( n77175 , n77174 );
buf ( n77176 , n77175 );
nand ( n77177 , n76976 , n77176 );
buf ( n77178 , n77177 );
nand ( n77179 , n76973 , n77178 );
not ( n77180 , n77179 );
not ( n77181 , n77180 );
or ( n77182 , n77181 , C0 );
buf ( n77183 , n76264 );
not ( n77184 , n77183 );
buf ( n77185 , n75614 );
not ( n77186 , n77185 );
or ( n77187 , n77184 , n77186 );
buf ( n77188 , n75614 );
buf ( n77189 , n76264 );
or ( n77190 , n77188 , n77189 );
nand ( n77191 , n77187 , n77190 );
buf ( n77192 , n77191 );
buf ( n77193 , n77192 );
not ( n77194 , n77193 );
buf ( n77195 , n75589 );
not ( n77196 , n77195 );
and ( n77197 , n77194 , n77196 );
buf ( n77198 , n77192 );
buf ( n77199 , n75589 );
and ( n77200 , n77198 , n77199 );
nor ( n77201 , n77197 , n77200 );
buf ( n77202 , n77201 );
buf ( n77203 , n77202 );
not ( n77204 , n77203 );
buf ( n77205 , n77204 );
buf ( n77206 , C0 );
buf ( n77207 , n77206 );
buf ( n77208 , n77205 );
or ( n77209 , n77207 , n77208 );
buf ( n77210 , n75683 );
not ( n77211 , n77210 );
buf ( n77212 , n76262 );
not ( n77213 , n77212 );
buf ( n77214 , n75693 );
not ( n77215 , n77214 );
and ( n77216 , n77213 , n77215 );
buf ( n77217 , n75693 );
buf ( n77218 , n76262 );
and ( n77219 , n77217 , n77218 );
nor ( n77220 , n77216 , n77219 );
buf ( n77221 , n77220 );
buf ( n77222 , n77221 );
not ( n77223 , n77222 );
or ( n77224 , n77211 , n77223 );
buf ( n77225 , n75683 );
buf ( n77226 , n77221 );
or ( n77227 , n77225 , n77226 );
nand ( n77228 , n77224 , n77227 );
buf ( n77229 , n77228 );
buf ( n77230 , n77229 );
buf ( n77231 , n48865 );
not ( n77232 , n77231 );
buf ( n77233 , n75607 );
not ( n77234 , n77233 );
or ( n77235 , n77232 , n77234 );
buf ( n77236 , n48808 );
not ( n77237 , n77236 );
buf ( n77238 , n60330 );
not ( n77239 , n77238 );
or ( n77240 , n77237 , n77239 );
buf ( n77241 , n60327 );
buf ( n77242 , n75377 );
nand ( n77243 , n77241 , n77242 );
buf ( n77244 , n77243 );
buf ( n77245 , n77244 );
nand ( n77246 , n77240 , n77245 );
buf ( n77247 , n77246 );
buf ( n77248 , n77247 );
buf ( n77249 , n48852 );
nand ( n77250 , n77248 , n77249 );
buf ( n77251 , n77250 );
buf ( n77252 , n77251 );
nand ( n77253 , n77235 , n77252 );
buf ( n77254 , n77253 );
buf ( n77255 , n77254 );
xor ( n77256 , n77230 , n77255 );
buf ( n77257 , n75661 );
not ( n77258 , n77257 );
buf ( n77259 , n75669 );
not ( n77260 , n77259 );
buf ( n77261 , n75640 );
not ( n77262 , n77261 );
and ( n77263 , n77260 , n77262 );
buf ( n77264 , n75669 );
buf ( n77265 , n75640 );
and ( n77266 , n77264 , n77265 );
nor ( n77267 , n77263 , n77266 );
buf ( n77268 , n77267 );
buf ( n77269 , n77268 );
not ( n77270 , n77269 );
and ( n77271 , n77258 , n77270 );
buf ( n77272 , n75661 );
buf ( n77273 , n77268 );
and ( n77274 , n77272 , n77273 );
nor ( n77275 , n77271 , n77274 );
buf ( n77276 , n77275 );
buf ( n77277 , n77276 );
not ( n77278 , n77277 );
buf ( n77279 , n77278 );
buf ( n77280 , n77279 );
not ( n77281 , n77280 );
buf ( n77282 , n52780 );
not ( n77283 , n77282 );
buf ( n77284 , n66463 );
not ( n77285 , n77284 );
or ( n77286 , n77283 , n77285 );
buf ( n77287 , n68062 );
buf ( n77288 , n52789 );
nand ( n77289 , n77287 , n77288 );
buf ( n77290 , n77289 );
buf ( n77291 , n77290 );
nand ( n77292 , n77286 , n77291 );
buf ( n77293 , n77292 );
buf ( n77294 , n77293 );
not ( n77295 , n77294 );
buf ( n77296 , n66459 );
not ( n77297 , n77296 );
or ( n77298 , n77295 , n77297 );
buf ( n77299 , n42333 );
not ( n77300 , n77299 );
buf ( n77301 , n75539 );
nand ( n77302 , n77300 , n77301 );
buf ( n77303 , n77302 );
buf ( n77304 , n77303 );
nand ( n77305 , n77298 , n77304 );
buf ( n77306 , n77305 );
buf ( n77307 , n77306 );
not ( n77308 , n77307 );
or ( n77309 , n77281 , n77308 );
buf ( n77310 , n77306 );
buf ( n77311 , n77279 );
or ( n77312 , n77310 , n77311 );
xor ( n77313 , n76217 , n76227 );
xor ( n77314 , n77313 , n76253 );
buf ( n77315 , n77314 );
buf ( n77316 , n77315 );
buf ( n77317 , n67149 );
not ( n77318 , n77317 );
buf ( n77319 , n76245 );
not ( n77320 , n77319 );
or ( n77321 , n77318 , n77320 );
buf ( n77322 , n45746 );
not ( n77323 , n77322 );
buf ( n77324 , n44946 );
not ( n77325 , n77324 );
or ( n77326 , n77323 , n77325 );
buf ( n77327 , n74500 );
buf ( n77328 , n45747 );
nand ( n77329 , n77327 , n77328 );
buf ( n77330 , n77329 );
buf ( n77331 , n77330 );
nand ( n77332 , n77326 , n77331 );
buf ( n77333 , n77332 );
buf ( n77334 , n77333 );
buf ( n77335 , n71048 );
nand ( n77336 , n77334 , n77335 );
buf ( n77337 , n77336 );
buf ( n77338 , n77337 );
nand ( n77339 , n77321 , n77338 );
buf ( n77340 , n77339 );
buf ( n77341 , n77340 );
not ( n77342 , n77341 );
buf ( n77343 , n67149 );
not ( n77344 , n77343 );
buf ( n77345 , n77333 );
not ( n77346 , n77345 );
or ( n77347 , n77344 , n77346 );
buf ( n77348 , n45746 );
not ( n77349 , n77348 );
buf ( n77350 , n74414 );
not ( n77351 , n77350 );
or ( n77352 , n77349 , n77351 );
buf ( n77353 , n74417 );
buf ( n77354 , n45747 );
nand ( n77355 , n77353 , n77354 );
buf ( n77356 , n77355 );
buf ( n77357 , n77356 );
nand ( n77358 , n77352 , n77357 );
buf ( n77359 , n77358 );
buf ( n77360 , n77359 );
buf ( n77361 , n71048 );
nand ( n77362 , n77360 , n77361 );
buf ( n77363 , n77362 );
buf ( n77364 , n77363 );
nand ( n77365 , n77347 , n77364 );
buf ( n77366 , n77365 );
buf ( n77367 , n77366 );
xor ( n77368 , n75726 , n75771 );
xor ( n77369 , n77368 , n75999 );
xor ( n77370 , n76008 , n76156 );
xor ( n77371 , n77369 , n77370 );
buf ( n77372 , n77371 );
or ( n77373 , n77367 , n77372 );
buf ( n77374 , n66601 );
buf ( n77375 , n64129 );
and ( n77376 , n77374 , n77375 );
buf ( n77377 , n66604 );
buf ( n77378 , n64133 );
and ( n77379 , n77377 , n77378 );
nor ( n77380 , n77376 , n77379 );
buf ( n77381 , n77380 );
buf ( n77382 , n77381 );
buf ( n77383 , n64141 );
or ( n77384 , n77382 , n77383 );
buf ( n77385 , n75802 );
buf ( n77386 , n63010 );
or ( n77387 , n77385 , n77386 );
nand ( n77388 , n77384 , n77387 );
buf ( n77389 , n77388 );
xor ( n77390 , n75956 , n75959 );
xor ( n77391 , n77390 , n75981 );
and ( n77392 , n77389 , n77391 );
xor ( n77393 , n75909 , n75926 );
xor ( n77394 , n77393 , n75952 );
buf ( n77395 , n77394 );
buf ( n77396 , n70348 );
buf ( n77397 , n60261 );
and ( n77398 , n77396 , n77397 );
buf ( n77399 , n70351 );
buf ( n77400 , n60090 );
and ( n77401 , n77399 , n77400 );
nor ( n77402 , n77398 , n77401 );
buf ( n77403 , n77402 );
buf ( n77404 , n77403 );
buf ( n77405 , n60270 );
or ( n77406 , n77404 , n77405 );
buf ( n77407 , n75976 );
buf ( n77408 , n60100 );
or ( n77409 , n77407 , n77408 );
nand ( n77410 , n77406 , n77409 );
buf ( n77411 , n77410 );
xor ( n77412 , n77395 , n77411 );
buf ( n77413 , n62691 );
not ( n77414 , n77413 );
buf ( n77415 , n76125 );
not ( n77416 , n77415 );
or ( n77417 , n77414 , n77416 );
buf ( n77418 , n68235 );
buf ( n77419 , n62684 );
or ( n77420 , n77418 , n77419 );
buf ( n77421 , n68232 );
buf ( n77422 , n60096 );
or ( n77423 , n77421 , n77422 );
nand ( n77424 , n77420 , n77423 );
buf ( n77425 , n77424 );
buf ( n77426 , n77425 );
not ( n77427 , n77426 );
buf ( n77428 , n77427 );
buf ( n77429 , n77428 );
buf ( n77430 , n62935 );
or ( n77431 , n77429 , n77430 );
nand ( n77432 , n77417 , n77431 );
buf ( n77433 , n77432 );
and ( n77434 , n77412 , n77433 );
and ( n77435 , n77395 , n77411 );
or ( n77436 , n77434 , n77435 );
xor ( n77437 , n75956 , n75959 );
xor ( n77438 , n77437 , n75981 );
and ( n77439 , n77436 , n77438 );
and ( n77440 , n77389 , n77436 );
or ( n77441 , n77392 , n77439 , n77440 );
xor ( n77442 , n75775 , n75791 );
xor ( n77443 , n77442 , n75813 );
and ( n77444 , n77441 , n77443 );
xor ( n77445 , n76056 , n76059 );
xor ( n77446 , n77445 , n76109 );
buf ( n77447 , n77446 );
buf ( n77448 , n58913 );
buf ( n77449 , n56789 );
buf ( n77450 , n71307 );
and ( n77451 , n77449 , n77450 );
buf ( n77452 , n56786 );
buf ( n77453 , n71310 );
and ( n77454 , n77452 , n77453 );
nor ( n77455 , n77451 , n77454 );
buf ( n77456 , n77455 );
buf ( n77457 , n77456 );
or ( n77458 , n77448 , n77457 );
buf ( n77459 , n76099 );
buf ( n77460 , n58884 );
or ( n77461 , n77459 , n77460 );
nand ( n77462 , n77458 , n77461 );
buf ( n77463 , n77462 );
buf ( n77464 , n55162 );
buf ( n77465 , n623 );
and ( n77466 , n77464 , n77465 );
buf ( n77467 , n55162 );
not ( n77468 , n77467 );
buf ( n77469 , n77468 );
buf ( n77470 , n77469 );
buf ( n77471 , n75821 );
and ( n77472 , n77470 , n77471 );
buf ( n77473 , n16469 );
nor ( n77474 , n77472 , n77473 );
buf ( n77475 , n77474 );
buf ( n77476 , n77475 );
buf ( n77477 , n55118 );
nor ( n77478 , n77466 , n77476 , n77477 );
buf ( n77479 , n77478 );
xor ( n77480 , n77463 , n77479 );
buf ( n77481 , n56799 );
buf ( n77482 , n56777 );
buf ( n77483 , n71818 );
and ( n77484 , n77482 , n77483 );
buf ( n77485 , n56804 );
buf ( n77486 , n71821 );
and ( n77487 , n77485 , n77486 );
nor ( n77488 , n77484 , n77487 );
buf ( n77489 , n77488 );
buf ( n77490 , n77489 );
or ( n77491 , n77481 , n77490 );
buf ( n77492 , n75941 );
buf ( n77493 , n58982 );
or ( n77494 , n77492 , n77493 );
nand ( n77495 , n77491 , n77494 );
buf ( n77496 , n77495 );
and ( n77497 , n77480 , n77496 );
and ( n77498 , n77463 , n77479 );
or ( n77499 , n77497 , n77498 );
buf ( n77500 , n77499 );
xor ( n77501 , n75932 , n75949 );
buf ( n77502 , n77501 );
buf ( n77503 , n77502 );
xor ( n77504 , n77500 , n77503 );
buf ( n77505 , n60101 );
not ( n77506 , n77505 );
buf ( n77507 , n70527 );
buf ( n77508 , n15265 );
and ( n77509 , n77507 , n77508 );
buf ( n77510 , n70530 );
buf ( n77511 , n60090 );
and ( n77512 , n77510 , n77511 );
nor ( n77513 , n77509 , n77512 );
buf ( n77514 , n77513 );
buf ( n77515 , n77514 );
not ( n77516 , n77515 );
buf ( n77517 , n77516 );
buf ( n77518 , n77517 );
not ( n77519 , n77518 );
or ( n77520 , n77506 , n77519 );
buf ( n77521 , n77403 );
buf ( n77522 , n60100 );
or ( n77523 , n77521 , n77522 );
nand ( n77524 , n77520 , n77523 );
buf ( n77525 , n77524 );
buf ( n77526 , n77525 );
and ( n77527 , n77504 , n77526 );
and ( n77528 , n77500 , n77503 );
or ( n77529 , n77527 , n77528 );
buf ( n77530 , n77529 );
xor ( n77531 , n77447 , n77530 );
buf ( n77532 , n63022 );
not ( n77533 , n77532 );
buf ( n77534 , n77381 );
not ( n77535 , n77534 );
buf ( n77536 , n77535 );
buf ( n77537 , n77536 );
not ( n77538 , n77537 );
or ( n77539 , n77533 , n77538 );
buf ( n77540 , n66690 );
buf ( n77541 , n64129 );
and ( n77542 , n77540 , n77541 );
buf ( n77543 , n66693 );
buf ( n77544 , n64133 );
and ( n77545 , n77543 , n77544 );
nor ( n77546 , n77542 , n77545 );
buf ( n77547 , n77546 );
buf ( n77548 , n77547 );
buf ( n77549 , n64141 );
or ( n77550 , n77548 , n77549 );
nand ( n77551 , n77539 , n77550 );
buf ( n77552 , n77551 );
and ( n77553 , n77531 , n77552 );
and ( n77554 , n77447 , n77530 );
or ( n77555 , n77553 , n77554 );
buf ( n77556 , n77555 );
buf ( n77557 , n64068 );
buf ( n77558 , n66742 );
and ( n77559 , n77557 , n77558 );
buf ( n77560 , n66579 );
buf ( n77561 , n63000 );
and ( n77562 , n77560 , n77561 );
nor ( n77563 , n77559 , n77562 );
buf ( n77564 , n77563 );
buf ( n77565 , n77564 );
buf ( n77566 , n64230 );
or ( n77567 , n77565 , n77566 );
buf ( n77568 , n76023 );
buf ( n77569 , n64227 );
or ( n77570 , n77568 , n77569 );
nand ( n77571 , n77567 , n77570 );
buf ( n77572 , n77571 );
buf ( n77573 , n77572 );
xor ( n77574 , n77556 , n77573 );
xor ( n77575 , n76036 , n76114 );
xor ( n77576 , n77575 , n76134 );
buf ( n77577 , n77576 );
buf ( n77578 , n77577 );
and ( n77579 , n77574 , n77578 );
and ( n77580 , n77556 , n77573 );
or ( n77581 , n77579 , n77580 );
buf ( n77582 , n77581 );
xor ( n77583 , n75775 , n75791 );
xor ( n77584 , n77583 , n75813 );
and ( n77585 , n77582 , n77584 );
and ( n77586 , n77441 , n77582 );
or ( n77587 , n77444 , n77585 , n77586 );
xor ( n77588 , n76015 , n76149 );
xor ( n77589 , n77588 , n76153 );
and ( n77590 , n77587 , n77589 );
xor ( n77591 , n75956 , n75959 );
xor ( n77592 , n77591 , n75981 );
xor ( n77593 , n77389 , n77436 );
xor ( n77594 , n77592 , n77593 );
buf ( n77595 , n55187 );
buf ( n77596 , n623 );
or ( n77597 , n77595 , n77596 );
buf ( n77598 , n55180 );
buf ( n77599 , n72427 );
buf ( n77600 , n623 );
and ( n77601 , n77598 , n77599 , n77600 );
buf ( n77602 , n55170 );
nor ( n77603 , n77601 , n77602 );
buf ( n77604 , n77603 );
buf ( n77605 , n77604 );
nand ( n77606 , n77597 , n77605 );
buf ( n77607 , n77606 );
buf ( n77608 , n56626 );
buf ( n77609 , n16469 );
buf ( n77610 , n74115 );
and ( n77611 , n77609 , n77610 );
buf ( n77612 , n16472 );
buf ( n77613 , n74118 );
and ( n77614 , n77612 , n77613 );
nor ( n77615 , n77611 , n77614 );
buf ( n77616 , n77615 );
buf ( n77617 , n77616 );
or ( n77618 , n77608 , n77617 );
buf ( n77619 , n76076 );
buf ( n77620 , n56614 );
or ( n77621 , n77619 , n77620 );
nand ( n77622 , n77618 , n77621 );
buf ( n77623 , n77622 );
xor ( n77624 , n77607 , n77623 );
buf ( n77625 , n55166 );
buf ( n77626 , n75821 );
nor ( n77627 , n77625 , n77626 );
buf ( n77628 , n77627 );
buf ( n77629 , n77628 );
buf ( n77630 , n58894 );
buf ( n77631 , n71804 );
or ( n77632 , n77630 , n77631 );
buf ( n77633 , n56789 );
buf ( n77634 , n71801 );
or ( n77635 , n77633 , n77634 );
nand ( n77636 , n77632 , n77635 );
buf ( n77637 , n77636 );
buf ( n77638 , n77637 );
not ( n77639 , n77638 );
buf ( n77640 , n58916 );
not ( n77641 , n77640 );
or ( n77642 , n77639 , n77641 );
buf ( n77643 , n77456 );
buf ( n77644 , n58884 );
or ( n77645 , n77643 , n77644 );
nand ( n77646 , n77642 , n77645 );
buf ( n77647 , n77646 );
buf ( n77648 , n77647 );
and ( n77649 , n77629 , n77648 );
buf ( n77650 , n77649 );
and ( n77651 , n77624 , n77650 );
and ( n77652 , n77607 , n77623 );
or ( n77653 , n77651 , n77652 );
xor ( n77654 , n76067 , n76084 );
xor ( n77655 , n77654 , n76104 );
buf ( n77656 , n77655 );
xor ( n77657 , n77653 , n77656 );
buf ( n77658 , n62691 );
not ( n77659 , n77658 );
buf ( n77660 , n77425 );
not ( n77661 , n77660 );
or ( n77662 , n77659 , n77661 );
buf ( n77663 , n70333 );
buf ( n77664 , n60096 );
and ( n77665 , n77663 , n77664 );
buf ( n77666 , n70336 );
buf ( n77667 , n62663 );
and ( n77668 , n77666 , n77667 );
nor ( n77669 , n77665 , n77668 );
buf ( n77670 , n77669 );
buf ( n77671 , n77670 );
buf ( n77672 , n62935 );
or ( n77673 , n77671 , n77672 );
nand ( n77674 , n77662 , n77673 );
buf ( n77675 , n77674 );
and ( n77676 , n77657 , n77675 );
and ( n77677 , n77653 , n77656 );
or ( n77678 , n77676 , n77677 );
xor ( n77679 , n77395 , n77411 );
xor ( n77680 , n77679 , n77433 );
and ( n77681 , n77678 , n77680 );
buf ( n77682 , n1664 );
not ( n77683 , n77682 );
buf ( n77684 , n77564 );
not ( n77685 , n77684 );
buf ( n77686 , n77685 );
buf ( n77687 , n77686 );
not ( n77688 , n77687 );
or ( n77689 , n77683 , n77688 );
buf ( n77690 , n64211 );
buf ( n77691 , n63003 );
and ( n77692 , n77690 , n77691 );
buf ( n77693 , n66610 );
buf ( n77694 , n64223 );
and ( n77695 , n77693 , n77694 );
nor ( n77696 , n77692 , n77695 );
buf ( n77697 , n77696 );
buf ( n77698 , n77697 );
buf ( n77699 , n64230 );
or ( n77700 , n77698 , n77699 );
nand ( n77701 , n77689 , n77700 );
buf ( n77702 , n77701 );
xor ( n77703 , n77395 , n77411 );
xor ( n77704 , n77703 , n77433 );
and ( n77705 , n77702 , n77704 );
and ( n77706 , n77678 , n77702 );
or ( n77707 , n77681 , n77705 , n77706 );
xor ( n77708 , n77594 , n77707 );
xor ( n77709 , n77556 , n77573 );
xor ( n77710 , n77709 , n77578 );
buf ( n77711 , n77710 );
and ( n77712 , n77708 , n77711 );
and ( n77713 , n77594 , n77707 );
or ( n77714 , n77712 , n77713 );
buf ( n77715 , n77714 );
xor ( n77716 , n76032 , n76139 );
xor ( n77717 , n77716 , n76145 );
buf ( n77718 , n77717 );
buf ( n77719 , n77718 );
xor ( n77720 , n77715 , n77719 );
xor ( n77721 , n75775 , n75791 );
xor ( n77722 , n77721 , n75813 );
xor ( n77723 , n77441 , n77582 );
xor ( n77724 , n77722 , n77723 );
buf ( n77725 , n77724 );
and ( n77726 , n77720 , n77725 );
and ( n77727 , n77715 , n77719 );
or ( n77728 , n77726 , n77727 );
buf ( n77729 , n77728 );
xor ( n77730 , n76015 , n76149 );
xor ( n77731 , n77730 , n76153 );
and ( n77732 , n77729 , n77731 );
and ( n77733 , n77587 , n77729 );
or ( n77734 , n77590 , n77732 , n77733 );
buf ( n77735 , n77734 );
nand ( n77736 , n77373 , n77735 );
buf ( n77737 , n77736 );
buf ( n77738 , n77737 );
buf ( n77739 , n77366 );
buf ( n77740 , n77371 );
nand ( n77741 , n77739 , n77740 );
buf ( n77742 , n77741 );
buf ( n77743 , n77742 );
and ( n77744 , n77738 , n77743 );
buf ( n77745 , n77744 );
buf ( n77746 , n77745 );
nand ( n77747 , n77342 , n77746 );
buf ( n77748 , n77747 );
buf ( n77749 , n77748 );
not ( n77750 , n77749 );
xor ( n77751 , n77046 , n77071 );
xor ( n77752 , n77751 , n77101 );
buf ( n77753 , n77752 );
buf ( n77754 , n77753 );
not ( n77755 , n77754 );
or ( n77756 , n77750 , n77755 );
buf ( n77757 , n77745 );
not ( n77758 , n77757 );
buf ( n77759 , n77340 );
nand ( n77760 , n77758 , n77759 );
buf ( n77761 , n77760 );
buf ( n77762 , n77761 );
nand ( n77763 , n77756 , n77762 );
buf ( n77764 , n77763 );
buf ( n77765 , n77764 );
xor ( n77766 , n77316 , n77765 );
buf ( n77767 , n56289 );
not ( n77768 , n77767 );
buf ( n77769 , n68606 );
not ( n77770 , n77769 );
or ( n77771 , n77768 , n77770 );
buf ( n77772 , n25226 );
buf ( n77773 , n52094 );
nand ( n77774 , n77772 , n77773 );
buf ( n77775 , n77774 );
buf ( n77776 , n77775 );
nand ( n77777 , n77771 , n77776 );
buf ( n77778 , n77777 );
buf ( n77779 , n77778 );
not ( n77780 , n77779 );
buf ( n77781 , n70268 );
not ( n77782 , n77781 );
or ( n77783 , n77780 , n77782 );
buf ( n77784 , n75649 );
buf ( n77785 , n42665 );
nand ( n77786 , n77784 , n77785 );
buf ( n77787 , n77786 );
buf ( n77788 , n77787 );
nand ( n77789 , n77783 , n77788 );
buf ( n77790 , n77789 );
buf ( n77791 , n77790 );
and ( n77792 , n77766 , n77791 );
and ( n77793 , n77316 , n77765 );
or ( n77794 , n77792 , n77793 );
buf ( n77795 , n77794 );
buf ( n77796 , n77795 );
nand ( n77797 , n77312 , n77796 );
buf ( n77798 , n77797 );
buf ( n77799 , n77798 );
nand ( n77800 , n77309 , n77799 );
buf ( n77801 , n77800 );
buf ( n77802 , n77801 );
and ( n77803 , n77256 , n77802 );
and ( n77804 , n77230 , n77255 );
or ( n77805 , n77803 , n77804 );
buf ( n77806 , n77805 );
buf ( n77807 , n77806 );
nand ( n77808 , n77209 , n77807 );
buf ( n77809 , n77808 );
buf ( n77810 , n77809 );
nand ( n77811 , C1 , n77810 );
buf ( n77812 , n77811 );
nand ( n77813 , n77182 , n77812 );
buf ( n77814 , n77813 );
buf ( n77815 , C1 );
nand ( n77816 , n77814 , n77815 );
buf ( n77817 , n77816 );
buf ( n77818 , n77817 );
not ( n77819 , n77818 );
buf ( n77820 , n77819 );
buf ( n77821 , n77820 );
and ( n77822 , n76952 , n77821 );
not ( n77823 , n76952 );
buf ( n77824 , n77817 );
and ( n77825 , n77823 , n77824 );
nor ( n77826 , n77822 , n77825 );
buf ( n77827 , n77826 );
buf ( n77828 , n77827 );
buf ( n77829 , n54067 );
not ( n77830 , n77829 );
buf ( n77831 , n12481 );
not ( n77832 , n77831 );
or ( n77833 , n77830 , n77832 );
buf ( n77834 , n48356 );
buf ( n77835 , n56325 );
nand ( n77836 , n77834 , n77835 );
buf ( n77837 , n77836 );
buf ( n77838 , n77837 );
nand ( n77839 , n77833 , n77838 );
buf ( n77840 , n77839 );
buf ( n77841 , n77840 );
not ( n77842 , n77841 );
buf ( n77843 , n53628 );
not ( n77844 , n77843 );
or ( n77845 , n77842 , n77844 );
buf ( n77846 , n76324 );
buf ( n77847 , n43905 );
nand ( n77848 , n77846 , n77847 );
buf ( n77849 , n77848 );
buf ( n77850 , n77849 );
nand ( n77851 , n77845 , n77850 );
buf ( n77852 , n77851 );
buf ( n77853 , n77852 );
not ( n77854 , n77853 );
buf ( n77855 , n60545 );
not ( n77856 , n77855 );
buf ( n77857 , n76961 );
not ( n77858 , n77857 );
or ( n77859 , n77856 , n77858 );
buf ( n77860 , n48836 );
not ( n77861 , n77860 );
buf ( n77862 , n56545 );
not ( n77863 , n77862 );
or ( n77864 , n77861 , n77863 );
buf ( n77865 , n29754 );
buf ( n77866 , n72931 );
nand ( n77867 , n77865 , n77866 );
buf ( n77868 , n77867 );
buf ( n77869 , n77868 );
nand ( n77870 , n77864 , n77869 );
buf ( n77871 , n77870 );
buf ( n77872 , n77871 );
buf ( n77873 , n51488 );
nand ( n77874 , n77872 , n77873 );
buf ( n77875 , n77874 );
buf ( n77876 , n77875 );
nand ( n77877 , n77859 , n77876 );
buf ( n77878 , n77877 );
buf ( n77879 , n77878 );
not ( n77880 , n77879 );
buf ( n77881 , n77880 );
buf ( n77882 , n77881 );
nand ( n77883 , n77854 , n77882 );
buf ( n77884 , n77883 );
xor ( n77885 , n75552 , n75577 );
xor ( n77886 , n77885 , n75582 );
buf ( n77887 , n77886 );
and ( n77888 , n77884 , n77887 );
and ( n77889 , n77878 , n77852 );
nor ( n77890 , n77888 , n77889 );
buf ( n77891 , n77890 );
buf ( n77892 , n76310 );
buf ( n77893 , n76344 );
xor ( n77894 , n77892 , n77893 );
buf ( n77895 , n76336 );
xor ( n77896 , n77894 , n77895 );
buf ( n77897 , n77896 );
buf ( n77898 , n77897 );
xor ( n77899 , n77891 , n77898 );
buf ( n77900 , C1 );
and ( n77901 , n77899 , n77900 );
and ( n77902 , n77891 , n77898 );
or ( n77903 , n77901 , n77902 );
buf ( n77904 , n77903 );
buf ( n77905 , n77904 );
not ( n77906 , n77905 );
not ( n77907 , n77180 );
and ( n77908 , n77907 , C1 );
nor ( n77909 , C0 , n77908 );
and ( n77910 , n77909 , n77812 );
not ( n77911 , n77909 );
not ( n77912 , n77812 );
and ( n77913 , n77911 , n77912 );
nor ( n77914 , n77910 , n77913 );
buf ( n77915 , n77914 );
not ( n77916 , n77915 );
or ( n77917 , n77906 , n77916 );
buf ( n77918 , n77175 );
buf ( n77919 , n76968 );
xor ( n77920 , n77918 , n77919 );
buf ( n77921 , n76971 );
xnor ( n77922 , n77920 , n77921 );
buf ( n77923 , n77922 );
not ( n77924 , n77923 );
buf ( n77925 , n50995 );
not ( n77926 , n77925 );
buf ( n77927 , n25293 );
not ( n77928 , n77927 );
or ( n77929 , n77926 , n77928 );
buf ( n77930 , n25290 );
buf ( n77931 , n50992 );
nand ( n77932 , n77930 , n77931 );
buf ( n77933 , n77932 );
buf ( n77934 , n77933 );
nand ( n77935 , n77929 , n77934 );
buf ( n77936 , n77935 );
buf ( n77937 , n77936 );
not ( n77938 , n77937 );
buf ( n77939 , n42246 );
not ( n77940 , n77939 );
or ( n77941 , n77938 , n77940 );
buf ( n77942 , n77110 );
buf ( n77943 , n42309 );
nand ( n77944 , n77942 , n77943 );
buf ( n77945 , n77944 );
buf ( n77946 , n77945 );
nand ( n77947 , n77941 , n77946 );
buf ( n77948 , n77947 );
buf ( n77949 , n77948 );
buf ( n77950 , n47716 );
buf ( n77951 , n44524 );
and ( n77952 , n77950 , n77951 );
not ( n77953 , n77950 );
buf ( n77954 , n74492 );
and ( n77955 , n77953 , n77954 );
nor ( n77956 , n77952 , n77955 );
buf ( n77957 , n77956 );
buf ( n77958 , n77957 );
not ( n77959 , n77958 );
buf ( n77960 , n44517 );
not ( n77961 , n77960 );
or ( n77962 , n77959 , n77961 );
buf ( n77963 , n77058 );
buf ( n77964 , n44496 );
nand ( n77965 , n77963 , n77964 );
buf ( n77966 , n77965 );
buf ( n77967 , n77966 );
nand ( n77968 , n77962 , n77967 );
buf ( n77969 , n77968 );
buf ( n77970 , n77969 );
buf ( n77971 , n71232 );
buf ( n77972 , n15265 );
and ( n77973 , n77971 , n77972 );
buf ( n77974 , n71235 );
buf ( n77975 , n60090 );
and ( n77976 , n77974 , n77975 );
nor ( n77977 , n77973 , n77976 );
buf ( n77978 , n77977 );
buf ( n77979 , n77978 );
buf ( n77980 , n60270 );
or ( n77981 , n77979 , n77980 );
buf ( n77982 , n77514 );
buf ( n77983 , n60100 );
or ( n77984 , n77982 , n77983 );
nand ( n77985 , n77981 , n77984 );
buf ( n77986 , n77985 );
xor ( n77987 , n77463 , n77479 );
xor ( n77988 , n77987 , n77496 );
and ( n77989 , n77986 , n77988 );
buf ( n77990 , n77616 );
buf ( n77991 , n56614 );
or ( n77992 , n77990 , n77991 );
buf ( n77993 , n56634 );
nand ( n77994 , n77992 , n77993 );
buf ( n77995 , n77994 );
buf ( n77996 , n77995 );
buf ( n77997 , n56799 );
buf ( n77998 , n56777 );
buf ( n77999 , n72445 );
and ( n78000 , n77998 , n77999 );
buf ( n78001 , n56804 );
buf ( n78002 , n72448 );
and ( n78003 , n78001 , n78002 );
nor ( n78004 , n78000 , n78003 );
buf ( n78005 , n78004 );
buf ( n78006 , n78005 );
or ( n78007 , n77997 , n78006 );
buf ( n78008 , n77489 );
buf ( n78009 , n56796 );
or ( n78010 , n78008 , n78009 );
nand ( n78011 , n78007 , n78010 );
buf ( n78012 , n78011 );
buf ( n78013 , n78012 );
xor ( n78014 , n77996 , n78013 );
buf ( n78015 , n71225 );
buf ( n78016 , n15265 );
and ( n78017 , n78015 , n78016 );
buf ( n78018 , n71228 );
buf ( n78019 , n60090 );
and ( n78020 , n78018 , n78019 );
nor ( n78021 , n78017 , n78020 );
buf ( n78022 , n78021 );
buf ( n78023 , n78022 );
not ( n78024 , n78023 );
buf ( n78025 , n78024 );
buf ( n78026 , n78025 );
not ( n78027 , n78026 );
buf ( n78028 , n60101 );
not ( n78029 , n78028 );
or ( n78030 , n78027 , n78029 );
buf ( n78031 , n77978 );
buf ( n78032 , n60100 );
or ( n78033 , n78031 , n78032 );
nand ( n78034 , n78030 , n78033 );
buf ( n78035 , n78034 );
buf ( n78036 , n78035 );
and ( n78037 , n78014 , n78036 );
and ( n78038 , n77996 , n78013 );
or ( n78039 , n78037 , n78038 );
buf ( n78040 , n78039 );
xor ( n78041 , n77463 , n77479 );
xor ( n78042 , n78041 , n77496 );
and ( n78043 , n78040 , n78042 );
and ( n78044 , n77986 , n78040 );
or ( n78045 , n77989 , n78043 , n78044 );
buf ( n78046 , n78045 );
buf ( n78047 , n68217 );
buf ( n78048 , n64129 );
and ( n78049 , n78047 , n78048 );
buf ( n78050 , n68220 );
buf ( n78051 , n64133 );
and ( n78052 , n78050 , n78051 );
nor ( n78053 , n78049 , n78052 );
buf ( n78054 , n78053 );
buf ( n78055 , n78054 );
buf ( n78056 , n64141 );
or ( n78057 , n78055 , n78056 );
buf ( n78058 , n77547 );
buf ( n78059 , n63010 );
or ( n78060 , n78058 , n78059 );
nand ( n78061 , n78057 , n78060 );
buf ( n78062 , n78061 );
buf ( n78063 , n78062 );
xor ( n78064 , n78046 , n78063 );
xor ( n78065 , n77500 , n77503 );
xor ( n78066 , n78065 , n77526 );
buf ( n78067 , n78066 );
buf ( n78068 , n78067 );
and ( n78069 , n78064 , n78068 );
and ( n78070 , n78046 , n78063 );
or ( n78071 , n78069 , n78070 );
buf ( n78072 , n78071 );
xor ( n78073 , n77447 , n77530 );
xor ( n78074 , n78073 , n77552 );
and ( n78075 , n78072 , n78074 );
buf ( n78076 , n66601 );
buf ( n78077 , n63003 );
and ( n78078 , n78076 , n78077 );
buf ( n78079 , n66604 );
buf ( n78080 , n63000 );
and ( n78081 , n78079 , n78080 );
nor ( n78082 , n78078 , n78081 );
buf ( n78083 , n78082 );
buf ( n78084 , n78083 );
buf ( n78085 , n64230 );
or ( n78086 , n78084 , n78085 );
buf ( n78087 , n77697 );
buf ( n78088 , n64227 );
or ( n78089 , n78087 , n78088 );
nand ( n78090 , n78086 , n78089 );
buf ( n78091 , n78090 );
xor ( n78092 , n77653 , n77656 );
xor ( n78093 , n78092 , n77675 );
and ( n78094 , n78091 , n78093 );
buf ( n78095 , n70348 );
buf ( n78096 , n62681 );
and ( n78097 , n78095 , n78096 );
buf ( n78098 , n70351 );
buf ( n78099 , n62663 );
and ( n78100 , n78098 , n78099 );
nor ( n78101 , n78097 , n78100 );
buf ( n78102 , n78101 );
buf ( n78103 , n78102 );
buf ( n78104 , n62935 );
or ( n78105 , n78103 , n78104 );
buf ( n78106 , n77670 );
buf ( n78107 , n62676 );
or ( n78108 , n78106 , n78107 );
nand ( n78109 , n78105 , n78108 );
buf ( n78110 , n78109 );
xor ( n78111 , n77607 , n77623 );
xor ( n78112 , n78111 , n77650 );
and ( n78113 , n78110 , n78112 );
buf ( n78114 , n63013 );
not ( n78115 , n78114 );
buf ( n78116 , n68232 );
buf ( n78117 , n64129 );
and ( n78118 , n78116 , n78117 );
buf ( n78119 , n68235 );
buf ( n78120 , n64133 );
and ( n78121 , n78119 , n78120 );
nor ( n78122 , n78118 , n78121 );
buf ( n78123 , n78122 );
not ( n78124 , n78123 );
buf ( n78125 , n78124 );
not ( n78126 , n78125 );
or ( n78127 , n78115 , n78126 );
buf ( n78128 , n78054 );
buf ( n78129 , n63010 );
or ( n78130 , n78128 , n78129 );
nand ( n78131 , n78127 , n78130 );
buf ( n78132 , n78131 );
xor ( n78133 , n77607 , n77623 );
xor ( n78134 , n78133 , n77650 );
and ( n78135 , n78132 , n78134 );
and ( n78136 , n78110 , n78132 );
or ( n78137 , n78113 , n78135 , n78136 );
xor ( n78138 , n77653 , n77656 );
xor ( n78139 , n78138 , n77675 );
and ( n78140 , n78137 , n78139 );
and ( n78141 , n78091 , n78137 );
or ( n78142 , n78094 , n78140 , n78141 );
xor ( n78143 , n77447 , n77530 );
xor ( n78144 , n78143 , n77552 );
and ( n78145 , n78142 , n78144 );
and ( n78146 , n78072 , n78142 );
or ( n78147 , n78075 , n78145 , n78146 );
xor ( n78148 , n77594 , n77707 );
xor ( n78149 , n78148 , n77711 );
and ( n78150 , n78147 , n78149 );
xor ( n78151 , n78046 , n78063 );
xor ( n78152 , n78151 , n78068 );
buf ( n78153 , n78152 );
buf ( n78154 , n66690 );
buf ( n78155 , n63003 );
and ( n78156 , n78154 , n78155 );
buf ( n78157 , n66693 );
buf ( n78158 , n63000 );
and ( n78159 , n78157 , n78158 );
nor ( n78160 , n78156 , n78159 );
buf ( n78161 , n78160 );
buf ( n78162 , n78161 );
buf ( n78163 , n64230 );
or ( n78164 , n78162 , n78163 );
buf ( n78165 , n78083 );
buf ( n78166 , n64227 );
or ( n78167 , n78165 , n78166 );
nand ( n78168 , n78164 , n78167 );
buf ( n78169 , n78168 );
buf ( n78170 , n78169 );
buf ( n78171 , n60270 );
buf ( n78172 , n15265 );
buf ( n78173 , n71307 );
and ( n78174 , n78172 , n78173 );
buf ( n78175 , n71310 );
buf ( n78176 , n60090 );
and ( n78177 , n78175 , n78176 );
nor ( n78178 , n78174 , n78177 );
buf ( n78179 , n78178 );
buf ( n78180 , n78179 );
or ( n78181 , n78171 , n78180 );
buf ( n78182 , n78022 );
buf ( n78183 , n60100 );
or ( n78184 , n78182 , n78183 );
nand ( n78185 , n78181 , n78184 );
buf ( n78186 , n78185 );
buf ( n78187 , n16808 );
buf ( n78188 , n623 );
and ( n78189 , n78187 , n78188 );
buf ( n78190 , n7201 );
buf ( n78191 , n75821 );
and ( n78192 , n78190 , n78191 );
buf ( n78193 , n56777 );
nor ( n78194 , n78192 , n78193 );
buf ( n78195 , n78194 );
buf ( n78196 , n78195 );
buf ( n78197 , n16469 );
nor ( n78198 , n78189 , n78196 , n78197 );
buf ( n78199 , n78198 );
xor ( n78200 , n78186 , n78199 );
buf ( n78201 , n56799 );
buf ( n78202 , n56777 );
buf ( n78203 , n74115 );
and ( n78204 , n78202 , n78203 );
buf ( n78205 , n56804 );
buf ( n78206 , n74118 );
and ( n78207 , n78205 , n78206 );
nor ( n78208 , n78204 , n78207 );
buf ( n78209 , n78208 );
buf ( n78210 , n78209 );
or ( n78211 , n78201 , n78210 );
buf ( n78212 , n78005 );
buf ( n78213 , n58982 );
or ( n78214 , n78212 , n78213 );
nand ( n78215 , n78211 , n78214 );
buf ( n78216 , n78215 );
and ( n78217 , n78200 , n78216 );
and ( n78218 , n78186 , n78199 );
or ( n78219 , n78217 , n78218 );
buf ( n78220 , n78219 );
xor ( n78221 , n77629 , n77648 );
buf ( n78222 , n78221 );
buf ( n78223 , n78222 );
xor ( n78224 , n78220 , n78223 );
buf ( n78225 , n62679 );
not ( n78226 , n78225 );
buf ( n78227 , n70530 );
buf ( n78228 , n62684 );
or ( n78229 , n78227 , n78228 );
buf ( n78230 , n70527 );
buf ( n78231 , n62681 );
or ( n78232 , n78230 , n78231 );
nand ( n78233 , n78229 , n78232 );
buf ( n78234 , n78233 );
buf ( n78235 , n78234 );
not ( n78236 , n78235 );
or ( n78237 , n78226 , n78236 );
buf ( n78238 , n78102 );
buf ( n78239 , n62676 );
or ( n78240 , n78238 , n78239 );
nand ( n78241 , n78237 , n78240 );
buf ( n78242 , n78241 );
buf ( n78243 , n78242 );
and ( n78244 , n78224 , n78243 );
and ( n78245 , n78220 , n78223 );
or ( n78246 , n78244 , n78245 );
buf ( n78247 , n78246 );
buf ( n78248 , n78247 );
xor ( n78249 , n78170 , n78248 );
xor ( n78250 , n77463 , n77479 );
xor ( n78251 , n78250 , n77496 );
xor ( n78252 , n77986 , n78040 );
xor ( n78253 , n78251 , n78252 );
buf ( n78254 , n78253 );
and ( n78255 , n78249 , n78254 );
and ( n78256 , n78170 , n78248 );
or ( n78257 , n78255 , n78256 );
buf ( n78258 , n78257 );
xor ( n78259 , n78153 , n78258 );
xor ( n78260 , n77653 , n77656 );
xor ( n78261 , n78260 , n77675 );
xor ( n78262 , n78091 , n78137 );
xor ( n78263 , n78261 , n78262 );
and ( n78264 , n78259 , n78263 );
and ( n78265 , n78153 , n78258 );
or ( n78266 , n78264 , n78265 );
buf ( n78267 , n78266 );
xor ( n78268 , n77395 , n77411 );
xor ( n78269 , n78268 , n77433 );
xor ( n78270 , n77678 , n77702 );
xor ( n78271 , n78269 , n78270 );
buf ( n78272 , n78271 );
xor ( n78273 , n78267 , n78272 );
xor ( n78274 , n77447 , n77530 );
xor ( n78275 , n78274 , n77552 );
xor ( n78276 , n78072 , n78142 );
xor ( n78277 , n78275 , n78276 );
buf ( n78278 , n78277 );
and ( n78279 , n78273 , n78278 );
and ( n78280 , n78267 , n78272 );
or ( n78281 , n78279 , n78280 );
buf ( n78282 , n78281 );
xor ( n78283 , n77594 , n77707 );
xor ( n78284 , n78283 , n77711 );
and ( n78285 , n78282 , n78284 );
and ( n78286 , n78147 , n78282 );
or ( n78287 , n78150 , n78285 , n78286 );
not ( n78288 , n78287 );
buf ( n78289 , n47716 );
not ( n78290 , n78289 );
buf ( n78291 , n44491 );
not ( n78292 , n78291 );
or ( n78293 , n78290 , n78292 );
buf ( n78294 , n44494 );
buf ( n78295 , n47713 );
nand ( n78296 , n78294 , n78295 );
buf ( n78297 , n78296 );
buf ( n78298 , n78297 );
nand ( n78299 , n78293 , n78298 );
buf ( n78300 , n78299 );
buf ( n78301 , n78300 );
not ( n78302 , n78301 );
buf ( n78303 , n45741 );
not ( n78304 , n78303 );
or ( n78305 , n78302 , n78304 );
buf ( n78306 , n45746 );
not ( n78307 , n78306 );
buf ( n78308 , n46384 );
not ( n78309 , n78308 );
or ( n78310 , n78307 , n78309 );
buf ( n78311 , n44491 );
buf ( n78312 , n46384 );
not ( n78313 , n78312 );
buf ( n78314 , n78313 );
buf ( n78315 , n78314 );
nand ( n78316 , n78311 , n78315 );
buf ( n78317 , n78316 );
buf ( n78318 , n78317 );
nand ( n78319 , n78310 , n78318 );
buf ( n78320 , n78319 );
buf ( n78321 , n78320 );
buf ( n78322 , n46246 );
nand ( n78323 , n78321 , n78322 );
buf ( n78324 , n78323 );
buf ( n78325 , n78324 );
nand ( n78326 , n78305 , n78325 );
buf ( n78327 , n78326 );
not ( n78328 , n78327 );
or ( n78329 , n78288 , n78328 );
buf ( n78330 , n78327 );
buf ( n78331 , n78287 );
or ( n78332 , n78330 , n78331 );
xor ( n78333 , n77715 , n77719 );
xor ( n78334 , n78333 , n77725 );
buf ( n78335 , n78334 );
buf ( n78336 , n78335 );
nand ( n78337 , n78332 , n78336 );
buf ( n78338 , n78337 );
nand ( n78339 , n78329 , n78338 );
not ( n78340 , n78339 );
xor ( n78341 , n76015 , n76149 );
xor ( n78342 , n78341 , n76153 );
xor ( n78343 , n77587 , n77729 );
xor ( n78344 , n78342 , n78343 );
buf ( n78345 , n78344 );
not ( n78346 , n78345 );
buf ( n78347 , n78346 );
buf ( n78348 , n77359 );
buf ( n78349 , n67149 );
and ( n78350 , n78348 , n78349 );
buf ( n78351 , n78320 );
not ( n78352 , n78351 );
buf ( n78353 , n45742 );
nor ( n78354 , n78352 , n78353 );
buf ( n78355 , n78354 );
buf ( n78356 , n78355 );
nor ( n78357 , n78350 , n78356 );
buf ( n78358 , n78357 );
nand ( n78359 , n78347 , n78358 );
not ( n78360 , n78359 );
or ( n78361 , n78340 , n78360 );
buf ( n78362 , n78358 );
not ( n78363 , n78362 );
buf ( n78364 , n78344 );
nand ( n78365 , n78363 , n78364 );
buf ( n78366 , n78365 );
nand ( n78367 , n78361 , n78366 );
buf ( n78368 , n78367 );
xor ( n78369 , n77970 , n78368 );
buf ( n78370 , n50060 );
not ( n78371 , n78370 );
buf ( n78372 , n77077 );
not ( n78373 , n78372 );
or ( n78374 , n78371 , n78373 );
buf ( n78375 , n42228 );
buf ( n78376 , n67438 );
nand ( n78377 , n78375 , n78376 );
buf ( n78378 , n78377 );
buf ( n78379 , n78378 );
nand ( n78380 , n78374 , n78379 );
buf ( n78381 , n78380 );
buf ( n78382 , n78381 );
not ( n78383 , n78382 );
buf ( n78384 , n41596 );
not ( n78385 , n78384 );
or ( n78386 , n78383 , n78385 );
buf ( n78387 , n77088 );
buf ( n78388 , n41574 );
nand ( n78389 , n78387 , n78388 );
buf ( n78390 , n78389 );
buf ( n78391 , n78390 );
nand ( n78392 , n78386 , n78391 );
buf ( n78393 , n78392 );
buf ( n78394 , n78393 );
and ( n78395 , n78369 , n78394 );
and ( n78396 , n77970 , n78368 );
or ( n78397 , n78395 , n78396 );
buf ( n78398 , n78397 );
buf ( n78399 , n78398 );
xor ( n78400 , n77949 , n78399 );
buf ( n78401 , n46912 );
not ( n78402 , n78401 );
buf ( n78403 , n77141 );
not ( n78404 , n78403 );
or ( n78405 , n78402 , n78404 );
buf ( n78406 , n46875 );
buf ( n78407 , n42856 );
and ( n78408 , n78406 , n78407 );
not ( n78409 , n78406 );
buf ( n78410 , n72235 );
and ( n78411 , n78409 , n78410 );
nor ( n78412 , n78408 , n78411 );
buf ( n78413 , n78412 );
buf ( n78414 , n78413 );
buf ( n78415 , n46907 );
nand ( n78416 , n78414 , n78415 );
buf ( n78417 , n78416 );
buf ( n78418 , n78417 );
nand ( n78419 , n78405 , n78418 );
buf ( n78420 , n78419 );
buf ( n78421 , n78420 );
and ( n78422 , n78400 , n78421 );
and ( n78423 , n77949 , n78399 );
or ( n78424 , n78422 , n78423 );
buf ( n78425 , n78424 );
buf ( n78426 , n78425 );
buf ( n78427 , n66463 );
not ( n78428 , n78427 );
buf ( n78429 , n41634 );
not ( n78430 , n78429 );
or ( n78431 , n78428 , n78430 );
buf ( n78432 , n12481 );
nand ( n78433 , n78431 , n78432 );
buf ( n78434 , n78433 );
buf ( n78435 , n78434 );
buf ( n78436 , n61434 );
buf ( n78437 , n42366 );
buf ( n78438 , n25010 );
nand ( n78439 , n78437 , n78438 );
buf ( n78440 , n78439 );
buf ( n78441 , n78440 );
and ( n78442 , n78435 , n78436 , n78441 );
buf ( n78443 , n78442 );
buf ( n78444 , n78443 );
xor ( n78445 , n78426 , n78444 );
xor ( n78446 , n77106 , n77123 );
xor ( n78447 , n78446 , n77149 );
buf ( n78448 , n78447 );
buf ( n78449 , n78448 );
and ( n78450 , n78445 , n78449 );
and ( n78451 , n78426 , n78444 );
or ( n78452 , n78450 , n78451 );
buf ( n78453 , n78452 );
buf ( n78454 , n78453 );
xor ( n78455 , n77036 , n77040 );
xor ( n78456 , n78455 , n77154 );
buf ( n78457 , n78456 );
buf ( n78458 , n78457 );
xor ( n78459 , n78454 , n78458 );
buf ( n78460 , n60545 );
not ( n78461 , n78460 );
buf ( n78462 , n77871 );
not ( n78463 , n78462 );
or ( n78464 , n78461 , n78463 );
buf ( n78465 , n48836 );
not ( n78466 , n78465 );
buf ( n78467 , n58632 );
not ( n78468 , n78467 );
or ( n78469 , n78466 , n78468 );
buf ( n78470 , n13653 );
buf ( n78471 , n72931 );
nand ( n78472 , n78470 , n78471 );
buf ( n78473 , n78472 );
buf ( n78474 , n78473 );
nand ( n78475 , n78469 , n78474 );
buf ( n78476 , n78475 );
buf ( n78477 , n78476 );
buf ( n78478 , n51488 );
nand ( n78479 , n78477 , n78478 );
buf ( n78480 , n78479 );
buf ( n78481 , n78480 );
nand ( n78482 , n78464 , n78481 );
buf ( n78483 , n78482 );
buf ( n78484 , n78483 );
and ( n78485 , n78459 , n78484 );
and ( n78486 , n78454 , n78458 );
or ( n78487 , n78485 , n78486 );
buf ( n78488 , n78487 );
buf ( n78489 , n78488 );
buf ( n78490 , n77165 );
buf ( n78491 , n77169 );
and ( n78492 , n78490 , n78491 );
not ( n78493 , n78490 );
buf ( n78494 , n77016 );
and ( n78495 , n78493 , n78494 );
nor ( n78496 , n78492 , n78495 );
buf ( n78497 , n78496 );
xor ( n78498 , n78497 , n77158 );
buf ( n78499 , n78498 );
not ( n78500 , n78499 );
buf ( n78501 , n78500 );
buf ( n78502 , n78501 );
nor ( n78503 , n43904 , n56325 );
buf ( n78504 , n78503 );
buf ( n78505 , n48865 );
not ( n78506 , n78505 );
buf ( n78507 , n77247 );
not ( n78508 , n78507 );
or ( n78509 , n78506 , n78508 );
and ( n78510 , n13662 , n75377 );
not ( n78511 , n13662 );
and ( n78512 , n78511 , n48808 );
or ( n78513 , n78510 , n78512 );
buf ( n78514 , n78513 );
buf ( n78515 , n48852 );
nand ( n78516 , n78514 , n78515 );
buf ( n78517 , n78516 );
buf ( n78518 , n78517 );
nand ( n78519 , n78509 , n78518 );
buf ( n78520 , n78519 );
buf ( n78521 , n78520 );
xor ( n78522 , n78504 , n78521 );
buf ( n78523 , n50979 );
buf ( n78524 , n58361 );
buf ( n78525 , n61434 );
and ( n78526 , n78524 , n78525 );
not ( n78527 , n78524 );
buf ( n78528 , n62598 );
and ( n78529 , n78527 , n78528 );
nor ( n78530 , n78526 , n78529 );
buf ( n78531 , n78530 );
buf ( n78532 , n78531 );
or ( n78533 , n78523 , n78532 );
buf ( n78534 , n77006 );
buf ( n78535 , n62579 );
or ( n78536 , n78534 , n78535 );
nand ( n78537 , n78533 , n78536 );
buf ( n78538 , n78537 );
buf ( n78539 , n78538 );
and ( n78540 , n78522 , n78539 );
and ( n78541 , n78504 , n78521 );
or ( n78542 , n78540 , n78541 );
buf ( n78543 , n78542 );
buf ( n78544 , n78543 );
not ( n78545 , n78544 );
buf ( n78546 , n78545 );
buf ( n78547 , n78546 );
nand ( n78548 , n78502 , n78547 );
buf ( n78549 , n78548 );
buf ( n78550 , n78549 );
and ( n78551 , n78489 , n78550 );
buf ( n78552 , n78546 );
buf ( n78553 , n78501 );
nor ( n78554 , n78552 , n78553 );
buf ( n78555 , n78554 );
buf ( n78556 , n78555 );
nor ( n78557 , n78551 , n78556 );
buf ( n78558 , n78557 );
not ( n78559 , n78558 );
or ( n78560 , n77924 , n78559 );
xor ( n78561 , n77276 , n77306 );
xor ( n78562 , n78561 , n77795 );
not ( n78563 , n78562 );
xor ( n78564 , n77340 , n77745 );
xnor ( n78565 , n78564 , n77753 );
buf ( n78566 , n78565 );
buf ( n78567 , n77371 );
buf ( n78568 , n77734 );
xnor ( n78569 , n78567 , n78568 );
buf ( n78570 , n78569 );
buf ( n78571 , n78570 );
not ( n78572 , n78571 );
buf ( n78573 , n77366 );
not ( n78574 , n78573 );
or ( n78575 , n78572 , n78574 );
buf ( n78576 , n77366 );
buf ( n78577 , n78570 );
or ( n78578 , n78576 , n78577 );
nand ( n78579 , n78575 , n78578 );
buf ( n78580 , n78579 );
buf ( n78581 , n78580 );
buf ( n78582 , n46912 );
not ( n78583 , n78582 );
buf ( n78584 , n78413 );
not ( n78585 , n78584 );
or ( n78586 , n78583 , n78585 );
buf ( n78587 , n46875 );
not ( n78588 , n78587 );
buf ( n78589 , n74460 );
not ( n78590 , n78589 );
or ( n78591 , n78588 , n78590 );
buf ( n78592 , n42844 );
buf ( n78593 , n46887 );
nand ( n78594 , n78592 , n78593 );
buf ( n78595 , n78594 );
buf ( n78596 , n78595 );
nand ( n78597 , n78591 , n78596 );
buf ( n78598 , n78597 );
buf ( n78599 , n78598 );
buf ( n78600 , n46907 );
nand ( n78601 , n78599 , n78600 );
buf ( n78602 , n78601 );
buf ( n78603 , n78602 );
nand ( n78604 , n78586 , n78603 );
buf ( n78605 , n78604 );
buf ( n78606 , n78605 );
xor ( n78607 , n78581 , n78606 );
buf ( n78608 , n71078 );
not ( n78609 , n78608 );
buf ( n78610 , n74492 );
not ( n78611 , n78610 );
or ( n78612 , n78609 , n78611 );
buf ( n78613 , n44524 );
buf ( n78614 , n48320 );
nand ( n78615 , n78613 , n78614 );
buf ( n78616 , n78615 );
buf ( n78617 , n78616 );
nand ( n78618 , n78612 , n78617 );
buf ( n78619 , n78618 );
buf ( n78620 , n78619 );
not ( n78621 , n78620 );
buf ( n78622 , n74488 );
not ( n78623 , n78622 );
or ( n78624 , n78621 , n78623 );
buf ( n78625 , n77957 );
buf ( n78626 , n44496 );
nand ( n78627 , n78625 , n78626 );
buf ( n78628 , n78627 );
buf ( n78629 , n78628 );
nand ( n78630 , n78624 , n78629 );
buf ( n78631 , n78630 );
buf ( n78632 , n78631 );
buf ( n78633 , n46912 );
not ( n78634 , n78633 );
buf ( n78635 , n78598 );
not ( n78636 , n78635 );
or ( n78637 , n78634 , n78636 );
buf ( n78638 , n46875 );
not ( n78639 , n78638 );
buf ( n78640 , n44946 );
not ( n78641 , n78640 );
or ( n78642 , n78639 , n78641 );
buf ( n78643 , n74500 );
buf ( n78644 , n46887 );
nand ( n78645 , n78643 , n78644 );
buf ( n78646 , n78645 );
buf ( n78647 , n78646 );
nand ( n78648 , n78642 , n78647 );
buf ( n78649 , n78648 );
buf ( n78650 , n78649 );
buf ( n78651 , n46907 );
nand ( n78652 , n78650 , n78651 );
buf ( n78653 , n78652 );
buf ( n78654 , n78653 );
nand ( n78655 , n78637 , n78654 );
buf ( n78656 , n78655 );
buf ( n78657 , n78656 );
xor ( n78658 , n78632 , n78657 );
buf ( n78659 , n50995 );
not ( n78660 , n78659 );
buf ( n78661 , n77077 );
not ( n78662 , n78661 );
or ( n78663 , n78660 , n78662 );
buf ( n78664 , n42228 );
buf ( n78665 , n50992 );
nand ( n78666 , n78664 , n78665 );
buf ( n78667 , n78666 );
buf ( n78668 , n78667 );
nand ( n78669 , n78663 , n78668 );
buf ( n78670 , n78669 );
buf ( n78671 , n78670 );
not ( n78672 , n78671 );
buf ( n78673 , n67354 );
not ( n78674 , n78673 );
or ( n78675 , n78672 , n78674 );
buf ( n78676 , n78381 );
buf ( n78677 , n41574 );
nand ( n78678 , n78676 , n78677 );
buf ( n78679 , n78678 );
buf ( n78680 , n78679 );
nand ( n78681 , n78675 , n78680 );
buf ( n78682 , n78681 );
buf ( n78683 , n78682 );
and ( n78684 , n78658 , n78683 );
and ( n78685 , n78632 , n78657 );
or ( n78686 , n78684 , n78685 );
buf ( n78687 , n78686 );
buf ( n78688 , n78687 );
and ( n78689 , n78607 , n78688 );
and ( n78690 , n78581 , n78606 );
or ( n78691 , n78689 , n78690 );
buf ( n78692 , n78691 );
buf ( n78693 , n78692 );
xor ( n78694 , n78566 , n78693 );
buf ( n78695 , n74651 );
buf ( n78696 , n52789 );
buf ( n78697 , n25226 );
and ( n78698 , n78696 , n78697 );
not ( n78699 , n78696 );
buf ( n78700 , n62510 );
and ( n78701 , n78699 , n78700 );
nor ( n78702 , n78698 , n78701 );
buf ( n78703 , n78702 );
buf ( n78704 , n78703 );
or ( n78705 , n78695 , n78704 );
buf ( n78706 , n77778 );
not ( n78707 , n78706 );
buf ( n78708 , n78707 );
buf ( n78709 , n78708 );
buf ( n78710 , n74674 );
or ( n78711 , n78709 , n78710 );
nand ( n78712 , n78705 , n78711 );
buf ( n78713 , n78712 );
buf ( n78714 , n78713 );
and ( n78715 , n78694 , n78714 );
and ( n78716 , n78566 , n78693 );
or ( n78717 , n78715 , n78716 );
buf ( n78718 , n78717 );
not ( n78719 , n78718 );
buf ( n78720 , n78513 );
buf ( n78721 , n48865 );
and ( n78722 , n78720 , n78721 );
buf ( n78723 , n48808 );
not ( n78724 , n78723 );
buf ( n78725 , n70855 );
not ( n78726 , n78725 );
or ( n78727 , n78724 , n78726 );
buf ( n78728 , n29463 );
buf ( n78729 , n75377 );
nand ( n78730 , n78728 , n78729 );
buf ( n78731 , n78730 );
buf ( n78732 , n78731 );
nand ( n78733 , n78727 , n78732 );
buf ( n78734 , n78733 );
buf ( n78735 , n78734 );
not ( n78736 , n78735 );
buf ( n78737 , n48849 );
nor ( n78738 , n78736 , n78737 );
buf ( n78739 , n78738 );
buf ( n78740 , n78739 );
nor ( n78741 , n78722 , n78740 );
buf ( n78742 , n78741 );
buf ( n78743 , n78742 );
buf ( n78744 , n53539 );
not ( n78745 , n78744 );
buf ( n78746 , n69798 );
not ( n78747 , n78746 );
or ( n78748 , n78745 , n78747 );
buf ( n78749 , n69804 );
buf ( n78750 , n53548 );
nand ( n78751 , n78749 , n78750 );
buf ( n78752 , n78751 );
buf ( n78753 , n78752 );
nand ( n78754 , n78748 , n78753 );
buf ( n78755 , n78754 );
not ( n78756 , n78755 );
not ( n78757 , n66459 );
or ( n78758 , n78756 , n78757 );
buf ( n78759 , n77293 );
buf ( n78760 , n66482 );
nand ( n78761 , n78759 , n78760 );
buf ( n78762 , n78761 );
nand ( n78763 , n78758 , n78762 );
not ( n78764 , n78763 );
buf ( n78765 , n78764 );
nand ( n78766 , n78743 , n78765 );
buf ( n78767 , n78766 );
not ( n78768 , n78767 );
or ( n78769 , n78719 , n78768 );
not ( n78770 , n78742 );
nand ( n78771 , n78770 , n78763 );
nand ( n78772 , n78769 , n78771 );
nand ( n78773 , n78563 , n78772 );
not ( n78774 , n78562 );
not ( n78775 , n78772 );
not ( n78776 , n78775 );
or ( n78777 , n78774 , n78776 );
xor ( n78778 , n77316 , n77765 );
xor ( n78779 , n78778 , n77791 );
buf ( n78780 , n78779 );
buf ( n78781 , n78780 );
buf ( n78782 , n48865 );
not ( n78783 , n78782 );
buf ( n78784 , n78734 );
not ( n78785 , n78784 );
or ( n78786 , n78783 , n78785 );
buf ( n78787 , n48808 );
not ( n78788 , n78787 );
buf ( n78789 , n28430 );
not ( n78790 , n78789 );
buf ( n78791 , n78790 );
buf ( n78792 , n78791 );
not ( n78793 , n78792 );
or ( n78794 , n78788 , n78793 );
buf ( n78795 , n28430 );
buf ( n78796 , n75377 );
nand ( n78797 , n78795 , n78796 );
buf ( n78798 , n78797 );
buf ( n78799 , n78798 );
nand ( n78800 , n78794 , n78799 );
buf ( n78801 , n78800 );
buf ( n78802 , n78801 );
buf ( n78803 , n48852 );
nand ( n78804 , n78802 , n78803 );
buf ( n78805 , n78804 );
buf ( n78806 , n78805 );
nand ( n78807 , n78786 , n78806 );
buf ( n78808 , n78807 );
buf ( n78809 , n78808 );
not ( n78810 , n78809 );
buf ( n78811 , n78810 );
buf ( n78812 , n78811 );
not ( n78813 , n78812 );
buf ( n78814 , n62579 );
not ( n78815 , n78814 );
buf ( n78816 , n12481 );
nand ( n78817 , n78815 , n78816 );
buf ( n78818 , n78817 );
buf ( n78819 , n78818 );
not ( n78820 , n78819 );
or ( n78821 , n78813 , n78820 );
xor ( n78822 , n77949 , n78399 );
xor ( n78823 , n78822 , n78421 );
buf ( n78824 , n78823 );
buf ( n78825 , n78824 );
nand ( n78826 , n78821 , n78825 );
buf ( n78827 , n78826 );
buf ( n78828 , n78827 );
buf ( n78829 , n78818 );
not ( n78830 , n78829 );
buf ( n78831 , n78830 );
buf ( n78832 , n78831 );
buf ( n78833 , n78808 );
nand ( n78834 , n78832 , n78833 );
buf ( n78835 , n78834 );
buf ( n78836 , n78835 );
nand ( n78837 , n78828 , n78836 );
buf ( n78838 , n78837 );
buf ( n78839 , n78838 );
xor ( n78840 , n78781 , n78839 );
xor ( n78841 , n78426 , n78444 );
xor ( n78842 , n78841 , n78449 );
buf ( n78843 , n78842 );
buf ( n78844 , n78843 );
and ( n78845 , n78840 , n78844 );
and ( n78846 , n78781 , n78839 );
or ( n78847 , n78845 , n78846 );
buf ( n78848 , n78847 );
nand ( n78849 , n78777 , n78848 );
nand ( n78850 , n78773 , n78849 );
buf ( n78851 , n78850 );
xor ( n78852 , n77230 , n77255 );
xor ( n78853 , n78852 , n77802 );
buf ( n78854 , n78853 );
buf ( n78855 , n78854 );
buf ( n78856 , C0 );
buf ( n78857 , n78856 );
and ( n78858 , n78851 , n78855 );
or ( n78859 , C0 , n78858 );
buf ( n78860 , n78859 );
nand ( n78861 , n78560 , n78860 );
buf ( n78862 , n77923 );
not ( n78863 , n78862 );
buf ( n78864 , n78863 );
buf ( n78865 , n78864 );
buf ( n78866 , n78558 );
not ( n78867 , n78866 );
buf ( n78868 , n78867 );
buf ( n78869 , n78868 );
nand ( n78870 , n78865 , n78869 );
buf ( n78871 , n78870 );
nand ( n78872 , n78861 , n78871 );
buf ( n78873 , n78872 );
nand ( n78874 , n77917 , n78873 );
buf ( n78875 , n78874 );
buf ( n78876 , n77914 );
buf ( n78877 , n77904 );
or ( n78878 , n78876 , n78877 );
buf ( n78879 , n78878 );
and ( n78880 , n78875 , n78879 );
buf ( n78881 , n78880 );
xor ( n78882 , n77828 , n78881 );
xor ( n78883 , n76272 , C0 );
xor ( n78884 , n78883 , n76276 );
buf ( n78885 , n78884 );
xor ( n78886 , n76281 , n76362 );
xor ( n78887 , n78886 , n76367 );
buf ( n78888 , n78887 );
buf ( n78889 , n78888 );
xor ( n78890 , n78885 , n78889 );
xor ( n78891 , n75522 , n75526 );
xor ( n78892 , n78891 , n76268 );
buf ( n78893 , n78892 );
buf ( n78894 , n78893 );
not ( n78895 , n78894 );
xor ( n78896 , n76302 , n76305 );
xor ( n78897 , n78896 , n76357 );
buf ( n78898 , n78897 );
buf ( n78899 , n78898 );
not ( n78900 , n78899 );
or ( n78901 , n78895 , n78900 );
xor ( n78902 , n76927 , n76929 );
xor ( n78903 , n78902 , n76934 );
buf ( n78904 , n78903 );
buf ( n78905 , n78904 );
buf ( n78906 , n78893 );
not ( n78907 , n78906 );
buf ( n78908 , n78898 );
not ( n78909 , n78908 );
buf ( n78910 , n78909 );
buf ( n78911 , n78910 );
nand ( n78912 , n78907 , n78911 );
buf ( n78913 , n78912 );
buf ( n78914 , n78913 );
nand ( n78915 , n78905 , n78914 );
buf ( n78916 , n78915 );
buf ( n78917 , n78916 );
nand ( n78918 , n78901 , n78917 );
buf ( n78919 , n78918 );
buf ( n78920 , n78919 );
xnor ( n78921 , n78890 , n78920 );
buf ( n78922 , n78921 );
buf ( n78923 , n78922 );
xor ( n78924 , n78882 , n78923 );
buf ( n78925 , n78924 );
buf ( n78926 , n78925 );
buf ( n78927 , C1 );
buf ( n78928 , n78927 );
buf ( n78929 , n77887 );
buf ( n78930 , n77852 );
xor ( n78931 , n78929 , n78930 );
buf ( n78932 , n77881 );
xor ( n78933 , n78931 , n78932 );
buf ( n78934 , n78933 );
buf ( n78935 , n78934 );
nand ( n78936 , n78928 , n78935 );
buf ( n78937 , n78936 );
buf ( n78938 , n78937 );
xor ( n78939 , n78504 , n78521 );
xor ( n78940 , n78939 , n78539 );
buf ( n78941 , n78940 );
buf ( n78942 , n78941 );
buf ( n78943 , C0 );
buf ( n78944 , n78943 );
xor ( n78945 , n78942 , n78944 );
buf ( n78946 , n50979 );
buf ( n78947 , n12481 );
buf ( n78948 , n41660 );
and ( n78949 , n78947 , n78948 );
not ( n78950 , n78947 );
buf ( n78951 , n59403 );
and ( n78952 , n78950 , n78951 );
nor ( n78953 , n78949 , n78952 );
buf ( n78954 , n78953 );
buf ( n78955 , n78954 );
or ( n78956 , n78946 , n78955 );
buf ( n78957 , n78531 );
buf ( n78958 , n62579 );
or ( n78959 , n78957 , n78958 );
nand ( n78960 , n78956 , n78959 );
buf ( n78961 , n78960 );
buf ( n78962 , n78961 );
buf ( n78963 , n48865 );
not ( n78964 , n78963 );
buf ( n78965 , n78801 );
not ( n78966 , n78965 );
or ( n78967 , n78964 , n78966 );
buf ( n78968 , n48808 );
not ( n78969 , n78968 );
buf ( n78970 , n72213 );
not ( n78971 , n78970 );
or ( n78972 , n78969 , n78971 );
buf ( n78973 , n43056 );
buf ( n78974 , n75377 );
nand ( n78975 , n78973 , n78974 );
buf ( n78976 , n78975 );
buf ( n78977 , n78976 );
nand ( n78978 , n78972 , n78977 );
buf ( n78979 , n78978 );
buf ( n78980 , n78979 );
buf ( n78981 , n48852 );
nand ( n78982 , n78980 , n78981 );
buf ( n78983 , n78982 );
buf ( n78984 , n78983 );
nand ( n78985 , n78967 , n78984 );
buf ( n78986 , n78985 );
buf ( n78987 , n78986 );
xor ( n78988 , n78581 , n78606 );
xor ( n78989 , n78988 , n78688 );
buf ( n78990 , n78989 );
buf ( n78991 , n78990 );
xor ( n78992 , n78987 , n78991 );
and ( n78993 , n78358 , n78344 );
not ( n78994 , n78358 );
and ( n78995 , n78994 , n78347 );
or ( n78996 , n78993 , n78995 );
xor ( n78997 , n78996 , n78339 );
xor ( n78998 , n78335 , n78287 );
xor ( n78999 , n78998 , n78327 );
buf ( n79000 , n78999 );
buf ( n79001 , n46912 );
not ( n79002 , n79001 );
buf ( n79003 , n78649 );
not ( n79004 , n79003 );
or ( n79005 , n79002 , n79004 );
buf ( n79006 , n46875 );
not ( n79007 , n79006 );
buf ( n79008 , n74414 );
not ( n79009 , n79008 );
or ( n79010 , n79007 , n79009 );
buf ( n79011 , n46114 );
buf ( n79012 , n46887 );
nand ( n79013 , n79011 , n79012 );
buf ( n79014 , n79013 );
buf ( n79015 , n79014 );
nand ( n79016 , n79010 , n79015 );
buf ( n79017 , n79016 );
buf ( n79018 , n79017 );
buf ( n79019 , n46907 );
nand ( n79020 , n79018 , n79019 );
buf ( n79021 , n79020 );
buf ( n79022 , n79021 );
nand ( n79023 , n79005 , n79022 );
buf ( n79024 , n79023 );
buf ( n79025 , n79024 );
xor ( n79026 , n79000 , n79025 );
buf ( n79027 , n50060 );
not ( n79028 , n79027 );
buf ( n79029 , n25385 );
not ( n79030 , n79029 );
buf ( n79031 , n79030 );
buf ( n79032 , n79031 );
not ( n79033 , n79032 );
or ( n79034 , n79028 , n79033 );
buf ( n79035 , n44503 );
buf ( n79036 , n67438 );
nand ( n79037 , n79035 , n79036 );
buf ( n79038 , n79037 );
buf ( n79039 , n79038 );
nand ( n79040 , n79034 , n79039 );
buf ( n79041 , n79040 );
buf ( n79042 , n79041 );
not ( n79043 , n79042 );
buf ( n79044 , n74488 );
not ( n79045 , n79044 );
or ( n79046 , n79043 , n79045 );
buf ( n79047 , n78619 );
buf ( n79048 , n44496 );
nand ( n79049 , n79047 , n79048 );
buf ( n79050 , n79049 );
buf ( n79051 , n79050 );
nand ( n79052 , n79046 , n79051 );
buf ( n79053 , n79052 );
buf ( n79054 , n79053 );
and ( n79055 , n79026 , n79054 );
and ( n79056 , n79000 , n79025 );
or ( n79057 , n79055 , n79056 );
buf ( n79058 , n79057 );
xor ( n79059 , n78997 , n79058 );
buf ( n79060 , n48865 );
not ( n79061 , n79060 );
buf ( n79062 , n78979 );
not ( n79063 , n79062 );
or ( n79064 , n79061 , n79063 );
buf ( n79065 , n48808 );
buf ( n79066 , n42856 );
and ( n79067 , n79065 , n79066 );
not ( n79068 , n79065 );
buf ( n79069 , n72235 );
and ( n79070 , n79068 , n79069 );
nor ( n79071 , n79067 , n79070 );
buf ( n79072 , n79071 );
buf ( n79073 , n79072 );
buf ( n79074 , n48852 );
nand ( n79075 , n79073 , n79074 );
buf ( n79076 , n79075 );
buf ( n79077 , n79076 );
nand ( n79078 , n79064 , n79077 );
buf ( n79079 , n79078 );
and ( n79080 , n79059 , n79079 );
and ( n79081 , n78997 , n79058 );
or ( n79082 , n79080 , n79081 );
buf ( n79083 , n79082 );
and ( n79084 , n78992 , n79083 );
and ( n79085 , n78987 , n78991 );
or ( n79086 , n79084 , n79085 );
buf ( n79087 , n79086 );
buf ( n79088 , n79087 );
xor ( n79089 , n77970 , n78368 );
xor ( n79090 , n79089 , n78394 );
buf ( n79091 , n79090 );
buf ( n79092 , n79091 );
buf ( n79093 , n56289 );
buf ( n79094 , n25306 );
and ( n79095 , n79093 , n79094 );
not ( n79096 , n79093 );
buf ( n79097 , n25293 );
and ( n79098 , n79096 , n79097 );
nor ( n79099 , n79095 , n79098 );
buf ( n79100 , n79099 );
buf ( n79101 , n79100 );
not ( n79102 , n79101 );
buf ( n79103 , n42246 );
not ( n79104 , n79103 );
or ( n79105 , n79102 , n79104 );
buf ( n79106 , n77936 );
buf ( n79107 , n42309 );
nand ( n79108 , n79106 , n79107 );
buf ( n79109 , n79108 );
buf ( n79110 , n79109 );
nand ( n79111 , n79105 , n79110 );
buf ( n79112 , n79111 );
buf ( n79113 , n79112 );
xor ( n79114 , n79092 , n79113 );
buf ( n79115 , n63913 );
not ( n79116 , n24926 );
not ( n79117 , n25226 );
or ( n79118 , n79116 , n79117 );
buf ( n79119 , n24926 );
buf ( n79120 , n25226 );
nor ( n79121 , n79119 , n79120 );
buf ( n79122 , n79121 );
or ( n79123 , n79122 , n56325 );
nand ( n79124 , n79118 , n79123 );
buf ( n79125 , n79124 );
nor ( n79126 , n79115 , n79125 );
buf ( n79127 , n79126 );
buf ( n79128 , n79127 );
and ( n79129 , n79114 , n79128 );
and ( n79130 , n79092 , n79113 );
or ( n79131 , n79129 , n79130 );
buf ( n79132 , n79131 );
buf ( n79133 , n79132 );
xor ( n79134 , n79088 , n79133 );
buf ( n79135 , n42375 );
buf ( n79136 , n55841 );
not ( n79137 , n79136 );
buf ( n79138 , n42342 );
not ( n79139 , n79138 );
or ( n79140 , n79137 , n79139 );
buf ( n79141 , n24951 );
buf ( n79142 , n55840 );
nand ( n79143 , n79141 , n79142 );
buf ( n79144 , n79143 );
buf ( n79145 , n79144 );
nand ( n79146 , n79140 , n79145 );
buf ( n79147 , n79146 );
buf ( n79148 , n79147 );
not ( n79149 , n79148 );
buf ( n79150 , n79149 );
buf ( n79151 , n79150 );
or ( n79152 , n79135 , n79151 );
buf ( n79153 , n78755 );
not ( n79154 , n79153 );
buf ( n79155 , n79154 );
buf ( n79156 , n79155 );
buf ( n79157 , n42333 );
or ( n79158 , n79156 , n79157 );
nand ( n79159 , n79152 , n79158 );
buf ( n79160 , n79159 );
buf ( n79161 , n79160 );
and ( n79162 , n79134 , n79161 );
and ( n79163 , n79088 , n79133 );
or ( n79164 , n79162 , n79163 );
buf ( n79165 , n79164 );
buf ( n79166 , n79165 );
xor ( n79167 , n78962 , n79166 );
buf ( n79168 , n62125 );
not ( n79169 , n79168 );
buf ( n79170 , n78476 );
not ( n79171 , n79170 );
or ( n79172 , n79169 , n79171 );
buf ( n79173 , n48836 );
not ( n79174 , n79173 );
buf ( n79175 , n41733 );
not ( n79176 , n79175 );
or ( n79177 , n79174 , n79176 );
buf ( n79178 , n60327 );
buf ( n79179 , n72931 );
nand ( n79180 , n79178 , n79179 );
buf ( n79181 , n79180 );
buf ( n79182 , n79181 );
nand ( n79183 , n79177 , n79182 );
buf ( n79184 , n79183 );
buf ( n79185 , n79184 );
buf ( n79186 , n51488 );
nand ( n79187 , n79185 , n79186 );
buf ( n79188 , n79187 );
buf ( n79189 , n79188 );
nand ( n79190 , n79172 , n79189 );
buf ( n79191 , n79190 );
buf ( n79192 , n79191 );
and ( n79193 , n79167 , n79192 );
and ( n79194 , n78962 , n79166 );
or ( n79195 , n79193 , n79194 );
buf ( n79196 , n79195 );
buf ( n79197 , n79196 );
and ( n79198 , n78945 , n79197 );
or ( n79199 , n79198 , C0 );
buf ( n79200 , n79199 );
buf ( n79201 , n79200 );
and ( n79202 , n78938 , n79201 );
buf ( n79203 , C0 );
buf ( n79204 , n79203 );
nor ( n79205 , n79202 , n79204 );
buf ( n79206 , n79205 );
not ( n79207 , n79206 );
xor ( n79208 , n77891 , n77898 );
xor ( n79209 , n79208 , n77900 );
buf ( n79210 , n79209 );
not ( n79211 , n79210 );
or ( n79212 , n79207 , n79211 );
or ( n79213 , n79210 , n79206 );
xor ( n79214 , n77206 , n77806 );
xnor ( n79215 , n79214 , n77202 );
not ( n79216 , n79215 );
nand ( n79217 , n79213 , n79216 );
nand ( n79218 , n79212 , n79217 );
buf ( n79219 , n78893 );
buf ( n79220 , n78910 );
and ( n79221 , n79219 , n79220 );
not ( n79222 , n79219 );
buf ( n79223 , n78898 );
and ( n79224 , n79222 , n79223 );
nor ( n79225 , n79221 , n79224 );
buf ( n79226 , n79225 );
xor ( n79227 , n79226 , n78904 );
xor ( n79228 , n79218 , n79227 );
xor ( n79229 , n77904 , n78872 );
xnor ( n79230 , n79229 , n77914 );
and ( n79231 , n79228 , n79230 );
and ( n79232 , n79218 , n79227 );
or ( n79233 , n79231 , n79232 );
buf ( n79234 , n79233 );
nand ( n79235 , n78926 , n79234 );
buf ( n79236 , n79235 );
not ( n79237 , n79236 );
xor ( n79238 , n79218 , n79227 );
xor ( n79239 , n79238 , n79230 );
buf ( n79240 , n79239 );
not ( n79241 , n79240 );
buf ( n79242 , n79241 );
buf ( n79243 , n79242 );
buf ( n79244 , n78864 );
not ( n79245 , n79244 );
buf ( n79246 , n78558 );
not ( n79247 , n79246 );
or ( n79248 , n79245 , n79247 );
buf ( n79249 , n77923 );
buf ( n79250 , n78868 );
nand ( n79251 , n79249 , n79250 );
buf ( n79252 , n79251 );
buf ( n79253 , n79252 );
nand ( n79254 , n79248 , n79253 );
buf ( n79255 , n79254 );
buf ( n79256 , n79255 );
buf ( n79257 , n78860 );
buf ( n79258 , n79257 );
buf ( n79259 , n79258 );
buf ( n79260 , n79259 );
xnor ( n79261 , n79256 , n79260 );
buf ( n79262 , n79261 );
not ( n79263 , n79262 );
not ( n79264 , n79210 );
xor ( n79265 , n79215 , n79264 );
xnor ( n79266 , n79265 , n79206 );
not ( n79267 , n79266 );
not ( n79268 , n79267 );
or ( n79269 , n79263 , n79268 );
buf ( n79270 , n78543 );
buf ( n79271 , n78498 );
xor ( n79272 , n79270 , n79271 );
buf ( n79273 , n78488 );
xor ( n79274 , n79272 , n79273 );
buf ( n79275 , n79274 );
not ( n79276 , n79275 );
xor ( n79277 , n78454 , n78458 );
xor ( n79278 , n79277 , n78484 );
buf ( n79279 , n79278 );
buf ( n79280 , n79279 );
not ( n79281 , n78848 );
not ( n79282 , n78562 );
not ( n79283 , n78772 );
and ( n79284 , n79282 , n79283 );
and ( n79285 , n78562 , n78772 );
nor ( n79286 , n79284 , n79285 );
not ( n79287 , n79286 );
or ( n79288 , n79281 , n79287 );
or ( n79289 , n79286 , n78848 );
nand ( n79290 , n79288 , n79289 );
buf ( n79291 , n79290 );
buf ( n79292 , C0 );
buf ( n79293 , n79292 );
and ( n79294 , n79280 , n79291 );
or ( n79295 , C0 , n79294 );
buf ( n79296 , n79295 );
not ( n79297 , n79296 );
or ( n79298 , n79276 , n79297 );
not ( n79299 , n79275 );
not ( n79300 , n79299 );
not ( n79301 , n79296 );
not ( n79302 , n79301 );
or ( n79303 , n79300 , n79302 );
xor ( n79304 , n78851 , n78855 );
xor ( n79305 , n79304 , n78857 );
buf ( n79306 , n79305 );
nand ( n79307 , n79303 , n79306 );
nand ( n79308 , n79298 , n79307 );
nand ( n79309 , n79269 , n79308 );
buf ( n79310 , n79309 );
buf ( n79311 , n79262 );
not ( n79312 , n79311 );
buf ( n79313 , n79266 );
nand ( n79314 , n79312 , n79313 );
buf ( n79315 , n79314 );
buf ( n79316 , n79315 );
and ( n79317 , n79310 , n79316 );
buf ( n79318 , n79317 );
buf ( n79319 , n79318 );
not ( n79320 , n79319 );
buf ( n79321 , n79320 );
buf ( n79322 , n79321 );
nand ( n79323 , n79243 , n79322 );
buf ( n79324 , n79323 );
buf ( n79325 , n79324 );
not ( n79326 , n79266 );
not ( n79327 , n79275 );
not ( n79328 , n79296 );
or ( n79329 , n79327 , n79328 );
nand ( n79330 , n79329 , n79307 );
not ( n79331 , n79330 );
not ( n79332 , n79262 );
or ( n79333 , n79331 , n79332 );
or ( n79334 , n79262 , n79308 );
nand ( n79335 , n79333 , n79334 );
or ( n79336 , n79326 , n79335 );
not ( n79337 , n79266 );
nand ( n79338 , n79337 , n79335 );
nand ( n79339 , n79336 , n79338 );
xnor ( n79340 , n78927 , n78934 );
xor ( n79341 , n79200 , n79340 );
not ( n79342 , n79341 );
xnor ( n79343 , n78742 , n78718 );
buf ( n79344 , n79343 );
buf ( n79345 , n78763 );
and ( n79346 , n79344 , n79345 );
not ( n79347 , n79344 );
buf ( n79348 , n78764 );
and ( n79349 , n79347 , n79348 );
nor ( n79350 , n79346 , n79349 );
buf ( n79351 , n79350 );
buf ( n79352 , n79351 );
xor ( n79353 , n78566 , n78693 );
xor ( n79354 , n79353 , n78714 );
buf ( n79355 , n79354 );
buf ( n79356 , n79355 );
buf ( n79357 , n60545 );
not ( n79358 , n79357 );
buf ( n79359 , n79184 );
not ( n79360 , n79359 );
or ( n79361 , n79358 , n79360 );
buf ( n79362 , n48836 );
not ( n79363 , n79362 );
buf ( n79364 , n41721 );
not ( n79365 , n79364 );
or ( n79366 , n79363 , n79365 );
buf ( n79367 , n13662 );
buf ( n79368 , n72931 );
nand ( n79369 , n79367 , n79368 );
buf ( n79370 , n79369 );
buf ( n79371 , n79370 );
nand ( n79372 , n79366 , n79371 );
buf ( n79373 , n79372 );
buf ( n79374 , n79373 );
buf ( n79375 , n51488 );
nand ( n79376 , n79374 , n79375 );
buf ( n79377 , n79376 );
buf ( n79378 , n79377 );
nand ( n79379 , n79361 , n79378 );
buf ( n79380 , n79379 );
buf ( n79381 , n79380 );
xor ( n79382 , n79356 , n79381 );
xor ( n79383 , n78632 , n78657 );
xor ( n79384 , n79383 , n78683 );
buf ( n79385 , n79384 );
buf ( n79386 , n79385 );
buf ( n79387 , n52780 );
not ( n79388 , n79387 );
buf ( n79389 , n25303 );
not ( n79390 , n79389 );
or ( n79391 , n79388 , n79390 );
buf ( n79392 , n52789 );
buf ( n79393 , n25290 );
nand ( n79394 , n79392 , n79393 );
buf ( n79395 , n79394 );
buf ( n79396 , n79395 );
nand ( n79397 , n79391 , n79396 );
buf ( n79398 , n79397 );
buf ( n79399 , n79398 );
not ( n79400 , n79399 );
buf ( n79401 , n42246 );
not ( n79402 , n79401 );
or ( n79403 , n79400 , n79402 );
buf ( n79404 , n79100 );
buf ( n79405 , n42309 );
nand ( n79406 , n79404 , n79405 );
buf ( n79407 , n79406 );
buf ( n79408 , n79407 );
nand ( n79409 , n79403 , n79408 );
buf ( n79410 , n79409 );
buf ( n79411 , n79410 );
xor ( n79412 , n79386 , n79411 );
xor ( n79413 , n77594 , n77707 );
xor ( n79414 , n79413 , n77711 );
xor ( n79415 , n78147 , n78282 );
xor ( n79416 , n79414 , n79415 );
buf ( n79417 , n79416 );
buf ( n79418 , n71078 );
not ( n79419 , n79418 );
buf ( n79420 , n76179 );
not ( n79421 , n79420 );
or ( n79422 , n79419 , n79421 );
buf ( n79423 , n48320 );
buf ( n79424 , n45746 );
nand ( n79425 , n79423 , n79424 );
buf ( n79426 , n79425 );
buf ( n79427 , n79426 );
nand ( n79428 , n79422 , n79427 );
buf ( n79429 , n79428 );
buf ( n79430 , n79429 );
not ( n79431 , n79430 );
buf ( n79432 , n45741 );
not ( n79433 , n79432 );
or ( n79434 , n79431 , n79433 );
buf ( n79435 , n78300 );
buf ( n79436 , n67149 );
nand ( n79437 , n79435 , n79436 );
buf ( n79438 , n79437 );
buf ( n79439 , n79438 );
nand ( n79440 , n79434 , n79439 );
buf ( n79441 , n79440 );
buf ( n79442 , n79441 );
xor ( n79443 , n79417 , n79442 );
buf ( n79444 , n46912 );
not ( n79445 , n79444 );
buf ( n79446 , n79017 );
not ( n79447 , n79446 );
or ( n79448 , n79445 , n79447 );
buf ( n79449 , n46875 );
not ( n79450 , n79449 );
buf ( n79451 , n46387 );
not ( n79452 , n79451 );
or ( n79453 , n79450 , n79452 );
buf ( n79454 , n78314 );
buf ( n79455 , n46887 );
nand ( n79456 , n79454 , n79455 );
buf ( n79457 , n79456 );
buf ( n79458 , n79457 );
nand ( n79459 , n79453 , n79458 );
buf ( n79460 , n79459 );
buf ( n79461 , n79460 );
buf ( n79462 , n46907 );
nand ( n79463 , n79461 , n79462 );
buf ( n79464 , n79463 );
buf ( n79465 , n79464 );
nand ( n79466 , n79448 , n79465 );
buf ( n79467 , n79466 );
buf ( n79468 , n79467 );
and ( n79469 , n79443 , n79468 );
and ( n79470 , n79417 , n79442 );
or ( n79471 , n79469 , n79470 );
buf ( n79472 , n79471 );
buf ( n79473 , n79472 );
buf ( n79474 , n56289 );
not ( n79475 , n79474 );
buf ( n79476 , n77077 );
not ( n79477 , n79476 );
or ( n79478 , n79475 , n79477 );
buf ( n79479 , n42228 );
buf ( n79480 , n52094 );
nand ( n79481 , n79479 , n79480 );
buf ( n79482 , n79481 );
buf ( n79483 , n79482 );
nand ( n79484 , n79478 , n79483 );
buf ( n79485 , n79484 );
buf ( n79486 , n79485 );
not ( n79487 , n79486 );
buf ( n79488 , n41596 );
not ( n79489 , n79488 );
or ( n79490 , n79487 , n79489 );
buf ( n79491 , n78670 );
buf ( n79492 , n41574 );
nand ( n79493 , n79491 , n79492 );
buf ( n79494 , n79493 );
buf ( n79495 , n79494 );
nand ( n79496 , n79490 , n79495 );
buf ( n79497 , n79496 );
buf ( n79498 , n79497 );
xor ( n79499 , n79473 , n79498 );
xor ( n79500 , n79000 , n79025 );
xor ( n79501 , n79500 , n79054 );
buf ( n79502 , n79501 );
buf ( n79503 , n79502 );
and ( n79504 , n79499 , n79503 );
and ( n79505 , n79473 , n79498 );
or ( n79506 , n79504 , n79505 );
buf ( n79507 , n79506 );
buf ( n79508 , n79507 );
and ( n79509 , n79412 , n79508 );
and ( n79510 , n79386 , n79411 );
or ( n79511 , n79509 , n79510 );
buf ( n79512 , n79511 );
buf ( n79513 , n79512 );
buf ( n79514 , n53539 );
not ( n79515 , n79514 );
buf ( n79516 , n62510 );
not ( n79517 , n79516 );
or ( n79518 , n79515 , n79517 );
buf ( n79519 , n25226 );
buf ( n79520 , n53548 );
nand ( n79521 , n79519 , n79520 );
buf ( n79522 , n79521 );
buf ( n79523 , n79522 );
nand ( n79524 , n79518 , n79523 );
buf ( n79525 , n79524 );
buf ( n79526 , n79525 );
not ( n79527 , n79526 );
buf ( n79528 , n73163 );
not ( n79529 , n79528 );
or ( n79530 , n79527 , n79529 );
buf ( n79531 , n78703 );
not ( n79532 , n79531 );
buf ( n79533 , n42665 );
nand ( n79534 , n79532 , n79533 );
buf ( n79535 , n79534 );
buf ( n79536 , n79535 );
nand ( n79537 , n79530 , n79536 );
buf ( n79538 , n79537 );
buf ( n79539 , n79538 );
xor ( n79540 , n79513 , n79539 );
xor ( n79541 , n79092 , n79113 );
xor ( n79542 , n79541 , n79128 );
buf ( n79543 , n79542 );
buf ( n79544 , n79543 );
and ( n79545 , n79540 , n79544 );
and ( n79546 , n79513 , n79539 );
or ( n79547 , n79545 , n79546 );
buf ( n79548 , n79547 );
buf ( n79549 , n79548 );
and ( n79550 , n79382 , n79549 );
and ( n79551 , n79356 , n79381 );
or ( n79552 , n79550 , n79551 );
buf ( n79553 , n79552 );
buf ( n79554 , n79553 );
buf ( n79555 , C0 );
buf ( n79556 , n79555 );
and ( n79557 , n79352 , n79554 );
or ( n79558 , C0 , n79557 );
buf ( n79559 , n79558 );
not ( n79560 , n79559 );
not ( n79561 , n79560 );
not ( n79562 , n79561 );
xor ( n79563 , n78781 , n78839 );
xor ( n79564 , n79563 , n78844 );
buf ( n79565 , n79564 );
buf ( n79566 , n79565 );
xnor ( n79567 , n78811 , n78824 );
buf ( n79568 , n79567 );
buf ( n79569 , n78831 );
and ( n79570 , n79568 , n79569 );
not ( n79571 , n79568 );
buf ( n79572 , n78818 );
and ( n79573 , n79571 , n79572 );
nor ( n79574 , n79570 , n79573 );
buf ( n79575 , n79574 );
buf ( n79576 , n79575 );
buf ( n79577 , C0 );
buf ( n79578 , n79577 );
xor ( n79579 , n79576 , n79578 );
buf ( n79580 , n12481 );
not ( n79581 , n79580 );
buf ( n79582 , n42331 );
nor ( n79583 , n79581 , n79582 );
buf ( n79584 , n79583 );
buf ( n79585 , n79584 );
buf ( n79586 , n50995 );
not ( n79587 , n79586 );
buf ( n79588 , n25382 );
not ( n79589 , n79588 );
or ( n79590 , n79587 , n79589 );
buf ( n79591 , n41570 );
buf ( n79592 , n50992 );
nand ( n79593 , n79591 , n79592 );
buf ( n79594 , n79593 );
buf ( n79595 , n79594 );
nand ( n79596 , n79590 , n79595 );
buf ( n79597 , n79596 );
buf ( n79598 , n79597 );
not ( n79599 , n79598 );
buf ( n79600 , n74488 );
not ( n79601 , n79600 );
or ( n79602 , n79599 , n79601 );
buf ( n79603 , n44496 );
buf ( n79604 , n79041 );
nand ( n79605 , n79603 , n79604 );
buf ( n79606 , n79605 );
buf ( n79607 , n79606 );
nand ( n79608 , n79602 , n79607 );
buf ( n79609 , n79608 );
buf ( n79610 , n79609 );
xor ( n79611 , n77607 , n77623 );
xor ( n79612 , n79611 , n77650 );
xor ( n79613 , n78110 , n78132 );
xor ( n79614 , n79612 , n79613 );
buf ( n79615 , n79614 );
not ( n79616 , n68273 );
not ( n79617 , n78124 );
or ( n79618 , n79616 , n79617 );
not ( n79619 , n64141 );
not ( n79620 , n64133 );
not ( n79621 , n70336 );
or ( n79622 , n79620 , n79621 );
nand ( n79623 , n64129 , n70333 );
nand ( n79624 , n79622 , n79623 );
nand ( n79625 , n79619 , n79624 );
nand ( n79626 , n79618 , n79625 );
buf ( n79627 , n56639 );
buf ( n79628 , n75821 );
nor ( n79629 , n79627 , n79628 );
buf ( n79630 , n79629 );
buf ( n79631 , n79630 );
buf ( n79632 , n60270 );
buf ( n79633 , n15265 );
buf ( n79634 , n71801 );
and ( n79635 , n79633 , n79634 );
buf ( n79636 , n60090 );
buf ( n79637 , n71804 );
and ( n79638 , n79636 , n79637 );
nor ( n79639 , n79635 , n79638 );
buf ( n79640 , n79639 );
buf ( n79641 , n79640 );
or ( n79642 , n79632 , n79641 );
buf ( n79643 , n78179 );
buf ( n79644 , n60100 );
or ( n79645 , n79643 , n79644 );
nand ( n79646 , n79642 , n79645 );
buf ( n79647 , n79646 );
buf ( n79648 , n79647 );
and ( n79649 , n79631 , n79648 );
buf ( n79650 , n79649 );
buf ( n79651 , n58913 );
buf ( n79652 , n58897 );
buf ( n79653 , n71818 );
and ( n79654 , n79652 , n79653 );
buf ( n79655 , n58894 );
buf ( n79656 , n71821 );
and ( n79657 , n79655 , n79656 );
nor ( n79658 , n79654 , n79657 );
buf ( n79659 , n79658 );
buf ( n79660 , n79659 );
or ( n79661 , n79651 , n79660 );
buf ( n79662 , n77637 );
not ( n79663 , n79662 );
buf ( n79664 , n79663 );
buf ( n79665 , n79664 );
buf ( n79666 , n58884 );
or ( n79667 , n79665 , n79666 );
nand ( n79668 , n79661 , n79667 );
buf ( n79669 , n79668 );
xor ( n79670 , n79650 , n79669 );
buf ( n79671 , n56634 );
buf ( n79672 , n623 );
or ( n79673 , n79671 , n79672 );
buf ( n79674 , n56629 );
buf ( n79675 , n56641 );
buf ( n79676 , n623 );
and ( n79677 , n79674 , n79675 , n79676 );
buf ( n79678 , n56644 );
nor ( n79679 , n79677 , n79678 );
buf ( n79680 , n79679 );
buf ( n79681 , n79680 );
nand ( n79682 , n79673 , n79681 );
buf ( n79683 , n79682 );
and ( n79684 , n79670 , n79683 );
and ( n79685 , n79650 , n79669 );
or ( n79686 , n79684 , n79685 );
xor ( n79687 , n79626 , n79686 );
xor ( n79688 , n77996 , n78013 );
xor ( n79689 , n79688 , n78036 );
buf ( n79690 , n79689 );
and ( n79691 , n79687 , n79690 );
and ( n79692 , n79626 , n79686 );
or ( n79693 , n79691 , n79692 );
buf ( n79694 , n79693 );
xor ( n79695 , n79615 , n79694 );
buf ( n79696 , n71232 );
buf ( n79697 , n60096 );
and ( n79698 , n79696 , n79697 );
buf ( n79699 , n71235 );
buf ( n79700 , n62663 );
and ( n79701 , n79699 , n79700 );
nor ( n79702 , n79698 , n79701 );
buf ( n79703 , n79702 );
buf ( n79704 , n79703 );
buf ( n79705 , n62935 );
or ( n79706 , n79704 , n79705 );
buf ( n79707 , n78234 );
not ( n79708 , n79707 );
buf ( n79709 , n79708 );
buf ( n79710 , n79709 );
buf ( n79711 , n62676 );
or ( n79712 , n79710 , n79711 );
nand ( n79713 , n79706 , n79712 );
buf ( n79714 , n79713 );
xor ( n79715 , n78186 , n78199 );
xor ( n79716 , n79715 , n78216 );
and ( n79717 , n79714 , n79716 );
buf ( n79718 , n71225 );
buf ( n79719 , n62681 );
and ( n79720 , n79718 , n79719 );
buf ( n79721 , n71228 );
buf ( n79722 , n62684 );
and ( n79723 , n79721 , n79722 );
nor ( n79724 , n79720 , n79723 );
buf ( n79725 , n79724 );
buf ( n79726 , n79725 );
buf ( n79727 , n62935 );
or ( n79728 , n79726 , n79727 );
buf ( n79729 , n79703 );
buf ( n79730 , n62676 );
or ( n79731 , n79729 , n79730 );
nand ( n79732 , n79728 , n79731 );
buf ( n79733 , n79732 );
buf ( n79734 , n79733 );
buf ( n79735 , n58897 );
buf ( n79736 , n72445 );
and ( n79737 , n79735 , n79736 );
buf ( n79738 , n58894 );
buf ( n79739 , n72448 );
and ( n79740 , n79738 , n79739 );
nor ( n79741 , n79737 , n79740 );
buf ( n79742 , n79741 );
buf ( n79743 , n79742 );
buf ( n79744 , n58913 );
or ( n79745 , n79743 , n79744 );
buf ( n79746 , n79659 );
buf ( n79747 , n58884 );
or ( n79748 , n79746 , n79747 );
nand ( n79749 , n79745 , n79748 );
buf ( n79750 , n79749 );
buf ( n79751 , n79750 );
xor ( n79752 , n79734 , n79751 );
buf ( n79753 , n78209 );
buf ( n79754 , n58982 );
or ( n79755 , n79753 , n79754 );
buf ( n79756 , n56807 );
nand ( n79757 , n79755 , n79756 );
buf ( n79758 , n79757 );
buf ( n79759 , n79758 );
and ( n79760 , n79752 , n79759 );
and ( n79761 , n79734 , n79751 );
or ( n79762 , n79760 , n79761 );
buf ( n79763 , n79762 );
xor ( n79764 , n78186 , n78199 );
xor ( n79765 , n79764 , n78216 );
and ( n79766 , n79763 , n79765 );
and ( n79767 , n79714 , n79763 );
or ( n79768 , n79717 , n79766 , n79767 );
buf ( n79769 , n79768 );
buf ( n79770 , n68217 );
buf ( n79771 , n66742 );
and ( n79772 , n79770 , n79771 );
buf ( n79773 , n68220 );
buf ( n79774 , n63000 );
and ( n79775 , n79773 , n79774 );
nor ( n79776 , n79772 , n79775 );
buf ( n79777 , n79776 );
buf ( n79778 , n79777 );
buf ( n79779 , n64230 );
or ( n79780 , n79778 , n79779 );
buf ( n79781 , n78161 );
buf ( n79782 , n64227 );
or ( n79783 , n79781 , n79782 );
nand ( n79784 , n79780 , n79783 );
buf ( n79785 , n79784 );
buf ( n79786 , n79785 );
xor ( n79787 , n79769 , n79786 );
xor ( n79788 , n78220 , n78223 );
xor ( n79789 , n79788 , n78243 );
buf ( n79790 , n79789 );
buf ( n79791 , n79790 );
and ( n79792 , n79787 , n79791 );
and ( n79793 , n79769 , n79786 );
or ( n79794 , n79792 , n79793 );
buf ( n79795 , n79794 );
buf ( n79796 , n79795 );
and ( n79797 , n79695 , n79796 );
and ( n79798 , n79615 , n79694 );
or ( n79799 , n79797 , n79798 );
buf ( n79800 , n79799 );
xor ( n79801 , n78153 , n78258 );
xor ( n79802 , n79801 , n78263 );
and ( n79803 , n79800 , n79802 );
buf ( n79804 , n70348 );
buf ( n79805 , n64129 );
and ( n79806 , n79804 , n79805 );
buf ( n79807 , n70351 );
buf ( n79808 , n64133 );
and ( n79809 , n79807 , n79808 );
nor ( n79810 , n79806 , n79809 );
buf ( n79811 , n79810 );
or ( n79812 , n79811 , n64141 );
nand ( n79813 , n79624 , n68273 );
nand ( n79814 , n79812 , n79813 );
xor ( n79815 , n79650 , n79669 );
xor ( n79816 , n79815 , n79683 );
and ( n79817 , n79814 , n79816 );
buf ( n79818 , n68232 );
buf ( n79819 , n66742 );
and ( n79820 , n79818 , n79819 );
buf ( n79821 , n68235 );
buf ( n79822 , n63000 );
and ( n79823 , n79821 , n79822 );
nor ( n79824 , n79820 , n79823 );
buf ( n79825 , n79824 );
buf ( n79826 , n79825 );
buf ( n79827 , n64230 );
or ( n79828 , n79826 , n79827 );
buf ( n79829 , n79777 );
buf ( n79830 , n64227 );
or ( n79831 , n79829 , n79830 );
nand ( n79832 , n79828 , n79831 );
buf ( n79833 , n79832 );
xor ( n79834 , n79650 , n79669 );
xor ( n79835 , n79834 , n79683 );
and ( n79836 , n79833 , n79835 );
and ( n79837 , n79814 , n79833 );
or ( n79838 , n79817 , n79836 , n79837 );
xor ( n79839 , n79626 , n79686 );
xor ( n79840 , n79839 , n79690 );
and ( n79841 , n79838 , n79840 );
xor ( n79842 , n79769 , n79786 );
xor ( n79843 , n79842 , n79791 );
buf ( n79844 , n79843 );
xor ( n79845 , n79626 , n79686 );
xor ( n79846 , n79845 , n79690 );
and ( n79847 , n79844 , n79846 );
and ( n79848 , n79838 , n79844 );
or ( n79849 , n79841 , n79847 , n79848 );
buf ( n79850 , n79849 );
xor ( n79851 , n78170 , n78248 );
xor ( n79852 , n79851 , n78254 );
buf ( n79853 , n79852 );
buf ( n79854 , n79853 );
xor ( n79855 , n79850 , n79854 );
xor ( n79856 , n79615 , n79694 );
xor ( n79857 , n79856 , n79796 );
buf ( n79858 , n79857 );
buf ( n79859 , n79858 );
and ( n79860 , n79855 , n79859 );
and ( n79861 , n79850 , n79854 );
or ( n79862 , n79860 , n79861 );
buf ( n79863 , n79862 );
xor ( n79864 , n78153 , n78258 );
xor ( n79865 , n79864 , n78263 );
and ( n79866 , n79863 , n79865 );
and ( n79867 , n79800 , n79863 );
or ( n79868 , n79803 , n79866 , n79867 );
buf ( n79869 , n79868 );
xor ( n79870 , n78267 , n78272 );
xor ( n79871 , n79870 , n78278 );
buf ( n79872 , n79871 );
buf ( n79873 , n79872 );
xor ( n79874 , n79869 , n79873 );
not ( n79875 , n50059 );
not ( n79876 , n79875 );
not ( n79877 , n76179 );
or ( n79878 , n79876 , n79877 );
buf ( n79879 , n44494 );
buf ( n79880 , n79875 );
not ( n79881 , n79880 );
buf ( n79882 , n79881 );
buf ( n79883 , n79882 );
nand ( n79884 , n79879 , n79883 );
buf ( n79885 , n79884 );
nand ( n79886 , n79878 , n79885 );
not ( n79887 , n79886 );
not ( n79888 , n45741 );
or ( n79889 , n79887 , n79888 );
buf ( n79890 , n46246 );
buf ( n79891 , n79429 );
nand ( n79892 , n79890 , n79891 );
buf ( n79893 , n79892 );
nand ( n79894 , n79889 , n79893 );
buf ( n79895 , n79894 );
and ( n79896 , n79874 , n79895 );
and ( n79897 , n79869 , n79873 );
or ( n79898 , n79896 , n79897 );
buf ( n79899 , n79898 );
buf ( n79900 , n79899 );
or ( n79901 , n79610 , n79900 );
xor ( n79902 , n79417 , n79442 );
xor ( n79903 , n79902 , n79468 );
buf ( n79904 , n79903 );
buf ( n79905 , n79904 );
nand ( n79906 , n79901 , n79905 );
buf ( n79907 , n79906 );
buf ( n79908 , n79907 );
buf ( n79909 , n79609 );
buf ( n79910 , n79899 );
nand ( n79911 , n79909 , n79910 );
buf ( n79912 , n79911 );
buf ( n79913 , n79912 );
nand ( n79914 , n79908 , n79913 );
buf ( n79915 , n79914 );
buf ( n79916 , n79915 );
buf ( n79917 , n48865 );
not ( n79918 , n79917 );
buf ( n79919 , n79072 );
not ( n79920 , n79919 );
or ( n79921 , n79918 , n79920 );
buf ( n79922 , n48852 );
buf ( n79923 , n48808 );
not ( n79924 , n79923 );
buf ( n79925 , n74460 );
not ( n79926 , n79925 );
or ( n79927 , n79924 , n79926 );
buf ( n79928 , n42844 );
buf ( n79929 , n72891 );
nand ( n79930 , n79928 , n79929 );
buf ( n79931 , n79930 );
buf ( n79932 , n79931 );
nand ( n79933 , n79927 , n79932 );
buf ( n79934 , n79933 );
buf ( n79935 , n79934 );
nand ( n79936 , n79922 , n79935 );
buf ( n79937 , n79936 );
buf ( n79938 , n79937 );
nand ( n79939 , n79921 , n79938 );
buf ( n79940 , n79939 );
buf ( n79941 , n79940 );
xor ( n79942 , n79916 , n79941 );
buf ( n79943 , n25226 );
not ( n79944 , n79943 );
not ( n79945 , n25257 );
not ( n79946 , n71123 );
or ( n79947 , n79945 , n79946 );
buf ( n79948 , n25257 );
buf ( n79949 , n71123 );
nor ( n79950 , n79948 , n79949 );
buf ( n79951 , n79950 );
or ( n79952 , n79951 , n56325 );
nand ( n79953 , n79947 , n79952 );
buf ( n79954 , n79953 );
nor ( n79955 , n79944 , n79954 );
buf ( n79956 , n79955 );
buf ( n79957 , n79956 );
and ( n79958 , n79942 , n79957 );
and ( n79959 , n79916 , n79941 );
or ( n79960 , n79958 , n79959 );
buf ( n79961 , n79960 );
buf ( n79962 , n79961 );
xor ( n79963 , n79585 , n79962 );
xor ( n79964 , n78997 , n79058 );
xor ( n79965 , n79964 , n79079 );
buf ( n79966 , n79965 );
and ( n79967 , n79963 , n79966 );
and ( n79968 , n79585 , n79962 );
or ( n79969 , n79967 , n79968 );
buf ( n79970 , n79969 );
buf ( n79971 , n79970 );
buf ( n79972 , n12481 );
buf ( n79973 , n42366 );
and ( n79974 , n79972 , n79973 );
not ( n79975 , n79972 );
buf ( n79976 , n63913 );
and ( n79977 , n79975 , n79976 );
nor ( n79978 , n79974 , n79977 );
buf ( n79979 , n79978 );
buf ( n79980 , n79979 );
not ( n79981 , n79980 );
buf ( n79982 , n66459 );
not ( n79983 , n79982 );
or ( n79984 , n79981 , n79983 );
buf ( n79985 , n79147 );
buf ( n79986 , n42336 );
nand ( n79987 , n79985 , n79986 );
buf ( n79988 , n79987 );
buf ( n79989 , n79988 );
nand ( n79990 , n79984 , n79989 );
buf ( n79991 , n79990 );
buf ( n79992 , n79991 );
xor ( n79993 , n79971 , n79992 );
buf ( n79994 , n60545 );
not ( n79995 , n79994 );
buf ( n79996 , n79373 );
not ( n79997 , n79996 );
or ( n79998 , n79995 , n79997 );
and ( n79999 , n48836 , n70855 );
not ( n80000 , n48836 );
and ( n80001 , n80000 , n29463 );
or ( n80002 , n79999 , n80001 );
buf ( n80003 , n80002 );
buf ( n80004 , n51488 );
nand ( n80005 , n80003 , n80004 );
buf ( n80006 , n80005 );
buf ( n80007 , n80006 );
nand ( n80008 , n79998 , n80007 );
buf ( n80009 , n80008 );
buf ( n80010 , n80009 );
and ( n80011 , n79993 , n80010 );
and ( n80012 , n79971 , n79992 );
or ( n80013 , n80011 , n80012 );
buf ( n80014 , n80013 );
buf ( n80015 , n80014 );
and ( n80016 , n79579 , n80015 );
or ( n80017 , n80016 , C0 );
buf ( n80018 , n80017 );
buf ( n80019 , n80018 );
buf ( n80020 , C0 );
buf ( n80021 , n80020 );
and ( n80022 , n79566 , n80019 );
or ( n80023 , C0 , n80022 );
buf ( n80024 , n80023 );
not ( n80025 , n80024 );
or ( n80026 , n79562 , n80025 );
not ( n80027 , n79560 );
not ( n80028 , n80024 );
not ( n80029 , n80028 );
or ( n80030 , n80027 , n80029 );
xor ( n80031 , n78942 , n78944 );
xor ( n80032 , n80031 , n79197 );
buf ( n80033 , n80032 );
nand ( n80034 , n80030 , n80033 );
nand ( n80035 , n80026 , n80034 );
nor ( n80036 , n79342 , n80035 );
and ( n80037 , n79306 , n79299 );
not ( n80038 , n79306 );
and ( n80039 , n80038 , n79275 );
or ( n80040 , n80037 , n80039 );
buf ( n80041 , n79296 );
not ( n80042 , n80041 );
and ( n80043 , n80040 , n80042 );
not ( n80044 , n80040 );
and ( n80045 , n80044 , n80041 );
nor ( n80046 , n80043 , n80045 );
or ( n80047 , n80036 , n80046 );
not ( n80048 , n79341 );
nand ( n80049 , n80048 , n80035 );
nand ( n80050 , n80047 , n80049 );
nand ( n80051 , n79339 , n80050 );
buf ( n80052 , n80051 );
not ( n80053 , n80052 );
buf ( n80054 , n79239 );
buf ( n80055 , n79318 );
nand ( n80056 , n80054 , n80055 );
buf ( n80057 , n80056 );
buf ( n80058 , n80057 );
nand ( n80059 , n80053 , n80058 );
buf ( n80060 , n80059 );
buf ( n80061 , n80060 );
nand ( n80062 , n79325 , n80061 );
buf ( n80063 , n80062 );
not ( n80064 , n80063 );
or ( n80065 , n79237 , n80064 );
buf ( n80066 , n78925 );
not ( n80067 , n80066 );
buf ( n80068 , n80067 );
buf ( n80069 , n80068 );
buf ( n80070 , n79233 );
not ( n80071 , n80070 );
buf ( n80072 , n80071 );
buf ( n80073 , n80072 );
nand ( n80074 , n80069 , n80073 );
buf ( n80075 , n80074 );
nand ( n80076 , n80065 , n80075 );
buf ( n80077 , n78884 );
buf ( n80078 , n80077 );
not ( n80079 , n80078 );
buf ( n80080 , n78888 );
not ( n80081 , n80080 );
or ( n80082 , n80079 , n80081 );
buf ( n80083 , n78888 );
buf ( n80084 , n80077 );
or ( n80085 , n80083 , n80084 );
buf ( n80086 , n78919 );
nand ( n80087 , n80085 , n80086 );
buf ( n80088 , n80087 );
buf ( n80089 , n80088 );
nand ( n80090 , n80082 , n80089 );
buf ( n80091 , n80090 );
xor ( n80092 , n76279 , n76371 );
xor ( n80093 , n80092 , n76375 );
buf ( n80094 , n80093 );
buf ( n80095 , n80094 );
not ( n80096 , n80095 );
buf ( n80097 , n80096 );
and ( n80098 , n80091 , n80097 );
not ( n80099 , n80091 );
and ( n80100 , n80099 , n80094 );
or ( n80101 , n80098 , n80100 );
buf ( n80102 , n80101 );
xor ( n80103 , n75311 , n75421 );
xor ( n80104 , n80103 , n75423 );
buf ( n80105 , n80104 );
buf ( n80106 , n80105 );
xor ( n80107 , n75109 , n75111 );
xor ( n80108 , n80107 , n75116 );
buf ( n80109 , n80108 );
buf ( n80110 , n80109 );
xor ( n80111 , n80106 , n80110 );
buf ( n80112 , n76941 );
not ( n80113 , n80112 );
buf ( n80114 , n77817 );
not ( n80115 , n80114 );
or ( n80116 , n80113 , n80115 );
buf ( n80117 , n76947 );
not ( n80118 , n80117 );
buf ( n80119 , n77820 );
not ( n80120 , n80119 );
or ( n80121 , n80118 , n80120 );
buf ( n80122 , n76937 );
nand ( n80123 , n80121 , n80122 );
buf ( n80124 , n80123 );
buf ( n80125 , n80124 );
nand ( n80126 , n80116 , n80125 );
buf ( n80127 , n80126 );
buf ( n80128 , n80127 );
xor ( n80129 , n80111 , n80128 );
buf ( n80130 , n80129 );
buf ( n80131 , n80130 );
not ( n80132 , n80131 );
buf ( n80133 , n80132 );
buf ( n80134 , n80133 );
and ( n80135 , n80102 , n80134 );
not ( n80136 , n80102 );
buf ( n80137 , n80130 );
and ( n80138 , n80136 , n80137 );
nor ( n80139 , n80135 , n80138 );
buf ( n80140 , n80139 );
xor ( n80141 , n77828 , n78881 );
and ( n80142 , n80141 , n78923 );
and ( n80143 , n77828 , n78881 );
or ( n80144 , n80142 , n80143 );
buf ( n80145 , n80144 );
nand ( n80146 , n80140 , n80145 );
nand ( n80147 , n80076 , n80146 );
buf ( n80148 , n80057 );
not ( n80149 , n80148 );
nor ( n80150 , n79339 , n80050 );
buf ( n80151 , n80150 );
nor ( n80152 , n80149 , n80151 );
buf ( n80153 , n80152 );
and ( n80154 , n80153 , n79236 );
xor ( n80155 , n79280 , n79291 );
xor ( n80156 , n80155 , n79293 );
buf ( n80157 , n80156 );
not ( n80158 , n80157 );
xor ( n80159 , n78962 , n79166 );
xor ( n80160 , n80159 , n79192 );
buf ( n80161 , n80160 );
buf ( n80162 , n80161 );
xor ( n80163 , n79088 , n79133 );
xor ( n80164 , n80163 , n79161 );
buf ( n80165 , n80164 );
buf ( n80166 , n80165 );
xor ( n80167 , n78987 , n78991 );
xor ( n80168 , n80167 , n79083 );
buf ( n80169 , n80168 );
buf ( n80170 , n80169 );
buf ( n80171 , n55841 );
not ( n80172 , n80171 );
buf ( n80173 , n62510 );
not ( n80174 , n80173 );
or ( n80175 , n80172 , n80174 );
buf ( n80176 , n25226 );
buf ( n80177 , n55840 );
nand ( n80178 , n80176 , n80177 );
buf ( n80179 , n80178 );
buf ( n80180 , n80179 );
nand ( n80181 , n80175 , n80180 );
buf ( n80182 , n80181 );
buf ( n80183 , n80182 );
not ( n80184 , n80183 );
buf ( n80185 , n73163 );
not ( n80186 , n80185 );
or ( n80187 , n80184 , n80186 );
buf ( n80188 , n79525 );
buf ( n80189 , n42665 );
nand ( n80190 , n80188 , n80189 );
buf ( n80191 , n80190 );
buf ( n80192 , n80191 );
nand ( n80193 , n80187 , n80192 );
buf ( n80194 , n80193 );
buf ( n80195 , n80194 );
buf ( n80196 , n60545 );
not ( n80197 , n80196 );
buf ( n80198 , n80002 );
not ( n80199 , n80198 );
or ( n80200 , n80197 , n80199 );
and ( n80201 , n28430 , n57174 );
not ( n80202 , n28430 );
and ( n80203 , n80202 , n48836 );
or ( n80204 , n80201 , n80203 );
buf ( n80205 , n80204 );
buf ( n80206 , n51488 );
nand ( n80207 , n80205 , n80206 );
buf ( n80208 , n80207 );
buf ( n80209 , n80208 );
nand ( n80210 , n80200 , n80209 );
buf ( n80211 , n80210 );
buf ( n80212 , n80211 );
xor ( n80213 , n80195 , n80212 );
buf ( n80214 , n53539 );
buf ( n80215 , n71123 );
and ( n80216 , n80214 , n80215 );
not ( n80217 , n80214 );
buf ( n80218 , n42257 );
and ( n80219 , n80217 , n80218 );
nor ( n80220 , n80216 , n80219 );
buf ( n80221 , n80220 );
buf ( n80222 , n80221 );
not ( n80223 , n80222 );
buf ( n80224 , n42246 );
not ( n80225 , n80224 );
or ( n80226 , n80223 , n80225 );
buf ( n80227 , n79398 );
buf ( n80228 , n42309 );
nand ( n80229 , n80227 , n80228 );
buf ( n80230 , n80229 );
buf ( n80231 , n80230 );
nand ( n80232 , n80226 , n80231 );
buf ( n80233 , n80232 );
buf ( n80234 , n80233 );
buf ( n80235 , n48865 );
not ( n80236 , n80235 );
buf ( n80237 , n79934 );
not ( n80238 , n80237 );
or ( n80239 , n80236 , n80238 );
buf ( n80240 , n48808 );
not ( n80241 , n80240 );
buf ( n80242 , n44946 );
not ( n80243 , n80242 );
or ( n80244 , n80241 , n80243 );
buf ( n80245 , n72891 );
buf ( n80246 , n74500 );
nand ( n80247 , n80245 , n80246 );
buf ( n80248 , n80247 );
buf ( n80249 , n80248 );
nand ( n80250 , n80244 , n80249 );
buf ( n80251 , n80250 );
buf ( n80252 , n80251 );
buf ( n80253 , n48852 );
nand ( n80254 , n80252 , n80253 );
buf ( n80255 , n80254 );
buf ( n80256 , n80255 );
nand ( n80257 , n80239 , n80256 );
buf ( n80258 , n80257 );
buf ( n80259 , n80258 );
buf ( n80260 , n46912 );
not ( n80261 , n80260 );
buf ( n80262 , n79460 );
not ( n80263 , n80262 );
or ( n80264 , n80261 , n80263 );
and ( n80265 , n47713 , n45723 );
not ( n80266 , n47713 );
buf ( n80267 , n45723 );
not ( n80268 , n80267 );
buf ( n80269 , n80268 );
and ( n80270 , n80266 , n80269 );
or ( n80271 , n80265 , n80270 );
nand ( n80272 , n80271 , n46907 );
buf ( n80273 , n80272 );
nand ( n80274 , n80264 , n80273 );
buf ( n80275 , n80274 );
buf ( n80276 , n80275 );
xor ( n80277 , n78153 , n78258 );
xor ( n80278 , n80277 , n78263 );
xor ( n80279 , n79800 , n79863 );
xor ( n80280 , n80278 , n80279 );
not ( n80281 , n46905 );
not ( n80282 , n80281 );
not ( n80283 , n80271 );
or ( n80284 , n80282 , n80283 );
and ( n80285 , n48320 , n45723 );
not ( n80286 , n48320 );
and ( n80287 , n80286 , n80269 );
or ( n80288 , n80285 , n80287 );
nand ( n80289 , n80288 , n46907 );
nand ( n80290 , n80284 , n80289 );
xor ( n80291 , n80280 , n80290 );
xor ( n80292 , n79626 , n79686 );
xor ( n80293 , n80292 , n79690 );
xor ( n80294 , n79838 , n79844 );
xor ( n80295 , n80293 , n80294 );
buf ( n80296 , n80295 );
xor ( n80297 , n78186 , n78199 );
xor ( n80298 , n80297 , n78216 );
xor ( n80299 , n79714 , n79763 );
xor ( n80300 , n80298 , n80299 );
buf ( n80301 , n80300 );
buf ( n80302 , n60270 );
buf ( n80303 , n15265 );
buf ( n80304 , n71818 );
and ( n80305 , n80303 , n80304 );
buf ( n80306 , n60090 );
buf ( n80307 , n71821 );
and ( n80308 , n80306 , n80307 );
nor ( n80309 , n80305 , n80308 );
buf ( n80310 , n80309 );
buf ( n80311 , n80310 );
or ( n80312 , n80302 , n80311 );
buf ( n80313 , n79640 );
buf ( n80314 , n60100 );
or ( n80315 , n80313 , n80314 );
nand ( n80316 , n80312 , n80315 );
buf ( n80317 , n80316 );
buf ( n80318 , n56781 );
buf ( n80319 , n623 );
and ( n80320 , n80318 , n80319 );
not ( n80321 , n56781 );
buf ( n80322 , n80321 );
buf ( n80323 , n75821 );
and ( n80324 , n80322 , n80323 );
buf ( n80325 , n58897 );
nor ( n80326 , n80324 , n80325 );
buf ( n80327 , n80326 );
buf ( n80328 , n80327 );
buf ( n80329 , n56777 );
nor ( n80330 , n80320 , n80328 , n80329 );
buf ( n80331 , n80330 );
xor ( n80332 , n80317 , n80331 );
buf ( n80333 , n58913 );
buf ( n80334 , n58897 );
buf ( n80335 , n74115 );
and ( n80336 , n80334 , n80335 );
buf ( n80337 , n58894 );
buf ( n80338 , n74118 );
and ( n80339 , n80337 , n80338 );
nor ( n80340 , n80336 , n80339 );
buf ( n80341 , n80340 );
buf ( n80342 , n80341 );
or ( n80343 , n80333 , n80342 );
buf ( n80344 , n79742 );
buf ( n80345 , n58884 );
or ( n80346 , n80344 , n80345 );
nand ( n80347 , n80343 , n80346 );
buf ( n80348 , n80347 );
and ( n80349 , n80332 , n80348 );
and ( n80350 , n80317 , n80331 );
or ( n80351 , n80349 , n80350 );
buf ( n80352 , n80351 );
xor ( n80353 , n79631 , n79648 );
buf ( n80354 , n80353 );
buf ( n80355 , n80354 );
xor ( n80356 , n80352 , n80355 );
buf ( n80357 , n70527 );
buf ( n80358 , n64129 );
and ( n80359 , n80357 , n80358 );
buf ( n80360 , n70530 );
buf ( n80361 , n63015 );
and ( n80362 , n80360 , n80361 );
nor ( n80363 , n80359 , n80362 );
buf ( n80364 , n80363 );
buf ( n80365 , n80364 );
buf ( n80366 , n64141 );
or ( n80367 , n80365 , n80366 );
buf ( n80368 , n79811 );
buf ( n80369 , n63010 );
or ( n80370 , n80368 , n80369 );
nand ( n80371 , n80367 , n80370 );
buf ( n80372 , n80371 );
buf ( n80373 , n80372 );
and ( n80374 , n80356 , n80373 );
and ( n80375 , n80352 , n80355 );
or ( n80376 , n80374 , n80375 );
buf ( n80377 , n80376 );
buf ( n80378 , n80377 );
xor ( n80379 , n80301 , n80378 );
xor ( n80380 , n79734 , n79751 );
xor ( n80381 , n80380 , n79759 );
buf ( n80382 , n80381 );
buf ( n80383 , n80382 );
buf ( n80384 , n58982 );
buf ( n80385 , n75821 );
nor ( n80386 , n80384 , n80385 );
buf ( n80387 , n80386 );
buf ( n80388 , n80387 );
buf ( n80389 , n60270 );
buf ( n80390 , n15265 );
buf ( n80391 , n72445 );
and ( n80392 , n80390 , n80391 );
buf ( n80393 , n60090 );
buf ( n80394 , n72448 );
and ( n80395 , n80393 , n80394 );
nor ( n80396 , n80392 , n80395 );
buf ( n80397 , n80396 );
buf ( n80398 , n80397 );
or ( n80399 , n80389 , n80398 );
buf ( n80400 , n80310 );
buf ( n80401 , n60100 );
or ( n80402 , n80400 , n80401 );
nand ( n80403 , n80399 , n80402 );
buf ( n80404 , n80403 );
buf ( n80405 , n80404 );
and ( n80406 , n80388 , n80405 );
buf ( n80407 , n80406 );
buf ( n80408 , n62935 );
buf ( n80409 , n71307 );
buf ( n80410 , n60096 );
and ( n80411 , n80409 , n80410 );
buf ( n80412 , n71310 );
buf ( n80413 , n62684 );
and ( n80414 , n80412 , n80413 );
nor ( n80415 , n80411 , n80414 );
buf ( n80416 , n80415 );
buf ( n80417 , n80416 );
or ( n80418 , n80408 , n80417 );
buf ( n80419 , n79725 );
buf ( n80420 , n62676 );
or ( n80421 , n80419 , n80420 );
nand ( n80422 , n80418 , n80421 );
buf ( n80423 , n80422 );
xor ( n80424 , n80407 , n80423 );
buf ( n80425 , n56807 );
buf ( n80426 , n623 );
or ( n80427 , n80425 , n80426 );
and ( n80428 , n56800 , n56777 , n623 );
not ( n80429 , n56815 );
nor ( n80430 , n80428 , n80429 );
buf ( n80431 , n80430 );
nand ( n80432 , n80427 , n80431 );
buf ( n80433 , n80432 );
and ( n80434 , n80424 , n80433 );
and ( n80435 , n80407 , n80423 );
or ( n80436 , n80434 , n80435 );
buf ( n80437 , n80436 );
xor ( n80438 , n80383 , n80437 );
buf ( n80439 , n70333 );
buf ( n80440 , n66742 );
and ( n80441 , n80439 , n80440 );
buf ( n80442 , n70336 );
buf ( n80443 , n63000 );
and ( n80444 , n80442 , n80443 );
nor ( n80445 , n80441 , n80444 );
buf ( n80446 , n80445 );
buf ( n80447 , n80446 );
buf ( n80448 , n64230 );
or ( n80449 , n80447 , n80448 );
buf ( n80450 , n79825 );
buf ( n80451 , n64227 );
or ( n80452 , n80450 , n80451 );
nand ( n80453 , n80449 , n80452 );
buf ( n80454 , n80453 );
buf ( n80455 , n80454 );
and ( n80456 , n80438 , n80455 );
and ( n80457 , n80383 , n80437 );
or ( n80458 , n80456 , n80457 );
buf ( n80459 , n80458 );
buf ( n80460 , n80459 );
and ( n80461 , n80379 , n80460 );
and ( n80462 , n80301 , n80378 );
or ( n80463 , n80461 , n80462 );
buf ( n80464 , n80463 );
buf ( n80465 , n80464 );
xor ( n80466 , n80296 , n80465 );
xor ( n80467 , n80352 , n80355 );
xor ( n80468 , n80467 , n80373 );
buf ( n80469 , n80468 );
buf ( n80470 , n71232 );
buf ( n80471 , n64129 );
and ( n80472 , n80470 , n80471 );
buf ( n80473 , n71235 );
buf ( n80474 , n63015 );
and ( n80475 , n80473 , n80474 );
nor ( n80476 , n80472 , n80475 );
buf ( n80477 , n80476 );
buf ( n80478 , n80477 );
buf ( n80479 , n64141 );
or ( n80480 , n80478 , n80479 );
buf ( n80481 , n80364 );
buf ( n80482 , n63010 );
or ( n80483 , n80481 , n80482 );
nand ( n80484 , n80480 , n80483 );
buf ( n80485 , n80484 );
xor ( n80486 , n80317 , n80331 );
xor ( n80487 , n80486 , n80348 );
and ( n80488 , n80485 , n80487 );
buf ( n80489 , n80341 );
buf ( n80490 , n58884 );
or ( n80491 , n80489 , n80490 );
buf ( n80492 , n58920 );
nand ( n80493 , n80491 , n80492 );
buf ( n80494 , n80493 );
buf ( n80495 , n80494 );
buf ( n80496 , n62681 );
buf ( n80497 , n71801 );
and ( n80498 , n80496 , n80497 );
buf ( n80499 , n62663 );
buf ( n80500 , n71804 );
and ( n80501 , n80499 , n80500 );
nor ( n80502 , n80498 , n80501 );
buf ( n80503 , n80502 );
buf ( n80504 , n80503 );
buf ( n80505 , n62935 );
or ( n80506 , n80504 , n80505 );
buf ( n80507 , n80416 );
buf ( n80508 , n62676 );
or ( n80509 , n80507 , n80508 );
nand ( n80510 , n80506 , n80509 );
buf ( n80511 , n80510 );
buf ( n80512 , n80511 );
xor ( n80513 , n80495 , n80512 );
buf ( n80514 , n71225 );
buf ( n80515 , n64129 );
and ( n80516 , n80514 , n80515 );
buf ( n80517 , n71228 );
buf ( n80518 , n63015 );
and ( n80519 , n80517 , n80518 );
nor ( n80520 , n80516 , n80519 );
buf ( n80521 , n80520 );
buf ( n80522 , n80521 );
buf ( n80523 , n64141 );
or ( n80524 , n80522 , n80523 );
buf ( n80525 , n80477 );
buf ( n80526 , n63010 );
or ( n80527 , n80525 , n80526 );
nand ( n80528 , n80524 , n80527 );
buf ( n80529 , n80528 );
buf ( n80530 , n80529 );
and ( n80531 , n80513 , n80530 );
and ( n80532 , n80495 , n80512 );
or ( n80533 , n80531 , n80532 );
buf ( n80534 , n80533 );
xor ( n80535 , n80317 , n80331 );
xor ( n80536 , n80535 , n80348 );
and ( n80537 , n80534 , n80536 );
and ( n80538 , n80485 , n80534 );
or ( n80539 , n80488 , n80537 , n80538 );
xor ( n80540 , n80469 , n80539 );
xor ( n80541 , n80383 , n80437 );
xor ( n80542 , n80541 , n80455 );
buf ( n80543 , n80542 );
and ( n80544 , n80540 , n80543 );
and ( n80545 , n80469 , n80539 );
or ( n80546 , n80544 , n80545 );
buf ( n80547 , n80546 );
xor ( n80548 , n79650 , n79669 );
xor ( n80549 , n80548 , n79683 );
xor ( n80550 , n79814 , n79833 );
xor ( n80551 , n80549 , n80550 );
buf ( n80552 , n80551 );
xor ( n80553 , n80547 , n80552 );
xor ( n80554 , n80301 , n80378 );
xor ( n80555 , n80554 , n80460 );
buf ( n80556 , n80555 );
buf ( n80557 , n80556 );
and ( n80558 , n80553 , n80557 );
and ( n80559 , n80547 , n80552 );
or ( n80560 , n80558 , n80559 );
buf ( n80561 , n80560 );
buf ( n80562 , n80561 );
and ( n80563 , n80466 , n80562 );
and ( n80564 , n80296 , n80465 );
or ( n80565 , n80563 , n80564 );
buf ( n80566 , n80565 );
buf ( n80567 , n80566 );
xor ( n80568 , n79850 , n79854 );
xor ( n80569 , n80568 , n79859 );
buf ( n80570 , n80569 );
buf ( n80571 , n80570 );
xor ( n80572 , n80567 , n80571 );
buf ( n80573 , n80281 );
not ( n80574 , n80573 );
buf ( n80575 , n80288 );
not ( n80576 , n80575 );
or ( n80577 , n80574 , n80576 );
buf ( n80578 , n46906 );
not ( n80579 , n80578 );
buf ( n80580 , n80579 );
buf ( n80581 , n80580 );
buf ( n80582 , n79875 );
not ( n80583 , n80582 );
buf ( n80584 , n80269 );
not ( n80585 , n80584 );
or ( n80586 , n80583 , n80585 );
buf ( n80587 , n45723 );
buf ( n80588 , n79882 );
nand ( n80589 , n80587 , n80588 );
buf ( n80590 , n80589 );
buf ( n80591 , n80590 );
nand ( n80592 , n80586 , n80591 );
buf ( n80593 , n80592 );
buf ( n80594 , n80593 );
nand ( n80595 , n80581 , n80594 );
buf ( n80596 , n80595 );
buf ( n80597 , n80596 );
nand ( n80598 , n80577 , n80597 );
buf ( n80599 , n80598 );
buf ( n80600 , n80599 );
and ( n80601 , n80572 , n80600 );
and ( n80602 , n80567 , n80571 );
or ( n80603 , n80601 , n80602 );
buf ( n80604 , n80603 );
and ( n80605 , n80291 , n80604 );
and ( n80606 , n80280 , n80290 );
or ( n80607 , n80605 , n80606 );
buf ( n80608 , n80607 );
xor ( n80609 , n80276 , n80608 );
buf ( n80610 , n48865 );
not ( n80611 , n80610 );
buf ( n80612 , n80251 );
not ( n80613 , n80612 );
or ( n80614 , n80611 , n80613 );
and ( n80615 , n25977 , n72891 );
not ( n80616 , n25977 );
and ( n80617 , n80616 , n48808 );
or ( n80618 , n80615 , n80617 );
buf ( n80619 , n80618 );
buf ( n80620 , n48852 );
nand ( n80621 , n80619 , n80620 );
buf ( n80622 , n80621 );
buf ( n80623 , n80622 );
nand ( n80624 , n80614 , n80623 );
buf ( n80625 , n80624 );
buf ( n80626 , n80625 );
and ( n80627 , n80609 , n80626 );
and ( n80628 , n80276 , n80608 );
or ( n80629 , n80627 , n80628 );
buf ( n80630 , n80629 );
buf ( n80631 , n80630 );
xor ( n80632 , n80259 , n80631 );
buf ( n80633 , n52780 );
not ( n80634 , n80633 );
buf ( n80635 , n72240 );
not ( n80636 , n80635 );
or ( n80637 , n80634 , n80636 );
buf ( n80638 , n42228 );
buf ( n80639 , n52789 );
nand ( n80640 , n80638 , n80639 );
buf ( n80641 , n80640 );
buf ( n80642 , n80641 );
nand ( n80643 , n80637 , n80642 );
buf ( n80644 , n80643 );
buf ( n80645 , n80644 );
not ( n80646 , n80645 );
buf ( n80647 , n41596 );
not ( n80648 , n80647 );
or ( n80649 , n80646 , n80648 );
buf ( n80650 , n79485 );
buf ( n80651 , n41574 );
nand ( n80652 , n80650 , n80651 );
buf ( n80653 , n80652 );
buf ( n80654 , n80653 );
nand ( n80655 , n80649 , n80654 );
buf ( n80656 , n80655 );
buf ( n80657 , n80656 );
and ( n80658 , n80632 , n80657 );
and ( n80659 , n80259 , n80631 );
or ( n80660 , n80658 , n80659 );
buf ( n80661 , n80660 );
buf ( n80662 , n80661 );
xor ( n80663 , n80234 , n80662 );
xor ( n80664 , n79473 , n79498 );
xor ( n80665 , n80664 , n79503 );
buf ( n80666 , n80665 );
buf ( n80667 , n80666 );
and ( n80668 , n80663 , n80667 );
and ( n80669 , n80234 , n80662 );
or ( n80670 , n80668 , n80669 );
buf ( n80671 , n80670 );
buf ( n80672 , n80671 );
and ( n80673 , n80213 , n80672 );
and ( n80674 , n80195 , n80212 );
or ( n80675 , n80673 , n80674 );
buf ( n80676 , n80675 );
buf ( n80677 , n80676 );
xor ( n80678 , n80170 , n80677 );
xor ( n80679 , n79513 , n79539 );
xor ( n80680 , n80679 , n79544 );
buf ( n80681 , n80680 );
buf ( n80682 , n80681 );
and ( n80683 , n80678 , n80682 );
and ( n80684 , n80170 , n80677 );
or ( n80685 , n80683 , n80684 );
buf ( n80686 , n80685 );
buf ( n80687 , n80686 );
xor ( n80688 , n80166 , n80687 );
xor ( n80689 , n79356 , n79381 );
xor ( n80690 , n80689 , n79549 );
buf ( n80691 , n80690 );
buf ( n80692 , n80691 );
and ( n80693 , n80688 , n80692 );
and ( n80694 , n80166 , n80687 );
or ( n80695 , n80693 , n80694 );
buf ( n80696 , n80695 );
buf ( n80697 , n80696 );
xor ( n80698 , n80162 , n80697 );
xor ( n80699 , n79352 , n79554 );
xor ( n80700 , n80699 , n79556 );
buf ( n80701 , n80700 );
buf ( n80702 , n80701 );
and ( n80703 , n80698 , n80702 );
and ( n80704 , n80162 , n80697 );
or ( n80705 , n80703 , n80704 );
buf ( n80706 , n80705 );
not ( n80707 , n80706 );
or ( n80708 , n80158 , n80707 );
not ( n80709 , n80157 );
not ( n80710 , n80709 );
not ( n80711 , n80706 );
not ( n80712 , n80711 );
or ( n80713 , n80710 , n80712 );
xor ( n80714 , n79560 , n80024 );
xnor ( n80715 , n80714 , n80033 );
nand ( n80716 , n80713 , n80715 );
nand ( n80717 , n80708 , n80716 );
not ( n80718 , n80717 );
not ( n80719 , n79561 );
not ( n80720 , n80024 );
or ( n80721 , n80719 , n80720 );
nand ( n80722 , n80721 , n80034 );
not ( n80723 , n80722 );
not ( n80724 , n79341 );
or ( n80725 , n80723 , n80724 );
or ( n80726 , n80035 , n79341 );
nand ( n80727 , n80725 , n80726 );
not ( n80728 , n80727 );
not ( n80729 , n80046 );
and ( n80730 , n80728 , n80729 );
and ( n80731 , n80046 , n80727 );
nor ( n80732 , n80730 , n80731 );
nand ( n80733 , n80718 , n80732 );
not ( n80734 , n80733 );
buf ( n80735 , C0 );
buf ( n80736 , n80735 );
xor ( n80737 , n79576 , n79578 );
xor ( n80738 , n80737 , n80015 );
buf ( n80739 , n80738 );
buf ( n80740 , n80739 );
xor ( n80741 , n80736 , n80740 );
xor ( n80742 , n79386 , n79411 );
xor ( n80743 , n80742 , n79508 );
buf ( n80744 , n80743 );
buf ( n80745 , n80744 );
buf ( n80746 , n60545 );
not ( n80747 , n80746 );
buf ( n80748 , n80204 );
not ( n80749 , n80748 );
or ( n80750 , n80747 , n80749 );
buf ( n80751 , n48836 );
not ( n80752 , n80751 );
buf ( n80753 , n43055 );
not ( n80754 , n80753 );
or ( n80755 , n80752 , n80754 );
buf ( n80756 , n43056 );
buf ( n80757 , n57174 );
nand ( n80758 , n80756 , n80757 );
buf ( n80759 , n80758 );
buf ( n80760 , n80759 );
nand ( n80761 , n80755 , n80760 );
buf ( n80762 , n80761 );
buf ( n80763 , n80762 );
buf ( n80764 , n51488 );
nand ( n80765 , n80763 , n80764 );
buf ( n80766 , n80765 );
buf ( n80767 , n80766 );
nand ( n80768 , n80750 , n80767 );
buf ( n80769 , n80768 );
buf ( n80770 , n80769 );
buf ( n80771 , n79899 );
buf ( n80772 , n79609 );
xor ( n80773 , n80771 , n80772 );
buf ( n80774 , n79904 );
xnor ( n80775 , n80773 , n80774 );
buf ( n80776 , n80775 );
buf ( n80777 , n80776 );
not ( n80778 , n80777 );
buf ( n80779 , n80778 );
not ( n80780 , n80779 );
not ( n80781 , n12481 );
nor ( n80782 , n80781 , n42664 );
not ( n80783 , n80782 );
or ( n80784 , n80780 , n80783 );
not ( n80785 , n80776 );
not ( n80786 , n42664 );
nand ( n80787 , n80786 , n12481 );
not ( n80788 , n80787 );
or ( n80789 , n80785 , n80788 );
xor ( n80790 , n79869 , n79873 );
xor ( n80791 , n80790 , n79895 );
buf ( n80792 , n80791 );
and ( n80793 , n56289 , n74492 );
not ( n80794 , n56289 );
and ( n80795 , n80794 , n41570 );
or ( n80796 , n80793 , n80795 );
buf ( n80797 , n80796 );
not ( n80798 , n80797 );
buf ( n80799 , n74487 );
not ( n80800 , n80799 );
or ( n80801 , n80798 , n80800 );
buf ( n80802 , n44495 );
not ( n80803 , n80802 );
buf ( n80804 , n79597 );
nand ( n80805 , n80803 , n80804 );
buf ( n80806 , n80805 );
buf ( n80807 , n80806 );
nand ( n80808 , n80801 , n80807 );
buf ( n80809 , n80808 );
xor ( n80810 , n80792 , n80809 );
not ( n80811 , n45741 );
buf ( n80812 , n50992 );
not ( n80813 , n80812 );
buf ( n80814 , n80813 );
buf ( n80815 , n80814 );
not ( n80816 , n80815 );
buf ( n80817 , n76179 );
not ( n80818 , n80817 );
or ( n80819 , n80816 , n80818 );
buf ( n80820 , n45746 );
buf ( n80821 , n50992 );
nand ( n80822 , n80820 , n80821 );
buf ( n80823 , n80822 );
buf ( n80824 , n80823 );
nand ( n80825 , n80819 , n80824 );
buf ( n80826 , n80825 );
not ( n80827 , n80826 );
or ( n80828 , n80811 , n80827 );
nand ( n80829 , n79886 , n67149 );
nand ( n80830 , n80828 , n80829 );
buf ( n80831 , n80830 );
not ( n80832 , n80831 );
buf ( n80833 , n48865 );
not ( n80834 , n80833 );
buf ( n80835 , n80618 );
not ( n80836 , n80835 );
or ( n80837 , n80834 , n80836 );
buf ( n80838 , n48852 );
buf ( n80839 , n48808 );
not ( n80840 , n80839 );
buf ( n80841 , n46384 );
not ( n80842 , n80841 );
or ( n80843 , n80840 , n80842 );
buf ( n80844 , n78314 );
buf ( n80845 , n72891 );
nand ( n80846 , n80844 , n80845 );
buf ( n80847 , n80846 );
buf ( n80848 , n80847 );
nand ( n80849 , n80843 , n80848 );
buf ( n80850 , n80849 );
buf ( n80851 , n80850 );
nand ( n80852 , n80838 , n80851 );
buf ( n80853 , n80852 );
buf ( n80854 , n80853 );
nand ( n80855 , n80837 , n80854 );
buf ( n80856 , n80855 );
buf ( n80857 , n80856 );
not ( n80858 , n80857 );
or ( n80859 , n80832 , n80858 );
buf ( n80860 , n80830 );
not ( n80861 , n80860 );
buf ( n80862 , n80861 );
buf ( n80863 , n80862 );
not ( n80864 , n80863 );
buf ( n80865 , n80856 );
not ( n80866 , n80865 );
buf ( n80867 , n80866 );
buf ( n80868 , n80867 );
not ( n80869 , n80868 );
or ( n80870 , n80864 , n80869 );
xor ( n80871 , n80280 , n80290 );
xor ( n80872 , n80871 , n80604 );
buf ( n80873 , n80872 );
nand ( n80874 , n80870 , n80873 );
buf ( n80875 , n80874 );
buf ( n80876 , n80875 );
nand ( n80877 , n80859 , n80876 );
buf ( n80878 , n80877 );
and ( n80879 , n80810 , n80878 );
and ( n80880 , n80792 , n80809 );
or ( n80881 , n80879 , n80880 );
nand ( n80882 , n80789 , n80881 );
nand ( n80883 , n80784 , n80882 );
buf ( n80884 , n80883 );
xor ( n80885 , n80770 , n80884 );
buf ( n80886 , n70268 );
not ( n80887 , n80886 );
buf ( n80888 , n12481 );
not ( n80889 , n80888 );
buf ( n80890 , n62510 );
not ( n80891 , n80890 );
or ( n80892 , n80889 , n80891 );
buf ( n80893 , n25226 );
buf ( n80894 , n56325 );
nand ( n80895 , n80893 , n80894 );
buf ( n80896 , n80895 );
buf ( n80897 , n80896 );
nand ( n80898 , n80892 , n80897 );
buf ( n80899 , n80898 );
buf ( n80900 , n80899 );
not ( n80901 , n80900 );
or ( n80902 , n80887 , n80901 );
buf ( n80903 , n80182 );
buf ( n80904 , n42665 );
nand ( n80905 , n80903 , n80904 );
buf ( n80906 , n80905 );
buf ( n80907 , n80906 );
nand ( n80908 , n80902 , n80907 );
buf ( n80909 , n80908 );
buf ( n80910 , n80909 );
and ( n80911 , n80885 , n80910 );
and ( n80912 , n80770 , n80884 );
or ( n80913 , n80911 , n80912 );
buf ( n80914 , n80913 );
buf ( n80915 , n80914 );
xor ( n80916 , n80745 , n80915 );
xor ( n80917 , n79585 , n79962 );
xor ( n80918 , n80917 , n79966 );
buf ( n80919 , n80918 );
buf ( n80920 , n80919 );
and ( n80921 , n80916 , n80920 );
and ( n80922 , n80745 , n80915 );
or ( n80923 , n80921 , n80922 );
buf ( n80924 , n80923 );
buf ( n80925 , n80924 );
xor ( n80926 , n79971 , n79992 );
xor ( n80927 , n80926 , n80010 );
buf ( n80928 , n80927 );
buf ( n80929 , n80928 );
buf ( n80930 , C0 );
buf ( n80931 , n80930 );
and ( n80932 , n80925 , n80929 );
or ( n80933 , C0 , n80932 );
buf ( n80934 , n80933 );
buf ( n80935 , n80934 );
and ( n80936 , n80741 , n80935 );
or ( n80937 , n80936 , C0 );
buf ( n80938 , n80937 );
buf ( n80939 , n80938 );
xor ( n80940 , n79566 , n80019 );
xor ( n80941 , n80940 , n80021 );
buf ( n80942 , n80941 );
buf ( n80943 , n80942 );
xor ( n80944 , n80939 , n80943 );
xor ( n80945 , n80162 , n80697 );
xor ( n80946 , n80945 , n80702 );
buf ( n80947 , n80946 );
buf ( n80948 , n80947 );
and ( n80949 , n80944 , n80948 );
and ( n80950 , n80939 , n80943 );
or ( n80951 , n80949 , n80950 );
buf ( n80952 , n80951 );
buf ( n80953 , n80952 );
xor ( n80954 , n80157 , n80711 );
xnor ( n80955 , n80954 , n80715 );
buf ( n80956 , n80955 );
xor ( n80957 , n80953 , n80956 );
xor ( n80958 , n79916 , n79941 );
xor ( n80959 , n80958 , n79957 );
buf ( n80960 , n80959 );
buf ( n80961 , n80960 );
buf ( n80962 , n52456 );
not ( n80963 , n80962 );
buf ( n80964 , n80762 );
not ( n80965 , n80964 );
or ( n80966 , n80963 , n80965 );
buf ( n80967 , n48836 );
not ( n80968 , n80967 );
buf ( n80969 , n72235 );
not ( n80970 , n80969 );
or ( n80971 , n80968 , n80970 );
buf ( n80972 , n42856 );
buf ( n80973 , n57174 );
nand ( n80974 , n80972 , n80973 );
buf ( n80975 , n80974 );
buf ( n80976 , n80975 );
nand ( n80977 , n80971 , n80976 );
buf ( n80978 , n80977 );
buf ( n80979 , n80978 );
buf ( n80980 , n51488 );
nand ( n80981 , n80979 , n80980 );
buf ( n80982 , n80981 );
buf ( n80983 , n80982 );
nand ( n80984 , n80966 , n80983 );
buf ( n80985 , n80984 );
buf ( n80986 , n80985 );
buf ( n80987 , n53539 );
not ( n80988 , n80987 );
buf ( n80989 , n41586 );
not ( n80990 , n80989 );
or ( n80991 , n80988 , n80990 );
buf ( n80992 , n42228 );
buf ( n80993 , n53548 );
nand ( n80994 , n80992 , n80993 );
buf ( n80995 , n80994 );
buf ( n80996 , n80995 );
nand ( n80997 , n80991 , n80996 );
buf ( n80998 , n80997 );
buf ( n80999 , n80998 );
not ( n81000 , n80999 );
buf ( n81001 , n67354 );
not ( n81002 , n81001 );
or ( n81003 , n81000 , n81002 );
buf ( n81004 , n41571 );
not ( n81005 , n81004 );
buf ( n81006 , n80644 );
nand ( n81007 , n81005 , n81006 );
buf ( n81008 , n81007 );
buf ( n81009 , n81008 );
nand ( n81010 , n81003 , n81009 );
buf ( n81011 , n81010 );
not ( n81012 , n81011 );
buf ( n81013 , n75152 );
buf ( n81014 , n42228 );
buf ( n81015 , n24883 );
or ( n81016 , n81014 , n81015 );
buf ( n81017 , n12481 );
nand ( n81018 , n81016 , n81017 );
buf ( n81019 , n81018 );
buf ( n81020 , n81019 );
not ( n81021 , n24884 );
nand ( n81022 , n81021 , n42228 );
buf ( n81023 , n81022 );
nand ( n81024 , n81013 , n81020 , n81023 );
buf ( n81025 , n81024 );
nand ( n81026 , n81012 , n81025 );
not ( n81027 , n81026 );
xor ( n81028 , n80276 , n80608 );
xor ( n81029 , n81028 , n80626 );
buf ( n81030 , n81029 );
not ( n81031 , n81030 );
or ( n81032 , n81027 , n81031 );
buf ( n81033 , n81025 );
not ( n81034 , n81033 );
buf ( n81035 , n81034 );
buf ( n81036 , n81035 );
buf ( n81037 , n81011 );
nand ( n81038 , n81036 , n81037 );
buf ( n81039 , n81038 );
nand ( n81040 , n81032 , n81039 );
buf ( n81041 , n81040 );
xor ( n81042 , n80986 , n81041 );
buf ( n81043 , n55841 );
not ( n81044 , n81043 );
buf ( n81045 , n25303 );
not ( n81046 , n81045 );
or ( n81047 , n81044 , n81046 );
buf ( n81048 , n75152 );
buf ( n81049 , n55840 );
nand ( n81050 , n81048 , n81049 );
buf ( n81051 , n81050 );
buf ( n81052 , n81051 );
nand ( n81053 , n81047 , n81052 );
buf ( n81054 , n81053 );
buf ( n81055 , n81054 );
not ( n81056 , n81055 );
buf ( n81057 , n42246 );
not ( n81058 , n81057 );
or ( n81059 , n81056 , n81058 );
buf ( n81060 , n80221 );
buf ( n81061 , n42309 );
nand ( n81062 , n81060 , n81061 );
buf ( n81063 , n81062 );
buf ( n81064 , n81063 );
nand ( n81065 , n81059 , n81064 );
buf ( n81066 , n81065 );
buf ( n81067 , n81066 );
and ( n81068 , n81042 , n81067 );
and ( n81069 , n80986 , n81041 );
or ( n81070 , n81068 , n81069 );
buf ( n81071 , n81070 );
buf ( n81072 , n81071 );
xor ( n81073 , n80961 , n81072 );
xor ( n81074 , n80234 , n80662 );
xor ( n81075 , n81074 , n80667 );
buf ( n81076 , n81075 );
buf ( n81077 , n81076 );
and ( n81078 , n81073 , n81077 );
and ( n81079 , n80961 , n81072 );
or ( n81080 , n81078 , n81079 );
buf ( n81081 , n81080 );
buf ( n81082 , n81081 );
xor ( n81083 , n80195 , n80212 );
xor ( n81084 , n81083 , n80672 );
buf ( n81085 , n81084 );
buf ( n81086 , n81085 );
buf ( n81087 , C0 );
buf ( n81088 , n81087 );
and ( n81089 , n81082 , n81086 );
or ( n81090 , C0 , n81089 );
buf ( n81091 , n81090 );
buf ( n81092 , n81091 );
xor ( n81093 , n80170 , n80677 );
xor ( n81094 , n81093 , n80682 );
buf ( n81095 , n81094 );
buf ( n81096 , n81095 );
buf ( n81097 , C0 );
buf ( n81098 , n81097 );
and ( n81099 , n81092 , n81096 );
or ( n81100 , C0 , n81099 );
buf ( n81101 , n81100 );
buf ( n81102 , n81101 );
xor ( n81103 , n80166 , n80687 );
xor ( n81104 , n81103 , n80692 );
buf ( n81105 , n81104 );
buf ( n81106 , n81105 );
xor ( n81107 , n81102 , n81106 );
xor ( n81108 , n80736 , n80740 );
xor ( n81109 , n81108 , n80935 );
buf ( n81110 , n81109 );
buf ( n81111 , n81110 );
and ( n81112 , n81107 , n81111 );
and ( n81113 , n81102 , n81106 );
or ( n81114 , n81112 , n81113 );
buf ( n81115 , n81114 );
buf ( n81116 , n81115 );
xor ( n81117 , n80939 , n80943 );
xor ( n81118 , n81117 , n80948 );
buf ( n81119 , n81118 );
buf ( n81120 , n81119 );
xor ( n81121 , n81116 , n81120 );
buf ( n81122 , C0 );
buf ( n81123 , n81122 );
xor ( n81124 , n80770 , n80884 );
xor ( n81125 , n81124 , n80910 );
buf ( n81126 , n81125 );
buf ( n81127 , n81126 );
or ( n81128 , n81123 , n81127 );
xor ( n81129 , n80259 , n80631 );
xor ( n81130 , n81129 , n80657 );
buf ( n81131 , n81130 );
buf ( n81132 , n81131 );
not ( n81133 , n81132 );
not ( n81134 , n52456 );
not ( n81135 , n80978 );
or ( n81136 , n81134 , n81135 );
buf ( n81137 , n48836 );
not ( n81138 , n81137 );
buf ( n81139 , n74460 );
not ( n81140 , n81139 );
or ( n81141 , n81138 , n81140 );
buf ( n81142 , n42844 );
buf ( n81143 , n57174 );
nand ( n81144 , n81142 , n81143 );
buf ( n81145 , n81144 );
buf ( n81146 , n81145 );
nand ( n81147 , n81141 , n81146 );
buf ( n81148 , n81147 );
buf ( n81149 , n81148 );
buf ( n81150 , n51488 );
nand ( n81151 , n81149 , n81150 );
buf ( n81152 , n81151 );
nand ( n81153 , n81136 , n81152 );
not ( n81154 , n81153 );
xor ( n81155 , n80792 , n80809 );
xor ( n81156 , n81155 , n80878 );
not ( n81157 , n81156 );
or ( n81158 , n81154 , n81157 );
not ( n81159 , n81153 );
not ( n81160 , n81159 );
not ( n81161 , n81156 );
not ( n81162 , n81161 );
or ( n81163 , n81160 , n81162 );
xor ( n81164 , n80296 , n80465 );
xor ( n81165 , n81164 , n80562 );
buf ( n81166 , n81165 );
buf ( n81167 , n81166 );
buf ( n81168 , n80814 );
not ( n81169 , n81168 );
buf ( n81170 , n80269 );
not ( n81171 , n81170 );
or ( n81172 , n81169 , n81171 );
buf ( n81173 , n45723 );
buf ( n81174 , n50992 );
nand ( n81175 , n81173 , n81174 );
buf ( n81176 , n81175 );
buf ( n81177 , n81176 );
nand ( n81178 , n81172 , n81177 );
buf ( n81179 , n81178 );
buf ( n81180 , n81179 );
not ( n81181 , n81180 );
buf ( n81182 , n80580 );
not ( n81183 , n81182 );
or ( n81184 , n81181 , n81183 );
buf ( n81185 , n80593 );
buf ( n81186 , n46912 );
nand ( n81187 , n81185 , n81186 );
buf ( n81188 , n81187 );
buf ( n81189 , n81188 );
nand ( n81190 , n81184 , n81189 );
buf ( n81191 , n81190 );
buf ( n81192 , n81191 );
xor ( n81193 , n81167 , n81192 );
buf ( n81194 , n48865 );
not ( n81195 , n81194 );
not ( n81196 , n24713 );
buf ( n81197 , n81196 );
not ( n81198 , n81197 );
buf ( n81199 , n47713 );
not ( n81200 , n81199 );
or ( n81201 , n81198 , n81200 );
buf ( n81202 , n81196 );
not ( n81203 , n81202 );
buf ( n81204 , n81203 );
buf ( n81205 , n81204 );
buf ( n81206 , n25938 );
nand ( n81207 , n81205 , n81206 );
buf ( n81208 , n81207 );
buf ( n81209 , n81208 );
nand ( n81210 , n81201 , n81209 );
buf ( n81211 , n81210 );
buf ( n81212 , n81211 );
not ( n81213 , n81212 );
or ( n81214 , n81195 , n81213 );
buf ( n81215 , n48808 );
buf ( n81216 , n71078 );
and ( n81217 , n81215 , n81216 );
not ( n81218 , n81215 );
buf ( n81219 , n48320 );
and ( n81220 , n81218 , n81219 );
nor ( n81221 , n81217 , n81220 );
buf ( n81222 , n81221 );
buf ( n81223 , n81222 );
buf ( n81224 , n48852 );
nand ( n81225 , n81223 , n81224 );
buf ( n81226 , n81225 );
buf ( n81227 , n81226 );
nand ( n81228 , n81214 , n81227 );
buf ( n81229 , n81228 );
buf ( n81230 , n81229 );
and ( n81231 , n81193 , n81230 );
and ( n81232 , n81167 , n81192 );
or ( n81233 , n81231 , n81232 );
buf ( n81234 , n81233 );
buf ( n81235 , n81234 );
buf ( n81236 , n60545 );
not ( n81237 , n81236 );
buf ( n81238 , n48836 );
not ( n81239 , n81238 );
buf ( n81240 , n74503 );
not ( n81241 , n81240 );
or ( n81242 , n81239 , n81241 );
buf ( n81243 , n74500 );
buf ( n81244 , n61847 );
nand ( n81245 , n81243 , n81244 );
buf ( n81246 , n81245 );
buf ( n81247 , n81246 );
nand ( n81248 , n81242 , n81247 );
buf ( n81249 , n81248 );
buf ( n81250 , n81249 );
not ( n81251 , n81250 );
or ( n81252 , n81237 , n81251 );
buf ( n81253 , n48836 );
not ( n81254 , n81253 );
buf ( n81255 , n72310 );
not ( n81256 , n81255 );
or ( n81257 , n81254 , n81256 );
buf ( n81258 , n46114 );
buf ( n81259 , n61847 );
nand ( n81260 , n81258 , n81259 );
buf ( n81261 , n81260 );
buf ( n81262 , n81261 );
nand ( n81263 , n81257 , n81262 );
buf ( n81264 , n81263 );
buf ( n81265 , n81264 );
buf ( n81266 , n51488 );
nand ( n81267 , n81265 , n81266 );
buf ( n81268 , n81267 );
buf ( n81269 , n81268 );
nand ( n81270 , n81252 , n81269 );
buf ( n81271 , n81270 );
buf ( n81272 , n81271 );
xor ( n81273 , n81235 , n81272 );
buf ( n81274 , n41582 );
not ( n81275 , n81274 );
buf ( n81276 , n81275 );
buf ( n81277 , n81276 );
buf ( n81278 , n25385 );
or ( n81279 , n81277 , n81278 );
buf ( n81280 , n12481 );
nand ( n81281 , n81279 , n81280 );
buf ( n81282 , n81281 );
buf ( n81283 , n81282 );
buf ( n81284 , n42228 );
buf ( n81285 , n81276 );
buf ( n81286 , n25385 );
nand ( n81287 , n81285 , n81286 );
buf ( n81288 , n81287 );
buf ( n81289 , n81288 );
and ( n81290 , n81283 , n81284 , n81289 );
buf ( n81291 , n81290 );
buf ( n81292 , n81291 );
and ( n81293 , n81273 , n81292 );
and ( n81294 , n81235 , n81272 );
or ( n81295 , n81293 , n81294 );
buf ( n81296 , n81295 );
not ( n81297 , n81296 );
xor ( n81298 , n80567 , n80571 );
xor ( n81299 , n81298 , n80600 );
buf ( n81300 , n81299 );
buf ( n81301 , n81300 );
buf ( n81302 , n48865 );
not ( n81303 , n81302 );
buf ( n81304 , n80850 );
not ( n81305 , n81304 );
or ( n81306 , n81303 , n81305 );
buf ( n81307 , n81211 );
buf ( n81308 , n48852 );
nand ( n81309 , n81307 , n81308 );
buf ( n81310 , n81309 );
buf ( n81311 , n81310 );
nand ( n81312 , n81306 , n81311 );
buf ( n81313 , n81312 );
buf ( n81314 , n81313 );
xor ( n81315 , n81301 , n81314 );
buf ( n81316 , n56289 );
not ( n81317 , n81316 );
buf ( n81318 , n44491 );
not ( n81319 , n81318 );
or ( n81320 , n81317 , n81319 );
buf ( n81321 , n44494 );
buf ( n81322 , n52094 );
nand ( n81323 , n81321 , n81322 );
buf ( n81324 , n81323 );
buf ( n81325 , n81324 );
nand ( n81326 , n81320 , n81325 );
buf ( n81327 , n81326 );
buf ( n81328 , n81327 );
not ( n81329 , n81328 );
buf ( n81330 , n45741 );
not ( n81331 , n81330 );
or ( n81332 , n81329 , n81331 );
buf ( n81333 , n80826 );
buf ( n81334 , n67149 );
nand ( n81335 , n81333 , n81334 );
buf ( n81336 , n81335 );
buf ( n81337 , n81336 );
nand ( n81338 , n81332 , n81337 );
buf ( n81339 , n81338 );
buf ( n81340 , n81339 );
and ( n81341 , n81315 , n81340 );
and ( n81342 , n81301 , n81314 );
or ( n81343 , n81341 , n81342 );
buf ( n81344 , n81343 );
not ( n81345 , n81344 );
buf ( n81346 , n52789 );
buf ( n81347 , n25385 );
and ( n81348 , n81346 , n81347 );
not ( n81349 , n81346 );
buf ( n81350 , n79031 );
and ( n81351 , n81349 , n81350 );
nor ( n81352 , n81348 , n81351 );
buf ( n81353 , n81352 );
buf ( n81354 , n81353 );
not ( n81355 , n81354 );
buf ( n81356 , n81355 );
buf ( n81357 , n81356 );
not ( n81358 , n81357 );
buf ( n81359 , n74488 );
not ( n81360 , n81359 );
or ( n81361 , n81358 , n81360 );
buf ( n81362 , n80796 );
buf ( n81363 , n44496 );
nand ( n81364 , n81362 , n81363 );
buf ( n81365 , n81364 );
buf ( n81366 , n81365 );
nand ( n81367 , n81361 , n81366 );
buf ( n81368 , n81367 );
not ( n81369 , n81368 );
nand ( n81370 , n81345 , n81369 );
not ( n81371 , n81370 );
or ( n81372 , n81297 , n81371 );
not ( n81373 , n81369 );
nand ( n81374 , n81373 , n81344 );
nand ( n81375 , n81372 , n81374 );
nand ( n81376 , n81163 , n81375 );
nand ( n81377 , n81158 , n81376 );
buf ( n81378 , n81377 );
not ( n81379 , n81378 );
or ( n81380 , n81133 , n81379 );
buf ( n81381 , n81377 );
buf ( n81382 , n81131 );
or ( n81383 , n81381 , n81382 );
and ( n81384 , n80881 , n80776 );
not ( n81385 , n80881 );
and ( n81386 , n81385 , n80779 );
or ( n81387 , n81384 , n81386 );
buf ( n81388 , n81387 );
buf ( n81389 , n80782 );
and ( n81390 , n81388 , n81389 );
not ( n81391 , n81388 );
buf ( n81392 , n80787 );
and ( n81393 , n81391 , n81392 );
nor ( n81394 , n81390 , n81393 );
buf ( n81395 , n81394 );
buf ( n81396 , n81395 );
nand ( n81397 , n81383 , n81396 );
buf ( n81398 , n81397 );
buf ( n81399 , n81398 );
nand ( n81400 , n81380 , n81399 );
buf ( n81401 , n81400 );
buf ( n81402 , n81401 );
nand ( n81403 , n81128 , n81402 );
buf ( n81404 , n81403 );
buf ( n81405 , n81404 );
buf ( n81406 , C1 );
buf ( n81407 , n81406 );
nand ( n81408 , n81405 , n81407 );
buf ( n81409 , n81408 );
buf ( n81410 , n81409 );
xor ( n81411 , n80745 , n80915 );
xor ( n81412 , n81411 , n80920 );
buf ( n81413 , n81412 );
buf ( n81414 , n81413 );
buf ( n81415 , C0 );
buf ( n81416 , n81415 );
and ( n81417 , n81410 , n81414 );
or ( n81418 , C0 , n81417 );
buf ( n81419 , n81418 );
buf ( n81420 , n81419 );
xor ( n81421 , n80925 , n80929 );
xor ( n81422 , n81421 , n80931 );
buf ( n81423 , n81422 );
buf ( n81424 , n81423 );
xor ( n81425 , n81420 , n81424 );
xor ( n81426 , n81092 , n81096 );
xor ( n81427 , n81426 , n81098 );
buf ( n81428 , n81427 );
buf ( n81429 , n81428 );
and ( n81430 , n81425 , n81429 );
and ( n81431 , n81420 , n81424 );
or ( n81432 , n81430 , n81431 );
buf ( n81433 , n81432 );
buf ( n81434 , n81433 );
xor ( n81435 , n81102 , n81106 );
xor ( n81436 , n81435 , n81111 );
buf ( n81437 , n81436 );
buf ( n81438 , n81437 );
xor ( n81439 , n81434 , n81438 );
xor ( n81440 , n81082 , n81086 );
xor ( n81441 , n81440 , n81088 );
buf ( n81442 , n81441 );
buf ( n81443 , n81442 );
xor ( n81444 , n80961 , n81072 );
xor ( n81445 , n81444 , n81077 );
buf ( n81446 , n81445 );
buf ( n81447 , n81446 );
buf ( n81448 , C0 );
or ( n81449 , n81447 , n81448 );
buf ( n81450 , C0 );
xor ( n81451 , n80986 , n81041 );
xor ( n81452 , n81451 , n81067 );
buf ( n81453 , n81452 );
buf ( n81454 , n81450 );
buf ( n81455 , n81453 );
or ( n81456 , n81454 , n81455 );
buf ( n81457 , n80862 );
buf ( n81458 , n80856 );
xor ( n81459 , n81457 , n81458 );
buf ( n81460 , n80872 );
xnor ( n81461 , n81459 , n81460 );
buf ( n81462 , n81461 );
buf ( n81463 , n81462 );
buf ( n81464 , n55841 );
not ( n81465 , n81464 );
buf ( n81466 , n74530 );
not ( n81467 , n81466 );
or ( n81468 , n81465 , n81467 );
buf ( n81469 , n42228 );
buf ( n81470 , n55840 );
nand ( n81471 , n81469 , n81470 );
buf ( n81472 , n81471 );
buf ( n81473 , n81472 );
nand ( n81474 , n81468 , n81473 );
buf ( n81475 , n81474 );
buf ( n81476 , n81475 );
not ( n81477 , n81476 );
buf ( n81478 , n67354 );
not ( n81479 , n81478 );
or ( n81480 , n81477 , n81479 );
buf ( n81481 , n80998 );
buf ( n81482 , n41574 );
nand ( n81483 , n81481 , n81482 );
buf ( n81484 , n81483 );
buf ( n81485 , n81484 );
nand ( n81486 , n81480 , n81485 );
buf ( n81487 , n81486 );
buf ( n81488 , n81487 );
xor ( n81489 , n81463 , n81488 );
buf ( n81490 , n42306 );
buf ( n81491 , n56325 );
nor ( n81492 , n81490 , n81491 );
buf ( n81493 , n81492 );
buf ( n81494 , n81493 );
and ( n81495 , n81489 , n81494 );
and ( n81496 , n81463 , n81488 );
or ( n81497 , n81495 , n81496 );
buf ( n81498 , n81497 );
buf ( n81499 , n81498 );
buf ( n81500 , n12481 );
buf ( n81501 , n25306 );
and ( n81502 , n81500 , n81501 );
not ( n81503 , n81500 );
buf ( n81504 , n42257 );
and ( n81505 , n81503 , n81504 );
nor ( n81506 , n81502 , n81505 );
buf ( n81507 , n81506 );
buf ( n81508 , n81507 );
not ( n81509 , n81508 );
buf ( n81510 , n42246 );
not ( n81511 , n81510 );
or ( n81512 , n81509 , n81511 );
buf ( n81513 , n81054 );
buf ( n81514 , n42309 );
nand ( n81515 , n81513 , n81514 );
buf ( n81516 , n81515 );
buf ( n81517 , n81516 );
nand ( n81518 , n81512 , n81517 );
buf ( n81519 , n81518 );
buf ( n81520 , n81519 );
xor ( n81521 , n81499 , n81520 );
buf ( n81522 , n81030 );
buf ( n81523 , n81011 );
xor ( n81524 , n81522 , n81523 );
buf ( n81525 , n81035 );
xor ( n81526 , n81524 , n81525 );
buf ( n81527 , n81526 );
buf ( n81528 , n81527 );
and ( n81529 , n81521 , n81528 );
and ( n81530 , n81499 , n81520 );
or ( n81531 , n81529 , n81530 );
buf ( n81532 , n81531 );
buf ( n81533 , n81532 );
nand ( n81534 , n81456 , n81533 );
buf ( n81535 , n81534 );
buf ( n81536 , n81535 );
nand ( n81537 , C1 , n81536 );
buf ( n81538 , n81537 );
buf ( n81539 , n81538 );
nand ( n81540 , n81449 , n81539 );
buf ( n81541 , n81540 );
buf ( n81542 , n81541 );
buf ( n81543 , C1 );
buf ( n81544 , n81543 );
nand ( n81545 , n81542 , n81544 );
buf ( n81546 , n81545 );
buf ( n81547 , n81546 );
xor ( n81548 , n81443 , n81547 );
xor ( n81549 , n81410 , n81414 );
xor ( n81550 , n81549 , n81416 );
buf ( n81551 , n81550 );
buf ( n81552 , n81551 );
and ( n81553 , n81548 , n81552 );
and ( n81554 , n81443 , n81547 );
or ( n81555 , n81553 , n81554 );
buf ( n81556 , n81555 );
buf ( n81557 , n81556 );
xor ( n81558 , n81420 , n81424 );
xor ( n81559 , n81558 , n81429 );
buf ( n81560 , n81559 );
buf ( n81561 , n81560 );
xor ( n81562 , n81557 , n81561 );
buf ( n81563 , n81401 );
buf ( n81564 , n81122 );
xor ( n81565 , n81563 , n81564 );
buf ( n81566 , n81126 );
xnor ( n81567 , n81565 , n81566 );
buf ( n81568 , n81567 );
buf ( n81569 , n81568 );
buf ( n81570 , n81131 );
buf ( n81571 , n81377 );
xor ( n81572 , n81570 , n81571 );
buf ( n81573 , n81395 );
xnor ( n81574 , n81572 , n81573 );
buf ( n81575 , n81574 );
buf ( n81576 , n81575 );
buf ( n81577 , C1 );
buf ( n81578 , n81577 );
xor ( n81579 , n81159 , n81156 );
xor ( n81580 , n81579 , n81375 );
buf ( n81581 , n81580 );
xor ( n81582 , n81578 , n81581 );
buf ( n81583 , C1 );
nand ( n81584 , n52456 , n81148 );
nand ( n81585 , n81249 , n51488 );
and ( n81586 , n81584 , n81585 );
nand ( n81587 , n81583 , n81586 );
buf ( n81588 , n44516 );
not ( n81589 , n81588 );
buf ( n81590 , n53548 );
buf ( n81591 , n41570 );
and ( n81592 , n81590 , n81591 );
not ( n81593 , n81590 );
buf ( n81594 , n79031 );
and ( n81595 , n81593 , n81594 );
nor ( n81596 , n81592 , n81595 );
buf ( n81597 , n81596 );
buf ( n81598 , n81597 );
not ( n81599 , n81598 );
and ( n81600 , n81589 , n81599 );
buf ( n81601 , n81353 );
buf ( n81602 , n44495 );
nor ( n81603 , n81601 , n81602 );
buf ( n81604 , n81603 );
buf ( n81605 , n81604 );
nor ( n81606 , n81600 , n81605 );
buf ( n81607 , n81606 );
buf ( n81608 , n81607 );
not ( n81609 , n81608 );
buf ( n81610 , n81609 );
not ( n81611 , n81610 );
buf ( n81612 , n70348 );
buf ( n81613 , n63003 );
and ( n81614 , n81612 , n81613 );
buf ( n81615 , n70351 );
buf ( n81616 , n64223 );
and ( n81617 , n81615 , n81616 );
nor ( n81618 , n81614 , n81617 );
buf ( n81619 , n81618 );
buf ( n81620 , n81619 );
buf ( n81621 , n64230 );
or ( n81622 , n81620 , n81621 );
buf ( n81623 , n80446 );
buf ( n81624 , n64227 );
or ( n81625 , n81623 , n81624 );
nand ( n81626 , n81622 , n81625 );
buf ( n81627 , n81626 );
xor ( n81628 , n80407 , n80423 );
xor ( n81629 , n81628 , n80433 );
and ( n81630 , n81627 , n81629 );
buf ( n81631 , n62935 );
buf ( n81632 , n60096 );
buf ( n81633 , n71818 );
and ( n81634 , n81632 , n81633 );
buf ( n81635 , n62663 );
buf ( n81636 , n71821 );
and ( n81637 , n81635 , n81636 );
nor ( n81638 , n81634 , n81637 );
buf ( n81639 , n81638 );
buf ( n81640 , n81639 );
or ( n81641 , n81631 , n81640 );
buf ( n81642 , n80503 );
buf ( n81643 , n62676 );
or ( n81644 , n81642 , n81643 );
nand ( n81645 , n81641 , n81644 );
buf ( n81646 , n81645 );
buf ( n81647 , n81646 );
buf ( n81648 , n58875 );
buf ( n81649 , n623 );
and ( n81650 , n81648 , n81649 );
buf ( n81651 , n15117 );
buf ( n81652 , n75821 );
and ( n81653 , n81651 , n81652 );
buf ( n81654 , n15265 );
nor ( n81655 , n81653 , n81654 );
buf ( n81656 , n81655 );
buf ( n81657 , n81656 );
buf ( n81658 , n58897 );
nor ( n81659 , n81650 , n81657 , n81658 );
buf ( n81660 , n81659 );
buf ( n81661 , n81660 );
xor ( n81662 , n81647 , n81661 );
buf ( n81663 , n60270 );
buf ( n81664 , n60261 );
buf ( n81665 , n74115 );
and ( n81666 , n81664 , n81665 );
buf ( n81667 , n60090 );
buf ( n81668 , n74118 );
and ( n81669 , n81667 , n81668 );
nor ( n81670 , n81666 , n81669 );
buf ( n81671 , n81670 );
buf ( n81672 , n81671 );
or ( n81673 , n81663 , n81672 );
buf ( n81674 , n80397 );
buf ( n81675 , n60100 );
or ( n81676 , n81674 , n81675 );
nand ( n81677 , n81673 , n81676 );
buf ( n81678 , n81677 );
buf ( n81679 , n81678 );
and ( n81680 , n81662 , n81679 );
and ( n81681 , n81647 , n81661 );
or ( n81682 , n81680 , n81681 );
buf ( n81683 , n81682 );
buf ( n81684 , n81683 );
xor ( n81685 , n80388 , n80405 );
buf ( n81686 , n81685 );
buf ( n81687 , n81686 );
xor ( n81688 , n81684 , n81687 );
buf ( n81689 , n71307 );
buf ( n81690 , n64129 );
and ( n81691 , n81689 , n81690 );
buf ( n81692 , n71310 );
buf ( n81693 , n63015 );
and ( n81694 , n81692 , n81693 );
nor ( n81695 , n81691 , n81694 );
buf ( n81696 , n81695 );
buf ( n81697 , n81696 );
buf ( n81698 , n64141 );
or ( n81699 , n81697 , n81698 );
buf ( n81700 , n80521 );
buf ( n81701 , n63010 );
or ( n81702 , n81700 , n81701 );
nand ( n81703 , n81699 , n81702 );
buf ( n81704 , n81703 );
buf ( n81705 , n81704 );
buf ( n81706 , n58890 );
buf ( n81707 , n75821 );
nor ( n81708 , n81706 , n81707 );
buf ( n81709 , n81708 );
buf ( n81710 , n81709 );
buf ( n81711 , n71801 );
buf ( n81712 , n62668 );
and ( n81713 , n81711 , n81712 );
buf ( n81714 , n71804 );
buf ( n81715 , n63015 );
and ( n81716 , n81714 , n81715 );
nor ( n81717 , n81713 , n81716 );
buf ( n81718 , n81717 );
buf ( n81719 , n81718 );
buf ( n81720 , n64141 );
or ( n81721 , n81719 , n81720 );
buf ( n81722 , n81696 );
buf ( n81723 , n63010 );
or ( n81724 , n81722 , n81723 );
nand ( n81725 , n81721 , n81724 );
buf ( n81726 , n81725 );
buf ( n81727 , n81726 );
and ( n81728 , n81710 , n81727 );
buf ( n81729 , n81728 );
buf ( n81730 , n81729 );
xor ( n81731 , n81705 , n81730 );
buf ( n81732 , n58920 );
buf ( n81733 , n623 );
or ( n81734 , n81732 , n81733 );
buf ( n81735 , n58916 );
buf ( n81736 , n58897 );
buf ( n81737 , n623 );
and ( n81738 , n81735 , n81736 , n81737 );
buf ( n81739 , n58900 );
nor ( n81740 , n81738 , n81739 );
buf ( n81741 , n81740 );
buf ( n81742 , n81741 );
nand ( n81743 , n81734 , n81742 );
buf ( n81744 , n81743 );
buf ( n81745 , n81744 );
and ( n81746 , n81731 , n81745 );
and ( n81747 , n81705 , n81730 );
or ( n81748 , n81746 , n81747 );
buf ( n81749 , n81748 );
buf ( n81750 , n81749 );
and ( n81751 , n81688 , n81750 );
and ( n81752 , n81684 , n81687 );
or ( n81753 , n81751 , n81752 );
buf ( n81754 , n81753 );
xor ( n81755 , n80407 , n80423 );
xor ( n81756 , n81755 , n80433 );
and ( n81757 , n81754 , n81756 );
and ( n81758 , n81627 , n81754 );
or ( n81759 , n81630 , n81757 , n81758 );
xor ( n81760 , n80469 , n80539 );
xor ( n81761 , n81760 , n80543 );
and ( n81762 , n81759 , n81761 );
xor ( n81763 , n80495 , n80512 );
xor ( n81764 , n81763 , n80530 );
buf ( n81765 , n81764 );
buf ( n81766 , n70527 );
buf ( n81767 , n63003 );
and ( n81768 , n81766 , n81767 );
buf ( n81769 , n70530 );
buf ( n81770 , n63000 );
and ( n81771 , n81769 , n81770 );
nor ( n81772 , n81768 , n81771 );
buf ( n81773 , n81772 );
buf ( n81774 , n81773 );
buf ( n81775 , n64230 );
or ( n81776 , n81774 , n81775 );
buf ( n81777 , n81619 );
buf ( n81778 , n64227 );
or ( n81779 , n81777 , n81778 );
nand ( n81780 , n81776 , n81779 );
buf ( n81781 , n81780 );
xor ( n81782 , n81765 , n81781 );
buf ( n81783 , n71232 );
buf ( n81784 , n63003 );
and ( n81785 , n81783 , n81784 );
buf ( n81786 , n71235 );
buf ( n81787 , n63000 );
and ( n81788 , n81786 , n81787 );
nor ( n81789 , n81785 , n81788 );
buf ( n81790 , n81789 );
buf ( n81791 , n81790 );
buf ( n81792 , n64230 );
or ( n81793 , n81791 , n81792 );
buf ( n81794 , n81773 );
buf ( n81795 , n64227 );
or ( n81796 , n81794 , n81795 );
nand ( n81797 , n81793 , n81796 );
buf ( n81798 , n81797 );
buf ( n81799 , n81798 );
xor ( n81800 , n81647 , n81661 );
xor ( n81801 , n81800 , n81679 );
buf ( n81802 , n81801 );
buf ( n81803 , n81802 );
xor ( n81804 , n81799 , n81803 );
buf ( n81805 , n81671 );
buf ( n81806 , n60100 );
or ( n81807 , n81805 , n81806 );
buf ( n81808 , n60102 );
nand ( n81809 , n81807 , n81808 );
buf ( n81810 , n81809 );
buf ( n81811 , n81810 );
buf ( n81812 , n62935 );
buf ( n81813 , n62681 );
buf ( n81814 , n72445 );
and ( n81815 , n81813 , n81814 );
buf ( n81816 , n62663 );
buf ( n81817 , n72448 );
and ( n81818 , n81816 , n81817 );
nor ( n81819 , n81815 , n81818 );
buf ( n81820 , n81819 );
buf ( n81821 , n81820 );
or ( n81822 , n81812 , n81821 );
buf ( n81823 , n81639 );
buf ( n81824 , n62676 );
or ( n81825 , n81823 , n81824 );
nand ( n81826 , n81822 , n81825 );
buf ( n81827 , n81826 );
buf ( n81828 , n81827 );
xor ( n81829 , n81811 , n81828 );
xor ( n81830 , n81710 , n81727 );
buf ( n81831 , n81830 );
buf ( n81832 , n81831 );
and ( n81833 , n81829 , n81832 );
and ( n81834 , n81811 , n81828 );
or ( n81835 , n81833 , n81834 );
buf ( n81836 , n81835 );
buf ( n81837 , n81836 );
and ( n81838 , n81804 , n81837 );
and ( n81839 , n81799 , n81803 );
or ( n81840 , n81838 , n81839 );
buf ( n81841 , n81840 );
and ( n81842 , n81782 , n81841 );
and ( n81843 , n81765 , n81781 );
or ( n81844 , n81842 , n81843 );
buf ( n81845 , n81844 );
xor ( n81846 , n80317 , n80331 );
xor ( n81847 , n81846 , n80348 );
xor ( n81848 , n80485 , n80534 );
xor ( n81849 , n81847 , n81848 );
buf ( n81850 , n81849 );
xor ( n81851 , n81845 , n81850 );
xor ( n81852 , n80407 , n80423 );
xor ( n81853 , n81852 , n80433 );
xor ( n81854 , n81627 , n81754 );
xor ( n81855 , n81853 , n81854 );
buf ( n81856 , n81855 );
and ( n81857 , n81851 , n81856 );
and ( n81858 , n81845 , n81850 );
or ( n81859 , n81857 , n81858 );
buf ( n81860 , n81859 );
xor ( n81861 , n80469 , n80539 );
xor ( n81862 , n81861 , n80543 );
and ( n81863 , n81860 , n81862 );
and ( n81864 , n81759 , n81860 );
or ( n81865 , n81762 , n81863 , n81864 );
buf ( n81866 , n81865 );
xor ( n81867 , n80547 , n80552 );
xor ( n81868 , n81867 , n80557 );
buf ( n81869 , n81868 );
buf ( n81870 , n81869 );
xor ( n81871 , n81866 , n81870 );
buf ( n81872 , n56289 );
not ( n81873 , n81872 );
buf ( n81874 , n80269 );
not ( n81875 , n81874 );
or ( n81876 , n81873 , n81875 );
buf ( n81877 , n45723 );
buf ( n81878 , n52094 );
nand ( n81879 , n81877 , n81878 );
buf ( n81880 , n81879 );
buf ( n81881 , n81880 );
nand ( n81882 , n81876 , n81881 );
buf ( n81883 , n81882 );
buf ( n81884 , n81883 );
not ( n81885 , n81884 );
buf ( n81886 , n80580 );
not ( n81887 , n81886 );
or ( n81888 , n81885 , n81887 );
buf ( n81889 , n81179 );
buf ( n81890 , n80281 );
nand ( n81891 , n81889 , n81890 );
buf ( n81892 , n81891 );
buf ( n81893 , n81892 );
nand ( n81894 , n81888 , n81893 );
buf ( n81895 , n81894 );
buf ( n81896 , n81895 );
and ( n81897 , n81871 , n81896 );
and ( n81898 , n81866 , n81870 );
or ( n81899 , n81897 , n81898 );
buf ( n81900 , n81899 );
not ( n81901 , n81900 );
buf ( n81902 , n45727 );
not ( n81903 , n81902 );
buf ( n81904 , n81327 );
not ( n81905 , n81904 );
or ( n81906 , n81903 , n81905 );
buf ( n81907 , n45741 );
buf ( n81908 , n52780 );
not ( n81909 , n81908 );
buf ( n81910 , n44491 );
not ( n81911 , n81910 );
or ( n81912 , n81909 , n81911 );
buf ( n81913 , n45746 );
buf ( n81914 , n52789 );
nand ( n81915 , n81913 , n81914 );
buf ( n81916 , n81915 );
buf ( n81917 , n81916 );
nand ( n81918 , n81912 , n81917 );
buf ( n81919 , n81918 );
buf ( n81920 , n81919 );
nand ( n81921 , n81907 , n81920 );
buf ( n81922 , n81921 );
buf ( n81923 , n81922 );
nand ( n81924 , n81906 , n81923 );
buf ( n81925 , n81924 );
buf ( n81926 , n81925 );
not ( n81927 , n81926 );
buf ( n81928 , n81927 );
nand ( n81929 , n81901 , n81928 );
not ( n81930 , n81929 );
xor ( n81931 , n81167 , n81192 );
xor ( n81932 , n81931 , n81230 );
buf ( n81933 , n81932 );
not ( n81934 , n81933 );
or ( n81935 , n81930 , n81934 );
buf ( n81936 , n81900 );
buf ( n81937 , n81925 );
nand ( n81938 , n81936 , n81937 );
buf ( n81939 , n81938 );
nand ( n81940 , n81935 , n81939 );
not ( n81941 , n81940 );
or ( n81942 , n81611 , n81941 );
buf ( n81943 , n81940 );
not ( n81944 , n81943 );
buf ( n81945 , n81944 );
not ( n81946 , n81945 );
not ( n81947 , n81607 );
or ( n81948 , n81946 , n81947 );
xor ( n81949 , n81301 , n81314 );
xor ( n81950 , n81949 , n81340 );
buf ( n81951 , n81950 );
nand ( n81952 , n81948 , n81951 );
nand ( n81953 , n81942 , n81952 );
and ( n81954 , n81587 , n81953 );
nor ( n81955 , C0 , n81954 );
buf ( n81956 , n81955 );
and ( n81957 , n81582 , n81956 );
and ( n81958 , n81578 , n81581 );
or ( n81959 , n81957 , n81958 );
buf ( n81960 , n81959 );
buf ( n81961 , n81960 );
xor ( n81962 , n81576 , n81961 );
buf ( n81963 , C1 );
buf ( n81964 , n81963 );
and ( n81965 , n81962 , n81964 );
and ( n81966 , n81576 , n81961 );
or ( n81967 , n81965 , n81966 );
buf ( n81968 , n81967 );
buf ( n81969 , n81968 );
or ( n81970 , n81569 , n81969 );
buf ( n81971 , n81538 );
buf ( n81972 , n81446 );
xor ( n81973 , n81971 , n81972 );
buf ( n81974 , C0 );
xnor ( n81975 , n81973 , n81974 );
buf ( n81976 , n81975 );
buf ( n81977 , n81976 );
buf ( n81978 , n81968 );
buf ( n81979 , n81568 );
and ( n81980 , n81978 , n81979 );
buf ( n81981 , n81980 );
buf ( n81982 , n81981 );
or ( n81983 , n81977 , n81982 );
nand ( n81984 , n81970 , n81983 );
buf ( n81985 , n81984 );
buf ( n81986 , n81985 );
xor ( n81987 , n81443 , n81547 );
xor ( n81988 , n81987 , n81552 );
buf ( n81989 , n81988 );
buf ( n81990 , n81989 );
xor ( n81991 , n81986 , n81990 );
xor ( n81992 , C1 , n81453 );
xor ( n81993 , n81992 , n81532 );
buf ( n81994 , n81993 );
not ( n81995 , n81994 );
xor ( n81996 , n81576 , n81961 );
xor ( n81997 , n81996 , n81964 );
buf ( n81998 , n81997 );
buf ( n81999 , n81998 );
not ( n82000 , n81999 );
or ( n82001 , n81995 , n82000 );
buf ( n82002 , C0 );
not ( n82003 , n81475 );
not ( n82004 , n41574 );
or ( n82005 , n82003 , n82004 );
nand ( n82006 , n74530 , n12481 );
not ( n82007 , n82006 );
buf ( n82008 , n42228 );
buf ( n82009 , n56325 );
nand ( n82010 , n82008 , n82009 );
buf ( n82011 , n82010 );
not ( n82012 , n82011 );
or ( n82013 , n82007 , n82012 );
nand ( n82014 , n82013 , n67354 );
nand ( n82015 , n82005 , n82014 );
buf ( n82016 , n82015 );
buf ( n82017 , n81222 );
not ( n82018 , n82017 );
buf ( n82019 , n48865 );
not ( n82020 , n82019 );
or ( n82021 , n82018 , n82020 );
buf ( n82022 , n81196 );
not ( n82023 , n82022 );
buf ( n82024 , n25900 );
not ( n82025 , n82024 );
buf ( n82026 , n82025 );
buf ( n82027 , n82026 );
not ( n82028 , n82027 );
or ( n82029 , n82023 , n82028 );
buf ( n82030 , n81204 );
buf ( n82031 , n25900 );
nand ( n82032 , n82030 , n82031 );
buf ( n82033 , n82032 );
buf ( n82034 , n82033 );
nand ( n82035 , n82029 , n82034 );
buf ( n82036 , n82035 );
buf ( n82037 , n82036 );
buf ( n82038 , n48852 );
nand ( n82039 , n82037 , n82038 );
buf ( n82040 , n82039 );
buf ( n82041 , n82040 );
nand ( n82042 , n82021 , n82041 );
buf ( n82043 , n82042 );
buf ( n82044 , n82043 );
xor ( n82045 , n80469 , n80539 );
xor ( n82046 , n82045 , n80543 );
xor ( n82047 , n81759 , n81860 );
xor ( n82048 , n82046 , n82047 );
buf ( n82049 , n82048 );
buf ( n82050 , n48865 );
not ( n82051 , n82050 );
buf ( n82052 , n82036 );
not ( n82053 , n82052 );
or ( n82054 , n82051 , n82053 );
buf ( n82055 , n48852 );
buf ( n82056 , n80814 );
not ( n82057 , n82056 );
buf ( n82058 , n46903 );
not ( n82059 , n82058 );
or ( n82060 , n82057 , n82059 );
buf ( n82061 , n50992 );
buf ( n82062 , n24714 );
nand ( n82063 , n82061 , n82062 );
buf ( n82064 , n82063 );
buf ( n82065 , n82064 );
nand ( n82066 , n82060 , n82065 );
buf ( n82067 , n82066 );
buf ( n82068 , n82067 );
nand ( n82069 , n82055 , n82068 );
buf ( n82070 , n82069 );
buf ( n82071 , n82070 );
nand ( n82072 , n82054 , n82071 );
buf ( n82073 , n82072 );
buf ( n82074 , n82073 );
xor ( n82075 , n82049 , n82074 );
xor ( n82076 , n81684 , n81687 );
xor ( n82077 , n82076 , n81750 );
buf ( n82078 , n82077 );
xor ( n82079 , n81765 , n81781 );
xor ( n82080 , n82079 , n81841 );
and ( n82081 , n82078 , n82080 );
buf ( n82082 , n71225 );
buf ( n82083 , n63003 );
and ( n82084 , n82082 , n82083 );
buf ( n82085 , n71228 );
buf ( n82086 , n64223 );
and ( n82087 , n82085 , n82086 );
nor ( n82088 , n82084 , n82087 );
buf ( n82089 , n82088 );
buf ( n82090 , n82089 );
buf ( n82091 , n64230 );
or ( n82092 , n82090 , n82091 );
buf ( n82093 , n81790 );
buf ( n82094 , n64227 );
or ( n82095 , n82093 , n82094 );
nand ( n82096 , n82092 , n82095 );
buf ( n82097 , n82096 );
buf ( n82098 , n60084 );
buf ( n82099 , n623 );
and ( n82100 , n82098 , n82099 );
buf ( n82101 , n60087 );
buf ( n82102 , n75821 );
and ( n82103 , n82101 , n82102 );
buf ( n82104 , n62681 );
nor ( n82105 , n82103 , n82104 );
buf ( n82106 , n82105 );
buf ( n82107 , n82106 );
buf ( n82108 , n15265 );
nor ( n82109 , n82100 , n82107 , n82108 );
buf ( n82110 , n82109 );
buf ( n82111 , n82110 );
buf ( n82112 , n64141 );
buf ( n82113 , n62668 );
buf ( n82114 , n71818 );
and ( n82115 , n82113 , n82114 );
buf ( n82116 , n71821 );
buf ( n82117 , n63015 );
and ( n82118 , n82116 , n82117 );
nor ( n82119 , n82115 , n82118 );
buf ( n82120 , n82119 );
buf ( n82121 , n82120 );
or ( n82122 , n82112 , n82121 );
buf ( n82123 , n81718 );
buf ( n82124 , n63010 );
or ( n82125 , n82123 , n82124 );
nand ( n82126 , n82122 , n82125 );
buf ( n82127 , n82126 );
buf ( n82128 , n82127 );
xor ( n82129 , n82111 , n82128 );
buf ( n82130 , n64141 );
buf ( n82131 , n62668 );
buf ( n82132 , n72445 );
and ( n82133 , n82131 , n82132 );
buf ( n82134 , n63015 );
buf ( n82135 , n72448 );
and ( n82136 , n82134 , n82135 );
nor ( n82137 , n82133 , n82136 );
buf ( n82138 , n82137 );
buf ( n82139 , n82138 );
or ( n82140 , n82130 , n82139 );
buf ( n82141 , n82120 );
buf ( n82142 , n63010 );
or ( n82143 , n82141 , n82142 );
nand ( n82144 , n82140 , n82143 );
buf ( n82145 , n82144 );
buf ( n82146 , n82145 );
buf ( n82147 , n60100 );
buf ( n82148 , n75821 );
nor ( n82149 , n82147 , n82148 );
buf ( n82150 , n82149 );
buf ( n82151 , n82150 );
and ( n82152 , n82146 , n82151 );
buf ( n82153 , n82152 );
buf ( n82154 , n82153 );
and ( n82155 , n82129 , n82154 );
and ( n82156 , n82111 , n82128 );
or ( n82157 , n82155 , n82156 );
buf ( n82158 , n82157 );
xor ( n82159 , n82097 , n82158 );
xor ( n82160 , n81811 , n81828 );
xor ( n82161 , n82160 , n81832 );
buf ( n82162 , n82161 );
and ( n82163 , n82159 , n82162 );
and ( n82164 , n82097 , n82158 );
or ( n82165 , n82163 , n82164 );
buf ( n82166 , n82165 );
xor ( n82167 , n81705 , n81730 );
xor ( n82168 , n82167 , n81745 );
buf ( n82169 , n82168 );
buf ( n82170 , n82169 );
xor ( n82171 , n82166 , n82170 );
xor ( n82172 , n81799 , n81803 );
xor ( n82173 , n82172 , n81837 );
buf ( n82174 , n82173 );
buf ( n82175 , n82174 );
and ( n82176 , n82171 , n82175 );
and ( n82177 , n82166 , n82170 );
or ( n82178 , n82176 , n82177 );
buf ( n82179 , n82178 );
xor ( n82180 , n81765 , n81781 );
xor ( n82181 , n82180 , n81841 );
and ( n82182 , n82179 , n82181 );
and ( n82183 , n82078 , n82179 );
or ( n82184 , n82081 , n82182 , n82183 );
buf ( n82185 , n82184 );
xor ( n82186 , n81845 , n81850 );
xor ( n82187 , n82186 , n81856 );
buf ( n82188 , n82187 );
buf ( n82189 , n82188 );
xor ( n82190 , n82185 , n82189 );
buf ( n82191 , n48848 );
not ( n82192 , n82191 );
nand ( n82193 , n52084 , n52087 , n52088 , n52091 );
buf ( n82194 , n82193 );
not ( n82195 , n82194 );
buf ( n82196 , n46903 );
not ( n82197 , n82196 );
or ( n82198 , n82195 , n82197 );
buf ( n82199 , n52093 );
buf ( n82200 , n24714 );
nand ( n82201 , n82199 , n82200 );
buf ( n82202 , n82201 );
buf ( n82203 , n82202 );
nand ( n82204 , n82198 , n82203 );
buf ( n82205 , n82204 );
buf ( n82206 , n82205 );
not ( n82207 , n82206 );
or ( n82208 , n82192 , n82207 );
buf ( n82209 , n82067 );
buf ( n82210 , n48865 );
nand ( n82211 , n82209 , n82210 );
buf ( n82212 , n82211 );
buf ( n82213 , n82212 );
nand ( n82214 , n82208 , n82213 );
buf ( n82215 , n82214 );
buf ( n82216 , n82215 );
and ( n82217 , n82190 , n82216 );
and ( n82218 , n82185 , n82189 );
or ( n82219 , n82217 , n82218 );
buf ( n82220 , n82219 );
buf ( n82221 , n82220 );
and ( n82222 , n82075 , n82221 );
and ( n82223 , n82049 , n82074 );
or ( n82224 , n82222 , n82223 );
buf ( n82225 , n82224 );
buf ( n82226 , n82225 );
xor ( n82227 , n82044 , n82226 );
xor ( n82228 , n81866 , n81870 );
xor ( n82229 , n82228 , n81896 );
buf ( n82230 , n82229 );
buf ( n82231 , n82230 );
and ( n82232 , n82227 , n82231 );
and ( n82233 , n82044 , n82226 );
or ( n82234 , n82232 , n82233 );
buf ( n82235 , n82234 );
buf ( n82236 , n82235 );
buf ( n82237 , n52456 );
not ( n82238 , n82237 );
buf ( n82239 , n81264 );
not ( n82240 , n82239 );
or ( n82241 , n82238 , n82240 );
buf ( n82242 , n48836 );
not ( n82243 , n82242 );
buf ( n82244 , n46384 );
not ( n82245 , n82244 );
or ( n82246 , n82243 , n82245 );
buf ( n82247 , n25951 );
buf ( n82248 , n61847 );
nand ( n82249 , n82247 , n82248 );
buf ( n82250 , n82249 );
buf ( n82251 , n82250 );
nand ( n82252 , n82246 , n82251 );
buf ( n82253 , n82252 );
buf ( n82254 , n82253 );
buf ( n82255 , n51488 );
nand ( n82256 , n82254 , n82255 );
buf ( n82257 , n82256 );
buf ( n82258 , n82257 );
nand ( n82259 , n82241 , n82258 );
buf ( n82260 , n82259 );
buf ( n82261 , n82260 );
xor ( n82262 , n82236 , n82261 );
buf ( n82263 , n41571 );
buf ( n82264 , n56325 );
nor ( n82265 , n82263 , n82264 );
buf ( n82266 , n82265 );
buf ( n82267 , n82266 );
and ( n82268 , n82262 , n82267 );
and ( n82269 , n82236 , n82261 );
or ( n82270 , n82268 , n82269 );
buf ( n82271 , n82270 );
buf ( n82272 , n82271 );
xor ( n82273 , n82016 , n82272 );
not ( n82274 , n55841 );
not ( n82275 , n74492 );
or ( n82276 , n82274 , n82275 );
buf ( n82277 , n44503 );
buf ( n82278 , n55840 );
nand ( n82279 , n82277 , n82278 );
buf ( n82280 , n82279 );
nand ( n82281 , n82276 , n82280 );
not ( n82282 , n82281 );
not ( n82283 , n74488 );
or ( n82284 , n82282 , n82283 );
buf ( n82285 , n81597 );
not ( n82286 , n82285 );
buf ( n82287 , n44496 );
nand ( n82288 , n82286 , n82287 );
buf ( n82289 , n82288 );
nand ( n82290 , n82284 , n82289 );
buf ( n82291 , n82290 );
buf ( n82292 , n52456 );
not ( n82293 , n82292 );
buf ( n82294 , n82253 );
not ( n82295 , n82294 );
or ( n82296 , n82293 , n82295 );
and ( n82297 , n47713 , n48836 );
not ( n82298 , n47713 );
and ( n82299 , n82298 , n61847 );
or ( n82300 , n82297 , n82299 );
buf ( n82301 , n82300 );
buf ( n82302 , n51488 );
nand ( n82303 , n82301 , n82302 );
buf ( n82304 , n82303 );
buf ( n82305 , n82304 );
nand ( n82306 , n82296 , n82305 );
buf ( n82307 , n82306 );
buf ( n82308 , n82307 );
buf ( n82309 , n53539 );
not ( n82310 , n82309 );
buf ( n82311 , n76179 );
not ( n82312 , n82311 );
or ( n82313 , n82310 , n82312 );
buf ( n82314 , n44494 );
buf ( n82315 , n53548 );
nand ( n82316 , n82314 , n82315 );
buf ( n82317 , n82316 );
buf ( n82318 , n82317 );
nand ( n82319 , n82313 , n82318 );
buf ( n82320 , n82319 );
buf ( n82321 , n82320 );
not ( n82322 , n82321 );
buf ( n82323 , n45741 );
not ( n82324 , n82323 );
or ( n82325 , n82322 , n82324 );
buf ( n82326 , n81919 );
buf ( n82327 , n67149 );
nand ( n82328 , n82326 , n82327 );
buf ( n82329 , n82328 );
buf ( n82330 , n82329 );
nand ( n82331 , n82325 , n82330 );
buf ( n82332 , n82331 );
buf ( n82333 , n82332 );
xor ( n82334 , n82308 , n82333 );
buf ( n82335 , n25382 );
nor ( n82336 , n45746 , n24833 );
or ( n82337 , n82336 , n56325 );
buf ( n82338 , n45746 );
buf ( n82339 , n24833 );
nand ( n82340 , n82338 , n82339 );
buf ( n82341 , n82340 );
nand ( n82342 , n82337 , n82341 );
buf ( n82343 , n82342 );
nor ( n82344 , n82335 , n82343 );
buf ( n82345 , n82344 );
buf ( n82346 , n82345 );
and ( n82347 , n82334 , n82346 );
and ( n82348 , n82308 , n82333 );
or ( n82349 , n82347 , n82348 );
buf ( n82350 , n82349 );
buf ( n82351 , n82350 );
or ( n82352 , n82291 , n82351 );
xor ( n82353 , n81900 , n81928 );
xor ( n82354 , n82353 , n81933 );
buf ( n82355 , n82354 );
not ( n82356 , n82355 );
buf ( n82357 , n82356 );
buf ( n82358 , n82357 );
nand ( n82359 , n82352 , n82358 );
buf ( n82360 , n82359 );
buf ( n82361 , n82360 );
buf ( n82362 , n82290 );
buf ( n82363 , n82350 );
nand ( n82364 , n82362 , n82363 );
buf ( n82365 , n82364 );
buf ( n82366 , n82365 );
nand ( n82367 , n82361 , n82366 );
buf ( n82368 , n82367 );
buf ( n82369 , n82368 );
and ( n82370 , n82273 , n82369 );
and ( n82371 , n82016 , n82272 );
or ( n82372 , n82370 , n82371 );
buf ( n82373 , n82372 );
not ( n82374 , n82373 );
not ( n82375 , n81344 );
not ( n82376 , n81369 );
and ( n82377 , n82375 , n82376 );
and ( n82378 , n81344 , n81369 );
nor ( n82379 , n82377 , n82378 );
not ( n82380 , n81296 );
and ( n82381 , n82379 , n82380 );
not ( n82382 , n82379 );
and ( n82383 , n82382 , n81296 );
nor ( n82384 , n82381 , n82383 );
not ( n82385 , n82384 );
nand ( n82386 , n82374 , n82385 );
not ( n82387 , n82386 );
xor ( n82388 , n81463 , n81488 );
xor ( n82389 , n82388 , n81494 );
buf ( n82390 , n82389 );
not ( n82391 , n82390 );
or ( n82392 , n82387 , n82391 );
not ( n82393 , n82385 );
nand ( n82394 , n82393 , n82373 );
nand ( n82395 , n82392 , n82394 );
buf ( n82396 , n82002 );
buf ( n82397 , n82395 );
or ( n82398 , n82396 , n82397 );
xor ( n82399 , n81499 , n81520 );
xor ( n82400 , n82399 , n81528 );
buf ( n82401 , n82400 );
buf ( n82402 , n82401 );
nand ( n82403 , n82398 , n82402 );
buf ( n82404 , n82403 );
nand ( n82405 , C1 , n82404 );
buf ( n82406 , n82405 );
nand ( n82407 , n82001 , n82406 );
buf ( n82408 , n82407 );
buf ( n82409 , n82408 );
not ( n82410 , n81998 );
buf ( n82411 , n81993 );
not ( n82412 , n82411 );
buf ( n82413 , n82412 );
nand ( n82414 , n82410 , n82413 );
buf ( n82415 , n82414 );
nand ( n82416 , n82409 , n82415 );
buf ( n82417 , n82416 );
buf ( n82418 , n82417 );
not ( n82419 , n82418 );
buf ( n82420 , n81976 );
not ( n82421 , n82420 );
xor ( n82422 , n81978 , n81979 );
buf ( n82423 , n82422 );
buf ( n82424 , n82423 );
not ( n82425 , n82424 );
and ( n82426 , n82421 , n82425 );
buf ( n82427 , n81976 );
buf ( n82428 , n82423 );
and ( n82429 , n82427 , n82428 );
nor ( n82430 , n82426 , n82429 );
buf ( n82431 , n82430 );
buf ( n82432 , n82431 );
nand ( n82433 , n82419 , n82432 );
buf ( n82434 , n82433 );
not ( n82435 , n82434 );
buf ( n82436 , n82395 );
buf ( n82437 , n82401 );
xor ( n82438 , n82436 , n82437 );
buf ( n82439 , n82002 );
xnor ( n82440 , n82438 , n82439 );
buf ( n82441 , n82440 );
buf ( n82442 , n82441 );
xor ( n82443 , n81578 , n81581 );
xor ( n82444 , n82443 , n81956 );
buf ( n82445 , n82444 );
buf ( n82446 , n82445 );
or ( n82447 , n82442 , n82446 );
buf ( n82448 , n82447 );
buf ( n82449 , n82448 );
buf ( n82450 , n82445 );
not ( n82451 , n82450 );
buf ( n82452 , n82441 );
not ( n82453 , n82452 );
or ( n82454 , n82451 , n82453 );
xor ( n82455 , n81235 , n81272 );
xor ( n82456 , n82455 , n81292 );
buf ( n82457 , n82456 );
buf ( n82458 , n82457 );
buf ( n82459 , C0 );
buf ( n82460 , n82459 );
xor ( n82461 , n82458 , n82460 );
buf ( n82462 , n81940 );
buf ( n82463 , n81951 );
xor ( n82464 , n82462 , n82463 );
buf ( n82465 , n81610 );
xor ( n82466 , n82464 , n82465 );
buf ( n82467 , n82466 );
buf ( n82468 , n82467 );
and ( n82469 , n82461 , n82468 );
or ( n82470 , n82469 , C0 );
buf ( n82471 , n82470 );
buf ( n82472 , n82471 );
not ( n82473 , n81586 );
not ( n82474 , n82473 );
not ( n82475 , n81953 );
or ( n82476 , n82474 , n82475 );
or ( n82477 , n81953 , n82473 );
nand ( n82478 , n82476 , n82477 );
not ( n82479 , n82478 );
not ( n82480 , n82479 );
or ( n82481 , C0 , n82480 );
nand ( n82482 , n82481 , C1 );
buf ( n82483 , n82482 );
buf ( n82484 , C0 );
buf ( n82485 , n82484 );
and ( n82486 , n82472 , n82483 );
or ( n82487 , C0 , n82486 );
buf ( n82488 , n82487 );
buf ( n82489 , n82488 );
nand ( n82490 , n82454 , n82489 );
buf ( n82491 , n82490 );
buf ( n82492 , n82491 );
and ( n82493 , n82449 , n82492 );
buf ( n82494 , n82493 );
buf ( n82495 , n82494 );
and ( n82496 , n82405 , n81993 );
not ( n82497 , n82405 );
and ( n82498 , n82497 , n82413 );
or ( n82499 , n82496 , n82498 );
xor ( n82500 , n82499 , n81998 );
buf ( n82501 , n82500 );
and ( n82502 , n82495 , n82501 );
buf ( n82503 , n82502 );
xnor ( n82504 , n82445 , n82488 );
xnor ( n82505 , n82504 , n82441 );
buf ( n82506 , n82505 );
buf ( n82507 , C0 );
buf ( n82508 , n82507 );
xor ( n82509 , n82044 , n82226 );
xor ( n82510 , n82509 , n82231 );
buf ( n82511 , n82510 );
buf ( n82512 , n82511 );
and ( n82513 , n52780 , n80269 );
not ( n82514 , n52780 );
and ( n82515 , n82514 , n45723 );
or ( n82516 , n82513 , n82515 );
buf ( n82517 , n82516 );
not ( n82518 , n82517 );
buf ( n82519 , n82518 );
or ( n82520 , n82519 , n46906 );
buf ( n82521 , n81883 );
not ( n82522 , n82521 );
buf ( n82523 , n82522 );
or ( n82524 , n82523 , n46905 );
nand ( n82525 , n82520 , n82524 );
buf ( n82526 , n82525 );
xor ( n82527 , n82049 , n82074 );
xor ( n82528 , n82527 , n82221 );
buf ( n82529 , n82528 );
buf ( n82530 , n82529 );
xor ( n82531 , n82526 , n82530 );
buf ( n82532 , n60545 );
not ( n82533 , n82532 );
buf ( n82534 , n82300 );
not ( n82535 , n82534 );
or ( n82536 , n82533 , n82535 );
and ( n82537 , n48836 , n48320 );
not ( n82538 , n48836 );
and ( n82539 , n82538 , n71078 );
or ( n82540 , n82537 , n82539 );
buf ( n82541 , n82540 );
buf ( n82542 , n51488 );
nand ( n82543 , n82541 , n82542 );
buf ( n82544 , n82543 );
buf ( n82545 , n82544 );
nand ( n82546 , n82536 , n82545 );
buf ( n82547 , n82546 );
buf ( n82548 , n82547 );
and ( n82549 , n82531 , n82548 );
and ( n82550 , n82526 , n82530 );
or ( n82551 , n82549 , n82550 );
buf ( n82552 , n82551 );
buf ( n82553 , n82552 );
buf ( n82554 , C0 );
buf ( n82555 , n82554 );
and ( n82556 , n82512 , n82553 );
or ( n82557 , C0 , n82556 );
buf ( n82558 , n82557 );
buf ( n82559 , n82558 );
xor ( n82560 , n82508 , n82559 );
xor ( n82561 , n82236 , n82261 );
xor ( n82562 , n82561 , n82267 );
buf ( n82563 , n82562 );
buf ( n82564 , n82563 );
and ( n82565 , n82560 , n82564 );
or ( n82566 , n82565 , C0 );
buf ( n82567 , n82566 );
buf ( n82568 , n82567 );
xor ( n82569 , n82016 , n82272 );
xor ( n82570 , n82569 , n82369 );
buf ( n82571 , n82570 );
buf ( n82572 , n82571 );
buf ( n82573 , C0 );
buf ( n82574 , n82573 );
and ( n82575 , n82568 , n82572 );
or ( n82576 , C0 , n82575 );
buf ( n82577 , n82576 );
buf ( n82578 , n82577 );
xor ( n82579 , n82384 , n82374 );
not ( n82580 , n82390 );
xor ( n82581 , n82579 , n82580 );
buf ( n82582 , n82581 );
xor ( n82583 , n82578 , n82582 );
xor ( n82584 , n82472 , n82483 );
xor ( n82585 , n82584 , n82485 );
buf ( n82586 , n82585 );
buf ( n82587 , n82586 );
and ( n82588 , n82583 , n82587 );
and ( n82589 , n82578 , n82582 );
or ( n82590 , n82588 , n82589 );
buf ( n82591 , n82590 );
buf ( n82592 , n82591 );
nor ( n82593 , n82506 , n82592 );
buf ( n82594 , n82593 );
xor ( n82595 , n81765 , n81781 );
xor ( n82596 , n82595 , n81841 );
xor ( n82597 , n82078 , n82179 );
xor ( n82598 , n82596 , n82597 );
buf ( n82599 , n82598 );
buf ( n82600 , n52777 );
not ( n82601 , n82600 );
buf ( n82602 , n46903 );
not ( n82603 , n82602 );
or ( n82604 , n82601 , n82603 );
buf ( n82605 , n81196 );
buf ( n82606 , n52777 );
not ( n82607 , n82606 );
buf ( n82608 , n82607 );
buf ( n82609 , n82608 );
nand ( n82610 , n82605 , n82609 );
buf ( n82611 , n82610 );
buf ( n82612 , n82611 );
nand ( n82613 , n82604 , n82612 );
buf ( n82614 , n82613 );
buf ( n82615 , n82614 );
not ( n82616 , n82615 );
buf ( n82617 , n48848 );
not ( n82618 , n82617 );
or ( n82619 , n82616 , n82618 );
buf ( n82620 , n82205 );
buf ( n82621 , n48865 );
nand ( n82622 , n82620 , n82621 );
buf ( n82623 , n82622 );
buf ( n82624 , n82623 );
nand ( n82625 , n82619 , n82624 );
buf ( n82626 , n82625 );
buf ( n82627 , n82626 );
xor ( n82628 , n82599 , n82627 );
buf ( n82629 , n71307 );
buf ( n82630 , n63003 );
and ( n82631 , n82629 , n82630 );
buf ( n82632 , n71310 );
buf ( n82633 , n64223 );
and ( n82634 , n82632 , n82633 );
nor ( n82635 , n82631 , n82634 );
buf ( n82636 , n82635 );
buf ( n82637 , n82636 );
buf ( n82638 , n64230 );
or ( n82639 , n82637 , n82638 );
buf ( n82640 , n82089 );
buf ( n82641 , n64227 );
or ( n82642 , n82640 , n82641 );
nand ( n82643 , n82639 , n82642 );
buf ( n82644 , n82643 );
buf ( n82645 , n82644 );
buf ( n82646 , n62935 );
buf ( n82647 , n62681 );
buf ( n82648 , n74115 );
and ( n82649 , n82647 , n82648 );
buf ( n82650 , n62684 );
buf ( n82651 , n74118 );
and ( n82652 , n82650 , n82651 );
nor ( n82653 , n82649 , n82652 );
buf ( n82654 , n82653 );
buf ( n82655 , n82654 );
or ( n82656 , n82646 , n82655 );
buf ( n82657 , n81820 );
buf ( n82658 , n62676 );
or ( n82659 , n82657 , n82658 );
nand ( n82660 , n82656 , n82659 );
buf ( n82661 , n82660 );
buf ( n82662 , n82661 );
xor ( n82663 , n82645 , n82662 );
buf ( n82664 , n60102 );
buf ( n82665 , n623 );
or ( n82666 , n82664 , n82665 );
buf ( n82667 , n60101 );
buf ( n82668 , n60261 );
buf ( n82669 , n623 );
and ( n82670 , n82667 , n82668 , n82669 );
buf ( n82671 , n60108 );
not ( n82672 , n82671 );
buf ( n82673 , n82672 );
buf ( n82674 , n82673 );
nor ( n82675 , n82670 , n82674 );
buf ( n82676 , n82675 );
buf ( n82677 , n82676 );
nand ( n82678 , n82666 , n82677 );
buf ( n82679 , n82678 );
buf ( n82680 , n82679 );
and ( n82681 , n82663 , n82680 );
and ( n82682 , n82645 , n82662 );
or ( n82683 , n82681 , n82682 );
buf ( n82684 , n82683 );
xor ( n82685 , n82097 , n82158 );
xor ( n82686 , n82685 , n82162 );
and ( n82687 , n82684 , n82686 );
buf ( n82688 , n82654 );
buf ( n82689 , n62676 );
or ( n82690 , n82688 , n82689 );
buf ( n82691 , n62687 );
nand ( n82692 , n82690 , n82691 );
buf ( n82693 , n82692 );
buf ( n82694 , n71801 );
buf ( n82695 , n63003 );
and ( n82696 , n82694 , n82695 );
buf ( n82697 , n71804 );
buf ( n82698 , n64223 );
and ( n82699 , n82697 , n82698 );
nor ( n82700 , n82696 , n82699 );
buf ( n82701 , n82700 );
buf ( n82702 , n82701 );
buf ( n82703 , n64230 );
or ( n82704 , n82702 , n82703 );
buf ( n82705 , n82636 );
buf ( n82706 , n64227 );
or ( n82707 , n82705 , n82706 );
nand ( n82708 , n82704 , n82707 );
buf ( n82709 , n82708 );
xor ( n82710 , n82693 , n82709 );
xor ( n82711 , n82146 , n82151 );
buf ( n82712 , n82711 );
and ( n82713 , n82710 , n82712 );
and ( n82714 , n82693 , n82709 );
or ( n82715 , n82713 , n82714 );
buf ( n82716 , n82715 );
xor ( n82717 , n82111 , n82128 );
xor ( n82718 , n82717 , n82154 );
buf ( n82719 , n82718 );
buf ( n82720 , n82719 );
xor ( n82721 , n82716 , n82720 );
xor ( n82722 , n82645 , n82662 );
xor ( n82723 , n82722 , n82680 );
buf ( n82724 , n82723 );
buf ( n82725 , n82724 );
and ( n82726 , n82721 , n82725 );
and ( n82727 , n82716 , n82720 );
or ( n82728 , n82726 , n82727 );
buf ( n82729 , n82728 );
xor ( n82730 , n82097 , n82158 );
xor ( n82731 , n82730 , n82162 );
and ( n82732 , n82729 , n82731 );
and ( n82733 , n82684 , n82729 );
or ( n82734 , n82687 , n82732 , n82733 );
buf ( n82735 , n82734 );
xor ( n82736 , n82166 , n82170 );
xor ( n82737 , n82736 , n82175 );
buf ( n82738 , n82737 );
buf ( n82739 , n82738 );
xor ( n82740 , n82735 , n82739 );
buf ( n82741 , n52456 );
not ( n82742 , n82741 );
buf ( n82743 , n24661 );
not ( n82744 , n82743 );
buf ( n82745 , n82744 );
and ( n82746 , n25879 , n82745 );
not ( n82747 , n25879 );
and ( n82748 , n82747 , n48836 );
or ( n82749 , n82746 , n82748 );
buf ( n82750 , n82749 );
not ( n82751 , n82750 );
or ( n82752 , n82742 , n82751 );
buf ( n82753 , n48836 );
buf ( n82754 , n82193 );
and ( n82755 , n82753 , n82754 );
not ( n82756 , n82753 );
buf ( n82757 , n82193 );
not ( n82758 , n82757 );
buf ( n82759 , n82758 );
buf ( n82760 , n82759 );
and ( n82761 , n82756 , n82760 );
nor ( n82762 , n82755 , n82761 );
buf ( n82763 , n82762 );
buf ( n82764 , n82763 );
buf ( n82765 , n51487 );
nand ( n82766 , n82764 , n82765 );
buf ( n82767 , n82766 );
buf ( n82768 , n82767 );
nand ( n82769 , n82752 , n82768 );
buf ( n82770 , n82769 );
buf ( n82771 , n82770 );
and ( n82772 , n82740 , n82771 );
and ( n82773 , n82735 , n82739 );
or ( n82774 , n82772 , n82773 );
buf ( n82775 , n82774 );
buf ( n82776 , n82775 );
xor ( n82777 , n82628 , n82776 );
buf ( n82778 , n82777 );
buf ( n82779 , n82778 );
buf ( n82780 , C0 );
buf ( n82781 , n82780 );
xor ( n82782 , n82779 , n82781 );
buf ( n82783 , n55841 );
not ( n82784 , n82783 );
buf ( n82785 , n45723 );
not ( n82786 , n82785 );
buf ( n82787 , n82786 );
buf ( n82788 , n82787 );
not ( n82789 , n82788 );
or ( n82790 , n82784 , n82789 );
buf ( n82791 , n45723 );
buf ( n82792 , n55840 );
nand ( n82793 , n82791 , n82792 );
buf ( n82794 , n82793 );
buf ( n82795 , n82794 );
nand ( n82796 , n82790 , n82795 );
buf ( n82797 , n82796 );
buf ( n82798 , n82797 );
not ( n82799 , n82798 );
buf ( n82800 , n80580 );
not ( n82801 , n82800 );
or ( n82802 , n82799 , n82801 );
buf ( n82803 , n53539 );
not ( n82804 , n82803 );
buf ( n82805 , n80269 );
not ( n82806 , n82805 );
or ( n82807 , n82804 , n82806 );
buf ( n82808 , n45723 );
buf ( n82809 , n53548 );
nand ( n82810 , n82808 , n82809 );
buf ( n82811 , n82810 );
buf ( n82812 , n82811 );
nand ( n82813 , n82807 , n82812 );
buf ( n82814 , n82813 );
buf ( n82815 , n82814 );
buf ( n82816 , n46912 );
nand ( n82817 , n82815 , n82816 );
buf ( n82818 , n82817 );
buf ( n82819 , n82818 );
nand ( n82820 , n82802 , n82819 );
buf ( n82821 , n82820 );
buf ( n82822 , n82821 );
and ( n82823 , n82782 , n82822 );
or ( n82824 , n82823 , C0 );
buf ( n82825 , n82824 );
buf ( n82826 , n82825 );
buf ( n82827 , n52456 );
not ( n82828 , n82827 );
buf ( n82829 , n82540 );
not ( n82830 , n82829 );
or ( n82831 , n82828 , n82830 );
buf ( n82832 , n51488 );
and ( n82833 , n25900 , n51493 );
not ( n82834 , n25900 );
and ( n82835 , n82834 , n48836 );
or ( n82836 , n82833 , n82835 );
buf ( n82837 , n82836 );
nand ( n82838 , n82832 , n82837 );
buf ( n82839 , n82838 );
buf ( n82840 , n82839 );
nand ( n82841 , n82831 , n82840 );
buf ( n82842 , n82841 );
buf ( n82843 , n82842 );
buf ( n82844 , n45746 );
buf ( n82845 , n45737 );
buf ( n82846 , n80269 );
nand ( n82847 , n82845 , n82846 );
buf ( n82848 , n82847 );
buf ( n82849 , n82848 );
buf ( n82850 , n12481 );
and ( n82851 , n82849 , n82850 );
and ( n82852 , n45724 , n45725 );
buf ( n82853 , n82852 );
buf ( n82854 , n82853 );
nor ( n82855 , n82851 , n82854 );
buf ( n82856 , n82855 );
buf ( n82857 , n82856 );
and ( n82858 , n82844 , n82857 );
buf ( n82859 , n82858 );
buf ( n82860 , n82859 );
xor ( n82861 , n82843 , n82860 );
buf ( n82862 , n52456 );
not ( n82863 , n82862 );
buf ( n82864 , n82836 );
not ( n82865 , n82864 );
or ( n82866 , n82863 , n82865 );
buf ( n82867 , n82749 );
buf ( n82868 , n51488 );
nand ( n82869 , n82867 , n82868 );
buf ( n82870 , n82869 );
buf ( n82871 , n82870 );
nand ( n82872 , n82866 , n82871 );
buf ( n82873 , n82872 );
buf ( n82874 , n82873 );
buf ( n82875 , n45727 );
buf ( n82876 , n12481 );
nand ( n82877 , n82875 , n82876 );
buf ( n82878 , n82877 );
buf ( n82879 , n82878 );
not ( n82880 , n82879 );
buf ( n82881 , n82880 );
buf ( n82882 , n82881 );
xor ( n82883 , n82874 , n82882 );
buf ( n82884 , n53539 );
not ( n82885 , n82884 );
buf ( n82886 , n46903 );
not ( n82887 , n82886 );
or ( n82888 , n82885 , n82887 );
buf ( n82889 , n53548 );
buf ( n82890 , n24714 );
nand ( n82891 , n82889 , n82890 );
buf ( n82892 , n82891 );
buf ( n82893 , n82892 );
nand ( n82894 , n82888 , n82893 );
buf ( n82895 , n82894 );
buf ( n82896 , n82895 );
not ( n82897 , n82896 );
buf ( n82898 , n48848 );
not ( n82899 , n82898 );
or ( n82900 , n82897 , n82899 );
buf ( n82901 , n48865 );
buf ( n82902 , n82614 );
nand ( n82903 , n82901 , n82902 );
buf ( n82904 , n82903 );
buf ( n82905 , n82904 );
nand ( n82906 , n82900 , n82905 );
buf ( n82907 , n82906 );
buf ( n82908 , n82907 );
xor ( n82909 , n82735 , n82739 );
xor ( n82910 , n82909 , n82771 );
buf ( n82911 , n82910 );
buf ( n82912 , n82911 );
xor ( n82913 , n82908 , n82912 );
buf ( n82914 , n45723 );
buf ( n82915 , n24750 );
buf ( n82916 , n81196 );
or ( n82917 , n82915 , n82916 );
buf ( n82918 , n12481 );
nand ( n82919 , n82917 , n82918 );
buf ( n82920 , n82919 );
buf ( n82921 , n82920 );
buf ( n82922 , n81196 );
buf ( n82923 , n24750 );
nand ( n82924 , n82922 , n82923 );
buf ( n82925 , n82924 );
buf ( n82926 , n82925 );
and ( n82927 , n82914 , n82921 , n82926 );
buf ( n82928 , n82927 );
buf ( n82929 , n82928 );
and ( n82930 , n82913 , n82929 );
and ( n82931 , n82908 , n82912 );
or ( n82932 , n82930 , n82931 );
buf ( n82933 , n82932 );
buf ( n82934 , n82933 );
and ( n82935 , n82883 , n82934 );
and ( n82936 , n82874 , n82882 );
or ( n82937 , n82935 , n82936 );
buf ( n82938 , n82937 );
buf ( n82939 , n82938 );
xor ( n82940 , n82861 , n82939 );
buf ( n82941 , n82940 );
buf ( n82942 , n82941 );
buf ( n82943 , C0 );
buf ( n82944 , n82943 );
and ( n82945 , n82826 , n82942 );
or ( n82946 , C0 , n82945 );
buf ( n82947 , n82946 );
buf ( n82948 , n82947 );
xor ( n82949 , n82185 , n82189 );
xor ( n82950 , n82949 , n82216 );
buf ( n82951 , n82950 );
buf ( n82952 , n82951 );
xor ( n82953 , n82599 , n82627 );
and ( n82954 , n82953 , n82776 );
and ( n82955 , n82599 , n82627 );
or ( n82956 , n82954 , n82955 );
buf ( n82957 , n82956 );
buf ( n82958 , n82957 );
xor ( n82959 , n82952 , n82958 );
buf ( n82960 , n80281 );
not ( n82961 , n82960 );
buf ( n82962 , n82516 );
not ( n82963 , n82962 );
or ( n82964 , n82961 , n82963 );
buf ( n82965 , n82814 );
buf ( n82966 , n80580 );
nand ( n82967 , n82965 , n82966 );
buf ( n82968 , n82967 );
buf ( n82969 , n82968 );
nand ( n82970 , n82964 , n82969 );
buf ( n82971 , n82970 );
buf ( n82972 , n82971 );
xor ( n82973 , n82959 , n82972 );
buf ( n82974 , n82973 );
buf ( n82975 , n82974 );
buf ( n82976 , C0 );
buf ( n82977 , n82976 );
xor ( n82978 , n82975 , n82977 );
buf ( n82979 , n67149 );
not ( n82980 , n82979 );
buf ( n82981 , n55841 );
not ( n82982 , n82981 );
buf ( n82983 , n76179 );
not ( n82984 , n82983 );
or ( n82985 , n82982 , n82984 );
buf ( n82986 , n44494 );
buf ( n82987 , n55840 );
nand ( n82988 , n82986 , n82987 );
buf ( n82989 , n82988 );
buf ( n82990 , n82989 );
nand ( n82991 , n82985 , n82990 );
buf ( n82992 , n82991 );
buf ( n82993 , n82992 );
not ( n82994 , n82993 );
or ( n82995 , n82980 , n82994 );
buf ( n82996 , n45741 );
buf ( n82997 , n12481 );
not ( n82998 , n82997 );
buf ( n82999 , n76179 );
not ( n83000 , n82999 );
or ( n83001 , n82998 , n83000 );
buf ( n83002 , n45746 );
buf ( n83003 , n56325 );
nand ( n83004 , n83002 , n83003 );
buf ( n83005 , n83004 );
buf ( n83006 , n83005 );
nand ( n83007 , n83001 , n83006 );
buf ( n83008 , n83007 );
buf ( n83009 , n83008 );
nand ( n83010 , n82996 , n83009 );
buf ( n83011 , n83010 );
buf ( n83012 , n83011 );
nand ( n83013 , n82995 , n83012 );
buf ( n83014 , n83013 );
buf ( n83015 , n83014 );
and ( n83016 , n82978 , n83015 );
or ( n83017 , n83016 , C0 );
buf ( n83018 , n83017 );
buf ( n83019 , n83018 );
xor ( n83020 , n82948 , n83019 );
xor ( n83021 , n82952 , n82958 );
and ( n83022 , n83021 , n82972 );
and ( n83023 , n82952 , n82958 );
or ( n83024 , n83022 , n83023 );
buf ( n83025 , n83024 );
buf ( n83026 , n83025 );
buf ( n83027 , n82992 );
not ( n83028 , n83027 );
buf ( n83029 , n45741 );
not ( n83030 , n83029 );
or ( n83031 , n83028 , n83030 );
buf ( n83032 , n67149 );
buf ( n83033 , n82320 );
nand ( n83034 , n83032 , n83033 );
buf ( n83035 , n83034 );
buf ( n83036 , n83035 );
nand ( n83037 , n83031 , n83036 );
buf ( n83038 , n83037 );
buf ( n83039 , n83038 );
xor ( n83040 , n83026 , n83039 );
buf ( n83041 , n44495 );
buf ( n83042 , n56325 );
nor ( n83043 , n83041 , n83042 );
buf ( n83044 , n83043 );
buf ( n83045 , n83044 );
xor ( n83046 , n83040 , n83045 );
buf ( n83047 , n83046 );
buf ( n83048 , n83047 );
and ( n83049 , n83020 , n83048 );
and ( n83050 , n82948 , n83019 );
or ( n83051 , n83049 , n83050 );
buf ( n83052 , n83051 );
buf ( n83053 , n83052 );
xor ( n83054 , n83026 , n83039 );
and ( n83055 , n83054 , n83045 );
and ( n83056 , n83026 , n83039 );
or ( n83057 , n83055 , n83056 );
buf ( n83058 , n83057 );
buf ( n83059 , n83058 );
xor ( n83060 , n82308 , n82333 );
xor ( n83061 , n83060 , n82346 );
buf ( n83062 , n83061 );
buf ( n83063 , n83062 );
xor ( n83064 , n83059 , n83063 );
buf ( n83065 , n12481 );
not ( n83066 , n83065 );
buf ( n83067 , n79031 );
not ( n83068 , n83067 );
or ( n83069 , n83066 , n83068 );
buf ( n83070 , n41570 );
buf ( n83071 , n56325 );
nand ( n83072 , n83070 , n83071 );
buf ( n83073 , n83072 );
buf ( n83074 , n83073 );
nand ( n83075 , n83069 , n83074 );
buf ( n83076 , n83075 );
buf ( n83077 , n83076 );
not ( n83078 , n83077 );
buf ( n83079 , n74488 );
not ( n83080 , n83079 );
or ( n83081 , n83078 , n83080 );
nand ( n83082 , n82281 , n44496 );
buf ( n83083 , n83082 );
nand ( n83084 , n83081 , n83083 );
buf ( n83085 , n83084 );
buf ( n83086 , n83085 );
xor ( n83087 , n83064 , n83086 );
buf ( n83088 , n83087 );
buf ( n83089 , n83088 );
xor ( n83090 , n83053 , n83089 );
xor ( n83091 , n82843 , n82860 );
and ( n83092 , n83091 , n82939 );
and ( n83093 , n82843 , n82860 );
or ( n83094 , n83092 , n83093 );
buf ( n83095 , n83094 );
buf ( n83096 , n83095 );
xor ( n83097 , n82526 , n82530 );
xor ( n83098 , n83097 , n82548 );
buf ( n83099 , n83098 );
buf ( n83100 , n83099 );
buf ( n83101 , C0 );
buf ( n83102 , n83101 );
and ( n83103 , n83096 , n83100 );
or ( n83104 , C0 , n83103 );
buf ( n83105 , n83104 );
buf ( n83106 , n83105 );
xor ( n83107 , n82512 , n82553 );
xor ( n83108 , n83107 , n82555 );
buf ( n83109 , n83108 );
buf ( n83110 , n83109 );
xor ( n83111 , n83106 , n83110 );
buf ( n83112 , C0 );
xor ( n83113 , n83111 , n83112 );
buf ( n83114 , n83113 );
buf ( n83115 , n83114 );
and ( n83116 , n83090 , n83115 );
and ( n83117 , n83053 , n83089 );
or ( n83118 , n83116 , n83117 );
buf ( n83119 , n83118 );
buf ( n83120 , n83119 );
not ( n83121 , n83120 );
xor ( n83122 , n83059 , n83063 );
and ( n83123 , n83122 , n83086 );
and ( n83124 , n83059 , n83063 );
or ( n83125 , n83123 , n83124 );
buf ( n83126 , n83125 );
buf ( n83127 , n83126 );
buf ( n83128 , n82350 );
not ( n83129 , n83128 );
buf ( n83130 , n83129 );
buf ( n83131 , n83130 );
not ( n83132 , n83131 );
buf ( n83133 , n82357 );
not ( n83134 , n83133 );
or ( n83135 , n83132 , n83134 );
buf ( n83136 , n82350 );
buf ( n83137 , n82354 );
nand ( n83138 , n83136 , n83137 );
buf ( n83139 , n83138 );
buf ( n83140 , n83139 );
nand ( n83141 , n83135 , n83140 );
buf ( n83142 , n83141 );
buf ( n83143 , n83142 );
buf ( n83144 , n82290 );
and ( n83145 , n83143 , n83144 );
not ( n83146 , n83143 );
buf ( n83147 , n82290 );
not ( n83148 , n83147 );
buf ( n83149 , n83148 );
buf ( n83150 , n83149 );
and ( n83151 , n83146 , n83150 );
nor ( n83152 , n83145 , n83151 );
buf ( n83153 , n83152 );
buf ( n83154 , n83153 );
xor ( n83155 , n83127 , n83154 );
buf ( n83156 , C0 );
buf ( n83157 , n83156 );
xor ( n83158 , n83155 , n83157 );
buf ( n83159 , n83158 );
and ( n83160 , n83106 , n83110 );
or ( n83161 , C0 , n83160 );
buf ( n83162 , n83161 );
buf ( n83163 , n83162 );
xor ( n83164 , n82508 , n82559 );
xor ( n83165 , n83164 , n82564 );
buf ( n83166 , n83165 );
buf ( n83167 , n83166 );
not ( n83168 , n83167 );
buf ( n83169 , n83168 );
buf ( n83170 , n83169 );
and ( n83171 , n83163 , n83170 );
not ( n83172 , n83163 );
buf ( n83173 , n83166 );
and ( n83174 , n83172 , n83173 );
nor ( n83175 , n83171 , n83174 );
buf ( n83176 , n83175 );
xor ( n83177 , n83159 , n83176 );
buf ( n83178 , n83177 );
nand ( n83179 , n83121 , n83178 );
buf ( n83180 , n83179 );
not ( n83181 , n83180 );
xor ( n83182 , n82779 , n82781 );
xor ( n83183 , n83182 , n82822 );
buf ( n83184 , n83183 );
buf ( n83185 , n83184 );
buf ( n83186 , n62659 );
buf ( n83187 , n623 );
and ( n83188 , n83186 , n83187 );
buf ( n83189 , n62681 );
buf ( n83190 , n62662 );
buf ( n83191 , n75821 );
and ( n83192 , n83190 , n83191 );
buf ( n83193 , n62668 );
nor ( n83194 , n83192 , n83193 );
buf ( n83195 , n83194 );
buf ( n83196 , n83195 );
nor ( n83197 , n83188 , n83189 , n83196 );
buf ( n83198 , n83197 );
buf ( n83199 , n83198 );
buf ( n83200 , n71818 );
buf ( n83201 , n63003 );
and ( n83202 , n83200 , n83201 );
buf ( n83203 , n71821 );
buf ( n83204 , n64223 );
and ( n83205 , n83203 , n83204 );
nor ( n83206 , n83202 , n83205 );
buf ( n83207 , n83206 );
buf ( n83208 , n83207 );
buf ( n83209 , n64230 );
or ( n83210 , n83208 , n83209 );
buf ( n83211 , n82701 );
buf ( n83212 , n64227 );
or ( n83213 , n83211 , n83212 );
nand ( n83214 , n83210 , n83213 );
buf ( n83215 , n83214 );
buf ( n83216 , n83215 );
xor ( n83217 , n83199 , n83216 );
buf ( n83218 , n64141 );
buf ( n83219 , n62668 );
buf ( n83220 , n74115 );
and ( n83221 , n83219 , n83220 );
buf ( n83222 , n63015 );
buf ( n83223 , n74118 );
and ( n83224 , n83222 , n83223 );
nor ( n83225 , n83221 , n83224 );
buf ( n83226 , n83225 );
buf ( n83227 , n83226 );
or ( n83228 , n83218 , n83227 );
buf ( n83229 , n82138 );
buf ( n83230 , n63010 );
or ( n83231 , n83229 , n83230 );
nand ( n83232 , n83228 , n83231 );
buf ( n83233 , n83232 );
buf ( n83234 , n83233 );
and ( n83235 , n83217 , n83234 );
and ( n83236 , n83199 , n83216 );
or ( n83237 , n83235 , n83236 );
buf ( n83238 , n83237 );
xor ( n83239 , n82693 , n82709 );
xor ( n83240 , n83239 , n82712 );
and ( n83241 , n83238 , n83240 );
buf ( n83242 , n62676 );
buf ( n83243 , n75821 );
nor ( n83244 , n83242 , n83243 );
buf ( n83245 , n83244 );
buf ( n83246 , n83245 );
buf ( n83247 , n83226 );
buf ( n83248 , n63010 );
or ( n83249 , n83247 , n83248 );
buf ( n83250 , n63018 );
nand ( n83251 , n83249 , n83250 );
buf ( n83252 , n83251 );
buf ( n83253 , n83252 );
and ( n83254 , n83246 , n83253 );
buf ( n83255 , n83254 );
buf ( n83256 , n83255 );
buf ( n83257 , n62687 );
buf ( n83258 , n623 );
or ( n83259 , n83257 , n83258 );
buf ( n83260 , n62679 );
buf ( n83261 , n62681 );
buf ( n83262 , n623 );
and ( n83263 , n83260 , n83261 , n83262 );
buf ( n83264 , n62695 );
not ( n83265 , n83264 );
buf ( n83266 , n83265 );
buf ( n83267 , n83266 );
nor ( n83268 , n83263 , n83267 );
buf ( n83269 , n83268 );
buf ( n83270 , n83269 );
nand ( n83271 , n83259 , n83270 );
buf ( n83272 , n83271 );
buf ( n83273 , n83272 );
xor ( n83274 , n83256 , n83273 );
xor ( n83275 , n83199 , n83216 );
xor ( n83276 , n83275 , n83234 );
buf ( n83277 , n83276 );
buf ( n83278 , n83277 );
and ( n83279 , n83274 , n83278 );
and ( n83280 , n83256 , n83273 );
or ( n83281 , n83279 , n83280 );
buf ( n83282 , n83281 );
xor ( n83283 , n82693 , n82709 );
xor ( n83284 , n83283 , n82712 );
and ( n83285 , n83282 , n83284 );
and ( n83286 , n83238 , n83282 );
or ( n83287 , n83241 , n83285 , n83286 );
xor ( n83288 , n82716 , n82720 );
xor ( n83289 , n83288 , n82725 );
buf ( n83290 , n83289 );
or ( n83291 , n83287 , n83290 );
not ( n83292 , n83291 );
not ( n83293 , n51487 );
not ( n83294 , n53539 );
not ( n83295 , n48839 );
or ( n83296 , n83294 , n83295 );
buf ( n83297 , n53548 );
buf ( n83298 , n48836 );
nand ( n83299 , n83297 , n83298 );
buf ( n83300 , n83299 );
nand ( n83301 , n83296 , n83300 );
not ( n83302 , n83301 );
or ( n83303 , n83293 , n83302 );
buf ( n83304 , n52777 );
buf ( n83305 , n48836 );
and ( n83306 , n83304 , n83305 );
not ( n83307 , n83304 );
buf ( n83308 , n82745 );
and ( n83309 , n83307 , n83308 );
nor ( n83310 , n83306 , n83309 );
buf ( n83311 , n83310 );
nand ( n83312 , n83311 , n52456 );
nand ( n83313 , n83303 , n83312 );
not ( n83314 , n83313 );
or ( n83315 , n83292 , n83314 );
nand ( n83316 , n83287 , n83290 );
nand ( n83317 , n83315 , n83316 );
not ( n83318 , n83317 );
buf ( n83319 , n52456 );
not ( n83320 , n83319 );
buf ( n83321 , n82763 );
not ( n83322 , n83321 );
or ( n83323 , n83320 , n83322 );
nand ( n83324 , n83311 , n51487 );
buf ( n83325 , n83324 );
nand ( n83326 , n83323 , n83325 );
buf ( n83327 , n83326 );
buf ( n83328 , n83327 );
xor ( n83329 , n82097 , n82158 );
xor ( n83330 , n83329 , n82162 );
xor ( n83331 , n82684 , n82729 );
xor ( n83332 , n83330 , n83331 );
buf ( n83333 , n83332 );
or ( n83334 , n83328 , n83333 );
buf ( n83335 , n83334 );
not ( n83336 , n83335 );
or ( n83337 , n83318 , n83336 );
buf ( n83338 , n83327 );
buf ( n83339 , n83332 );
nand ( n83340 , n83338 , n83339 );
buf ( n83341 , n83340 );
nand ( n83342 , n83337 , n83341 );
buf ( n83343 , n83342 );
not ( n83344 , n83343 );
buf ( n83345 , n12481 );
not ( n83346 , n83345 );
buf ( n83347 , n82787 );
not ( n83348 , n83347 );
or ( n83349 , n83346 , n83348 );
buf ( n83350 , n45723 );
buf ( n83351 , n56325 );
nand ( n83352 , n83350 , n83351 );
buf ( n83353 , n83352 );
buf ( n83354 , n83353 );
nand ( n83355 , n83349 , n83354 );
buf ( n83356 , n83355 );
buf ( n83357 , n83356 );
not ( n83358 , n83357 );
buf ( n83359 , n80580 );
not ( n83360 , n83359 );
or ( n83361 , n83358 , n83360 );
buf ( n83362 , n82797 );
buf ( n83363 , n80281 );
nand ( n83364 , n83362 , n83363 );
buf ( n83365 , n83364 );
buf ( n83366 , n83365 );
nand ( n83367 , n83361 , n83366 );
buf ( n83368 , n83367 );
buf ( n83369 , n83368 );
not ( n83370 , n83369 );
or ( n83371 , n83344 , n83370 );
buf ( n83372 , n83342 );
buf ( n83373 , n83368 );
or ( n83374 , n83372 , n83373 );
not ( n83375 , n48848 );
buf ( n83376 , n55840 );
buf ( n83377 , n81196 );
and ( n83378 , n83376 , n83377 );
not ( n83379 , n83376 );
buf ( n83380 , n46903 );
and ( n83381 , n83379 , n83380 );
nor ( n83382 , n83378 , n83381 );
buf ( n83383 , n83382 );
not ( n83384 , n83383 );
not ( n83385 , n83384 );
or ( n83386 , n83375 , n83385 );
nand ( n83387 , n82895 , n48865 );
nand ( n83388 , n83386 , n83387 );
not ( n83389 , n83388 );
buf ( n83390 , n83389 );
not ( n83391 , n83390 );
or ( n83392 , n83391 , C0 );
buf ( n83393 , n48831 );
buf ( n83394 , n82745 );
nand ( n83395 , n83393 , n83394 );
buf ( n83396 , n83395 );
and ( n83397 , n12481 , n83396 );
buf ( n83398 , n82745 );
not ( n83399 , n83398 );
buf ( n83400 , n83399 );
and ( n83401 , n48834 , n83400 );
nor ( n83402 , n83397 , n83401 , n46903 );
buf ( n83403 , n83402 );
xor ( n83404 , n83287 , n83290 );
and ( n83405 , n83313 , n83404 );
not ( n83406 , n83313 );
not ( n83407 , n83404 );
and ( n83408 , n83406 , n83407 );
nor ( n83409 , n83405 , n83408 );
buf ( n83410 , n83409 );
buf ( n83411 , C0 );
buf ( n83412 , n83411 );
and ( n83413 , n83403 , n83410 );
or ( n83414 , C0 , n83413 );
buf ( n83415 , n83414 );
buf ( n83416 , n83415 );
nand ( n83417 , n83392 , n83416 );
buf ( n83418 , n83417 );
buf ( n83419 , n83418 );
nand ( n83420 , C1 , n83419 );
buf ( n83421 , n83420 );
buf ( n83422 , n83421 );
nand ( n83423 , n83374 , n83422 );
buf ( n83424 , n83423 );
buf ( n83425 , n83424 );
nand ( n83426 , n83371 , n83425 );
buf ( n83427 , n83426 );
buf ( n83428 , n83427 );
not ( n83429 , n83428 );
xor ( n83430 , n82874 , n82882 );
xor ( n83431 , n83430 , n82934 );
buf ( n83432 , n83431 );
buf ( n83433 , n83432 );
not ( n83434 , n83433 );
buf ( n83435 , n83434 );
buf ( n83436 , n83435 );
nand ( n83437 , n83429 , n83436 );
buf ( n83438 , n83437 );
buf ( n83439 , n83438 );
and ( n83440 , n83185 , n83439 );
buf ( n83441 , n83427 );
not ( n83442 , n83441 );
buf ( n83443 , n83435 );
nor ( n83444 , n83442 , n83443 );
buf ( n83445 , n83444 );
buf ( n83446 , n83445 );
nor ( n83447 , n83440 , n83446 );
buf ( n83448 , n83447 );
buf ( n83449 , n83448 );
not ( n83450 , n83449 );
xor ( n83451 , n82826 , n82942 );
xor ( n83452 , n83451 , n82944 );
buf ( n83453 , n83452 );
buf ( n83454 , n83453 );
not ( n83455 , n83454 );
buf ( n83456 , n83455 );
buf ( n83457 , n83456 );
not ( n83458 , n83457 );
or ( n83459 , n83450 , n83458 );
xor ( n83460 , n82975 , n82977 );
xor ( n83461 , n83460 , n83015 );
buf ( n83462 , n83461 );
buf ( n83463 , n83462 );
nand ( n83464 , n83459 , n83463 );
buf ( n83465 , n83464 );
buf ( n83466 , n83465 );
buf ( n83467 , n83448 );
not ( n83468 , n83467 );
buf ( n83469 , n83453 );
nand ( n83470 , n83468 , n83469 );
buf ( n83471 , n83470 );
buf ( n83472 , n83471 );
nand ( n83473 , n83466 , n83472 );
buf ( n83474 , n83473 );
buf ( n83475 , n83474 );
buf ( n83476 , n83342 );
buf ( n83477 , n83368 );
xor ( n83478 , n83476 , n83477 );
buf ( n83479 , n83421 );
xnor ( n83480 , n83478 , n83479 );
buf ( n83481 , n83480 );
buf ( n83482 , n83481 );
buf ( n83483 , C1 );
buf ( n83484 , n83483 );
xor ( n83485 , n83482 , n83484 );
buf ( n83486 , C0 );
buf ( n83487 , n83486 );
xor ( n83488 , n82908 , n82912 );
xor ( n83489 , n83488 , n82929 );
buf ( n83490 , n83489 );
buf ( n83491 , n83490 );
xor ( n83492 , n83487 , n83491 );
buf ( n83493 , n56325 );
not ( n83494 , n83493 );
buf ( n83495 , n80281 );
nand ( n83496 , n83494 , n83495 );
buf ( n83497 , n83496 );
buf ( n83498 , n83497 );
buf ( n83499 , n83332 );
buf ( n83500 , n83327 );
xor ( n83501 , n83499 , n83500 );
buf ( n83502 , n83317 );
xnor ( n83503 , n83501 , n83502 );
buf ( n83504 , n83503 );
buf ( n83505 , n83504 );
nand ( n83506 , n83498 , n83505 );
buf ( n83507 , n83506 );
buf ( n83508 , n83507 );
not ( n83509 , n83508 );
xor ( n83510 , n82693 , n82709 );
xor ( n83511 , n83510 , n82712 );
xor ( n83512 , n83238 , n83282 );
xor ( n83513 , n83511 , n83512 );
buf ( n83514 , n83513 );
not ( n83515 , n83514 );
buf ( n83516 , n83515 );
buf ( n83517 , n83516 );
not ( n83518 , n83517 );
not ( n83519 , n51487 );
buf ( n83520 , n55841 );
not ( n83521 , n83520 );
buf ( n83522 , n48839 );
not ( n83523 , n83522 );
or ( n83524 , n83521 , n83523 );
buf ( n83525 , n83400 );
buf ( n83526 , n55840 );
nand ( n83527 , n83525 , n83526 );
buf ( n83528 , n83527 );
buf ( n83529 , n83528 );
nand ( n83530 , n83524 , n83529 );
buf ( n83531 , n83530 );
not ( n83532 , n83531 );
or ( n83533 , n83519 , n83532 );
nand ( n83534 , n83301 , n52456 );
nand ( n83535 , n83533 , n83534 );
buf ( n83536 , n83535 );
not ( n83537 , n83536 );
buf ( n83538 , n83537 );
buf ( n83539 , n83538 );
not ( n83540 , n83539 );
or ( n83541 , n83518 , n83540 );
buf ( n83542 , n51482 );
buf ( n83543 , C0 );
nor ( n83544 , n83542 , n83543 );
buf ( n83545 , n83544 );
buf ( n83546 , n83545 );
buf ( n83547 , n56325 );
or ( n83548 , n83546 , n83547 );
buf ( n83549 , C1 );
buf ( n83550 , n83549 );
nand ( n83551 , n83548 , n83550 );
buf ( n83552 , n83551 );
not ( n83553 , n83552 );
nand ( n83554 , n83553 , n48836 );
not ( n83555 , n83554 );
xor ( n83556 , n83246 , n83253 );
buf ( n83557 , n83556 );
buf ( n83558 , n83557 );
buf ( n83559 , n63003 );
buf ( n83560 , n72445 );
and ( n83561 , n83559 , n83560 );
buf ( n83562 , n64223 );
buf ( n83563 , n72448 );
and ( n83564 , n83562 , n83563 );
nor ( n83565 , n83561 , n83564 );
buf ( n83566 , n83565 );
buf ( n83567 , n83566 );
buf ( n83568 , n64230 );
or ( n83569 , n83567 , n83568 );
buf ( n83570 , n83207 );
buf ( n83571 , n64227 );
or ( n83572 , n83570 , n83571 );
nand ( n83573 , n83569 , n83572 );
buf ( n83574 , n83573 );
buf ( n83575 , n83574 );
xor ( n83576 , n83558 , n83575 );
buf ( n83577 , n63003 );
buf ( n83578 , n74115 );
and ( n83579 , n83577 , n83578 );
buf ( n83580 , n64223 );
buf ( n83581 , n74118 );
and ( n83582 , n83580 , n83581 );
nor ( n83583 , n83579 , n83582 );
buf ( n83584 , n83583 );
buf ( n83585 , n83584 );
buf ( n83586 , n64230 );
or ( n83587 , n83585 , n83586 );
buf ( n83588 , n83566 );
buf ( n83589 , n64227 );
or ( n83590 , n83588 , n83589 );
nand ( n83591 , n83587 , n83590 );
buf ( n83592 , n83591 );
buf ( n83593 , n83592 );
buf ( n83594 , n6932 );
buf ( n83595 , n623 );
and ( n83596 , n83594 , n83595 );
buf ( n83597 , n62668 );
buf ( n83598 , n62990 );
buf ( n83599 , n75821 );
and ( n83600 , n83598 , n83599 );
buf ( n83601 , n63003 );
nor ( n83602 , n83600 , n83601 );
buf ( n83603 , n83602 );
buf ( n83604 , n83603 );
nor ( n83605 , n83596 , n83597 , n83604 );
buf ( n83606 , n83605 );
buf ( n83607 , n83606 );
xor ( n83608 , n83593 , n83607 );
buf ( n83609 , n63018 );
buf ( n83610 , n623 );
or ( n83611 , n83609 , n83610 );
buf ( n83612 , n63013 );
buf ( n83613 , n64129 );
buf ( n83614 , n623 );
and ( n83615 , n83612 , n83613 , n83614 );
buf ( n83616 , n63026 );
not ( n83617 , n83616 );
buf ( n83618 , n83617 );
buf ( n83619 , n83618 );
nor ( n83620 , n83615 , n83619 );
buf ( n83621 , n83620 );
buf ( n83622 , n83621 );
nand ( n83623 , n83611 , n83622 );
buf ( n83624 , n83623 );
buf ( n83625 , n83624 );
and ( n83626 , n83608 , n83625 );
and ( n83627 , n83593 , n83607 );
or ( n83628 , n83626 , n83627 );
buf ( n83629 , n83628 );
buf ( n83630 , n83629 );
and ( n83631 , n83576 , n83630 );
and ( n83632 , n83558 , n83575 );
or ( n83633 , n83631 , n83632 );
buf ( n83634 , n83633 );
buf ( n83635 , n83634 );
not ( n83636 , n83635 );
buf ( n83637 , n83636 );
not ( n83638 , n83637 );
and ( n83639 , n83555 , n83638 );
buf ( n83640 , n83637 );
buf ( n83641 , n83554 );
nand ( n83642 , n83640 , n83641 );
buf ( n83643 , n83642 );
xor ( n83644 , n83256 , n83273 );
xor ( n83645 , n83644 , n83278 );
buf ( n83646 , n83645 );
and ( n83647 , n83643 , n83646 );
nor ( n83648 , n83639 , n83647 );
buf ( n83649 , n83648 );
not ( n83650 , n83649 );
buf ( n83651 , n83650 );
buf ( n83652 , n83651 );
nand ( n83653 , n83541 , n83652 );
buf ( n83654 , n83653 );
buf ( n83655 , n83535 );
buf ( n83656 , n83513 );
nand ( n83657 , n83655 , n83656 );
buf ( n83658 , n83657 );
nand ( n83659 , n83654 , n83658 );
buf ( n83660 , n56325 );
buf ( n83661 , n81196 );
xnor ( n83662 , n83660 , n83661 );
buf ( n83663 , n83662 );
not ( n83664 , n83663 );
not ( n83665 , n48848 );
or ( n83666 , n83664 , n83665 );
buf ( n83667 , n83383 );
not ( n83668 , n83667 );
buf ( n83669 , n48865 );
nand ( n83670 , n83668 , n83669 );
buf ( n83671 , n83670 );
nand ( n83672 , n83666 , n83671 );
xor ( n83673 , n83659 , n83672 );
buf ( n83674 , n48862 );
buf ( n83675 , n12481 );
nand ( n83676 , n83674 , n83675 );
buf ( n83677 , n83676 );
not ( n83678 , n83535 );
not ( n83679 , n83516 );
not ( n83680 , n83651 );
or ( n83681 , n83679 , n83680 );
buf ( n83682 , n83513 );
buf ( n83683 , n83648 );
nand ( n83684 , n83682 , n83683 );
buf ( n83685 , n83684 );
nand ( n83686 , n83681 , n83685 );
not ( n83687 , n83686 );
or ( n83688 , n83678 , n83687 );
nand ( n83689 , n83651 , n83516 );
not ( n83690 , n83535 );
nand ( n83691 , n83689 , n83690 , n83685 );
nand ( n83692 , n83688 , n83691 );
buf ( n83693 , n83692 );
not ( n83694 , n83693 );
buf ( n83695 , n83694 );
buf ( n83696 , n83695 );
buf ( n83697 , n83677 );
nand ( n83698 , C1 , n83697 );
buf ( n83699 , n83698 );
buf ( n83700 , n83699 );
nand ( n83701 , n83696 , n83700 );
buf ( n83702 , n83701 );
nand ( n83703 , C1 , n83702 );
and ( n83704 , n83673 , n83703 );
and ( n83705 , n83659 , n83672 );
or ( n83706 , n83704 , n83705 );
buf ( n83707 , n83706 );
not ( n83708 , n83707 );
or ( n83709 , n83509 , n83708 );
buf ( n83710 , n83497 );
not ( n83711 , n83710 );
buf ( n83712 , n83711 );
buf ( n83713 , n83712 );
buf ( n83714 , n83504 );
not ( n83715 , n83714 );
buf ( n83716 , n83715 );
buf ( n83717 , n83716 );
nand ( n83718 , n83713 , n83717 );
buf ( n83719 , n83718 );
buf ( n83720 , n83719 );
nand ( n83721 , n83709 , n83720 );
buf ( n83722 , n83721 );
buf ( n83723 , n83722 );
xnor ( n83724 , n83492 , n83723 );
buf ( n83725 , n83724 );
buf ( n83726 , n83725 );
xor ( n83727 , n83485 , n83726 );
buf ( n83728 , n83727 );
buf ( n83729 , n83728 );
buf ( n83730 , n83388 );
not ( n83731 , n83730 );
or ( n83732 , n83731 , C0 );
buf ( n83733 , C1 );
buf ( n83734 , n83733 );
nand ( n83735 , n83732 , n83734 );
buf ( n83736 , n83735 );
buf ( n83737 , n83736 );
buf ( n83738 , n83415 );
xnor ( n83739 , n83737 , n83738 );
buf ( n83740 , n83739 );
buf ( n83741 , n83740 );
buf ( n83742 , C1 );
buf ( n83743 , n83742 );
xor ( n83744 , n83741 , n83743 );
xor ( n83745 , n83403 , n83410 );
xor ( n83746 , n83745 , n83412 );
buf ( n83747 , n83746 );
buf ( n83748 , n83747 );
not ( n83749 , n83748 );
buf ( n83750 , C0 );
buf ( n83751 , C1 );
buf ( n83752 , n83751 );
nand ( n83753 , n83749 , n83752 );
buf ( n83754 , n83753 );
buf ( n83755 , n83754 );
xor ( n83756 , n83659 , n83672 );
xor ( n83757 , n83756 , n83703 );
buf ( n83758 , n83757 );
and ( n83759 , n83755 , n83758 );
buf ( n83760 , C0 );
buf ( n83761 , n83760 );
nor ( n83762 , n83759 , n83761 );
buf ( n83763 , n83762 );
buf ( n83764 , n83763 );
and ( n83765 , n83744 , n83764 );
and ( n83766 , n83741 , n83743 );
or ( n83767 , n83765 , n83766 );
buf ( n83768 , n83767 );
buf ( n83769 , n83768 );
or ( n83770 , n83729 , n83769 );
buf ( n83771 , n83770 );
not ( n83772 , n83771 );
xor ( n83773 , n83558 , n83575 );
xor ( n83774 , n83773 , n83630 );
buf ( n83775 , n83774 );
buf ( n83776 , n83775 );
buf ( n83777 , n63022 );
buf ( n83778 , n623 );
nand ( n83779 , n83777 , n83778 );
buf ( n83780 , n83779 );
buf ( n83781 , n83780 );
not ( n83782 , n83781 );
buf ( n83783 , n83584 );
buf ( n83784 , n64227 );
or ( n83785 , n83783 , n83784 );
buf ( n83786 , n64230 );
nand ( n83787 , n83785 , n83786 );
buf ( n83788 , n83787 );
buf ( n83789 , n83788 );
nand ( n83790 , n83782 , n83789 );
buf ( n83791 , n83790 );
buf ( n83792 , n83791 );
not ( n83793 , n83792 );
or ( n83794 , n83793 , C0 );
xor ( n83795 , n83593 , n83607 );
xor ( n83796 , n83795 , n83625 );
buf ( n83797 , n83796 );
buf ( n83798 , n83797 );
nand ( n83799 , n83794 , n83798 );
buf ( n83800 , n83799 );
buf ( n83801 , n83800 );
buf ( n83802 , C1 );
buf ( n83803 , n83802 );
nand ( n83804 , n83801 , n83803 );
buf ( n83805 , n83804 );
buf ( n83806 , n83805 );
xor ( n83807 , n83776 , n83806 );
not ( n83808 , n51464 );
and ( n83809 , n83808 , C1 );
or ( n83810 , C0 , n83809 );
and ( n83811 , n51463 , n83810 );
not ( n83812 , n51463 );
not ( n83813 , n23615 );
and ( n83814 , n83813 , C1 );
or ( n83815 , C0 , n83814 );
and ( n83816 , n83812 , n83815 );
or ( n83817 , n83811 , n83816 );
nor ( n83818 , n83817 , n56325 );
buf ( n83819 , n83818 );
and ( n83820 , n83807 , n83819 );
and ( n83821 , n83776 , n83806 );
or ( n83822 , n83820 , n83821 );
buf ( n83823 , n83822 );
buf ( n83824 , n83823 );
buf ( n83825 , C0 );
buf ( n83826 , n83825 );
xor ( n83827 , n83824 , n83826 );
not ( n83828 , n83634 );
not ( n83829 , n83646 );
or ( n83830 , n83828 , n83829 );
or ( n83831 , n83646 , n83634 );
nand ( n83832 , n83830 , n83831 );
and ( n83833 , n83554 , n83832 );
not ( n83834 , n83554 );
not ( n83835 , n83832 );
and ( n83836 , n83834 , n83835 );
nor ( n83837 , n83833 , n83836 );
buf ( n83838 , n83837 );
and ( n83839 , n83827 , n83838 );
or ( n83840 , n83839 , C0 );
buf ( n83841 , n83840 );
buf ( n83842 , n83841 );
not ( n83843 , n52456 );
not ( n83844 , n83531 );
or ( n83845 , n83843 , n83844 );
and ( n83846 , n56325 , n82745 );
not ( n83847 , n56325 );
and ( n83848 , n83847 , n48836 );
nor ( n83849 , n83846 , n83848 );
nand ( n83850 , n83849 , n51487 );
nand ( n83851 , n83845 , n83850 );
buf ( n83852 , n83851 );
buf ( n83853 , C0 );
buf ( n83854 , n83853 );
buf ( n83855 , n83788 );
not ( n83856 , n83855 );
buf ( n83857 , n83780 );
not ( n83858 , n83857 );
or ( n83859 , n83856 , n83858 );
buf ( n83860 , n83780 );
buf ( n83861 , n83788 );
or ( n83862 , n83860 , n83861 );
nand ( n83863 , n83859 , n83862 );
buf ( n83864 , n83863 );
buf ( n83865 , n83864 );
buf ( n83866 , n63003 );
buf ( n83867 , n64227 );
buf ( n83868 , n75821 );
nor ( n83869 , n83867 , n83868 );
buf ( n83870 , n83869 );
buf ( n83871 , n83870 );
nor ( n83872 , n83866 , n83871 );
buf ( n83873 , n83872 );
buf ( n83874 , n83873 );
buf ( n83875 , n64230 );
buf ( n83876 , n623 );
or ( n83877 , n83875 , n83876 );
buf ( n83878 , n64235 );
nand ( n83879 , n83877 , n83878 );
buf ( n83880 , n83879 );
buf ( n83881 , n83880 );
buf ( n83882 , C0 );
buf ( n83883 , C0 );
buf ( n83884 , n83883 );
and ( n83885 , n83874 , n83881 );
or ( n83886 , C0 , n83885 );
buf ( n83887 , n83886 );
buf ( n83888 , n83887 );
buf ( n83889 , C0 );
buf ( n83890 , n83889 );
and ( n83891 , n83865 , n83888 );
or ( n83892 , C0 , n83891 );
buf ( n83893 , n83892 );
buf ( n83894 , n83893 );
buf ( n83895 , n83791 );
not ( n83896 , n83895 );
buf ( n83897 , n83797 );
not ( n83898 , n83897 );
or ( n83899 , n83896 , n83898 );
buf ( n83900 , n83797 );
buf ( n83901 , n83791 );
or ( n83902 , n83900 , n83901 );
nand ( n83903 , n83899 , n83902 );
buf ( n83904 , n83903 );
buf ( n83905 , n83904 );
not ( n83906 , n83905 );
or ( n83907 , C0 , n83906 );
nand ( n83908 , n83907 , C1 );
buf ( n83909 , n83908 );
buf ( n83910 , n83909 );
buf ( n83911 , C0 );
buf ( n83912 , n83911 );
and ( n83913 , n83894 , n83910 );
or ( n83914 , C0 , n83913 );
buf ( n83915 , n83914 );
buf ( n83916 , n83915 );
xor ( n83917 , n83854 , n83916 );
xor ( n83918 , n83776 , n83806 );
xor ( n83919 , n83918 , n83819 );
buf ( n83920 , n83919 );
buf ( n83921 , n83920 );
and ( n83922 , n83917 , n83921 );
or ( n83923 , n83922 , C0 );
buf ( n83924 , n83923 );
buf ( n83925 , n83924 );
xor ( n83926 , n83852 , n83925 );
xor ( n83927 , n83824 , n83826 );
xor ( n83928 , n83927 , n83838 );
buf ( n83929 , n83928 );
buf ( n83930 , n83929 );
and ( n83931 , n83926 , n83930 );
and ( n83932 , n83852 , n83925 );
or ( n83933 , n83931 , n83932 );
buf ( n83934 , n83933 );
buf ( n83935 , n83934 );
xor ( n83936 , n83842 , n83935 );
buf ( n83937 , n83695 );
not ( n83938 , n83937 );
buf ( n83939 , n83677 );
and ( n83940 , C1 , n83939 );
nor ( n83941 , C0 , n83940 );
buf ( n83942 , n83941 );
buf ( n83943 , n83942 );
not ( n83944 , n83943 );
buf ( n83945 , n83944 );
buf ( n83946 , n83945 );
not ( n83947 , n83946 );
or ( n83948 , n83938 , n83947 );
buf ( n83949 , n83692 );
buf ( n83950 , n83942 );
nand ( n83951 , n83949 , n83950 );
buf ( n83952 , n83951 );
buf ( n83953 , n83952 );
nand ( n83954 , n83948 , n83953 );
buf ( n83955 , n83954 );
buf ( n83956 , n83955 );
and ( n83957 , n83936 , n83956 );
or ( n83958 , n83957 , C0 );
buf ( n83959 , n83958 );
buf ( n83960 , n83959 );
xor ( n83961 , n83894 , n83910 );
xor ( n83962 , n83961 , n83912 );
buf ( n83963 , n83962 );
buf ( n83964 , n83963 );
xor ( n83965 , n83865 , n83888 );
xor ( n83966 , n83965 , n83890 );
buf ( n83967 , n83966 );
buf ( n83968 , n83967 );
buf ( n83969 , C0 );
buf ( n83970 , n83969 );
xor ( n83971 , n83874 , n83881 );
xor ( n83972 , n83971 , n83884 );
buf ( n83973 , n83972 );
buf ( n83974 , n83973 );
buf ( n83975 , C0 );
buf ( n83976 , n83975 );
buf ( n83977 , C0 );
buf ( n83978 , n83977 );
buf ( n83979 , C0 );
buf ( n83980 , n83979 );
buf ( n83981 , C0 );
buf ( n83982 , n83981 );
buf ( n83983 , C0 );
buf ( n83984 , n83983 );
buf ( n83985 , C0 );
xor ( n83986 , n83854 , n83916 );
xor ( n83987 , n83986 , n83921 );
buf ( n83988 , n83987 );
buf ( n83989 , n83988 );
buf ( n83990 , C0 );
buf ( n83991 , n83990 );
nor ( n83992 , n83989 , n83991 );
buf ( n83993 , n83992 );
buf ( n83994 , C1 );
xor ( n83995 , n83852 , n83925 );
xor ( n83996 , n83995 , n83930 );
buf ( n83997 , n83996 );
buf ( n83998 , n83997 );
xor ( n83999 , n83842 , n83935 );
xor ( n84000 , n83999 , n83956 );
buf ( n84001 , n84000 );
buf ( n84002 , n84001 );
buf ( n84003 , C0 );
buf ( n84004 , n84003 );
xor ( n84005 , n83960 , n84004 );
buf ( n84006 , n83750 );
buf ( n84007 , n83747 );
xor ( n84008 , n84006 , n84007 );
buf ( n84009 , n83757 );
xor ( n84010 , n84008 , n84009 );
buf ( n84011 , n84010 );
buf ( n84012 , n84011 );
and ( n84013 , n84005 , n84012 );
or ( n84014 , n84013 , C0 );
buf ( n84015 , n84014 );
not ( n84016 , n84015 );
xor ( n84017 , n83741 , n83743 );
xor ( n84018 , n84017 , n83764 );
buf ( n84019 , n84018 );
buf ( n84020 , n84019 );
buf ( n84021 , n83504 );
not ( n84022 , n84021 );
buf ( n84023 , n83712 );
not ( n84024 , n84023 );
or ( n84025 , n84022 , n84024 );
buf ( n84026 , n83497 );
buf ( n84027 , n83716 );
nand ( n84028 , n84026 , n84027 );
buf ( n84029 , n84028 );
buf ( n84030 , n84029 );
nand ( n84031 , n84025 , n84030 );
buf ( n84032 , n84031 );
xnor ( n84033 , n84032 , n83706 );
buf ( n84034 , n84033 );
nand ( n84035 , n84020 , n84034 );
buf ( n84036 , n84035 );
not ( n84037 , n84036 );
or ( n84038 , n84016 , n84037 );
buf ( n84039 , n84019 );
buf ( n84040 , n84033 );
or ( n84041 , n84039 , n84040 );
buf ( n84042 , n84041 );
nand ( n84043 , n84038 , n84042 );
buf ( n84044 , n84043 );
buf ( n84045 , n83728 );
buf ( n84046 , n83768 );
nand ( n84047 , n84045 , n84046 );
buf ( n84048 , n84047 );
buf ( n84049 , n84048 );
nand ( n84050 , n84044 , n84049 );
buf ( n84051 , n84050 );
not ( n84052 , n84051 );
or ( n84053 , n83772 , n84052 );
buf ( n84054 , n83432 );
buf ( n84055 , n83427 );
xor ( n84056 , n84054 , n84055 );
buf ( n84057 , n83184 );
xor ( n84058 , n84056 , n84057 );
buf ( n84059 , n84058 );
buf ( n84060 , n84059 );
not ( n84061 , n84060 );
buf ( n84062 , n83486 );
buf ( n84063 , n83490 );
or ( n84064 , n84062 , n84063 );
buf ( n84065 , n83722 );
nand ( n84066 , n84064 , n84065 );
buf ( n84067 , n84066 );
buf ( n84068 , n84067 );
buf ( n84069 , C1 );
buf ( n84070 , n84069 );
nand ( n84071 , n84068 , n84070 );
buf ( n84072 , n84071 );
xor ( n84073 , C1 , n84072 );
buf ( n84074 , n84073 );
not ( n84075 , n84074 );
and ( n84076 , n84061 , n84075 );
buf ( n84077 , n84059 );
buf ( n84078 , n84073 );
and ( n84079 , n84077 , n84078 );
nor ( n84080 , n84076 , n84079 );
buf ( n84081 , n84080 );
xor ( n84082 , n83482 , n83484 );
and ( n84083 , n84082 , n83726 );
and ( n84084 , n83482 , n83484 );
or ( n84085 , n84083 , n84084 );
buf ( n84086 , n84085 );
nand ( n84087 , n84081 , n84086 );
nand ( n84088 , n84053 , n84087 );
buf ( n84089 , n84088 );
buf ( n84090 , n84081 );
buf ( n84091 , n84086 );
or ( n84092 , n84090 , n84091 );
buf ( n84093 , n84092 );
buf ( n84094 , n84093 );
nand ( n84095 , n84089 , n84094 );
buf ( n84096 , n84095 );
not ( n84097 , n84096 );
buf ( n84098 , n83462 );
not ( n84099 , n84098 );
buf ( n84100 , n83448 );
not ( n84101 , n84100 );
and ( n84102 , n84099 , n84101 );
buf ( n84103 , n83462 );
buf ( n84104 , n83448 );
and ( n84105 , n84103 , n84104 );
nor ( n84106 , n84102 , n84105 );
buf ( n84107 , n84106 );
buf ( n84108 , n84107 );
not ( n84109 , n84108 );
buf ( n84110 , n83453 );
not ( n84111 , n84110 );
and ( n84112 , n84109 , n84111 );
buf ( n84113 , n84107 );
buf ( n84114 , n83453 );
and ( n84115 , n84113 , n84114 );
nor ( n84116 , n84112 , n84115 );
buf ( n84117 , n84116 );
buf ( n84118 , n84117 );
buf ( n84119 , n84059 );
buf ( n84120 , n84072 );
not ( n84121 , n84120 );
buf ( n84122 , C1 );
nand ( n84123 , n84121 , n84122 );
buf ( n84124 , n84123 );
buf ( n84125 , n84124 );
nand ( n84126 , n84119 , n84125 );
buf ( n84127 , n84126 );
buf ( n84128 , n84127 );
buf ( n84129 , C1 );
buf ( n84130 , n84129 );
and ( n84131 , n84128 , n84130 );
buf ( n84132 , n84131 );
buf ( n84133 , n84132 );
nand ( n84134 , n84118 , n84133 );
buf ( n84135 , n84134 );
not ( n84136 , n84135 );
or ( n84137 , n84097 , n84136 );
buf ( n84138 , n84117 );
not ( n84139 , n84138 );
buf ( n84140 , n84139 );
buf ( n84141 , n84140 );
buf ( n84142 , n84132 );
not ( n84143 , n84142 );
buf ( n84144 , n84143 );
buf ( n84145 , n84144 );
nand ( n84146 , n84141 , n84145 );
buf ( n84147 , n84146 );
nand ( n84148 , n84137 , n84147 );
buf ( n84149 , n84148 );
xor ( n84150 , n83475 , n84149 );
buf ( n84151 , C0 );
buf ( n84152 , n84151 );
xor ( n84153 , n83096 , n83100 );
xor ( n84154 , n84153 , n83102 );
buf ( n84155 , n84154 );
buf ( n84156 , n84155 );
xor ( n84157 , n84152 , n84156 );
xor ( n84158 , n82948 , n83019 );
xor ( n84159 , n84158 , n83048 );
buf ( n84160 , n84159 );
buf ( n84161 , n84160 );
xor ( n84162 , n84157 , n84161 );
buf ( n84163 , n84162 );
buf ( n84164 , n84163 );
and ( n84165 , n84150 , n84164 );
and ( n84166 , n83475 , n84149 );
or ( n84167 , n84165 , n84166 );
buf ( n84168 , n84167 );
buf ( n84169 , n84168 );
not ( n84170 , n84169 );
buf ( n84171 , n84170 );
buf ( n84172 , n84171 );
xor ( n84173 , n83053 , n83089 );
xor ( n84174 , n84173 , n83115 );
buf ( n84175 , n84174 );
buf ( n84176 , n84175 );
xor ( n84177 , n84152 , n84156 );
and ( n84178 , n84177 , n84161 );
or ( n84179 , n84178 , C0 );
buf ( n84180 , n84179 );
buf ( n84181 , n84180 );
nor ( n84182 , n84176 , n84181 );
buf ( n84183 , n84182 );
buf ( n84184 , n84183 );
or ( n84185 , n84172 , n84184 );
buf ( n84186 , n84175 );
buf ( n84187 , n84180 );
nand ( n84188 , n84186 , n84187 );
buf ( n84189 , n84188 );
buf ( n84190 , n84189 );
nand ( n84191 , n84185 , n84190 );
buf ( n84192 , n84191 );
not ( n84193 , n84192 );
or ( n84194 , n83181 , n84193 );
buf ( n84195 , n83177 );
not ( n84196 , n84195 );
buf ( n84197 , n83119 );
nand ( n84198 , n84196 , n84197 );
buf ( n84199 , n84198 );
nand ( n84200 , n84194 , n84199 );
not ( n84201 , n84200 );
buf ( n84202 , n83162 );
not ( n84203 , n84202 );
buf ( n84204 , n83169 );
nand ( n84205 , n84203 , n84204 );
buf ( n84206 , n84205 );
buf ( n84207 , n84206 );
not ( n84208 , n84207 );
buf ( n84209 , n83159 );
not ( n84210 , n84209 );
or ( n84211 , n84208 , n84210 );
buf ( n84212 , n83166 );
buf ( n84213 , n83162 );
nand ( n84214 , n84212 , n84213 );
buf ( n84215 , n84214 );
buf ( n84216 , n84215 );
nand ( n84217 , n84211 , n84216 );
buf ( n84218 , n84217 );
buf ( n84219 , n84218 );
not ( n84220 , n84219 );
and ( n84221 , n83127 , n83154 );
or ( n84222 , C0 , n84221 );
buf ( n84223 , n84222 );
buf ( n84224 , n84223 );
xor ( n84225 , n82458 , n82460 );
xor ( n84226 , n84225 , n82468 );
buf ( n84227 , n84226 );
buf ( n84228 , n84227 );
and ( n84229 , n84224 , n84228 );
not ( n84230 , n84224 );
buf ( n84231 , n84227 );
not ( n84232 , n84231 );
buf ( n84233 , n84232 );
buf ( n84234 , n84233 );
and ( n84235 , n84230 , n84234 );
or ( n84236 , n84229 , n84235 );
buf ( n84237 , n84236 );
buf ( n84238 , n84237 );
not ( n84239 , n84238 );
xor ( n84240 , n82568 , n82572 );
xor ( n84241 , n84240 , n82574 );
buf ( n84242 , n84241 );
buf ( n84243 , n84242 );
not ( n84244 , n84243 );
and ( n84245 , n84239 , n84244 );
buf ( n84246 , n84237 );
buf ( n84247 , n84242 );
and ( n84248 , n84246 , n84247 );
nor ( n84249 , n84245 , n84248 );
buf ( n84250 , n84249 );
buf ( n84251 , n84250 );
nand ( n84252 , n84220 , n84251 );
buf ( n84253 , n84252 );
not ( n84254 , n84253 );
or ( n84255 , n84201 , n84254 );
buf ( n84256 , n84250 );
not ( n84257 , n84256 );
buf ( n84258 , n84218 );
nand ( n84259 , n84257 , n84258 );
buf ( n84260 , n84259 );
nand ( n84261 , n84255 , n84260 );
buf ( n84262 , n84227 );
not ( n84263 , n84262 );
buf ( n84264 , n84223 );
not ( n84265 , n84264 );
or ( n84266 , n84263 , n84265 );
buf ( n84267 , n84242 );
buf ( n84268 , n84223 );
not ( n84269 , n84268 );
buf ( n84270 , n84233 );
nand ( n84271 , n84269 , n84270 );
buf ( n84272 , n84271 );
buf ( n84273 , n84272 );
nand ( n84274 , n84267 , n84273 );
buf ( n84275 , n84274 );
buf ( n84276 , n84275 );
nand ( n84277 , n84266 , n84276 );
buf ( n84278 , n84277 );
not ( n84279 , n84278 );
xor ( n84280 , n82578 , n82582 );
xor ( n84281 , n84280 , n82587 );
buf ( n84282 , n84281 );
not ( n84283 , n84282 );
nand ( n84284 , n84279 , n84283 );
and ( n84285 , n84261 , n84284 );
and ( n84286 , n84282 , n84278 );
nor ( n84287 , n84285 , n84286 );
or ( n84288 , n82594 , n84287 );
buf ( n84289 , n82505 );
buf ( n84290 , n82591 );
nand ( n84291 , n84289 , n84290 );
buf ( n84292 , n84291 );
nand ( n84293 , n84288 , n84292 );
not ( n84294 , n84293 );
or ( n84295 , n82503 , n84294 );
buf ( n84296 , n82500 );
buf ( n84297 , n82494 );
or ( n84298 , n84296 , n84297 );
buf ( n84299 , n84298 );
nand ( n84300 , n84295 , n84299 );
not ( n84301 , n84300 );
or ( n84302 , n82435 , n84301 );
buf ( n84303 , n82431 );
not ( n84304 , n84303 );
buf ( n84305 , n82417 );
nand ( n84306 , n84304 , n84305 );
buf ( n84307 , n84306 );
nand ( n84308 , n84302 , n84307 );
buf ( n84309 , n84308 );
and ( n84310 , n81991 , n84309 );
and ( n84311 , n81986 , n81990 );
or ( n84312 , n84310 , n84311 );
buf ( n84313 , n84312 );
buf ( n84314 , n84313 );
and ( n84315 , n81562 , n84314 );
and ( n84316 , n81557 , n81561 );
or ( n84317 , n84315 , n84316 );
buf ( n84318 , n84317 );
buf ( n84319 , n84318 );
and ( n84320 , n81439 , n84319 );
and ( n84321 , n81434 , n81438 );
or ( n84322 , n84320 , n84321 );
buf ( n84323 , n84322 );
buf ( n84324 , n84323 );
and ( n84325 , n81121 , n84324 );
and ( n84326 , n81116 , n81120 );
or ( n84327 , n84325 , n84326 );
buf ( n84328 , n84327 );
buf ( n84329 , n84328 );
and ( n84330 , n80957 , n84329 );
and ( n84331 , n80953 , n80956 );
or ( n84332 , n84330 , n84331 );
buf ( n84333 , n84332 );
not ( n84334 , n84333 );
or ( n84335 , n80734 , n84334 );
not ( n84336 , n80732 );
nand ( n84337 , n84336 , n80717 );
nand ( n84338 , n84335 , n84337 );
nand ( n84339 , n80154 , n84338 , n80146 );
or ( n84340 , n80140 , n80145 );
nand ( n84341 , n80147 , n84339 , n84340 );
xor ( n84342 , n75105 , n75120 );
xor ( n84343 , n84342 , n75427 );
buf ( n84344 , n84343 );
buf ( n84345 , n84344 );
xor ( n84346 , n80106 , n80110 );
and ( n84347 , n84346 , n80128 );
and ( n84348 , n80106 , n80110 );
or ( n84349 , n84347 , n84348 );
buf ( n84350 , n84349 );
buf ( n84351 , n84350 );
xor ( n84352 , n84345 , n84351 );
xor ( n84353 , n76388 , n76392 );
buf ( n84354 , n84353 );
buf ( n84355 , n84354 );
buf ( n84356 , n76379 );
and ( n84357 , n84355 , n84356 );
not ( n84358 , n84355 );
buf ( n84359 , n76379 );
not ( n84360 , n84359 );
buf ( n84361 , n84360 );
buf ( n84362 , n84361 );
and ( n84363 , n84358 , n84362 );
nor ( n84364 , n84357 , n84363 );
buf ( n84365 , n84364 );
buf ( n84366 , n84365 );
xor ( n84367 , n84352 , n84366 );
buf ( n84368 , n84367 );
buf ( n84369 , n84368 );
buf ( n84370 , n80097 );
not ( n84371 , n84370 );
buf ( n84372 , n80133 );
not ( n84373 , n84372 );
or ( n84374 , n84371 , n84373 );
buf ( n84375 , n80091 );
nand ( n84376 , n84374 , n84375 );
buf ( n84377 , n84376 );
buf ( n84378 , n84377 );
buf ( n84379 , n80130 );
buf ( n84380 , n80094 );
nand ( n84381 , n84379 , n84380 );
buf ( n84382 , n84381 );
buf ( n84383 , n84382 );
nand ( n84384 , n84378 , n84383 );
buf ( n84385 , n84384 );
buf ( n84386 , n84385 );
nor ( n84387 , n84369 , n84386 );
buf ( n84388 , n84387 );
not ( n84389 , n84388 );
nand ( n84390 , n84341 , n84389 );
buf ( n84391 , n84390 );
xor ( n84392 , n84345 , n84351 );
and ( n84393 , n84392 , n84366 );
and ( n84394 , n84345 , n84351 );
or ( n84395 , n84393 , n84394 );
buf ( n84396 , n84395 );
buf ( n84397 , n84396 );
not ( n84398 , n84397 );
buf ( n84399 , n76397 );
not ( n84400 , n84399 );
buf ( n84401 , n74639 );
not ( n84402 , n84401 );
or ( n84403 , n84400 , n84402 );
buf ( n84404 , n74639 );
buf ( n84405 , n76397 );
or ( n84406 , n84404 , n84405 );
nand ( n84407 , n84403 , n84406 );
buf ( n84408 , n84407 );
xor ( n84409 , n75441 , n84408 );
buf ( n84410 , n84409 );
nand ( n84411 , n84398 , n84410 );
buf ( n84412 , n84411 );
buf ( n84413 , n84412 );
not ( n84414 , n84413 );
buf ( n84415 , n84414 );
buf ( n84416 , n84415 );
or ( n84417 , n84391 , n84416 );
buf ( n84418 , n84412 );
nand ( n84419 , n84368 , n84385 );
not ( n84420 , n84419 );
buf ( n84421 , n84420 );
and ( n84422 , n84418 , n84421 );
not ( n84423 , n84396 );
nor ( n84424 , n84423 , n84409 );
buf ( n84425 , n84424 );
nor ( n84426 , n84422 , n84425 );
buf ( n84427 , n84426 );
buf ( n84428 , n84427 );
nand ( n84429 , n84417 , n84428 );
buf ( n84430 , n84429 );
buf ( n84431 , n84430 );
and ( n84432 , n76906 , n84431 );
and ( n84433 , n76413 , n76905 );
or ( n84434 , n84432 , n84433 );
buf ( n84435 , n84434 );
buf ( n84436 , n84435 );
not ( n84437 , n84436 );
xor ( n84438 , n76663 , n76664 );
and ( n84439 , n84438 , n76671 );
or ( n84440 , n84439 , C0 );
buf ( n84441 , n84440 );
buf ( n84442 , n84441 );
buf ( n84443 , n76729 );
not ( n84444 , n84443 );
buf ( n84445 , n47050 );
not ( n84446 , n84445 );
or ( n84447 , n84444 , n84446 );
buf ( n84448 , n52780 );
buf ( n84449 , n42468 );
and ( n84450 , n84448 , n84449 );
not ( n84451 , n84448 );
buf ( n84452 , n47031 );
and ( n84453 , n84451 , n84452 );
nor ( n84454 , n84450 , n84453 );
buf ( n84455 , n84454 );
buf ( n84456 , n84455 );
buf ( n84457 , n52595 );
nand ( n84458 , n84456 , n84457 );
buf ( n84459 , n84458 );
buf ( n84460 , n84459 );
nand ( n84461 , n84447 , n84460 );
buf ( n84462 , n84461 );
buf ( n84463 , n84462 );
buf ( n84464 , n46912 );
not ( n84465 , n84464 );
buf ( n84466 , n46875 );
not ( n84467 , n84466 );
buf ( n84468 , n41915 );
not ( n84469 , n84468 );
or ( n84470 , n84467 , n84469 );
buf ( n84471 , n41912 );
buf ( n84472 , n46887 );
nand ( n84473 , n84471 , n84472 );
buf ( n84474 , n84473 );
buf ( n84475 , n84474 );
nand ( n84476 , n84470 , n84475 );
buf ( n84477 , n84476 );
buf ( n84478 , n84477 );
not ( n84479 , n84478 );
or ( n84480 , n84465 , n84479 );
buf ( n84481 , n76881 );
buf ( n84482 , n46907 );
nand ( n84483 , n84481 , n84482 );
buf ( n84484 , n84483 );
buf ( n84485 , n84484 );
nand ( n84486 , n84480 , n84485 );
buf ( n84487 , n84486 );
buf ( n84488 , n84487 );
xor ( n84489 , n84463 , n84488 );
xor ( n84490 , n76752 , n76809 );
and ( n84491 , n84490 , n76816 );
and ( n84492 , n76752 , n76809 );
or ( n84493 , n84491 , n84492 );
buf ( n84494 , n84493 );
buf ( n84495 , n84494 );
xor ( n84496 , n84489 , n84495 );
buf ( n84497 , n84496 );
buf ( n84498 , n84497 );
xor ( n84499 , n76737 , n76819 );
and ( n84500 , n84499 , n76837 );
and ( n84501 , n76737 , n76819 );
or ( n84502 , n84500 , n84501 );
buf ( n84503 , n84502 );
buf ( n84504 , n84503 );
buf ( n84505 , C1 );
buf ( n84506 , n84505 );
and ( n84507 , n84504 , n84506 );
nor ( n84508 , n84507 , C0 );
buf ( n84509 , n84508 );
buf ( n84510 , n84509 );
xor ( n84511 , n84498 , n84510 );
buf ( n84512 , n84511 );
buf ( n84513 , n84512 );
not ( n84514 , n84513 );
buf ( n84515 , n84514 );
buf ( n84516 , n84515 );
or ( n84517 , n84442 , n84516 );
xor ( n84518 , n76840 , n76844 );
and ( n84519 , n84518 , n76896 );
and ( n84520 , n76840 , n76844 );
or ( n84521 , n84519 , n84520 );
buf ( n84522 , n84521 );
buf ( n84523 , n84522 );
nand ( n84524 , n84517 , n84523 );
buf ( n84525 , n84524 );
buf ( n84526 , n84525 );
buf ( n84527 , n84441 );
buf ( n84528 , n84515 );
nand ( n84529 , n84527 , n84528 );
buf ( n84530 , n84529 );
buf ( n84531 , n84530 );
and ( n84532 , n84526 , n84531 );
buf ( n84533 , n84532 );
buf ( n84534 , n84533 );
xor ( n84535 , n76481 , n76483 );
and ( n84536 , n84535 , n76501 );
or ( n84537 , n84536 , C0 );
buf ( n84538 , n84537 );
not ( n84539 , n76856 );
not ( n84540 , n84539 );
not ( n84541 , n76865 );
or ( n84542 , n84540 , n84541 );
not ( n84543 , n76856 );
not ( n84544 , n76865 );
not ( n84545 , n84544 );
or ( n84546 , n84543 , n84545 );
nand ( n84547 , n84546 , n76887 );
nand ( n84548 , n84542 , n84547 );
buf ( n84549 , n67149 );
not ( n84550 , n84549 );
buf ( n84551 , n53492 );
not ( n84552 , n84551 );
buf ( n84553 , n46657 );
not ( n84554 , n84553 );
or ( n84555 , n84552 , n84554 );
buf ( n84556 , n28411 );
buf ( n84557 , n45747 );
nand ( n84558 , n84556 , n84557 );
buf ( n84559 , n84558 );
buf ( n84560 , n84559 );
nand ( n84561 , n84555 , n84560 );
buf ( n84562 , n84561 );
buf ( n84563 , n84562 );
not ( n84564 , n84563 );
or ( n84565 , n84550 , n84564 );
buf ( n84566 , n76427 );
buf ( n84567 , n46225 );
nand ( n84568 , n84566 , n84567 );
buf ( n84569 , n84568 );
buf ( n84570 , n84569 );
nand ( n84571 , n84565 , n84570 );
buf ( n84572 , n84571 );
not ( n84573 , n84572 );
not ( n84574 , n84573 );
not ( n84575 , n76549 );
not ( n84576 , n76565 );
or ( n84577 , n84575 , n84576 );
buf ( n84578 , n76549 );
buf ( n84579 , n76565 );
nor ( n84580 , n84578 , n84579 );
buf ( n84581 , n84580 );
or ( n84582 , n84581 , n76626 );
nand ( n84583 , n84577 , n84582 );
not ( n84584 , n84583 );
buf ( n84585 , n76455 );
not ( n84586 , n84585 );
buf ( n84587 , n50128 );
not ( n84588 , n84587 );
or ( n84589 , n84586 , n84588 );
buf ( n84590 , n48323 );
not ( n84591 , n84590 );
buf ( n84592 , n51804 );
not ( n84593 , n84592 );
or ( n84594 , n84591 , n84593 );
buf ( n84595 , n52673 );
buf ( n84596 , n48320 );
nand ( n84597 , n84595 , n84596 );
buf ( n84598 , n84597 );
buf ( n84599 , n84598 );
nand ( n84600 , n84594 , n84599 );
buf ( n84601 , n84600 );
buf ( n84602 , n84601 );
buf ( n84603 , n47872 );
nand ( n84604 , n84602 , n84603 );
buf ( n84605 , n84604 );
buf ( n84606 , n84605 );
nand ( n84607 , n84589 , n84606 );
buf ( n84608 , n84607 );
not ( n84609 , n84608 );
not ( n84610 , n84609 );
or ( n84611 , n84584 , n84610 );
not ( n84612 , n84583 );
nand ( n84613 , n84608 , n84612 );
nand ( n84614 , n84611 , n84613 );
not ( n84615 , n84614 );
or ( n84616 , n84574 , n84615 );
or ( n84617 , n84614 , n84573 );
nand ( n84618 , n84616 , n84617 );
and ( n84619 , n84548 , n84618 );
not ( n84620 , n84548 );
not ( n84621 , n84618 );
and ( n84622 , n84620 , n84621 );
nor ( n84623 , n84619 , n84622 );
xor ( n84624 , n76628 , n76653 );
and ( n84625 , n84624 , n76660 );
and ( n84626 , n76628 , n76653 );
or ( n84627 , n84625 , n84626 );
buf ( n84628 , n84627 );
and ( n84629 , n84623 , n84628 );
not ( n84630 , n84623 );
buf ( n84631 , n84628 );
not ( n84632 , n84631 );
buf ( n84633 , n84632 );
and ( n84634 , n84630 , n84633 );
nor ( n84635 , n84629 , n84634 );
xnor ( n84636 , n84538 , n84635 );
buf ( n84637 , n84636 );
xor ( n84638 , n76438 , n76463 );
and ( n84639 , n84638 , n76478 );
and ( n84640 , n76438 , n76463 );
or ( n84641 , n84639 , n84640 );
buf ( n84642 , n84641 );
buf ( n84643 , n84642 );
buf ( n84644 , n48836 );
not ( n84645 , n84644 );
buf ( n84646 , n43777 );
not ( n84647 , n84646 );
or ( n84648 , n84645 , n84647 );
buf ( n84649 , n42398 );
buf ( n84650 , n61847 );
nand ( n84651 , n84649 , n84650 );
buf ( n84652 , n84651 );
buf ( n84653 , n84652 );
nand ( n84654 , n84648 , n84653 );
buf ( n84655 , n84654 );
buf ( n84656 , n84655 );
buf ( n84657 , n62125 );
and ( n84658 , n84656 , n84657 );
buf ( n84659 , n76831 );
buf ( n84660 , n51489 );
nor ( n84661 , n84659 , n84660 );
buf ( n84662 , n84661 );
buf ( n84663 , n84662 );
nor ( n84664 , n84658 , n84663 );
buf ( n84665 , n84664 );
buf ( n84666 , n84665 );
not ( n84667 , n84666 );
buf ( n84668 , n84667 );
buf ( n84669 , n84668 );
xor ( n84670 , n84643 , n84669 );
not ( n84671 , n76473 );
not ( n84672 , n50608 );
or ( n84673 , n84671 , n84672 );
buf ( n84674 , n50995 );
not ( n84675 , n84674 );
buf ( n84676 , n50599 );
not ( n84677 , n84676 );
or ( n84678 , n84675 , n84677 );
buf ( n84679 , n50598 );
buf ( n84680 , n50998 );
nand ( n84681 , n84679 , n84680 );
buf ( n84682 , n84681 );
buf ( n84683 , n84682 );
nand ( n84684 , n84678 , n84683 );
buf ( n84685 , n84684 );
buf ( n84686 , n84685 );
not ( n84687 , n84686 );
buf ( n84688 , n84687 );
or ( n84689 , n84688 , n39980 );
nand ( n84690 , n84673 , n84689 );
buf ( n84691 , n38979 );
buf ( n84692 , n46615 );
not ( n84693 , n84692 );
buf ( n84694 , n84693 );
buf ( n84695 , n84694 );
nor ( n84696 , n84691 , n84695 );
buf ( n84697 , n84696 );
not ( n84698 , n84697 );
not ( n84699 , n56325 );
and ( n84700 , n84698 , n84699 );
not ( n84701 , n84694 );
not ( n84702 , n42468 );
or ( n84703 , n84701 , n84702 );
nand ( n84704 , n84703 , n42411 );
nor ( n84705 , n84700 , n84704 );
not ( n84706 , n76623 );
buf ( n84707 , n76584 );
buf ( n84708 , n76571 );
or ( n84709 , n84707 , n84708 );
buf ( n84710 , n84709 );
not ( n84711 , n84710 );
or ( n84712 , n84706 , n84711 );
buf ( n84713 , n76584 );
buf ( n84714 , n76571 );
nand ( n84715 , n84713 , n84714 );
buf ( n84716 , n84715 );
nand ( n84717 , n84712 , n84716 );
buf ( n84718 , n84717 );
xor ( n84719 , n70845 , n70873 );
xor ( n84720 , n84719 , n70899 );
buf ( n84721 , n84720 );
buf ( n84722 , n84721 );
xor ( n84723 , n84718 , n84722 );
buf ( n84724 , n76542 );
not ( n84725 , n84724 );
buf ( n84726 , n43935 );
not ( n84727 , n84726 );
or ( n84728 , n84725 , n84727 );
buf ( n84729 , n46390 );
not ( n84730 , n84729 );
buf ( n84731 , n25181 );
not ( n84732 , n84731 );
or ( n84733 , n84730 , n84732 );
buf ( n84734 , n54068 );
buf ( n84735 , n46393 );
nand ( n84736 , n84734 , n84735 );
buf ( n84737 , n84736 );
buf ( n84738 , n84737 );
nand ( n84739 , n84733 , n84738 );
buf ( n84740 , n84739 );
buf ( n84741 , n84740 );
buf ( n84742 , n43905 );
nand ( n84743 , n84741 , n84742 );
buf ( n84744 , n84743 );
buf ( n84745 , n84744 );
nand ( n84746 , n84728 , n84745 );
buf ( n84747 , n84746 );
buf ( n84748 , n84747 );
xor ( n84749 , n84723 , n84748 );
buf ( n84750 , n84749 );
nand ( n84751 , n84705 , n84750 );
and ( n84752 , n84690 , n84751 );
not ( n84753 , n84690 );
not ( n84754 , n84750 );
nand ( n84755 , n84705 , n84754 );
and ( n84756 , n84753 , n84755 );
or ( n84757 , n84752 , n84756 );
not ( n84758 , n84705 );
nand ( n84759 , n84758 , n84754 );
and ( n84760 , n84690 , n84759 );
not ( n84761 , n84690 );
not ( n84762 , n84705 );
nand ( n84763 , n84762 , n84750 );
and ( n84764 , n84761 , n84763 );
or ( n84765 , n84760 , n84764 );
nand ( n84766 , n84757 , n84765 );
buf ( n84767 , n84766 );
xnor ( n84768 , n84670 , n84767 );
buf ( n84769 , n84768 );
buf ( n84770 , n84769 );
and ( n84771 , n84637 , n84770 );
not ( n84772 , n84637 );
buf ( n84773 , n84769 );
not ( n84774 , n84773 );
buf ( n84775 , n84774 );
buf ( n84776 , n84775 );
and ( n84777 , n84772 , n84776 );
nor ( n84778 , n84771 , n84777 );
buf ( n84779 , n84778 );
not ( n84780 , n84779 );
buf ( n84781 , n12481 );
buf ( n84782 , n46623 );
and ( n84783 , n84781 , n84782 );
not ( n84784 , n84781 );
buf ( n84785 , n38412 );
and ( n84786 , n84784 , n84785 );
nor ( n84787 , n84783 , n84786 );
buf ( n84788 , n84787 );
not ( n84789 , n84788 );
not ( n84790 , n46620 );
or ( n84791 , n84789 , n84790 );
buf ( n84792 , n55841 );
not ( n84793 , n84792 );
buf ( n84794 , n45069 );
not ( n84795 , n84794 );
or ( n84796 , n84793 , n84795 );
buf ( n84797 , n46623 );
buf ( n84798 , n55840 );
nand ( n84799 , n84797 , n84798 );
buf ( n84800 , n84799 );
buf ( n84801 , n84800 );
nand ( n84802 , n84796 , n84801 );
buf ( n84803 , n84802 );
buf ( n84804 , n84803 );
buf ( n84805 , n38380 );
nand ( n84806 , n84804 , n84805 );
buf ( n84807 , n84806 );
nand ( n84808 , n84791 , n84807 );
buf ( n84809 , n84808 );
buf ( n84810 , n44496 );
not ( n84811 , n84810 );
buf ( n84812 , n65010 );
not ( n84813 , n84812 );
buf ( n84814 , n56342 );
not ( n84815 , n84814 );
or ( n84816 , n84813 , n84815 );
buf ( n84817 , n48172 );
buf ( n84818 , n44530 );
nand ( n84819 , n84817 , n84818 );
buf ( n84820 , n84819 );
buf ( n84821 , n84820 );
nand ( n84822 , n84816 , n84821 );
buf ( n84823 , n84822 );
buf ( n84824 , n84823 );
not ( n84825 , n84824 );
or ( n84826 , n84811 , n84825 );
buf ( n84827 , n76555 );
buf ( n84828 , n44517 );
nand ( n84829 , n84827 , n84828 );
buf ( n84830 , n84829 );
buf ( n84831 , n84830 );
nand ( n84832 , n84826 , n84831 );
buf ( n84833 , n84832 );
buf ( n84834 , n84833 );
xor ( n84835 , n76778 , n76799 );
and ( n84836 , n84835 , n76806 );
and ( n84837 , n76778 , n76799 );
or ( n84838 , n84836 , n84837 );
buf ( n84839 , n84838 );
buf ( n84840 , n84839 );
xor ( n84841 , n84834 , n84840 );
xor ( n84842 , n76597 , n76609 );
and ( n84843 , n84842 , n76622 );
and ( n84844 , n76597 , n76609 );
or ( n84845 , n84843 , n84844 );
buf ( n84846 , n84845 );
buf ( n84847 , n76791 );
not ( n84848 , n84847 );
buf ( n84849 , n59928 );
not ( n84850 , n84849 );
or ( n84851 , n84848 , n84850 );
nand ( n84852 , n70769 , n62582 );
buf ( n84853 , n84852 );
nand ( n84854 , n84851 , n84853 );
buf ( n84855 , n84854 );
buf ( n84856 , n84855 );
xor ( n84857 , n84846 , n84856 );
buf ( n84858 , n43868 );
not ( n84859 , n84858 );
buf ( n84860 , n70823 );
not ( n84861 , n84860 );
or ( n84862 , n84859 , n84861 );
buf ( n84863 , n76766 );
buf ( n84864 , n41596 );
nand ( n84865 , n84863 , n84864 );
buf ( n84866 , n84865 );
buf ( n84867 , n84866 );
nand ( n84868 , n84862 , n84867 );
buf ( n84869 , n84868 );
buf ( n84870 , n84869 );
xor ( n84871 , n84857 , n84870 );
buf ( n84872 , n84871 );
buf ( n84873 , n84872 );
xor ( n84874 , n84841 , n84873 );
buf ( n84875 , n84874 );
buf ( n84876 , n84875 );
xor ( n84877 , n84809 , n84876 );
buf ( n84878 , n48868 );
not ( n84879 , n84878 );
buf ( n84880 , n48808 );
not ( n84881 , n84880 );
buf ( n84882 , n44025 );
not ( n84883 , n84882 );
or ( n84884 , n84881 , n84883 );
buf ( n84885 , n28305 );
buf ( n84886 , n72891 );
nand ( n84887 , n84885 , n84886 );
buf ( n84888 , n84887 );
buf ( n84889 , n84888 );
nand ( n84890 , n84884 , n84889 );
buf ( n84891 , n84890 );
buf ( n84892 , n84891 );
not ( n84893 , n84892 );
or ( n84894 , n84879 , n84893 );
buf ( n84895 , n76645 );
buf ( n84896 , n48855 );
nand ( n84897 , n84895 , n84896 );
buf ( n84898 , n84897 );
buf ( n84899 , n84898 );
nand ( n84900 , n84894 , n84899 );
buf ( n84901 , n84900 );
buf ( n84902 , n84901 );
not ( n84903 , n84902 );
buf ( n84904 , n84903 );
buf ( n84905 , n84904 );
xor ( n84906 , n84877 , n84905 );
buf ( n84907 , n84906 );
buf ( n84908 , n84907 );
not ( n84909 , n84908 );
buf ( n84910 , n84909 );
not ( n84911 , n84910 );
or ( n84912 , C0 , n84911 );
buf ( n84913 , C1 );
nand ( n84914 , n84912 , n84913 );
buf ( n84915 , n76852 );
not ( n84916 , n84915 );
buf ( n84917 , n76888 );
not ( n84918 , n84917 );
buf ( n84919 , n84918 );
buf ( n84920 , n84919 );
not ( n84921 , n84920 );
or ( n84922 , n84916 , n84921 );
buf ( n84923 , n76855 );
not ( n84924 , n84923 );
buf ( n84925 , n76888 );
not ( n84926 , n84925 );
or ( n84927 , n84924 , n84926 );
buf ( n84928 , n76894 );
nand ( n84929 , n84927 , n84928 );
buf ( n84930 , n84929 );
buf ( n84931 , n84930 );
nand ( n84932 , n84922 , n84931 );
buf ( n84933 , n84932 );
buf ( n84934 , n84933 );
not ( n84935 , n84934 );
and ( n84936 , n84914 , n84935 );
not ( n84937 , n84914 );
and ( n84938 , n84937 , n84934 );
nor ( n84939 , n84936 , n84938 );
not ( n84940 , n84939 );
or ( n84941 , n84780 , n84940 );
buf ( n84942 , n76503 );
not ( n84943 , n84942 );
buf ( n84944 , n76520 );
nand ( n84945 , n84943 , n84944 );
buf ( n84946 , n84945 );
buf ( n84947 , n84946 );
not ( n84948 , n84947 );
buf ( n84949 , n76673 );
not ( n84950 , n84949 );
or ( n84951 , n84948 , n84950 );
buf ( n84952 , n76523 );
buf ( n84953 , n76503 );
nand ( n84954 , n84952 , n84953 );
buf ( n84955 , n84954 );
buf ( n84956 , n84955 );
nand ( n84957 , n84951 , n84956 );
buf ( n84958 , n84957 );
nand ( n84959 , n84941 , n84958 );
buf ( n84960 , n84959 );
not ( n84961 , n84939 );
buf ( n84962 , n84779 );
not ( n84963 , n84962 );
buf ( n84964 , n84963 );
nand ( n84965 , n84961 , n84964 );
buf ( n84966 , n84965 );
and ( n84967 , n84960 , n84966 );
buf ( n84968 , n84967 );
buf ( n84969 , n84968 );
xor ( n84970 , n84534 , n84969 );
not ( n84971 , n84769 );
not ( n84972 , n84635 );
and ( n84973 , n84971 , n84972 );
buf ( n84974 , n84769 );
buf ( n84975 , n84635 );
nand ( n84976 , n84974 , n84975 );
buf ( n84977 , n84976 );
and ( n84978 , n84977 , n84538 );
nor ( n84979 , n84973 , n84978 );
buf ( n84980 , n84628 );
not ( n84981 , n84980 );
buf ( n84982 , n84618 );
not ( n84983 , n84982 );
buf ( n84984 , n84548 );
nand ( n84985 , n84983 , n84984 );
buf ( n84986 , n84985 );
buf ( n84987 , n84986 );
not ( n84988 , n84987 );
or ( n84989 , n84981 , n84988 );
buf ( n84990 , n84548 );
not ( n84991 , n84990 );
buf ( n84992 , n84618 );
nand ( n84993 , n84991 , n84992 );
buf ( n84994 , n84993 );
buf ( n84995 , n84994 );
nand ( n84996 , n84989 , n84995 );
buf ( n84997 , n84996 );
buf ( n84998 , n84997 );
buf ( n84999 , n84497 );
not ( n85000 , n84999 );
buf ( n85001 , n85000 );
buf ( n85002 , n85001 );
not ( n85003 , n85002 );
or ( n85004 , n85003 , C0 );
buf ( n85005 , n84503 );
nand ( n85006 , n85004 , n85005 );
buf ( n85007 , n85006 );
buf ( n85008 , n85007 );
buf ( n85009 , C1 );
buf ( n85010 , n85009 );
nand ( n85011 , n85008 , n85010 );
buf ( n85012 , n85011 );
buf ( n85013 , n85012 );
xor ( n85014 , n84998 , n85013 );
buf ( n85015 , n84907 );
not ( n85016 , n85015 );
or ( n85017 , C0 , n85016 );
buf ( n85018 , n84933 );
nand ( n85019 , n85017 , n85018 );
buf ( n85020 , n85019 );
buf ( n85021 , n85020 );
buf ( n85022 , C1 );
buf ( n85023 , n85022 );
nand ( n85024 , n85021 , n85023 );
buf ( n85025 , n85024 );
buf ( n85026 , n85025 );
xor ( n85027 , n85014 , n85026 );
buf ( n85028 , n85027 );
xor ( n85029 , n84979 , n85028 );
xor ( n85030 , n84463 , n84488 );
and ( n85031 , n85030 , n84495 );
and ( n85032 , n84463 , n84488 );
or ( n85033 , n85031 , n85032 );
buf ( n85034 , n85033 );
buf ( n85035 , n85034 );
buf ( n85036 , n46912 );
not ( n85037 , n85036 );
buf ( n85038 , n46875 );
not ( n85039 , n85038 );
buf ( n85040 , n51250 );
not ( n85041 , n85040 );
or ( n85042 , n85039 , n85041 );
buf ( n85043 , n41822 );
buf ( n85044 , n46887 );
nand ( n85045 , n85043 , n85044 );
buf ( n85046 , n85045 );
buf ( n85047 , n85046 );
nand ( n85048 , n85042 , n85047 );
buf ( n85049 , n85048 );
buf ( n85050 , n85049 );
not ( n85051 , n85050 );
or ( n85052 , n85037 , n85051 );
buf ( n85053 , n84477 );
buf ( n85054 , n46907 );
nand ( n85055 , n85053 , n85054 );
buf ( n85056 , n85055 );
buf ( n85057 , n85056 );
nand ( n85058 , n85052 , n85057 );
buf ( n85059 , n85058 );
not ( n85060 , n85059 );
buf ( n85061 , n84455 );
not ( n85062 , n85061 );
buf ( n85063 , n44221 );
not ( n85064 , n85063 );
or ( n85065 , n85062 , n85064 );
buf ( n85066 , n56289 );
buf ( n85067 , n38994 );
and ( n85068 , n85066 , n85067 );
not ( n85069 , n85066 );
buf ( n85070 , n38979 );
and ( n85071 , n85069 , n85070 );
nor ( n85072 , n85068 , n85071 );
buf ( n85073 , n85072 );
buf ( n85074 , n85073 );
not ( n85075 , n85074 );
buf ( n85076 , n42448 );
nand ( n85077 , n85075 , n85076 );
buf ( n85078 , n85077 );
buf ( n85079 , n85078 );
nand ( n85080 , n85065 , n85079 );
buf ( n85081 , n85080 );
not ( n85082 , n85081 );
not ( n85083 , n85082 );
or ( n85084 , n85060 , n85083 );
not ( n85085 , n85059 );
nand ( n85086 , n85085 , n85081 );
nand ( n85087 , n85084 , n85086 );
buf ( n85088 , n44039 );
buf ( n85089 , n84803 );
not ( n85090 , n85089 );
buf ( n85091 , n85090 );
buf ( n85092 , n85091 );
or ( n85093 , n85088 , n85092 );
buf ( n85094 , n53539 );
buf ( n85095 , n42403 );
and ( n85096 , n85094 , n85095 );
not ( n85097 , n85094 );
buf ( n85098 , n47068 );
and ( n85099 , n85097 , n85098 );
nor ( n85100 , n85096 , n85099 );
buf ( n85101 , n85100 );
buf ( n85102 , n85101 );
buf ( n85103 , n52171 );
or ( n85104 , n85102 , n85103 );
nand ( n85105 , n85093 , n85104 );
buf ( n85106 , n85105 );
buf ( n85107 , n85106 );
and ( n85108 , n85087 , n85107 );
not ( n85109 , n85087 );
not ( n85110 , n85107 );
and ( n85111 , n85109 , n85110 );
nor ( n85112 , n85108 , n85111 );
buf ( n85113 , n85112 );
xor ( n85114 , n85035 , n85113 );
buf ( n85115 , C0 );
buf ( n85116 , n85115 );
xor ( n85117 , n85114 , n85116 );
buf ( n85118 , n85117 );
buf ( n85119 , n85118 );
not ( n85120 , n37410 );
nor ( n85121 , n85120 , n56325 );
xor ( n85122 , n84834 , n84840 );
and ( n85123 , n85122 , n84873 );
and ( n85124 , n84834 , n84840 );
or ( n85125 , n85123 , n85124 );
buf ( n85126 , n85125 );
xor ( n85127 , n85121 , n85126 );
buf ( n85128 , n84740 );
not ( n85129 , n85128 );
buf ( n85130 , n43935 );
not ( n85131 , n85130 );
or ( n85132 , n85129 , n85131 );
buf ( n85133 , n69726 );
buf ( n85134 , n53649 );
nand ( n85135 , n85133 , n85134 );
buf ( n85136 , n85135 );
buf ( n85137 , n85136 );
nand ( n85138 , n85132 , n85137 );
buf ( n85139 , n85138 );
buf ( n85140 , n85139 );
xor ( n85141 , n70743 , n70760 );
xor ( n85142 , n85141 , n70779 );
buf ( n85143 , n85142 );
buf ( n85144 , n85143 );
xor ( n85145 , n85140 , n85144 );
xor ( n85146 , n84846 , n84856 );
and ( n85147 , n85146 , n84870 );
and ( n85148 , n84846 , n84856 );
or ( n85149 , n85147 , n85148 );
buf ( n85150 , n85149 );
buf ( n85151 , n85150 );
xor ( n85152 , n85145 , n85151 );
buf ( n85153 , n85152 );
xor ( n85154 , n85127 , n85153 );
buf ( n85155 , n85154 );
buf ( n85156 , C0 );
buf ( n85157 , n85156 );
xor ( n85158 , n85155 , n85157 );
buf ( n85159 , n84808 );
not ( n85160 , n85159 );
buf ( n85161 , n84901 );
not ( n85162 , n85161 );
or ( n85163 , n85160 , n85162 );
buf ( n85164 , n84808 );
not ( n85165 , n85164 );
buf ( n85166 , n85165 );
buf ( n85167 , n85166 );
not ( n85168 , n85167 );
buf ( n85169 , n84904 );
not ( n85170 , n85169 );
or ( n85171 , n85168 , n85170 );
buf ( n85172 , n84875 );
nand ( n85173 , n85171 , n85172 );
buf ( n85174 , n85173 );
buf ( n85175 , n85174 );
nand ( n85176 , n85163 , n85175 );
buf ( n85177 , n85176 );
buf ( n85178 , n85177 );
xor ( n85179 , n85158 , n85178 );
buf ( n85180 , n85179 );
buf ( n85181 , n85180 );
xor ( n85182 , n85119 , n85181 );
not ( n85183 , n48855 );
not ( n85184 , n84891 );
or ( n85185 , n85183 , n85184 );
buf ( n85186 , n48808 );
not ( n85187 , n85186 );
buf ( n85188 , n41763 );
not ( n85189 , n85188 );
or ( n85190 , n85187 , n85189 );
buf ( n85191 , n41762 );
buf ( n85192 , n72891 );
nand ( n85193 , n85191 , n85192 );
buf ( n85194 , n85193 );
buf ( n85195 , n85194 );
nand ( n85196 , n85190 , n85195 );
buf ( n85197 , n85196 );
buf ( n85198 , n85197 );
buf ( n85199 , n48868 );
nand ( n85200 , n85198 , n85199 );
buf ( n85201 , n85200 );
nand ( n85202 , n85185 , n85201 );
not ( n85203 , n84583 );
not ( n85204 , n84608 );
or ( n85205 , n85203 , n85204 );
not ( n85206 , n84612 );
not ( n85207 , n84609 );
or ( n85208 , n85206 , n85207 );
nand ( n85209 , n85208 , n84572 );
nand ( n85210 , n85205 , n85209 );
xor ( n85211 , n85202 , n85210 );
not ( n85212 , n84759 );
not ( n85213 , n84690 );
or ( n85214 , n85212 , n85213 );
nand ( n85215 , n85214 , n84751 );
xor ( n85216 , n85211 , n85215 );
not ( n85217 , n84642 );
nand ( n85218 , n85217 , n84665 );
not ( n85219 , n85218 );
not ( n85220 , n84766 );
or ( n85221 , n85219 , n85220 );
buf ( n85222 , n84668 );
buf ( n85223 , n84642 );
nand ( n85224 , n85222 , n85223 );
buf ( n85225 , n85224 );
nand ( n85226 , n85221 , n85225 );
xor ( n85227 , n85216 , n85226 );
buf ( n85228 , n84601 );
not ( n85229 , n85228 );
buf ( n85230 , n50128 );
not ( n85231 , n85230 );
or ( n85232 , n85229 , n85231 );
buf ( n85233 , n47716 );
not ( n85234 , n85233 );
buf ( n85235 , n51804 );
not ( n85236 , n85235 );
or ( n85237 , n85234 , n85236 );
buf ( n85238 , n52673 );
buf ( n85239 , n47713 );
nand ( n85240 , n85238 , n85239 );
buf ( n85241 , n85240 );
buf ( n85242 , n85241 );
nand ( n85243 , n85237 , n85242 );
buf ( n85244 , n85243 );
buf ( n85245 , n85244 );
buf ( n85246 , n47872 );
nand ( n85247 , n85245 , n85246 );
buf ( n85248 , n85247 );
buf ( n85249 , n85248 );
nand ( n85250 , n85232 , n85249 );
buf ( n85251 , n85250 );
not ( n85252 , n39999 );
not ( n85253 , n84685 );
or ( n85254 , n85252 , n85253 );
buf ( n85255 , n70152 );
buf ( n85256 , n48975 );
nand ( n85257 , n85255 , n85256 );
buf ( n85258 , n85257 );
nand ( n85259 , n85254 , n85258 );
xor ( n85260 , n85251 , n85259 );
buf ( n85261 , n67149 );
not ( n85262 , n85261 );
buf ( n85263 , n64616 );
not ( n85264 , n85263 );
buf ( n85265 , n41873 );
not ( n85266 , n85265 );
or ( n85267 , n85264 , n85266 );
buf ( n85268 , n47063 );
buf ( n85269 , n45747 );
nand ( n85270 , n85268 , n85269 );
buf ( n85271 , n85270 );
buf ( n85272 , n85271 );
nand ( n85273 , n85267 , n85272 );
buf ( n85274 , n85273 );
buf ( n85275 , n85274 );
not ( n85276 , n85275 );
or ( n85277 , n85262 , n85276 );
buf ( n85278 , n84562 );
buf ( n85279 , n46225 );
nand ( n85280 , n85278 , n85279 );
buf ( n85281 , n85280 );
buf ( n85282 , n85281 );
nand ( n85283 , n85277 , n85282 );
buf ( n85284 , n85283 );
xor ( n85285 , n85260 , n85284 );
buf ( n85286 , n44496 );
not ( n85287 , n85286 );
buf ( n85288 , n70198 );
not ( n85289 , n85288 );
or ( n85290 , n85287 , n85289 );
buf ( n85291 , n84823 );
buf ( n85292 , n44517 );
nand ( n85293 , n85291 , n85292 );
buf ( n85294 , n85293 );
buf ( n85295 , n85294 );
nand ( n85296 , n85290 , n85295 );
buf ( n85297 , n85296 );
buf ( n85298 , n85297 );
xor ( n85299 , n70806 , n70831 );
xor ( n85300 , n85299 , n70904 );
buf ( n85301 , n85300 );
buf ( n85302 , n85301 );
xor ( n85303 , n85298 , n85302 );
xor ( n85304 , n84718 , n84722 );
and ( n85305 , n85304 , n84748 );
and ( n85306 , n84718 , n84722 );
or ( n85307 , n85305 , n85306 );
buf ( n85308 , n85307 );
buf ( n85309 , n85308 );
xor ( n85310 , n85303 , n85309 );
buf ( n85311 , n85310 );
xor ( n85312 , n85285 , n85311 );
not ( n85313 , n62125 );
not ( n85314 , n48836 );
not ( n85315 , n39672 );
or ( n85316 , n85314 , n85315 );
buf ( n85317 , n39685 );
not ( n85318 , n85317 );
buf ( n85319 , n61847 );
nand ( n85320 , n85318 , n85319 );
buf ( n85321 , n85320 );
nand ( n85322 , n85316 , n85321 );
not ( n85323 , n85322 );
or ( n85324 , n85313 , n85323 );
nand ( n85325 , n84655 , n51488 );
nand ( n85326 , n85324 , n85325 );
and ( n85327 , n85312 , n85326 );
not ( n85328 , n85312 );
not ( n85329 , n85326 );
and ( n85330 , n85328 , n85329 );
nor ( n85331 , n85327 , n85330 );
xor ( n85332 , n85227 , n85331 );
buf ( n85333 , n85332 );
xor ( n85334 , n85182 , n85333 );
buf ( n85335 , n85334 );
xor ( n85336 , n85029 , n85335 );
buf ( n85337 , n85336 );
xor ( n85338 , n84970 , n85337 );
buf ( n85339 , n85338 );
buf ( n85340 , n85339 );
xor ( n85341 , n84441 , n84512 );
xnor ( n85342 , n85341 , n84522 );
buf ( n85343 , n85342 );
xor ( n85344 , n76705 , n76711 );
and ( n85345 , n85344 , n76899 );
and ( n85346 , n76705 , n76711 );
or ( n85347 , n85345 , n85346 );
buf ( n85348 , n85347 );
buf ( n85349 , n85348 );
xor ( n85350 , n85343 , n85349 );
xor ( n85351 , n84939 , n84958 );
xnor ( n85352 , n85351 , n84964 );
buf ( n85353 , n85352 );
and ( n85354 , n85350 , n85353 );
and ( n85355 , n85343 , n85349 );
or ( n85356 , n85354 , n85355 );
buf ( n85357 , n85356 );
buf ( n85358 , n85357 );
not ( n85359 , n85358 );
buf ( n85360 , n85359 );
buf ( n85361 , n85360 );
nand ( n85362 , n85340 , n85361 );
buf ( n85363 , n85362 );
buf ( n85364 , n85363 );
not ( n85365 , n85364 );
xor ( n85366 , n85343 , n85349 );
xor ( n85367 , n85366 , n85353 );
buf ( n85368 , n85367 );
buf ( n85369 , n85368 );
buf ( n85370 , n85369 );
buf ( n85371 , n85370 );
buf ( n85372 , n85371 );
xor ( n85373 , n76677 , n76694 );
and ( n85374 , n85373 , n76902 );
and ( n85375 , n76677 , n76694 );
or ( n85376 , n85374 , n85375 );
buf ( n85377 , n85376 );
buf ( n85378 , n85377 );
nor ( n85379 , n85372 , n85378 );
buf ( n85380 , n85379 );
buf ( n85381 , n85380 );
nor ( n85382 , n85365 , n85381 );
buf ( n85383 , n85382 );
buf ( n85384 , n85383 );
buf ( n85385 , n67149 );
not ( n85386 , n85385 );
buf ( n85387 , n70928 );
not ( n85388 , n85387 );
or ( n85389 , n85386 , n85388 );
buf ( n85390 , n85274 );
buf ( n85391 , n46225 );
nand ( n85392 , n85390 , n85391 );
buf ( n85393 , n85392 );
buf ( n85394 , n85393 );
nand ( n85395 , n85389 , n85394 );
buf ( n85396 , n85395 );
not ( n85397 , n85396 );
xor ( n85398 , n85140 , n85144 );
and ( n85399 , n85398 , n85151 );
and ( n85400 , n85140 , n85144 );
or ( n85401 , n85399 , n85400 );
buf ( n85402 , n85401 );
not ( n85403 , n85402 );
not ( n85404 , n85403 );
or ( n85405 , n85397 , n85404 );
not ( n85406 , n85396 );
nand ( n85407 , n85402 , n85406 );
nand ( n85408 , n85405 , n85407 );
xor ( n85409 , n70784 , n70801 );
xor ( n85410 , n85409 , n70909 );
buf ( n85411 , n85410 );
and ( n85412 , n85408 , n85411 );
not ( n85413 , n85408 );
not ( n85414 , n85411 );
and ( n85415 , n85413 , n85414 );
nor ( n85416 , n85412 , n85415 );
buf ( n85417 , n85416 );
xor ( n85418 , n85202 , n85210 );
and ( n85419 , n85418 , n85215 );
and ( n85420 , n85202 , n85210 );
or ( n85421 , n85419 , n85420 );
buf ( n85422 , n85421 );
xor ( n85423 , n85417 , n85422 );
or ( n85424 , n85285 , n85311 );
not ( n85425 , n85424 );
not ( n85426 , n85326 );
or ( n85427 , n85425 , n85426 );
nand ( n85428 , n85285 , n85311 );
nand ( n85429 , n85427 , n85428 );
buf ( n85430 , n85429 );
xor ( n85431 , n85423 , n85430 );
buf ( n85432 , n85431 );
buf ( n85433 , n85432 );
buf ( n85434 , n44039 );
not ( n85435 , n85434 );
buf ( n85436 , n85101 );
not ( n85437 , n85436 );
and ( n85438 , n85435 , n85437 );
buf ( n85439 , n70951 );
buf ( n85440 , n38381 );
nor ( n85441 , n85439 , n85440 );
buf ( n85442 , n85441 );
buf ( n85443 , n85442 );
nor ( n85444 , n85438 , n85443 );
buf ( n85445 , n85444 );
not ( n85446 , n85445 );
not ( n85447 , n45053 );
not ( n85448 , n85073 );
and ( n85449 , n85447 , n85448 );
and ( n85450 , n70066 , n50104 );
nor ( n85451 , n85449 , n85450 );
not ( n85452 , n85451 );
xor ( n85453 , n85298 , n85302 );
and ( n85454 , n85453 , n85309 );
and ( n85455 , n85298 , n85302 );
or ( n85456 , n85454 , n85455 );
buf ( n85457 , n85456 );
xnor ( n85458 , n85452 , n85457 );
not ( n85459 , n85458 );
or ( n85460 , n85446 , n85459 );
or ( n85461 , n85458 , n85445 );
nand ( n85462 , n85460 , n85461 );
buf ( n85463 , n85462 );
buf ( n85464 , C1 );
buf ( n85465 , n85464 );
xor ( n85466 , n85463 , n85465 );
xor ( n85467 , n85251 , n85259 );
and ( n85468 , n85467 , n85284 );
and ( n85469 , n85251 , n85259 );
or ( n85470 , n85468 , n85469 );
and ( n85471 , n46907 , n85049 );
and ( n85472 , n28305 , n46890 );
not ( n85473 , n28305 );
and ( n85474 , n85473 , n46875 );
or ( n85475 , n85472 , n85474 );
and ( n85476 , n85475 , n46912 );
nor ( n85477 , n85471 , n85476 );
buf ( n85478 , n85477 );
not ( n85479 , n85478 );
buf ( n85480 , n85479 );
xor ( n85481 , n85470 , n85480 );
not ( n85482 , n48868 );
not ( n85483 , n70231 );
or ( n85484 , n85482 , n85483 );
buf ( n85485 , n85197 );
not ( n85486 , n85485 );
buf ( n85487 , n48858 );
nor ( n85488 , n85486 , n85487 );
buf ( n85489 , n85488 );
not ( n85490 , n85489 );
nand ( n85491 , n85484 , n85490 );
xnor ( n85492 , n85481 , n85491 );
buf ( n85493 , n85492 );
xor ( n85494 , n85466 , n85493 );
buf ( n85495 , n85494 );
buf ( n85496 , n85495 );
xor ( n85497 , n85433 , n85496 );
xor ( n85498 , n84998 , n85013 );
and ( n85499 , n85498 , n85026 );
and ( n85500 , n84998 , n85013 );
or ( n85501 , n85499 , n85500 );
buf ( n85502 , n85501 );
buf ( n85503 , n85502 );
xnor ( n85504 , n85497 , n85503 );
buf ( n85505 , n85504 );
buf ( n85506 , n85505 );
buf ( n85507 , n85028 );
not ( n85508 , n85507 );
buf ( n85509 , n84979 );
nand ( n85510 , n85508 , n85509 );
buf ( n85511 , n85510 );
buf ( n85512 , n85511 );
not ( n85513 , n85512 );
buf ( n85514 , n85335 );
not ( n85515 , n85514 );
or ( n85516 , n85513 , n85515 );
buf ( n85517 , n84979 );
not ( n85518 , n85517 );
buf ( n85519 , n85028 );
nand ( n85520 , n85518 , n85519 );
buf ( n85521 , n85520 );
buf ( n85522 , n85521 );
nand ( n85523 , n85516 , n85522 );
buf ( n85524 , n85523 );
buf ( n85525 , n85524 );
xor ( n85526 , n85506 , n85525 );
xor ( n85527 , n68618 , n68598 );
xnor ( n85528 , n85527 , n68644 );
buf ( n85529 , n85528 );
buf ( n85530 , n85244 );
not ( n85531 , n85530 );
buf ( n85532 , n42628 );
not ( n85533 , n85532 );
or ( n85534 , n85531 , n85533 );
buf ( n85535 , n69696 );
buf ( n85536 , n42564 );
nand ( n85537 , n85535 , n85536 );
buf ( n85538 , n85537 );
buf ( n85539 , n85538 );
nand ( n85540 , n85534 , n85539 );
buf ( n85541 , n85540 );
buf ( n85542 , n85541 );
xor ( n85543 , n85529 , n85542 );
buf ( n85544 , n69828 );
buf ( n85545 , n69758 );
xor ( n85546 , n85544 , n85545 );
buf ( n85547 , n69738 );
xnor ( n85548 , n85546 , n85547 );
buf ( n85549 , n85548 );
buf ( n85550 , n85549 );
xor ( n85551 , n85543 , n85550 );
buf ( n85552 , n85551 );
buf ( n85553 , n85552 );
buf ( n85554 , n70167 );
not ( n85555 , n85554 );
buf ( n85556 , n70205 );
not ( n85557 , n85556 );
or ( n85558 , n85555 , n85557 );
buf ( n85559 , n70205 );
buf ( n85560 , n70167 );
or ( n85561 , n85559 , n85560 );
nand ( n85562 , n85558 , n85561 );
buf ( n85563 , n85562 );
xnor ( n85564 , n70178 , n85563 );
buf ( n85565 , n85564 );
xor ( n85566 , n85553 , n85565 );
buf ( n85567 , n51290 );
buf ( n85568 , n56325 );
buf ( n85569 , n41795 );
and ( n85570 , n85568 , n85569 );
not ( n85571 , n85568 );
buf ( n85572 , n45270 );
and ( n85573 , n85571 , n85572 );
nor ( n85574 , n85570 , n85573 );
buf ( n85575 , n85574 );
buf ( n85576 , n85575 );
or ( n85577 , n85567 , n85576 );
buf ( n85578 , n55840 );
buf ( n85579 , n43434 );
and ( n85580 , n85578 , n85579 );
not ( n85581 , n85578 );
buf ( n85582 , n41772 );
and ( n85583 , n85581 , n85582 );
nor ( n85584 , n85580 , n85583 );
buf ( n85585 , n85584 );
buf ( n85586 , n85585 );
buf ( n85587 , n37416 );
or ( n85588 , n85586 , n85587 );
nand ( n85589 , n85577 , n85588 );
buf ( n85590 , n85589 );
buf ( n85591 , n85590 );
xor ( n85592 , n85566 , n85591 );
buf ( n85593 , n85592 );
buf ( n85594 , n85593 );
buf ( n85595 , C0 );
buf ( n85596 , n85595 );
xor ( n85597 , n85594 , n85596 );
and ( n85598 , n85035 , n85113 );
or ( n85599 , C0 , n85598 );
buf ( n85600 , n85599 );
buf ( n85601 , n85600 );
xor ( n85602 , n85597 , n85601 );
buf ( n85603 , n85602 );
buf ( n85604 , n85603 );
not ( n85605 , n85121 );
not ( n85606 , n85153 );
or ( n85607 , n85605 , n85606 );
nor ( n85608 , n85121 , n85153 );
not ( n85609 , n85126 );
or ( n85610 , n85608 , n85609 );
nand ( n85611 , n85607 , n85610 );
nand ( n85612 , n85082 , n85085 );
not ( n85613 , n85612 );
not ( n85614 , n85107 );
or ( n85615 , n85613 , n85614 );
nand ( n85616 , n85059 , n85081 );
nand ( n85617 , n85615 , n85616 );
xor ( n85618 , n85611 , n85617 );
not ( n85619 , n62125 );
buf ( n85620 , n48836 );
not ( n85621 , n85620 );
buf ( n85622 , n38851 );
not ( n85623 , n85622 );
or ( n85624 , n85621 , n85623 );
not ( n85625 , n44983 );
nand ( n85626 , n85625 , n61847 );
buf ( n85627 , n85626 );
nand ( n85628 , n85624 , n85627 );
buf ( n85629 , n85628 );
not ( n85630 , n85629 );
or ( n85631 , n85619 , n85630 );
nand ( n85632 , n85322 , n51488 );
nand ( n85633 , n85631 , n85632 );
xor ( n85634 , n85618 , n85633 );
buf ( n85635 , n85634 );
xor ( n85636 , n85155 , n85157 );
and ( n85637 , n85636 , n85178 );
or ( n85638 , n85637 , C0 );
buf ( n85639 , n85638 );
buf ( n85640 , n85639 );
xor ( n85641 , n85635 , n85640 );
xor ( n85642 , n85216 , n85226 );
and ( n85643 , n85642 , n85331 );
and ( n85644 , n85216 , n85226 );
or ( n85645 , n85643 , n85644 );
buf ( n85646 , n85645 );
xor ( n85647 , n85641 , n85646 );
buf ( n85648 , n85647 );
buf ( n85649 , n85648 );
xor ( n85650 , n85604 , n85649 );
xor ( n85651 , n85119 , n85181 );
and ( n85652 , n85651 , n85333 );
and ( n85653 , n85119 , n85181 );
or ( n85654 , n85652 , n85653 );
buf ( n85655 , n85654 );
buf ( n85656 , n85655 );
xor ( n85657 , n85650 , n85656 );
buf ( n85658 , n85657 );
buf ( n85659 , n85658 );
xnor ( n85660 , n85526 , n85659 );
buf ( n85661 , n85660 );
buf ( n85662 , n85661 );
xor ( n85663 , n84534 , n84969 );
and ( n85664 , n85663 , n85337 );
and ( n85665 , n84534 , n84969 );
or ( n85666 , n85664 , n85665 );
buf ( n85667 , n85666 );
buf ( n85668 , n85667 );
nand ( n85669 , n85662 , n85668 );
buf ( n85670 , n85669 );
buf ( n85671 , n85670 );
and ( n85672 , n85384 , n85671 );
buf ( n85673 , n85672 );
buf ( n85674 , n85673 );
not ( n85675 , n85674 );
or ( n85676 , n84437 , n85675 );
not ( n85677 , n85363 );
and ( n85678 , n85368 , n85377 );
not ( n85679 , n85678 );
or ( n85680 , n85677 , n85679 );
buf ( n85681 , n85339 );
buf ( n85682 , n85360 );
or ( n85683 , n85681 , n85682 );
buf ( n85684 , n85683 );
nand ( n85685 , n85680 , n85684 );
not ( n85686 , n85685 );
not ( n85687 , n85670 );
or ( n85688 , n85686 , n85687 );
buf ( n85689 , n85661 );
buf ( n85690 , n85667 );
or ( n85691 , n85689 , n85690 );
buf ( n85692 , n85691 );
nand ( n85693 , n85688 , n85692 );
buf ( n85694 , n85693 );
not ( n85695 , n85694 );
buf ( n85696 , n85695 );
buf ( n85697 , n85696 );
nand ( n85698 , n85676 , n85697 );
buf ( n85699 , n85698 );
buf ( n85700 , n85699 );
buf ( n85701 , n69708 );
buf ( n85702 , n69683 );
xor ( n85703 , n85701 , n85702 );
buf ( n85704 , n69839 );
xnor ( n85705 , n85703 , n85704 );
buf ( n85706 , n85705 );
buf ( n85707 , n85706 );
nand ( n85708 , n85403 , n85406 );
not ( n85709 , n85708 );
not ( n85710 , n85411 );
or ( n85711 , n85709 , n85710 );
nand ( n85712 , n85402 , n85396 );
nand ( n85713 , n85711 , n85712 );
buf ( n85714 , n85713 );
xor ( n85715 , n85707 , n85714 );
buf ( n85716 , n85452 );
not ( n85717 , n85716 );
buf ( n85718 , n85445 );
not ( n85719 , n85718 );
buf ( n85720 , n85719 );
buf ( n85721 , n85720 );
not ( n85722 , n85721 );
or ( n85723 , n85717 , n85722 );
buf ( n85724 , n85451 );
not ( n85725 , n85724 );
buf ( n85726 , n85445 );
not ( n85727 , n85726 );
or ( n85728 , n85725 , n85727 );
buf ( n85729 , n85457 );
nand ( n85730 , n85728 , n85729 );
buf ( n85731 , n85730 );
buf ( n85732 , n85731 );
nand ( n85733 , n85723 , n85732 );
buf ( n85734 , n85733 );
buf ( n85735 , n85734 );
and ( n85736 , n85715 , n85735 );
and ( n85737 , n85707 , n85714 );
or ( n85738 , n85736 , n85737 );
buf ( n85739 , n85738 );
buf ( n85740 , n85739 );
not ( n85741 , n70231 );
not ( n85742 , n48868 );
or ( n85743 , n85741 , n85742 );
not ( n85744 , n85477 );
nor ( n85745 , n85744 , n85489 );
nand ( n85746 , n85743 , n85745 );
not ( n85747 , n85746 );
not ( n85748 , n85470 );
or ( n85749 , n85747 , n85748 );
nand ( n85750 , n85480 , n85491 );
nand ( n85751 , n85749 , n85750 );
buf ( n85752 , n85751 );
buf ( n85753 , C0 );
buf ( n85754 , n85753 );
or ( n85755 , n85752 , n85754 );
xor ( n85756 , n85553 , n85565 );
and ( n85757 , n85756 , n85591 );
and ( n85758 , n85553 , n85565 );
or ( n85759 , n85757 , n85758 );
buf ( n85760 , n85759 );
buf ( n85761 , n85760 );
nand ( n85762 , n85755 , n85761 );
buf ( n85763 , n85762 );
buf ( n85764 , n85763 );
buf ( n85765 , C1 );
buf ( n85766 , n85765 );
and ( n85767 , n85764 , n85766 );
buf ( n85768 , n85767 );
buf ( n85769 , n85768 );
not ( n85770 , n85769 );
buf ( n85771 , n85770 );
buf ( n85772 , n85771 );
xor ( n85773 , n85740 , n85772 );
buf ( n85774 , n70138 );
buf ( n85775 , n70966 );
xor ( n85776 , n85774 , n85775 );
buf ( n85777 , n70243 );
xnor ( n85778 , n85776 , n85777 );
buf ( n85779 , n85778 );
buf ( n85780 , n85779 );
not ( n85781 , n85780 );
buf ( n85782 , n85781 );
buf ( n85783 , n85782 );
xnor ( n85784 , n85773 , n85783 );
buf ( n85785 , n85784 );
buf ( n85786 , n85785 );
not ( n85787 , n85786 );
buf ( n85788 , n85787 );
buf ( n85789 , n85788 );
not ( n85790 , n85789 );
buf ( n85791 , n69434 );
buf ( n85792 , n69465 );
xor ( n85793 , n85791 , n85792 );
buf ( n85794 , n69518 );
xnor ( n85795 , n85793 , n85794 );
buf ( n85796 , n85795 );
buf ( n85797 , n85796 );
not ( n85798 , n85797 );
buf ( n85799 , n85798 );
buf ( n85800 , n85799 );
not ( n85801 , n85800 );
buf ( n85802 , n69924 );
buf ( n85803 , n62125 );
and ( n85804 , n85802 , n85803 );
buf ( n85805 , n48836 );
not ( n85806 , n85805 );
buf ( n85807 , n42899 );
not ( n85808 , n85807 );
or ( n85809 , n85806 , n85808 );
buf ( n85810 , n42458 );
buf ( n85811 , n61847 );
nand ( n85812 , n85810 , n85811 );
buf ( n85813 , n85812 );
buf ( n85814 , n85813 );
nand ( n85815 , n85809 , n85814 );
buf ( n85816 , n85815 );
buf ( n85817 , n85816 );
not ( n85818 , n85817 );
buf ( n85819 , n51489 );
nor ( n85820 , n85818 , n85819 );
buf ( n85821 , n85820 );
buf ( n85822 , n85821 );
nor ( n85823 , n85804 , n85822 );
buf ( n85824 , n85823 );
buf ( n85825 , n85824 );
not ( n85826 , n85825 );
or ( n85827 , n85801 , n85826 );
buf ( n85828 , n85824 );
not ( n85829 , n85828 );
buf ( n85830 , n85829 );
buf ( n85831 , n85830 );
buf ( n85832 , n85796 );
nand ( n85833 , n85831 , n85832 );
buf ( n85834 , n85833 );
buf ( n85835 , n85834 );
nand ( n85836 , n85827 , n85835 );
buf ( n85837 , n85836 );
xor ( n85838 , n69842 , n69867 );
xor ( n85839 , n85838 , n69893 );
buf ( n85840 , n85839 );
xor ( n85841 , n85837 , n85840 );
buf ( n85842 , n85841 );
buf ( n85843 , C0 );
xor ( n85844 , n85529 , n85542 );
and ( n85845 , n85844 , n85550 );
and ( n85846 , n85529 , n85542 );
or ( n85847 , n85845 , n85846 );
buf ( n85848 , n85847 );
buf ( n85849 , n85848 );
buf ( n85850 , n46907 );
not ( n85851 , n85850 );
buf ( n85852 , n85475 );
not ( n85853 , n85852 );
or ( n85854 , n85851 , n85853 );
buf ( n85855 , n69624 );
not ( n85856 , n85855 );
buf ( n85857 , n46912 );
nand ( n85858 , n85856 , n85857 );
buf ( n85859 , n85858 );
buf ( n85860 , n85859 );
nand ( n85861 , n85854 , n85860 );
buf ( n85862 , n85861 );
buf ( n85863 , n85862 );
xor ( n85864 , n85849 , n85863 );
buf ( n85865 , n85585 );
not ( n85866 , n85865 );
buf ( n85867 , n85866 );
buf ( n85868 , n85867 );
not ( n85869 , n85868 );
buf ( n85870 , n37400 );
not ( n85871 , n85870 );
or ( n85872 , n85869 , n85871 );
buf ( n85873 , n69880 );
buf ( n85874 , n37413 );
nand ( n85875 , n85873 , n85874 );
buf ( n85876 , n85875 );
buf ( n85877 , n85876 );
nand ( n85878 , n85872 , n85877 );
buf ( n85879 , n85878 );
buf ( n85880 , n85879 );
and ( n85881 , n85864 , n85880 );
and ( n85882 , n85849 , n85863 );
or ( n85883 , n85881 , n85882 );
buf ( n85884 , n85883 );
xor ( n85885 , n85843 , n85884 );
not ( n85886 , n69657 );
not ( n85887 , n69630 );
or ( n85888 , n85886 , n85887 );
nand ( n85889 , n69654 , n69633 );
nand ( n85890 , n85888 , n85889 );
not ( n85891 , n69615 );
and ( n85892 , n85890 , n85891 );
not ( n85893 , n85890 );
and ( n85894 , n85893 , n69615 );
nor ( n85895 , n85892 , n85894 );
not ( n85896 , n85895 );
xor ( n85897 , n85885 , n85896 );
buf ( n85898 , n85897 );
xor ( n85899 , n85842 , n85898 );
xor ( n85900 , n70218 , n70225 );
xor ( n85901 , n85900 , n70239 );
buf ( n85902 , n85901 );
buf ( n85903 , C0 );
buf ( n85904 , n85903 );
buf ( n85905 , n85902 );
or ( n85906 , n85904 , n85905 );
xor ( n85907 , n85849 , n85863 );
xor ( n85908 , n85907 , n85880 );
buf ( n85909 , n85908 );
buf ( n85910 , n85909 );
nand ( n85911 , n85906 , n85910 );
buf ( n85912 , n85911 );
buf ( n85913 , n85912 );
nand ( n85914 , C1 , n85913 );
buf ( n85915 , n85914 );
buf ( n85916 , n85915 );
xor ( n85917 , n85899 , n85916 );
buf ( n85918 , n85917 );
buf ( n85919 , n85918 );
not ( n85920 , n85919 );
or ( n85921 , n85790 , n85920 );
buf ( n85922 , n85918 );
buf ( n85923 , n85788 );
or ( n85924 , n85922 , n85923 );
buf ( n85925 , n85909 );
buf ( n85926 , n85902 );
xor ( n85927 , n85925 , n85926 );
xor ( n85928 , n85927 , C1 );
buf ( n85929 , n85928 );
buf ( n85930 , n85929 );
not ( n85931 , n85930 );
buf ( n85932 , n85931 );
not ( n85933 , n85932 );
xor ( n85934 , n85594 , n85596 );
and ( n85935 , n85934 , n85601 );
or ( n85936 , n85935 , C0 );
buf ( n85937 , n85936 );
not ( n85938 , n85937 );
or ( n85939 , n85933 , n85938 );
buf ( n85940 , n85937 );
not ( n85941 , n85940 );
buf ( n85942 , n85941 );
not ( n85943 , n85942 );
not ( n85944 , n85929 );
or ( n85945 , n85943 , n85944 );
not ( n85946 , n85617 );
not ( n85947 , n85633 );
or ( n85948 , n85946 , n85947 );
or ( n85949 , n85633 , n85617 );
nand ( n85950 , n85949 , n85611 );
nand ( n85951 , n85948 , n85950 );
buf ( n85952 , n85951 );
xor ( n85953 , n85707 , n85714 );
xor ( n85954 , n85953 , n85735 );
buf ( n85955 , n85954 );
buf ( n85956 , n85955 );
xor ( n85957 , n85952 , n85956 );
buf ( n85958 , n85957 );
buf ( n85959 , n85958 );
buf ( n85960 , n70053 );
not ( n85961 , n85960 );
not ( n85962 , n70078 );
not ( n85963 , n68649 );
not ( n85964 , n70085 );
or ( n85965 , n85963 , n85964 );
or ( n85966 , n68649 , n70091 );
nand ( n85967 , n85965 , n85966 );
not ( n85968 , n85967 );
or ( n85969 , n85962 , n85968 );
or ( n85970 , n70078 , n70093 );
nand ( n85971 , n85969 , n85970 );
buf ( n85972 , n85971 );
not ( n85973 , n85972 );
or ( n85974 , n85961 , n85973 );
buf ( n85975 , n85971 );
buf ( n85976 , n70053 );
or ( n85977 , n85975 , n85976 );
nand ( n85978 , n85974 , n85977 );
buf ( n85979 , n85978 );
buf ( n85980 , n85979 );
buf ( n85981 , n51488 );
not ( n85982 , n85981 );
buf ( n85983 , n85629 );
not ( n85984 , n85983 );
or ( n85985 , n85982 , n85984 );
buf ( n85986 , n85816 );
buf ( n85987 , n62125 );
nand ( n85988 , n85986 , n85987 );
buf ( n85989 , n85988 );
buf ( n85990 , n85989 );
nand ( n85991 , n85985 , n85990 );
buf ( n85992 , n85991 );
buf ( n85993 , n85992 );
xor ( n85994 , n85980 , n85993 );
xor ( n85995 , n70914 , n70939 );
xor ( n85996 , n85995 , n70962 );
buf ( n85997 , n85996 );
buf ( n85998 , n85997 );
xor ( n85999 , n85994 , n85998 );
buf ( n86000 , n85999 );
buf ( n86001 , n86000 );
and ( n86002 , n85959 , n86001 );
not ( n86003 , n85959 );
buf ( n86004 , n86000 );
not ( n86005 , n86004 );
buf ( n86006 , n86005 );
buf ( n86007 , n86006 );
and ( n86008 , n86003 , n86007 );
nor ( n86009 , n86002 , n86008 );
buf ( n86010 , n86009 );
nand ( n86011 , n85945 , n86010 );
nand ( n86012 , n85939 , n86011 );
buf ( n86013 , n86012 );
nand ( n86014 , n85924 , n86013 );
buf ( n86015 , n86014 );
buf ( n86016 , n86015 );
nand ( n86017 , n85921 , n86016 );
buf ( n86018 , n86017 );
buf ( n86019 , n86018 );
xor ( n86020 , n70130 , n70134 );
xor ( n86021 , n86020 , n70973 );
buf ( n86022 , n86021 );
buf ( n86023 , n86022 );
buf ( n86024 , n70111 );
not ( n86025 , n86024 );
buf ( n86026 , n86025 );
not ( n86027 , n86026 );
and ( n86028 , n86027 , n70007 );
nor ( n86029 , C0 , n86028 );
nand ( n86030 , C1 , n70006 );
and ( n86031 , n86026 , n86030 );
not ( n86032 , n86026 );
and ( n86033 , n86032 , C1 );
or ( n86034 , n86031 , n86033 );
nand ( n86035 , n86029 , n86034 );
buf ( n86036 , n86035 );
xor ( n86037 , n86023 , n86036 );
xor ( n86038 , n85842 , n85898 );
and ( n86039 , n86038 , n85916 );
and ( n86040 , n85842 , n85898 );
or ( n86041 , n86039 , n86040 );
buf ( n86042 , n86041 );
buf ( n86043 , n86042 );
xor ( n86044 , n86037 , n86043 );
buf ( n86045 , n86044 );
buf ( n86046 , n86045 );
and ( n86047 , n86019 , n86046 );
not ( n86048 , n86019 );
buf ( n86049 , n86045 );
not ( n86050 , n86049 );
buf ( n86051 , n86050 );
buf ( n86052 , n86051 );
and ( n86053 , n86048 , n86052 );
nor ( n86054 , n86047 , n86053 );
buf ( n86055 , n86054 );
buf ( n86056 , n86055 );
buf ( n86057 , n85799 );
not ( n86058 , n86057 );
buf ( n86059 , n85830 );
not ( n86060 , n86059 );
or ( n86061 , n86058 , n86060 );
buf ( n86062 , n85796 );
not ( n86063 , n86062 );
buf ( n86064 , n85824 );
not ( n86065 , n86064 );
or ( n86066 , n86063 , n86065 );
buf ( n86067 , n85840 );
nand ( n86068 , n86066 , n86067 );
buf ( n86069 , n86068 );
buf ( n86070 , n86069 );
nand ( n86071 , n86061 , n86070 );
buf ( n86072 , n86071 );
buf ( n86073 , n86072 );
xor ( n86074 , n69926 , n69935 );
xor ( n86075 , n86074 , n69946 );
buf ( n86076 , n86075 );
xor ( n86077 , n86073 , n86076 );
xor ( n86078 , n69659 , n69897 );
xor ( n86079 , n86078 , n69901 );
buf ( n86080 , n86079 );
xnor ( n86081 , n86077 , n86080 );
buf ( n86082 , n86081 );
buf ( n86083 , n86082 );
not ( n86084 , n85771 );
not ( n86085 , n85782 );
or ( n86086 , n86084 , n86085 );
not ( n86087 , n85779 );
not ( n86088 , n85768 );
or ( n86089 , n86087 , n86088 );
nand ( n86090 , n86089 , n85739 );
nand ( n86091 , n86086 , n86090 );
not ( n86092 , n86091 );
not ( n86093 , n85896 );
or ( n86094 , n86093 , C1 );
not ( n86095 , n85895 );
or ( n86096 , C0 , n86095 );
nand ( n86097 , n86096 , n85884 );
nand ( n86098 , n86094 , n86097 );
not ( n86099 , n86098 );
not ( n86100 , n86099 );
buf ( n86101 , n70097 );
not ( n86102 , n86101 );
buf ( n86103 , n70026 );
not ( n86104 , n86103 );
or ( n86105 , n86102 , n86104 );
buf ( n86106 , n70097 );
not ( n86107 , n86106 );
buf ( n86108 , n70023 );
nand ( n86109 , n86107 , n86108 );
buf ( n86110 , n86109 );
buf ( n86111 , n86110 );
nand ( n86112 , n86105 , n86111 );
buf ( n86113 , n86112 );
buf ( n86114 , n86113 );
buf ( n86115 , n70046 );
and ( n86116 , n86114 , n86115 );
not ( n86117 , n86114 );
buf ( n86118 , n70104 );
and ( n86119 , n86117 , n86118 );
nor ( n86120 , n86116 , n86119 );
buf ( n86121 , n86120 );
buf ( n86122 , n86121 );
not ( n86123 , n86122 );
or ( n86124 , C0 , n86123 );
xor ( n86125 , n85980 , n85993 );
and ( n86126 , n86125 , n85998 );
and ( n86127 , n85980 , n85993 );
or ( n86128 , n86126 , n86127 );
buf ( n86129 , n86128 );
buf ( n86130 , n86129 );
nand ( n86131 , n86124 , n86130 );
buf ( n86132 , n86131 );
buf ( n86133 , n86121 );
not ( n86134 , n86133 );
buf ( n86135 , n86134 );
buf ( n86136 , C1 );
nand ( n86137 , n86132 , n86136 );
not ( n86138 , n86137 );
or ( n86139 , n86100 , n86138 );
or ( n86140 , n86137 , n86099 );
nand ( n86141 , n86139 , n86140 );
not ( n86142 , n86141 );
or ( n86143 , n86092 , n86142 );
not ( n86144 , n86091 );
not ( n86145 , n86144 );
or ( n86146 , n86145 , n86141 );
nand ( n86147 , n86143 , n86146 );
buf ( n86148 , n86147 );
xor ( n86149 , n86083 , n86148 );
buf ( n86150 , n85955 );
buf ( n86151 , n85951 );
or ( n86152 , n86150 , n86151 );
buf ( n86153 , n86152 );
buf ( n86154 , n86153 );
buf ( n86155 , n86000 );
and ( n86156 , n86154 , n86155 );
and ( n86157 , n85952 , n85956 );
buf ( n86158 , n86157 );
buf ( n86159 , n86158 );
nor ( n86160 , n86156 , n86159 );
buf ( n86161 , n86160 );
buf ( n86162 , n86161 );
and ( n86163 , n86129 , C1 );
or ( n86164 , n86163 , C0 );
buf ( n86165 , n86164 );
buf ( n86166 , n86135 );
xnor ( n86167 , n86165 , n86166 );
buf ( n86168 , n86167 );
buf ( n86169 , n86168 );
xor ( n86170 , n86162 , n86169 );
and ( n86171 , n85421 , n85416 );
or ( n86172 , n85429 , n86171 );
or ( n86173 , n85421 , n85416 );
nand ( n86174 , n86172 , n86173 );
buf ( n86175 , n86174 );
xor ( n86176 , n85463 , n85465 );
and ( n86177 , n86176 , n85493 );
and ( n86178 , n85463 , n85465 );
or ( n86179 , n86177 , n86178 );
buf ( n86180 , n86179 );
buf ( n86181 , n86180 );
xor ( n86182 , n86175 , n86181 );
xor ( n86183 , n85751 , n85753 );
xnor ( n86184 , n86183 , n85760 );
buf ( n86185 , n86184 );
and ( n86186 , n86182 , n86185 );
and ( n86187 , n86175 , n86181 );
or ( n86188 , n86186 , n86187 );
buf ( n86189 , n86188 );
buf ( n86190 , n86189 );
and ( n86191 , n86170 , n86190 );
and ( n86192 , n86162 , n86169 );
or ( n86193 , n86191 , n86192 );
buf ( n86194 , n86193 );
buf ( n86195 , n86194 );
xor ( n86196 , n86149 , n86195 );
buf ( n86197 , n86196 );
buf ( n86198 , n86197 );
and ( n86199 , n86056 , n86198 );
not ( n86200 , n86056 );
buf ( n86201 , n86197 );
not ( n86202 , n86201 );
buf ( n86203 , n86202 );
buf ( n86204 , n86203 );
and ( n86205 , n86200 , n86204 );
nor ( n86206 , n86199 , n86205 );
buf ( n86207 , n86206 );
buf ( n86208 , n86207 );
xor ( n86209 , n86162 , n86169 );
xor ( n86210 , n86209 , n86190 );
buf ( n86211 , n86210 );
buf ( n86212 , n86211 );
not ( n86213 , n85495 );
buf ( n86214 , n85432 );
not ( n86215 , n86214 );
buf ( n86216 , n86215 );
not ( n86217 , n86216 );
and ( n86218 , n86213 , n86217 );
buf ( n86219 , n85495 );
buf ( n86220 , n86216 );
nand ( n86221 , n86219 , n86220 );
buf ( n86222 , n86221 );
and ( n86223 , n86222 , n85502 );
nor ( n86224 , n86218 , n86223 );
buf ( n86225 , n86224 );
not ( n86226 , n86225 );
xor ( n86227 , n86175 , n86181 );
xor ( n86228 , n86227 , n86185 );
buf ( n86229 , n86228 );
buf ( n86230 , n86229 );
not ( n86231 , n86230 );
or ( n86232 , n86226 , n86231 );
xor ( n86233 , n85635 , n85640 );
and ( n86234 , n86233 , n85646 );
and ( n86235 , n85635 , n85640 );
or ( n86236 , n86234 , n86235 );
buf ( n86237 , n86236 );
buf ( n86238 , n86237 );
nand ( n86239 , n86232 , n86238 );
buf ( n86240 , n86239 );
buf ( n86241 , n86240 );
buf ( n86242 , n86224 );
not ( n86243 , n86242 );
buf ( n86244 , n86229 );
not ( n86245 , n86244 );
buf ( n86246 , n86245 );
buf ( n86247 , n86246 );
nand ( n86248 , n86243 , n86247 );
buf ( n86249 , n86248 );
buf ( n86250 , n86249 );
and ( n86251 , n86241 , n86250 );
buf ( n86252 , n86251 );
buf ( n86253 , n86252 );
xor ( n86254 , n86212 , n86253 );
buf ( n86255 , n85785 );
buf ( n86256 , n85918 );
xor ( n86257 , n86255 , n86256 );
buf ( n86258 , n86012 );
xor ( n86259 , n86257 , n86258 );
buf ( n86260 , n86259 );
buf ( n86261 , n86260 );
and ( n86262 , n86254 , n86261 );
and ( n86263 , n86212 , n86253 );
or ( n86264 , n86262 , n86263 );
buf ( n86265 , n86264 );
buf ( n86266 , n86265 );
nand ( n86267 , n86208 , n86266 );
buf ( n86268 , n86267 );
buf ( n86269 , n86268 );
buf ( n86270 , n85937 );
not ( n86271 , n86270 );
buf ( n86272 , n85929 );
not ( n86273 , n86272 );
or ( n86274 , n86271 , n86273 );
buf ( n86275 , n85932 );
buf ( n86276 , n85942 );
nand ( n86277 , n86275 , n86276 );
buf ( n86278 , n86277 );
buf ( n86279 , n86278 );
nand ( n86280 , n86274 , n86279 );
buf ( n86281 , n86280 );
buf ( n86282 , n86281 );
buf ( n86283 , n86010 );
xor ( n86284 , n86282 , n86283 );
buf ( n86285 , n86284 );
buf ( n86286 , n86285 );
xor ( n86287 , n85604 , n85649 );
and ( n86288 , n86287 , n85656 );
and ( n86289 , n85604 , n85649 );
or ( n86290 , n86288 , n86289 );
buf ( n86291 , n86290 );
buf ( n86292 , n86291 );
xor ( n86293 , n86286 , n86292 );
buf ( n86294 , n86237 );
buf ( n86295 , n86224 );
xor ( n86296 , n86294 , n86295 );
buf ( n86297 , n86246 );
xnor ( n86298 , n86296 , n86297 );
buf ( n86299 , n86298 );
buf ( n86300 , n86299 );
and ( n86301 , n86293 , n86300 );
and ( n86302 , n86286 , n86292 );
or ( n86303 , n86301 , n86302 );
buf ( n86304 , n86303 );
buf ( n86305 , n86304 );
not ( n86306 , n86305 );
xor ( n86307 , n86212 , n86253 );
xor ( n86308 , n86307 , n86261 );
buf ( n86309 , n86308 );
buf ( n86310 , n86309 );
nand ( n86311 , n86306 , n86310 );
buf ( n86312 , n86311 );
buf ( n86313 , n86312 );
not ( n86314 , n86313 );
xor ( n86315 , n86286 , n86292 );
xor ( n86316 , n86315 , n86300 );
buf ( n86317 , n86316 );
buf ( n86318 , n86317 );
buf ( n86319 , n85505 );
not ( n86320 , n86319 );
buf ( n86321 , n85524 );
not ( n86322 , n86321 );
or ( n86323 , n86320 , n86322 );
or ( n86324 , n85505 , n85524 );
nand ( n86325 , n86324 , n85658 );
buf ( n86326 , n86325 );
nand ( n86327 , n86323 , n86326 );
buf ( n86328 , n86327 );
buf ( n86329 , n86328 );
nor ( n86330 , n86318 , n86329 );
buf ( n86331 , n86330 );
buf ( n86332 , n86331 );
nor ( n86333 , n86314 , n86332 );
buf ( n86334 , n86333 );
buf ( n86335 , n86334 );
nand ( n86336 , n85700 , n86269 , n86335 );
buf ( n86337 , n86336 );
buf ( n86338 , n86337 );
not ( n86339 , n86312 );
buf ( n86340 , n86328 );
buf ( n86341 , n86317 );
and ( n86342 , n86340 , n86341 );
buf ( n86343 , n86342 );
not ( n86344 , n86343 );
or ( n86345 , n86339 , n86344 );
buf ( n86346 , n86309 );
not ( n86347 , n86346 );
buf ( n86348 , n86304 );
nand ( n86349 , n86347 , n86348 );
buf ( n86350 , n86349 );
nand ( n86351 , n86345 , n86350 );
buf ( n86352 , n86351 );
buf ( n86353 , n86268 );
nand ( n86354 , n86352 , n86353 );
buf ( n86355 , n86354 );
buf ( n86356 , n86355 );
buf ( n86357 , n86207 );
buf ( n86358 , n86265 );
or ( n86359 , n86357 , n86358 );
buf ( n86360 , n86359 );
buf ( n86361 , n86360 );
nand ( n86362 , n86338 , n86356 , n86361 );
buf ( n86363 , n86362 );
buf ( n86364 , n86363 );
xor ( n86365 , n69366 , n69562 );
xor ( n86366 , n86365 , n69964 );
buf ( n86367 , n86366 );
buf ( n86368 , n69536 );
buf ( n86369 , n69541 );
xor ( n86370 , n86368 , n86369 );
buf ( n86371 , n69556 );
xnor ( n86372 , n86370 , n86371 );
buf ( n86373 , n86372 );
buf ( n86374 , n86373 );
not ( n86375 , n86374 );
xor ( n86376 , n69910 , n69913 );
xor ( n86377 , n86376 , n69960 );
buf ( n86378 , n86377 );
buf ( n86379 , n86378 );
not ( n86380 , n86379 );
buf ( n86381 , n86380 );
buf ( n86382 , n86381 );
not ( n86383 , n86382 );
or ( n86384 , n86375 , n86383 );
not ( n86385 , n86072 );
not ( n86386 , n86079 );
or ( n86387 , n86385 , n86386 );
buf ( n86388 , n86079 );
buf ( n86389 , n86072 );
or ( n86390 , n86388 , n86389 );
buf ( n86391 , n86075 );
nand ( n86392 , n86390 , n86391 );
buf ( n86393 , n86392 );
nand ( n86394 , n86387 , n86393 );
xor ( n86395 , n69917 , n69950 );
xor ( n86396 , n86395 , n69955 );
buf ( n86397 , n86396 );
xor ( n86398 , n86394 , n86397 );
xor ( n86399 , n69991 , n69994 );
xor ( n86400 , n86399 , n70115 );
buf ( n86401 , n86400 );
and ( n86402 , n86398 , n86401 );
and ( n86403 , n86394 , n86397 );
or ( n86404 , n86402 , n86403 );
buf ( n86405 , n86404 );
nand ( n86406 , n86384 , n86405 );
buf ( n86407 , n86406 );
buf ( n86408 , n86407 );
buf ( n86409 , n86373 );
not ( n86410 , n86409 );
buf ( n86411 , n86378 );
nand ( n86412 , n86410 , n86411 );
buf ( n86413 , n86412 );
buf ( n86414 , n86413 );
nand ( n86415 , n86408 , n86414 );
buf ( n86416 , n86415 );
buf ( n86417 , n86416 );
xor ( n86418 , n86367 , n86417 );
xor ( n86419 , n69975 , n69979 );
xor ( n86420 , n86419 , n70992 );
buf ( n86421 , n86420 );
buf ( n86422 , n86421 );
xor ( n86423 , n86418 , n86422 );
buf ( n86424 , n86423 );
buf ( n86425 , n86424 );
not ( n86426 , n86425 );
buf ( n86427 , n86426 );
buf ( n86428 , n86427 );
xor ( n86429 , n70119 , n70123 );
xor ( n86430 , n86429 , n70987 );
buf ( n86431 , n86430 );
not ( n86432 , n86431 );
buf ( n86433 , n86432 );
not ( n86434 , n86433 );
buf ( n86435 , n86373 );
buf ( n86436 , n86404 );
xor ( n86437 , n86435 , n86436 );
buf ( n86438 , n86378 );
xor ( n86439 , n86437 , n86438 );
buf ( n86440 , n86439 );
buf ( n86441 , n86440 );
not ( n86442 , n86441 );
or ( n86443 , n86434 , n86442 );
xor ( n86444 , n70128 , n70977 );
xor ( n86445 , n86444 , n70982 );
buf ( n86446 , n86445 );
buf ( n86447 , n86446 );
not ( n86448 , n86098 );
not ( n86449 , n86091 );
or ( n86450 , n86448 , n86449 );
not ( n86451 , n86099 );
not ( n86452 , n86144 );
or ( n86453 , n86451 , n86452 );
nand ( n86454 , n86453 , n86137 );
nand ( n86455 , n86450 , n86454 );
buf ( n86456 , n86455 );
or ( n86457 , n86447 , n86456 );
buf ( n86458 , n86457 );
buf ( n86459 , n86458 );
xor ( n86460 , n86023 , n86036 );
and ( n86461 , n86460 , n86043 );
and ( n86462 , n86023 , n86036 );
or ( n86463 , n86461 , n86462 );
buf ( n86464 , n86463 );
buf ( n86465 , n86464 );
and ( n86466 , n86459 , n86465 );
buf ( n86467 , n86446 );
buf ( n86468 , n86455 );
and ( n86469 , n86467 , n86468 );
buf ( n86470 , n86469 );
buf ( n86471 , n86470 );
nor ( n86472 , n86466 , n86471 );
buf ( n86473 , n86472 );
not ( n86474 , n86473 );
buf ( n86475 , n86474 );
nand ( n86476 , n86443 , n86475 );
buf ( n86477 , n86476 );
buf ( n86478 , n86477 );
buf ( n86479 , n86440 );
not ( n86480 , n86479 );
buf ( n86481 , n86480 );
buf ( n86482 , n86481 );
buf ( n86483 , n86431 );
nand ( n86484 , n86482 , n86483 );
buf ( n86485 , n86484 );
buf ( n86486 , n86485 );
nand ( n86487 , n86478 , n86486 );
buf ( n86488 , n86487 );
buf ( n86489 , n86488 );
not ( n86490 , n86489 );
buf ( n86491 , n86490 );
buf ( n86492 , n86491 );
nand ( n86493 , n86428 , n86492 );
buf ( n86494 , n86493 );
buf ( n86495 , n86494 );
not ( n86496 , n86495 );
xor ( n86497 , n71002 , n71003 );
buf ( n86498 , n86497 );
buf ( n86499 , n86498 );
buf ( n86500 , n69357 );
and ( n86501 , n86499 , n86500 );
not ( n86502 , n86499 );
buf ( n86503 , n69357 );
not ( n86504 , n86503 );
buf ( n86505 , n86504 );
buf ( n86506 , n86505 );
and ( n86507 , n86502 , n86506 );
nor ( n86508 , n86501 , n86507 );
buf ( n86509 , n86508 );
buf ( n86510 , n86509 );
xor ( n86511 , n86367 , n86417 );
and ( n86512 , n86511 , n86422 );
and ( n86513 , n86367 , n86417 );
or ( n86514 , n86512 , n86513 );
buf ( n86515 , n86514 );
buf ( n86516 , n86515 );
nor ( n86517 , n86510 , n86516 );
buf ( n86518 , n86517 );
buf ( n86519 , n86518 );
nor ( n86520 , n86496 , n86519 );
buf ( n86521 , n86520 );
buf ( n86522 , n86521 );
buf ( n86523 , n86051 );
not ( n86524 , n86523 );
buf ( n86525 , n86197 );
not ( n86526 , n86525 );
or ( n86527 , n86524 , n86526 );
buf ( n86528 , n86018 );
nand ( n86529 , n86527 , n86528 );
buf ( n86530 , n86529 );
buf ( n86531 , n86530 );
buf ( n86532 , n86203 );
buf ( n86533 , n86045 );
nand ( n86534 , n86532 , n86533 );
buf ( n86535 , n86534 );
buf ( n86536 , n86535 );
nand ( n86537 , n86531 , n86536 );
buf ( n86538 , n86537 );
buf ( n86539 , n86538 );
xor ( n86540 , n86467 , n86468 );
buf ( n86541 , n86540 );
buf ( n86542 , n86541 );
buf ( n86543 , n86464 );
not ( n86544 , n86543 );
buf ( n86545 , n86544 );
buf ( n86546 , n86545 );
and ( n86547 , n86542 , n86546 );
not ( n86548 , n86542 );
buf ( n86549 , n86464 );
and ( n86550 , n86548 , n86549 );
nor ( n86551 , n86547 , n86550 );
buf ( n86552 , n86551 );
xor ( n86553 , n86394 , n86397 );
xor ( n86554 , n86553 , n86401 );
buf ( n86555 , n86554 );
not ( n86556 , n86555 );
buf ( n86557 , n86556 );
buf ( n86558 , n86557 );
not ( n86559 , n86558 );
xor ( n86560 , n86083 , n86148 );
and ( n86561 , n86560 , n86195 );
and ( n86562 , n86083 , n86148 );
or ( n86563 , n86561 , n86562 );
buf ( n86564 , n86563 );
buf ( n86565 , n86564 );
not ( n86566 , n86565 );
buf ( n86567 , n86566 );
buf ( n86568 , n86567 );
not ( n86569 , n86568 );
or ( n86570 , n86559 , n86569 );
buf ( n86571 , n86564 );
buf ( n86572 , n86554 );
nand ( n86573 , n86571 , n86572 );
buf ( n86574 , n86573 );
buf ( n86575 , n86574 );
nand ( n86576 , n86570 , n86575 );
buf ( n86577 , n86576 );
xnor ( n86578 , n86552 , n86577 );
buf ( n86579 , n86578 );
or ( n86580 , n86539 , n86579 );
buf ( n86581 , n86580 );
buf ( n86582 , n86581 );
not ( n86583 , n86432 );
not ( n86584 , n86473 );
or ( n86585 , n86583 , n86584 );
nand ( n86586 , n86474 , n86431 );
nand ( n86587 , n86585 , n86586 );
and ( n86588 , n86587 , n86481 );
not ( n86589 , n86587 );
not ( n86590 , n86481 );
and ( n86591 , n86589 , n86590 );
nor ( n86592 , n86588 , n86591 );
buf ( n86593 , n86592 );
not ( n86594 , n86552 );
not ( n86595 , n86557 );
and ( n86596 , n86594 , n86595 );
buf ( n86597 , n86552 );
buf ( n86598 , n86557 );
nand ( n86599 , n86597 , n86598 );
buf ( n86600 , n86599 );
and ( n86601 , n86600 , n86567 );
nor ( n86602 , n86596 , n86601 );
buf ( n86603 , n86602 );
nand ( n86604 , n86593 , n86603 );
buf ( n86605 , n86604 );
buf ( n86606 , n86605 );
and ( n86607 , n86582 , n86606 );
buf ( n86608 , n86607 );
buf ( n86609 , n86608 );
nand ( n86610 , n86364 , n86522 , n86609 );
buf ( n86611 , n86610 );
buf ( n86612 , n86611 );
not ( n86613 , n86494 );
not ( n86614 , n86605 );
buf ( n86615 , n86578 );
buf ( n86616 , n86538 );
and ( n86617 , n86615 , n86616 );
buf ( n86618 , n86617 );
not ( n86619 , n86618 );
or ( n86620 , n86614 , n86619 );
buf ( n86621 , n86592 );
not ( n86622 , n86621 );
buf ( n86623 , n86622 );
buf ( n86624 , n86623 );
buf ( n86625 , n86602 );
not ( n86626 , n86625 );
buf ( n86627 , n86626 );
buf ( n86628 , n86627 );
nand ( n86629 , n86624 , n86628 );
buf ( n86630 , n86629 );
nand ( n86631 , n86620 , n86630 );
not ( n86632 , n86631 );
or ( n86633 , n86613 , n86632 );
buf ( n86634 , n86509 );
buf ( n86635 , n86515 );
nand ( n86636 , n86634 , n86635 );
buf ( n86637 , n86636 );
buf ( n86638 , n86637 );
buf ( n86639 , n86424 );
buf ( n86640 , n86488 );
nand ( n86641 , n86639 , n86640 );
buf ( n86642 , n86641 );
buf ( n86643 , n86642 );
and ( n86644 , n86638 , n86643 );
buf ( n86645 , n86644 );
nand ( n86646 , n86633 , n86645 );
buf ( n86647 , n86518 );
not ( n86648 , n86647 );
buf ( n86649 , n86648 );
nand ( n86650 , n86646 , n86649 );
buf ( n86651 , n86650 );
nand ( n86652 , n86612 , n86651 );
buf ( n86653 , n86652 );
not ( n86654 , n86653 );
or ( n86655 , n71015 , n86654 );
not ( n86656 , n69350 );
buf ( n86657 , n69354 );
buf ( n86658 , n71008 );
nor ( n86659 , n86657 , n86658 );
buf ( n86660 , n86659 );
not ( n86661 , n86660 );
or ( n86662 , n86656 , n86661 );
buf ( n86663 , n69274 );
not ( n86664 , n86663 );
buf ( n86665 , n86664 );
buf ( n86666 , n86665 );
buf ( n86667 , n69347 );
not ( n86668 , n86667 );
buf ( n86669 , n86668 );
buf ( n86670 , n86669 );
nand ( n86671 , n86666 , n86670 );
buf ( n86672 , n86671 );
nand ( n86673 , n86662 , n86672 );
and ( n86674 , n86673 , n69270 );
nor ( n86675 , n67907 , n69269 );
nor ( n86676 , n86674 , n86675 );
nand ( n86677 , n86655 , n86676 );
not ( n86678 , n66005 );
not ( n86679 , n65910 );
and ( n86680 , n86678 , n86679 );
nor ( n86681 , n67864 , n66133 );
nor ( n86682 , n86680 , n86681 );
nand ( n86683 , n86682 , n67876 , n67871 );
not ( n86684 , n86683 );
nand ( n86685 , n86677 , n86684 , n67891 );
not ( n86686 , n67885 );
not ( n86687 , n67890 );
nand ( n86688 , n86686 , n86687 );
nand ( n86689 , n67892 , n86685 , n86688 );
nand ( n86690 , n53447 , n59133 , n63523 , n86689 );
not ( n86691 , n86690 );
buf ( n86692 , n49142 );
not ( n86693 , n86692 );
buf ( n86694 , n49684 );
not ( n86695 , n86694 );
or ( n86696 , n86693 , n86695 );
buf ( n86697 , n49684 );
buf ( n86698 , n49142 );
or ( n86699 , n86697 , n86698 );
buf ( n86700 , n49152 );
nand ( n86701 , n86699 , n86700 );
buf ( n86702 , n86701 );
buf ( n86703 , n86702 );
nand ( n86704 , n86696 , n86703 );
buf ( n86705 , n86704 );
buf ( n86706 , n86705 );
not ( n86707 , n86706 );
buf ( n86708 , n86707 );
buf ( n86709 , n86708 );
buf ( n86710 , n42312 );
not ( n86711 , n86710 );
buf ( n86712 , n42249 );
not ( n86713 , n86712 );
or ( n86714 , n86711 , n86713 );
buf ( n86715 , n49467 );
nand ( n86716 , n86714 , n86715 );
buf ( n86717 , n86716 );
buf ( n86718 , n86717 );
buf ( n86719 , n39986 );
not ( n86720 , n86719 );
buf ( n86721 , n40010 );
not ( n86722 , n86721 );
buf ( n86723 , n37268 );
not ( n86724 , n86723 );
or ( n86725 , n86722 , n86724 );
buf ( n86726 , n43142 );
buf ( n86727 , n40009 );
nand ( n86728 , n86726 , n86727 );
buf ( n86729 , n86728 );
buf ( n86730 , n86729 );
nand ( n86731 , n86725 , n86730 );
buf ( n86732 , n86731 );
buf ( n86733 , n86732 );
not ( n86734 , n86733 );
or ( n86735 , n86720 , n86734 );
buf ( n86736 , n49186 );
buf ( n86737 , n40002 );
nand ( n86738 , n86736 , n86737 );
buf ( n86739 , n86738 );
buf ( n86740 , n86739 );
nand ( n86741 , n86735 , n86740 );
buf ( n86742 , n86741 );
buf ( n86743 , n86742 );
xor ( n86744 , n86718 , n86743 );
buf ( n86745 , n42668 );
not ( n86746 , n86745 );
buf ( n86747 , n42672 );
not ( n86748 , n86747 );
buf ( n86749 , n36041 );
not ( n86750 , n86749 );
or ( n86751 , n86748 , n86750 );
buf ( n86752 , n36054 );
not ( n86753 , n86752 );
buf ( n86754 , n42671 );
nand ( n86755 , n86753 , n86754 );
buf ( n86756 , n86755 );
buf ( n86757 , n86756 );
nand ( n86758 , n86751 , n86757 );
buf ( n86759 , n86758 );
buf ( n86760 , n86759 );
not ( n86761 , n86760 );
or ( n86762 , n86746 , n86761 );
buf ( n86763 , n49366 );
buf ( n86764 , n42712 );
nand ( n86765 , n86763 , n86764 );
buf ( n86766 , n86765 );
buf ( n86767 , n86766 );
nand ( n86768 , n86762 , n86767 );
buf ( n86769 , n86768 );
buf ( n86770 , n86769 );
xor ( n86771 , n86744 , n86770 );
buf ( n86772 , n86771 );
buf ( n86773 , n86772 );
xor ( n86774 , n49357 , n49374 );
and ( n86775 , n86774 , n49446 );
and ( n86776 , n49357 , n49374 );
or ( n86777 , n86775 , n86776 );
buf ( n86778 , n86777 );
buf ( n86779 , n86778 );
xor ( n86780 , n86773 , n86779 );
xor ( n86781 , n49559 , n49570 );
and ( n86782 , n86781 , n49593 );
and ( n86783 , n49559 , n49570 );
or ( n86784 , n86782 , n86783 );
buf ( n86785 , n86784 );
buf ( n86786 , n86785 );
xor ( n86787 , n86780 , n86786 );
buf ( n86788 , n86787 );
buf ( n86789 , n86788 );
not ( n86790 , n49595 );
not ( n86791 , n49612 );
xor ( n86792 , n49670 , n49654 );
not ( n86793 , n86792 );
nand ( n86794 , n86793 , n49676 );
not ( n86795 , n49676 );
nand ( n86796 , n86795 , n86792 );
nand ( n86797 , n86791 , n86794 , n86796 );
not ( n86798 , n86797 );
or ( n86799 , n86790 , n86798 );
nand ( n86800 , n49612 , n49677 );
nand ( n86801 , n86799 , n86800 );
buf ( n86802 , n86801 );
xor ( n86803 , n86789 , n86802 );
xor ( n86804 , n49620 , n49645 );
and ( n86805 , n86804 , n49652 );
and ( n86806 , n49620 , n49645 );
or ( n86807 , n86805 , n86806 );
buf ( n86808 , n86807 );
buf ( n86809 , n86808 );
buf ( n86810 , n43909 );
not ( n86811 , n86810 );
buf ( n86812 , n25184 );
buf ( n86813 , n38436 );
and ( n86814 , n86812 , n86813 );
not ( n86815 , n86812 );
buf ( n86816 , n50871 );
and ( n86817 , n86815 , n86816 );
nor ( n86818 , n86814 , n86817 );
buf ( n86819 , n86818 );
buf ( n86820 , n86819 );
not ( n86821 , n86820 );
or ( n86822 , n86811 , n86821 );
buf ( n86823 , n49511 );
buf ( n86824 , n44586 );
nand ( n86825 , n86823 , n86824 );
buf ( n86826 , n86825 );
buf ( n86827 , n86826 );
nand ( n86828 , n86822 , n86827 );
buf ( n86829 , n86828 );
buf ( n86830 , n86829 );
xor ( n86831 , n86809 , n86830 );
xor ( n86832 , n49197 , n49203 );
and ( n86833 , n86832 , n49275 );
and ( n86834 , n49197 , n49203 );
or ( n86835 , n86833 , n86834 );
buf ( n86836 , n86835 );
buf ( n86837 , n86836 );
xor ( n86838 , n86831 , n86837 );
buf ( n86839 , n86838 );
buf ( n86840 , n86839 );
buf ( n86841 , n38758 );
not ( n86842 , n86841 );
buf ( n86843 , n45401 );
not ( n86844 , n86843 );
buf ( n86845 , n86844 );
buf ( n86846 , n86845 );
not ( n86847 , n86846 );
buf ( n86848 , n42973 );
not ( n86849 , n86848 );
or ( n86850 , n86847 , n86849 );
buf ( n86851 , n38480 );
buf ( n86852 , n38412 );
nand ( n86853 , n86851 , n86852 );
buf ( n86854 , n86853 );
buf ( n86855 , n86854 );
nand ( n86856 , n86850 , n86855 );
buf ( n86857 , n86856 );
buf ( n86858 , n86857 );
not ( n86859 , n86858 );
or ( n86860 , n86842 , n86859 );
buf ( n86861 , n49346 );
buf ( n86862 , n38775 );
nand ( n86863 , n86861 , n86862 );
buf ( n86864 , n86863 );
buf ( n86865 , n86864 );
nand ( n86866 , n86860 , n86865 );
buf ( n86867 , n86866 );
buf ( n86868 , n86867 );
buf ( n86869 , n49241 );
not ( n86870 , n86869 );
buf ( n86871 , n49218 );
not ( n86872 , n86871 );
or ( n86873 , n86870 , n86872 );
buf ( n86874 , n49269 );
nand ( n86875 , n86873 , n86874 );
buf ( n86876 , n86875 );
not ( n86877 , n49218 );
nand ( n86878 , n86877 , n49244 );
nand ( n86879 , n86876 , n86878 );
buf ( n86880 , n86879 );
xor ( n86881 , n86868 , n86880 );
buf ( n86882 , n39374 );
not ( n86883 , n86882 );
buf ( n86884 , n39000 );
not ( n86885 , n86884 );
buf ( n86886 , n39240 );
not ( n86887 , n86886 );
or ( n86888 , n86885 , n86887 );
buf ( n86889 , n37692 );
buf ( n86890 , n38997 );
nand ( n86891 , n86889 , n86890 );
buf ( n86892 , n86891 );
buf ( n86893 , n86892 );
nand ( n86894 , n86888 , n86893 );
buf ( n86895 , n86894 );
buf ( n86896 , n86895 );
not ( n86897 , n86896 );
or ( n86898 , n86883 , n86897 );
buf ( n86899 , n49637 );
buf ( n86900 , n38985 );
nand ( n86901 , n86899 , n86900 );
buf ( n86902 , n86901 );
buf ( n86903 , n86902 );
nand ( n86904 , n86898 , n86903 );
buf ( n86905 , n86904 );
buf ( n86906 , n86905 );
xor ( n86907 , n86881 , n86906 );
buf ( n86908 , n86907 );
buf ( n86909 , n86908 );
not ( n86910 , n41647 );
not ( n86911 , n36396 );
not ( n86912 , n41663 );
or ( n86913 , n86911 , n86912 );
nand ( n86914 , n41666 , n39891 );
nand ( n86915 , n86913 , n86914 );
not ( n86916 , n86915 );
or ( n86917 , n86910 , n86916 );
buf ( n86918 , n49582 );
buf ( n86919 , n41705 );
nand ( n86920 , n86918 , n86919 );
buf ( n86921 , n86920 );
nand ( n86922 , n86917 , n86921 );
buf ( n86923 , n86922 );
xor ( n86924 , n86909 , n86923 );
buf ( n86925 , n42339 );
not ( n86926 , n86925 );
and ( n86927 , n36565 , n42343 );
not ( n86928 , n36565 );
and ( n86929 , n86928 , n42350 );
or ( n86930 , n86927 , n86929 );
buf ( n86931 , n86930 );
not ( n86932 , n86931 );
or ( n86933 , n86926 , n86932 );
buf ( n86934 , n49660 );
buf ( n86935 , n42378 );
nand ( n86936 , n86934 , n86935 );
buf ( n86937 , n86936 );
buf ( n86938 , n86937 );
nand ( n86939 , n86933 , n86938 );
buf ( n86940 , n86939 );
buf ( n86941 , n86940 );
xor ( n86942 , n86924 , n86941 );
buf ( n86943 , n86942 );
buf ( n86944 , n86943 );
xor ( n86945 , n86840 , n86944 );
buf ( n86946 , n49654 );
buf ( n86947 , n86946 );
not ( n86948 , n86947 );
buf ( n86949 , n49670 );
not ( n86950 , n86949 );
or ( n86951 , n86948 , n86950 );
buf ( n86952 , n86946 );
buf ( n86953 , n49670 );
or ( n86954 , n86952 , n86953 );
buf ( n86955 , n49676 );
nand ( n86956 , n86954 , n86955 );
buf ( n86957 , n86956 );
buf ( n86958 , n86957 );
nand ( n86959 , n86951 , n86958 );
buf ( n86960 , n86959 );
buf ( n86961 , n86960 );
xor ( n86962 , n86945 , n86961 );
buf ( n86963 , n86962 );
buf ( n86964 , n86963 );
xor ( n86965 , n86803 , n86964 );
buf ( n86966 , n86965 );
not ( n86967 , n86966 );
not ( n86968 , n49158 );
nand ( n86969 , n49528 , n86968 );
not ( n86970 , n86969 );
not ( n86971 , n49683 );
or ( n86972 , n86970 , n86971 );
nand ( n86973 , n49527 , n49158 );
nand ( n86974 , n86972 , n86973 );
xor ( n86975 , n86967 , n86974 );
xor ( n86976 , n49164 , n49452 );
and ( n86977 , n86976 , n49525 );
and ( n86978 , n49164 , n49452 );
or ( n86979 , n86977 , n86978 );
buf ( n86980 , n86979 );
buf ( n86981 , n86980 );
xor ( n86982 , n49170 , n49278 );
and ( n86983 , n86982 , n49449 );
and ( n86984 , n49170 , n49278 );
or ( n86985 , n86983 , n86984 );
buf ( n86986 , n86985 );
buf ( n86987 , n86986 );
xor ( n86988 , n49459 , n49515 );
and ( n86989 , n86988 , n49522 );
and ( n86990 , n49459 , n49515 );
or ( n86991 , n86989 , n86990 );
buf ( n86992 , n86991 );
buf ( n86993 , n86992 );
xor ( n86994 , n86987 , n86993 );
buf ( n86995 , n49321 );
buf ( n86996 , n49263 );
not ( n86997 , n86996 );
buf ( n86998 , n43250 );
not ( n86999 , n86998 );
or ( n87000 , n86997 , n86999 );
buf ( n87001 , n32969 );
buf ( n87002 , n42152 );
not ( n87003 , n87002 );
buf ( n87004 , n36500 );
not ( n87005 , n87004 );
or ( n87006 , n87003 , n87005 );
buf ( n87007 , n39481 );
buf ( n87008 , n42160 );
nand ( n87009 , n87007 , n87008 );
buf ( n87010 , n87009 );
buf ( n87011 , n87010 );
nand ( n87012 , n87006 , n87011 );
buf ( n87013 , n87012 );
buf ( n87014 , n87013 );
nand ( n87015 , n87001 , n87014 );
buf ( n87016 , n87015 );
buf ( n87017 , n87016 );
nand ( n87018 , n87000 , n87017 );
buf ( n87019 , n87018 );
buf ( n87020 , n87019 );
xor ( n87021 , n86995 , n87020 );
buf ( n87022 , n49435 );
not ( n87023 , n87022 );
buf ( n87024 , n44776 );
not ( n87025 , n87024 );
or ( n87026 , n87023 , n87025 );
buf ( n87027 , n44679 );
not ( n87028 , n45370 );
not ( n87029 , n43104 );
or ( n87030 , n87028 , n87029 );
buf ( n87031 , n36929 );
buf ( n87032 , n42196 );
nand ( n87033 , n87031 , n87032 );
buf ( n87034 , n87033 );
nand ( n87035 , n87030 , n87034 );
buf ( n87036 , n87035 );
nand ( n87037 , n87027 , n87036 );
buf ( n87038 , n87037 );
buf ( n87039 , n87038 );
nand ( n87040 , n87026 , n87039 );
buf ( n87041 , n87040 );
buf ( n87042 , n87041 );
xor ( n87043 , n87021 , n87042 );
buf ( n87044 , n87043 );
buf ( n87045 , n87044 );
xor ( n87046 , n49401 , n49415 );
and ( n87047 , n87046 , n49443 );
and ( n87048 , n49401 , n49415 );
or ( n87049 , n87047 , n87048 );
buf ( n87050 , n87049 );
buf ( n87051 , n87050 );
xor ( n87052 , n87045 , n87051 );
buf ( n87053 , n38150 );
not ( n87054 , n87053 );
buf ( n87055 , n43434 );
not ( n87056 , n87055 );
buf ( n87057 , n39209 );
not ( n87058 , n87057 );
or ( n87059 , n87056 , n87058 );
buf ( n87060 , n37641 );
buf ( n87061 , n37329 );
nand ( n87062 , n87060 , n87061 );
buf ( n87063 , n87062 );
buf ( n87064 , n87063 );
nand ( n87065 , n87059 , n87064 );
buf ( n87066 , n87065 );
buf ( n87067 , n87066 );
not ( n87068 , n87067 );
or ( n87069 , n87054 , n87068 );
buf ( n87070 , n49293 );
buf ( n87071 , n37403 );
nand ( n87072 , n87070 , n87071 );
buf ( n87073 , n87072 );
buf ( n87074 , n87073 );
nand ( n87075 , n87069 , n87074 );
buf ( n87076 , n87075 );
buf ( n87077 , n87076 );
buf ( n87078 , n49395 );
not ( n87079 , n87078 );
buf ( n87080 , n87079 );
buf ( n87081 , n87080 );
not ( n87082 , n87081 );
buf ( n87083 , n38133 );
not ( n87084 , n87083 );
or ( n87085 , n87082 , n87084 );
and ( n87086 , n28306 , n43371 );
not ( n87087 , n28306 );
and ( n87088 , n87087 , n49391 );
or ( n87089 , n87086 , n87088 );
buf ( n87090 , n87089 );
buf ( n87091 , n38063 );
nand ( n87092 , n87090 , n87091 );
buf ( n87093 , n87092 );
buf ( n87094 , n87093 );
nand ( n87095 , n87085 , n87094 );
buf ( n87096 , n87095 );
buf ( n87097 , n87096 );
xor ( n87098 , n87077 , n87097 );
buf ( n87099 , n49412 );
not ( n87100 , n87099 );
buf ( n87101 , n36523 );
not ( n87102 , n87101 );
or ( n87103 , n87100 , n87102 );
buf ( n87104 , n36643 );
buf ( n87105 , n43996 );
not ( n87106 , n87105 );
buf ( n87107 , n52246 );
not ( n87108 , n87107 );
or ( n87109 , n87106 , n87108 );
buf ( n87110 , n41718 );
not ( n87111 , n87110 );
buf ( n87112 , n87111 );
buf ( n87113 , n87112 );
buf ( n87114 , n42075 );
nand ( n87115 , n87113 , n87114 );
buf ( n87116 , n87115 );
buf ( n87117 , n87116 );
nand ( n87118 , n87109 , n87117 );
buf ( n87119 , n87118 );
buf ( n87120 , n87119 );
nand ( n87121 , n87104 , n87120 );
buf ( n87122 , n87121 );
buf ( n87123 , n87122 );
nand ( n87124 , n87103 , n87123 );
buf ( n87125 , n87124 );
buf ( n87126 , n87125 );
xor ( n87127 , n87098 , n87126 );
buf ( n87128 , n87127 );
buf ( n87129 , n87128 );
xor ( n87130 , n87052 , n87129 );
buf ( n87131 , n87130 );
not ( n87132 , n42566 );
buf ( n87133 , n25160 );
not ( n87134 , n87133 );
buf ( n87135 , n39407 );
not ( n87136 , n87135 );
or ( n87137 , n87134 , n87136 );
buf ( n87138 , n52072 );
buf ( n87139 , n42581 );
nand ( n87140 , n87138 , n87139 );
buf ( n87141 , n87140 );
buf ( n87142 , n87141 );
nand ( n87143 , n87137 , n87142 );
buf ( n87144 , n87143 );
not ( n87145 , n87144 );
or ( n87146 , n87132 , n87145 );
nand ( n87147 , n49489 , n42631 );
nand ( n87148 , n87146 , n87147 );
not ( n87149 , n87148 );
xor ( n87150 , n49304 , n49325 );
and ( n87151 , n87150 , n49354 );
and ( n87152 , n49304 , n49325 );
or ( n87153 , n87151 , n87152 );
buf ( n87154 , n87153 );
not ( n87155 , n87154 );
not ( n87156 , n87155 );
or ( n87157 , n87149 , n87156 );
not ( n87158 , n87148 );
nand ( n87159 , n87154 , n87158 );
nand ( n87160 , n87157 , n87159 );
buf ( n87161 , n41976 );
not ( n87162 , n87161 );
buf ( n87163 , n38862 );
not ( n87164 , n87163 );
or ( n87165 , n87162 , n87164 );
buf ( n87166 , n38848 );
buf ( n87167 , n37472 );
nand ( n87168 , n87166 , n87167 );
buf ( n87169 , n87168 );
buf ( n87170 , n87169 );
nand ( n87171 , n87165 , n87170 );
buf ( n87172 , n87171 );
not ( n87173 , n87172 );
not ( n87174 , n44253 );
or ( n87175 , n87173 , n87174 );
nand ( n87176 , n41844 , n42434 );
or ( n87177 , n41844 , n42434 );
nand ( n87178 , n87176 , n87177 , n65307 );
nand ( n87179 , n87175 , n87178 );
not ( n87180 , n87179 );
buf ( n87181 , n49235 );
not ( n87182 , n87181 );
buf ( n87183 , n87182 );
not ( n87184 , n87183 );
not ( n87185 , n37872 );
or ( n87186 , n87184 , n87185 );
buf ( n87187 , n45617 );
buf ( n87188 , n41890 );
buf ( n87189 , n43777 );
and ( n87190 , n87188 , n87189 );
not ( n87191 , n87188 );
buf ( n87192 , n29290 );
and ( n87193 , n87191 , n87192 );
nor ( n87194 , n87190 , n87193 );
buf ( n87195 , n87194 );
buf ( n87196 , n87195 );
nand ( n87197 , n87187 , n87196 );
buf ( n87198 , n87197 );
nand ( n87199 , n87186 , n87198 );
xor ( n87200 , n87180 , n87199 );
buf ( n87201 , n42854 );
buf ( n87202 , n43108 );
buf ( n87203 , n37649 );
and ( n87204 , n87202 , n87203 );
not ( n87205 , n87202 );
buf ( n87206 , n36363 );
and ( n87207 , n87205 , n87206 );
nor ( n87208 , n87204 , n87207 );
buf ( n87209 , n87208 );
buf ( n87210 , n87209 );
or ( n87211 , n87201 , n87210 );
nand ( n87212 , C1 , n87211 );
buf ( n87213 , n87212 );
xnor ( n87214 , n87200 , n87213 );
not ( n87215 , n87214 );
xor ( n87216 , n87160 , n87215 );
or ( n87217 , n49494 , n49513 );
nand ( n87218 , n87217 , n49474 );
nand ( n87219 , n49513 , n49494 );
nand ( n87220 , n87218 , n87219 );
not ( n87221 , n87220 );
nand ( n87222 , n87216 , n87221 );
nand ( n87223 , n87131 , n87222 );
not ( n87224 , n87223 );
nor ( n87225 , n87222 , n87131 );
nor ( n87226 , n87216 , n87221 );
nor ( n87227 , n87225 , n87226 );
not ( n87228 , n87227 );
or ( n87229 , n87224 , n87228 );
not ( n87230 , n87216 );
nand ( n87231 , n87230 , n87131 , n87220 );
nand ( n87232 , n87229 , n87231 );
buf ( n87233 , n87232 );
xor ( n87234 , n86994 , n87233 );
buf ( n87235 , n87234 );
buf ( n87236 , n87235 );
xor ( n87237 , n86981 , n87236 );
xor ( n87238 , n49535 , n49541 );
and ( n87239 , n87238 , n49681 );
and ( n87240 , n49535 , n49541 );
or ( n87241 , n87239 , n87240 );
buf ( n87242 , n87241 );
buf ( n87243 , n87242 );
xor ( n87244 , n87237 , n87243 );
buf ( n87245 , n87244 );
xnor ( n87246 , n86975 , n87245 );
buf ( n87247 , n87246 );
not ( n87248 , n87247 );
buf ( n87249 , n87248 );
buf ( n87250 , n87249 );
nand ( n87251 , n86709 , n87250 );
buf ( n87252 , n87251 );
buf ( n87253 , n87252 );
xor ( n87254 , n86718 , n86743 );
and ( n87255 , n87254 , n86770 );
and ( n87256 , n86718 , n86743 );
or ( n87257 , n87255 , n87256 );
buf ( n87258 , n87257 );
buf ( n87259 , n87258 );
buf ( n87260 , n40002 );
not ( n87261 , n87260 );
buf ( n87262 , n86732 );
not ( n87263 , n87262 );
or ( n87264 , n87261 , n87263 );
buf ( n87265 , n39986 );
buf ( n87266 , n40010 );
buf ( n87267 , n38244 );
and ( n87268 , n87266 , n87267 );
not ( n87269 , n87266 );
buf ( n87270 , n43031 );
and ( n87271 , n87269 , n87270 );
nor ( n87272 , n87268 , n87271 );
buf ( n87273 , n87272 );
buf ( n87274 , n87273 );
nand ( n87275 , n87265 , n87274 );
buf ( n87276 , n87275 );
buf ( n87277 , n87276 );
nand ( n87278 , n87264 , n87277 );
buf ( n87279 , n87278 );
buf ( n87280 , n42712 );
not ( n87281 , n87280 );
buf ( n87282 , n86759 );
not ( n87283 , n87282 );
or ( n87284 , n87281 , n87283 );
not ( n87285 , n25227 );
not ( n87286 , n53159 );
or ( n87287 , n87285 , n87286 );
nand ( n87288 , n42672 , n41619 );
nand ( n87289 , n87287 , n87288 );
nand ( n87290 , n87289 , n42668 );
buf ( n87291 , n87290 );
nand ( n87292 , n87284 , n87291 );
buf ( n87293 , n87292 );
xor ( n87294 , n87279 , n87293 );
xor ( n87295 , n87077 , n87097 );
and ( n87296 , n87295 , n87126 );
and ( n87297 , n87077 , n87097 );
or ( n87298 , n87296 , n87297 );
buf ( n87299 , n87298 );
xor ( n87300 , n87294 , n87299 );
buf ( n87301 , n87300 );
xor ( n87302 , n87259 , n87301 );
buf ( n87303 , n42378 );
not ( n87304 , n87303 );
buf ( n87305 , n86930 );
not ( n87306 , n87305 );
or ( n87307 , n87304 , n87306 );
buf ( n87308 , n42350 );
buf ( n87309 , n36611 );
and ( n87310 , n87308 , n87309 );
not ( n87311 , n87308 );
buf ( n87312 , n45650 );
and ( n87313 , n87311 , n87312 );
nor ( n87314 , n87310 , n87313 );
buf ( n87315 , n87314 );
buf ( n87316 , n87315 );
not ( n87317 , n87316 );
buf ( n87318 , n42339 );
nand ( n87319 , n87317 , n87318 );
buf ( n87320 , n87319 );
buf ( n87321 , n87320 );
nand ( n87322 , n87307 , n87321 );
buf ( n87323 , n87322 );
buf ( n87324 , n87323 );
xor ( n87325 , n86868 , n86880 );
and ( n87326 , n87325 , n86906 );
and ( n87327 , n86868 , n86880 );
or ( n87328 , n87326 , n87327 );
buf ( n87329 , n87328 );
buf ( n87330 , n87329 );
xor ( n87331 , n87324 , n87330 );
buf ( n87332 , n44586 );
not ( n87333 , n87332 );
buf ( n87334 , n86819 );
not ( n87335 , n87334 );
or ( n87336 , n87333 , n87335 );
buf ( n87337 , n25184 );
not ( n87338 , n87337 );
buf ( n87339 , n38098 );
not ( n87340 , n87339 );
or ( n87341 , n87338 , n87340 );
nand ( n87342 , n40089 , n25183 );
buf ( n87343 , n87342 );
nand ( n87344 , n87341 , n87343 );
buf ( n87345 , n87344 );
buf ( n87346 , n87345 );
buf ( n87347 , n43909 );
nand ( n87348 , n87346 , n87347 );
buf ( n87349 , n87348 );
buf ( n87350 , n87349 );
nand ( n87351 , n87336 , n87350 );
buf ( n87352 , n87351 );
buf ( n87353 , n87352 );
xnor ( n87354 , n87331 , n87353 );
buf ( n87355 , n87354 );
buf ( n87356 , n87355 );
xnor ( n87357 , n87302 , n87356 );
buf ( n87358 , n87357 );
buf ( n87359 , n87358 );
xor ( n87360 , n86840 , n86944 );
and ( n87361 , n87360 , n86961 );
and ( n87362 , n86840 , n86944 );
or ( n87363 , n87361 , n87362 );
buf ( n87364 , n87363 );
buf ( n87365 , n87364 );
xor ( n87366 , n87359 , n87365 );
xor ( n87367 , n86909 , n86923 );
and ( n87368 , n87367 , n86941 );
and ( n87369 , n86909 , n86923 );
or ( n87370 , n87368 , n87369 );
buf ( n87371 , n87370 );
buf ( n87372 , n87371 );
not ( n87373 , n87372 );
buf ( n87374 , n87373 );
xor ( n87375 , n86809 , n86830 );
and ( n87376 , n87375 , n86837 );
and ( n87377 , n86809 , n86830 );
or ( n87378 , n87376 , n87377 );
buf ( n87379 , n87378 );
not ( n87380 , n87379 );
and ( n87381 , n87374 , n87380 );
not ( n87382 , n87374 );
and ( n87383 , n87382 , n87379 );
or ( n87384 , n87381 , n87383 );
buf ( n87385 , n87148 );
not ( n87386 , n87385 );
buf ( n87387 , n87214 );
not ( n87388 , n87387 );
or ( n87389 , n87386 , n87388 );
not ( n87390 , n87158 );
not ( n87391 , n87215 );
or ( n87392 , n87390 , n87391 );
nand ( n87393 , n87392 , n87154 );
buf ( n87394 , n87393 );
nand ( n87395 , n87389 , n87394 );
buf ( n87396 , n87395 );
not ( n87397 , n41705 );
not ( n87398 , n86915 );
or ( n87399 , n87397 , n87398 );
xor ( n87400 , n41666 , n36427 );
nand ( n87401 , n87400 , n41647 );
nand ( n87402 , n87399 , n87401 );
not ( n87403 , n87402 );
buf ( n87404 , n87119 );
not ( n87405 , n87404 );
buf ( n87406 , n50374 );
not ( n87407 , n87406 );
or ( n87408 , n87405 , n87407 );
buf ( n87409 , n36643 );
buf ( n87410 , n43368 );
not ( n87411 , n87410 );
buf ( n87412 , n52246 );
not ( n87413 , n87412 );
or ( n87414 , n87411 , n87413 );
buf ( n87415 , n39729 );
buf ( n87416 , n43365 );
nand ( n87417 , n87415 , n87416 );
buf ( n87418 , n87417 );
buf ( n87419 , n87418 );
nand ( n87420 , n87414 , n87419 );
buf ( n87421 , n87420 );
buf ( n87422 , n87421 );
nand ( n87423 , n87409 , n87422 );
buf ( n87424 , n87423 );
buf ( n87425 , n87424 );
nand ( n87426 , n87408 , n87425 );
buf ( n87427 , n87426 );
buf ( n87428 , n87427 );
buf ( n87429 , n87035 );
not ( n87430 , n87429 );
buf ( n87431 , n44670 );
not ( n87432 , n87431 );
buf ( n87433 , n87432 );
buf ( n87434 , n87433 );
not ( n87435 , n87434 );
or ( n87436 , n87430 , n87435 );
buf ( n87437 , n36929 );
not ( n87438 , n87437 );
buf ( n87439 , n41951 );
not ( n87440 , n87439 );
and ( n87441 , n87438 , n87440 );
buf ( n87442 , n43095 );
buf ( n87443 , n41951 );
and ( n87444 , n87442 , n87443 );
nor ( n87445 , n87441 , n87444 );
buf ( n87446 , n87445 );
buf ( n87447 , n87446 );
not ( n87448 , n87447 );
buf ( n87449 , n36912 );
nand ( n87450 , n87448 , n87449 );
buf ( n87451 , n87450 );
buf ( n87452 , n87451 );
nand ( n87453 , n87436 , n87452 );
buf ( n87454 , n87453 );
buf ( n87455 , n87454 );
xor ( n87456 , n87428 , n87455 );
buf ( n87457 , n87180 );
not ( n87458 , n87457 );
not ( n87459 , n87199 );
buf ( n87460 , n87459 );
not ( n87461 , n87460 );
or ( n87462 , n87458 , n87461 );
buf ( n87463 , n87213 );
nand ( n87464 , n87462 , n87463 );
buf ( n87465 , n87464 );
buf ( n87466 , n87465 );
buf ( n87467 , n87199 );
buf ( n87468 , n87179 );
nand ( n87469 , n87467 , n87468 );
buf ( n87470 , n87469 );
buf ( n87471 , n87470 );
nand ( n87472 , n87466 , n87471 );
buf ( n87473 , n87472 );
buf ( n87474 , n87473 );
xor ( n87475 , n87456 , n87474 );
buf ( n87476 , n87475 );
not ( n87477 , n87476 );
xor ( n87478 , n87403 , n87477 );
xnor ( n87479 , n87396 , n87478 );
buf ( n87480 , n87479 );
and ( n87481 , n87384 , n87480 );
not ( n87482 , n87384 );
not ( n87483 , n87480 );
and ( n87484 , n87482 , n87483 );
nor ( n87485 , n87481 , n87484 );
buf ( n87486 , n87485 );
xor ( n87487 , n87366 , n87486 );
buf ( n87488 , n87487 );
xor ( n87489 , n86981 , n87236 );
and ( n87490 , n87489 , n87243 );
and ( n87491 , n86981 , n87236 );
or ( n87492 , n87490 , n87491 );
buf ( n87493 , n87492 );
xor ( n87494 , n87488 , n87493 );
not ( n87495 , n87222 );
not ( n87496 , n87131 );
or ( n87497 , n87495 , n87496 );
not ( n87498 , n87226 );
nand ( n87499 , n87497 , n87498 );
buf ( n87500 , n87499 );
xor ( n87501 , n86773 , n86779 );
and ( n87502 , n87501 , n86786 );
and ( n87503 , n86773 , n86779 );
or ( n87504 , n87502 , n87503 );
buf ( n87505 , n87504 );
buf ( n87506 , n87505 );
xor ( n87507 , n87500 , n87506 );
buf ( n87508 , n38775 );
not ( n87509 , n87508 );
buf ( n87510 , n86857 );
not ( n87511 , n87510 );
or ( n87512 , n87509 , n87511 );
buf ( n87513 , n86845 );
not ( n87514 , n87513 );
buf ( n87515 , n37745 );
not ( n87516 , n87515 );
or ( n87517 , n87514 , n87516 );
buf ( n87518 , n43198 );
buf ( n87519 , n38412 );
nand ( n87520 , n87518 , n87519 );
buf ( n87521 , n87520 );
buf ( n87522 , n87521 );
nand ( n87523 , n87517 , n87522 );
buf ( n87524 , n87523 );
buf ( n87525 , n87524 );
buf ( n87526 , n38758 );
nand ( n87527 , n87525 , n87526 );
buf ( n87528 , n87527 );
buf ( n87529 , n87528 );
nand ( n87530 , n87512 , n87529 );
buf ( n87531 , n87530 );
buf ( n87532 , n87531 );
buf ( n87533 , n38985 );
not ( n87534 , n87533 );
buf ( n87535 , n86895 );
not ( n87536 , n87535 );
or ( n87537 , n87534 , n87536 );
buf ( n87538 , n39000 );
not ( n87539 , n87538 );
buf ( n87540 , n49178 );
not ( n87541 , n87540 );
or ( n87542 , n87539 , n87541 );
buf ( n87543 , n69992 );
buf ( n87544 , n38997 );
nand ( n87545 , n87543 , n87544 );
buf ( n87546 , n87545 );
buf ( n87547 , n87546 );
nand ( n87548 , n87542 , n87547 );
buf ( n87549 , n87548 );
buf ( n87550 , n87549 );
buf ( n87551 , n42448 );
nand ( n87552 , n87550 , n87551 );
buf ( n87553 , n87552 );
buf ( n87554 , n87553 );
nand ( n87555 , n87537 , n87554 );
buf ( n87556 , n87555 );
buf ( n87557 , n87556 );
xor ( n87558 , n87532 , n87557 );
xor ( n87559 , n86995 , n87020 );
and ( n87560 , n87559 , n87042 );
and ( n87561 , n86995 , n87020 );
or ( n87562 , n87560 , n87561 );
buf ( n87563 , n87562 );
buf ( n87564 , n87563 );
xor ( n87565 , n87558 , n87564 );
buf ( n87566 , n87565 );
buf ( n87567 , n87566 );
xor ( n87568 , n87045 , n87051 );
and ( n87569 , n87568 , n87129 );
and ( n87570 , n87045 , n87051 );
or ( n87571 , n87569 , n87570 );
buf ( n87572 , n87571 );
buf ( n87573 , n87572 );
xor ( n87574 , n87567 , n87573 );
buf ( n87575 , n38150 );
not ( n87576 , n87575 );
buf ( n87577 , n43434 );
not ( n87578 , n87577 );
buf ( n87579 , n49336 );
not ( n87580 , n87579 );
or ( n87581 , n87578 , n87580 );
buf ( n87582 , n44163 );
buf ( n87583 , n37329 );
nand ( n87584 , n87582 , n87583 );
buf ( n87585 , n87584 );
buf ( n87586 , n87585 );
nand ( n87587 , n87581 , n87586 );
buf ( n87588 , n87587 );
buf ( n87589 , n87588 );
not ( n87590 , n87589 );
or ( n87591 , n87576 , n87590 );
buf ( n87592 , n87066 );
buf ( n87593 , n37403 );
nand ( n87594 , n87592 , n87593 );
buf ( n87595 , n87594 );
buf ( n87596 , n87595 );
nand ( n87597 , n87591 , n87596 );
buf ( n87598 , n87597 );
and ( n87599 , n87089 , n43389 );
buf ( n87600 , n41762 );
not ( n87601 , n87600 );
buf ( n87602 , n43371 );
not ( n87603 , n87602 );
or ( n87604 , n87601 , n87603 );
buf ( n87605 , n38108 );
buf ( n87606 , n41975 );
nand ( n87607 , n87605 , n87606 );
buf ( n87608 , n87607 );
buf ( n87609 , n87608 );
nand ( n87610 , n87604 , n87609 );
buf ( n87611 , n87610 );
and ( n87612 , n87611 , n38060 );
nor ( n87613 , n87599 , n87612 );
xor ( n87614 , n87598 , n87613 );
not ( n87615 , n41905 );
not ( n87616 , n41894 );
not ( n87617 , n74977 );
or ( n87618 , n87616 , n87617 );
nand ( n87619 , n39671 , n41895 );
nand ( n87620 , n87618 , n87619 );
not ( n87621 , n87620 );
or ( n87622 , n87615 , n87621 );
nand ( n87623 , n87195 , n41862 );
nand ( n87624 , n87622 , n87623 );
buf ( n87625 , n87624 );
not ( n87626 , n87625 );
buf ( n87627 , n87626 );
and ( n87628 , n87614 , n87627 );
not ( n87629 , n87614 );
and ( n87630 , n87629 , n87624 );
nor ( n87631 , n87628 , n87630 );
buf ( n87632 , n87172 );
not ( n87633 , n87632 );
buf ( n87634 , n43766 );
not ( n87635 , n87634 );
or ( n87636 , n87633 , n87635 );
buf ( n87637 , n41976 );
not ( n87638 , n87637 );
buf ( n87639 , n42899 );
not ( n87640 , n87639 );
or ( n87641 , n87638 , n87640 );
buf ( n87642 , n42458 );
buf ( n87643 , n43780 );
nand ( n87644 , n87642 , n87643 );
buf ( n87645 , n87644 );
buf ( n87646 , n87645 );
nand ( n87647 , n87641 , n87646 );
buf ( n87648 , n87647 );
buf ( n87649 , n87648 );
buf ( n87650 , n41852 );
nand ( n87651 , n87649 , n87650 );
buf ( n87652 , n87651 );
buf ( n87653 , n87652 );
nand ( n87654 , n87636 , n87653 );
buf ( n87655 , n87654 );
buf ( n87656 , n87655 );
buf ( n87657 , n42055 );
not ( n87658 , n87657 );
buf ( n87659 , n37649 );
not ( n87660 , n87659 );
or ( n87661 , n87658 , n87660 );
buf ( n87662 , n38834 );
buf ( n87663 , n42052 );
nand ( n87664 , n87662 , n87663 );
buf ( n87665 , n87664 );
buf ( n87666 , n87665 );
nand ( n87667 , n87661 , n87666 );
buf ( n87668 , n87667 );
buf ( n87669 , n87668 );
not ( n87670 , n87669 );
buf ( n87671 , n87670 );
buf ( n87672 , n87671 );
buf ( n87673 , n42854 );
or ( n87674 , n87672 , n87673 );
nand ( n87675 , C1 , n87674 );
buf ( n87676 , n87675 );
buf ( n87677 , n87676 );
xor ( n87678 , n87656 , n87677 );
buf ( n87679 , n45288 );
not ( n87680 , n87679 );
buf ( n87681 , n87680 );
buf ( n87682 , n87681 );
buf ( n87683 , n87013 );
not ( n87684 , n87683 );
buf ( n87685 , n87684 );
buf ( n87686 , n87685 );
or ( n87687 , n87682 , n87686 );
buf ( n87688 , n42530 );
not ( n87689 , n87688 );
buf ( n87690 , n87689 );
buf ( n87691 , n87690 );
buf ( n87692 , n41882 );
not ( n87693 , n87692 );
buf ( n87694 , n39493 );
not ( n87695 , n87694 );
or ( n87696 , n87693 , n87695 );
buf ( n87697 , n51030 );
buf ( n87698 , n41879 );
nand ( n87699 , n87697 , n87698 );
buf ( n87700 , n87699 );
buf ( n87701 , n87700 );
nand ( n87702 , n87696 , n87701 );
buf ( n87703 , n87702 );
buf ( n87704 , n87703 );
not ( n87705 , n87704 );
buf ( n87706 , n87705 );
buf ( n87707 , n87706 );
or ( n87708 , n87691 , n87707 );
nand ( n87709 , n87687 , n87708 );
buf ( n87710 , n87709 );
buf ( n87711 , n87710 );
xor ( n87712 , n87678 , n87711 );
buf ( n87713 , n87712 );
buf ( n87714 , n87713 );
buf ( n87715 , n42566 );
not ( n87716 , n87715 );
buf ( n87717 , n25160 );
not ( n87718 , n87717 );
buf ( n87719 , n37971 );
not ( n87720 , n87719 );
or ( n87721 , n87718 , n87720 );
buf ( n87722 , n38447 );
buf ( n87723 , n42581 );
nand ( n87724 , n87722 , n87723 );
buf ( n87725 , n87724 );
buf ( n87726 , n87725 );
nand ( n87727 , n87721 , n87726 );
buf ( n87728 , n87727 );
buf ( n87729 , n87728 );
not ( n87730 , n87729 );
or ( n87731 , n87716 , n87730 );
buf ( n87732 , n87144 );
buf ( n87733 , n42631 );
nand ( n87734 , n87732 , n87733 );
buf ( n87735 , n87734 );
buf ( n87736 , n87735 );
nand ( n87737 , n87731 , n87736 );
buf ( n87738 , n87737 );
buf ( n87739 , n87738 );
xor ( n87740 , n87714 , n87739 );
buf ( n87741 , n87740 );
xor ( n87742 , n87631 , n87741 );
buf ( n87743 , n87742 );
not ( n87744 , n87743 );
buf ( n87745 , n87744 );
buf ( n87746 , n87745 );
xor ( n87747 , n87574 , n87746 );
buf ( n87748 , n87747 );
buf ( n87749 , n87748 );
xor ( n87750 , n87507 , n87749 );
buf ( n87751 , n87750 );
buf ( n87752 , n87751 );
xor ( n87753 , n86987 , n86993 );
and ( n87754 , n87753 , n87233 );
and ( n87755 , n86987 , n86993 );
or ( n87756 , n87754 , n87755 );
buf ( n87757 , n87756 );
buf ( n87758 , n87757 );
xor ( n87759 , n87752 , n87758 );
xor ( n87760 , n86789 , n86802 );
and ( n87761 , n87760 , n86964 );
and ( n87762 , n86789 , n86802 );
or ( n87763 , n87761 , n87762 );
buf ( n87764 , n87763 );
buf ( n87765 , n87764 );
xor ( n87766 , n87759 , n87765 );
buf ( n87767 , n87766 );
xnor ( n87768 , n87494 , n87767 );
not ( n87769 , n87245 );
nand ( n87770 , n87769 , n86967 );
buf ( n87771 , n86974 );
and ( n87772 , n87770 , n87771 );
not ( n87773 , n87245 );
nor ( n87774 , n87773 , n86967 );
nor ( n87775 , n87772 , n87774 );
nand ( n87776 , n87768 , n87775 );
buf ( n87777 , n87776 );
and ( n87778 , n87253 , n87777 );
buf ( n87779 , n87778 );
not ( n87780 , n87488 );
not ( n87781 , n87780 );
not ( n87782 , n87493 );
not ( n87783 , n87782 );
or ( n87784 , n87781 , n87783 );
nand ( n87785 , n87784 , n87767 );
nand ( n87786 , n87488 , n87493 );
nand ( n87787 , n87785 , n87786 );
xor ( n87788 , n87279 , n87293 );
and ( n87789 , n87788 , n87299 );
and ( n87790 , n87279 , n87293 );
or ( n87791 , n87789 , n87790 );
buf ( n87792 , n42668 );
not ( n87793 , n87792 );
buf ( n87794 , n87793 );
not ( n87795 , n87794 );
not ( n87796 , n42711 );
or ( n87797 , n87795 , n87796 );
nand ( n87798 , n87797 , n87289 );
not ( n87799 , n87315 );
not ( n87800 , n42375 );
and ( n87801 , n87799 , n87800 );
buf ( n87802 , n42343 );
not ( n87803 , n87802 );
buf ( n87804 , n36054 );
not ( n87805 , n87804 );
or ( n87806 , n87803 , n87805 );
buf ( n87807 , n52444 );
buf ( n87808 , n42350 );
nand ( n87809 , n87807 , n87808 );
buf ( n87810 , n87809 );
buf ( n87811 , n87810 );
nand ( n87812 , n87806 , n87811 );
buf ( n87813 , n87812 );
and ( n87814 , n87813 , n42339 );
nor ( n87815 , n87801 , n87814 );
and ( n87816 , n87798 , n87815 );
not ( n87817 , n87798 );
buf ( n87818 , n87815 );
not ( n87819 , n87818 );
buf ( n87820 , n87819 );
and ( n87821 , n87817 , n87820 );
or ( n87822 , n87816 , n87821 );
not ( n87823 , n39374 );
not ( n87824 , n39000 );
not ( n87825 , n37268 );
or ( n87826 , n87824 , n87825 );
buf ( n87827 , n43142 );
buf ( n87828 , n38997 );
nand ( n87829 , n87827 , n87828 );
buf ( n87830 , n87829 );
nand ( n87831 , n87826 , n87830 );
not ( n87832 , n87831 );
or ( n87833 , n87823 , n87832 );
not ( n87834 , n38988 );
nand ( n87835 , n87834 , n87549 );
nand ( n87836 , n87833 , n87835 );
and ( n87837 , n87822 , n87836 );
not ( n87838 , n87822 );
not ( n87839 , n87836 );
and ( n87840 , n87838 , n87839 );
nor ( n87841 , n87837 , n87840 );
xor ( n87842 , n87791 , n87841 );
not ( n87843 , n87352 );
not ( n87844 , n87323 );
or ( n87845 , n87843 , n87844 );
or ( n87846 , n87323 , n87352 );
nand ( n87847 , n87846 , n87329 );
nand ( n87848 , n87845 , n87847 );
xor ( n87849 , n87842 , n87848 );
buf ( n87850 , n87849 );
not ( n87851 , n87374 );
not ( n87852 , n87479 );
or ( n87853 , n87851 , n87852 );
nand ( n87854 , n87853 , n87379 );
buf ( n87855 , n87854 );
not ( n87856 , n87479 );
nand ( n87857 , n87856 , n87371 );
buf ( n87858 , n87857 );
nand ( n87859 , n87855 , n87858 );
buf ( n87860 , n87859 );
buf ( n87861 , n87860 );
xor ( n87862 , n87850 , n87861 );
xor ( n87863 , n87428 , n87455 );
and ( n87864 , n87863 , n87474 );
and ( n87865 , n87428 , n87455 );
or ( n87866 , n87864 , n87865 );
buf ( n87867 , n87866 );
buf ( n87868 , n87867 );
buf ( n87869 , n42566 );
not ( n87870 , n87869 );
buf ( n87871 , n25160 );
not ( n87872 , n87871 );
buf ( n87873 , n38435 );
not ( n87874 , n87873 );
or ( n87875 , n87872 , n87874 );
buf ( n87876 , n38436 );
buf ( n87877 , n42581 );
nand ( n87878 , n87876 , n87877 );
buf ( n87879 , n87878 );
buf ( n87880 , n87879 );
nand ( n87881 , n87875 , n87880 );
buf ( n87882 , n87881 );
buf ( n87883 , n87882 );
not ( n87884 , n87883 );
or ( n87885 , n87870 , n87884 );
buf ( n87886 , n87728 );
buf ( n87887 , n42631 );
nand ( n87888 , n87886 , n87887 );
buf ( n87889 , n87888 );
buf ( n87890 , n87889 );
nand ( n87891 , n87885 , n87890 );
buf ( n87892 , n87891 );
buf ( n87893 , n87892 );
xor ( n87894 , n87868 , n87893 );
buf ( n87895 , n87421 );
not ( n87896 , n87895 );
buf ( n87897 , n36523 );
not ( n87898 , n87897 );
or ( n87899 , n87896 , n87898 );
buf ( n87900 , n44141 );
buf ( n87901 , n42152 );
not ( n87902 , n87901 );
buf ( n87903 , n52246 );
not ( n87904 , n87903 );
or ( n87905 , n87902 , n87904 );
buf ( n87906 , n87112 );
buf ( n87907 , n42160 );
nand ( n87908 , n87906 , n87907 );
buf ( n87909 , n87908 );
buf ( n87910 , n87909 );
nand ( n87911 , n87905 , n87910 );
buf ( n87912 , n87911 );
buf ( n87913 , n87912 );
nand ( n87914 , n87900 , n87913 );
buf ( n87915 , n87914 );
buf ( n87916 , n87915 );
nand ( n87917 , n87899 , n87916 );
buf ( n87918 , n87917 );
buf ( n87919 , n87611 );
not ( n87920 , n87919 );
buf ( n87921 , n38133 );
not ( n87922 , n87921 );
or ( n87923 , n87920 , n87922 );
buf ( n87924 , n43777 );
buf ( n87925 , n44004 );
and ( n87926 , n87924 , n87925 );
not ( n87927 , n87924 );
buf ( n87928 , n44635 );
and ( n87929 , n87927 , n87928 );
nor ( n87930 , n87926 , n87929 );
buf ( n87931 , n87930 );
buf ( n87932 , n87931 );
not ( n87933 , n87932 );
buf ( n87934 , n43414 );
nand ( n87935 , n87933 , n87934 );
buf ( n87936 , n87935 );
buf ( n87937 , n87936 );
nand ( n87938 , n87923 , n87937 );
buf ( n87939 , n87938 );
not ( n87940 , n87939 );
xor ( n87941 , n87918 , n87940 );
buf ( n87942 , n38758 );
not ( n87943 , n87942 );
buf ( n87944 , n38413 );
not ( n87945 , n87944 );
buf ( n87946 , n39240 );
not ( n87947 , n87946 );
or ( n87948 , n87945 , n87947 );
buf ( n87949 , n37692 );
buf ( n87950 , n45401 );
nand ( n87951 , n87949 , n87950 );
buf ( n87952 , n87951 );
buf ( n87953 , n87952 );
nand ( n87954 , n87948 , n87953 );
buf ( n87955 , n87954 );
buf ( n87956 , n87955 );
not ( n87957 , n87956 );
or ( n87958 , n87943 , n87957 );
buf ( n87959 , n87524 );
buf ( n87960 , n38775 );
nand ( n87961 , n87959 , n87960 );
buf ( n87962 , n87961 );
buf ( n87963 , n87962 );
nand ( n87964 , n87958 , n87963 );
buf ( n87965 , n87964 );
xnor ( n87966 , n87941 , n87965 );
buf ( n87967 , n87966 );
xor ( n87968 , n87894 , n87967 );
buf ( n87969 , n87968 );
buf ( n87970 , n87969 );
xor ( n87971 , n87532 , n87557 );
and ( n87972 , n87971 , n87564 );
and ( n87973 , n87532 , n87557 );
or ( n87974 , n87972 , n87973 );
buf ( n87975 , n87974 );
not ( n87976 , n87975 );
not ( n87977 , n87976 );
buf ( n87978 , n43909 );
not ( n87979 , n87978 );
and ( n87980 , n36396 , n25183 );
not ( n87981 , n36396 );
and ( n87982 , n87981 , n25184 );
or ( n87983 , n87980 , n87982 );
buf ( n87984 , n87983 );
not ( n87985 , n87984 );
or ( n87986 , n87979 , n87985 );
buf ( n87987 , n87345 );
buf ( n87988 , n44586 );
nand ( n87989 , n87987 , n87988 );
buf ( n87990 , n87989 );
buf ( n87991 , n87990 );
nand ( n87992 , n87986 , n87991 );
buf ( n87993 , n87992 );
not ( n87994 , n87993 );
or ( n87995 , n87977 , n87994 );
not ( n87996 , n87993 );
nand ( n87997 , n87996 , n87975 );
nand ( n87998 , n87995 , n87997 );
buf ( n87999 , n41705 );
not ( n88000 , n87999 );
buf ( n88001 , n87400 );
not ( n88002 , n88001 );
or ( n88003 , n88000 , n88002 );
not ( n88004 , n41666 );
not ( n88005 , n39930 );
or ( n88006 , n88004 , n88005 );
not ( n88007 , n42277 );
nand ( n88008 , n88007 , n41663 );
nand ( n88009 , n88006 , n88008 );
buf ( n88010 , n88009 );
buf ( n88011 , n41647 );
nand ( n88012 , n88010 , n88011 );
buf ( n88013 , n88012 );
buf ( n88014 , n88013 );
nand ( n88015 , n88003 , n88014 );
buf ( n88016 , n88015 );
and ( n88017 , n87998 , n88016 );
not ( n88018 , n87998 );
not ( n88019 , n88016 );
and ( n88020 , n88018 , n88019 );
nor ( n88021 , n88017 , n88020 );
buf ( n88022 , n88021 );
xor ( n88023 , n87970 , n88022 );
not ( n88024 , n87402 );
not ( n88025 , n87476 );
or ( n88026 , n88024 , n88025 );
not ( n88027 , n87396 );
and ( n88028 , n87403 , n87477 );
or ( n88029 , n88027 , n88028 );
nand ( n88030 , n88026 , n88029 );
buf ( n88031 , n88030 );
xor ( n88032 , n88023 , n88031 );
buf ( n88033 , n88032 );
buf ( n88034 , n88033 );
xor ( n88035 , n87862 , n88034 );
buf ( n88036 , n88035 );
xor ( n88037 , n87752 , n87758 );
and ( n88038 , n88037 , n87765 );
and ( n88039 , n87752 , n87758 );
or ( n88040 , n88038 , n88039 );
buf ( n88041 , n88040 );
xor ( n88042 , n88036 , n88041 );
xor ( n88043 , n87500 , n87506 );
and ( n88044 , n88043 , n87749 );
and ( n88045 , n87500 , n87506 );
or ( n88046 , n88044 , n88045 );
buf ( n88047 , n88046 );
not ( n88048 , n88047 );
buf ( n88049 , n87566 );
not ( n88050 , n88049 );
buf ( n88051 , n88050 );
buf ( n88052 , n88051 );
not ( n88053 , n88052 );
buf ( n88054 , n87742 );
not ( n88055 , n88054 );
or ( n88056 , n88053 , n88055 );
buf ( n88057 , n87572 );
nand ( n88058 , n88056 , n88057 );
buf ( n88059 , n88058 );
buf ( n88060 , n88059 );
buf ( n88061 , n87745 );
buf ( n88062 , n87566 );
nand ( n88063 , n88061 , n88062 );
buf ( n88064 , n88063 );
buf ( n88065 , n88064 );
nand ( n88066 , n88060 , n88065 );
buf ( n88067 , n88066 );
buf ( n88068 , n88067 );
buf ( n88069 , n87355 );
buf ( n88070 , n87300 );
buf ( n88071 , n87258 );
nor ( n88072 , n88070 , n88071 );
buf ( n88073 , n88072 );
buf ( n88074 , n88073 );
or ( n88075 , n88069 , n88074 );
buf ( n88076 , n87300 );
buf ( n88077 , n87258 );
nand ( n88078 , n88076 , n88077 );
buf ( n88079 , n88078 );
buf ( n88080 , n88079 );
nand ( n88081 , n88075 , n88080 );
buf ( n88082 , n88081 );
buf ( n88083 , n88082 );
xor ( n88084 , n88068 , n88083 );
buf ( n88085 , n38150 );
not ( n88086 , n88085 );
buf ( n88087 , n37329 );
not ( n88088 , n88087 );
buf ( n88089 , n88088 );
buf ( n88090 , n88089 );
not ( n88091 , n88090 );
buf ( n88092 , n43678 );
not ( n88093 , n88092 );
or ( n88094 , n88091 , n88093 );
buf ( n88095 , n38480 );
buf ( n88096 , n37329 );
nand ( n88097 , n88095 , n88096 );
buf ( n88098 , n88097 );
buf ( n88099 , n88098 );
nand ( n88100 , n88094 , n88099 );
buf ( n88101 , n88100 );
buf ( n88102 , n88101 );
not ( n88103 , n88102 );
or ( n88104 , n88086 , n88103 );
buf ( n88105 , n87588 );
buf ( n88106 , n37403 );
nand ( n88107 , n88105 , n88106 );
buf ( n88108 , n88107 );
buf ( n88109 , n88108 );
nand ( n88110 , n88104 , n88109 );
buf ( n88111 , n88110 );
xor ( n88112 , n87656 , n87677 );
and ( n88113 , n88112 , n87711 );
and ( n88114 , n87656 , n87677 );
or ( n88115 , n88113 , n88114 );
buf ( n88116 , n88115 );
xor ( n88117 , n88111 , n88116 );
not ( n88118 , n87598 );
not ( n88119 , n87627 );
or ( n88120 , n88118 , n88119 );
buf ( n88121 , n87598 );
buf ( n88122 , n87627 );
nor ( n88123 , n88121 , n88122 );
buf ( n88124 , n88123 );
or ( n88125 , n88124 , n87613 );
nand ( n88126 , n88120 , n88125 );
xor ( n88127 , n88117 , n88126 );
buf ( n88128 , n87631 );
not ( n88129 , n88128 );
buf ( n88130 , n88129 );
not ( n88131 , n88130 );
buf ( n88132 , n87713 );
buf ( n88133 , n87738 );
or ( n88134 , n88132 , n88133 );
buf ( n88135 , n88134 );
not ( n88136 , n88135 );
or ( n88137 , n88131 , n88136 );
and ( n88138 , n87714 , n87739 );
buf ( n88139 , n88138 );
not ( n88140 , n88139 );
nand ( n88141 , n88137 , n88140 );
xor ( n88142 , n88127 , n88141 );
buf ( n88143 , n41844 );
buf ( n88144 , n88143 );
not ( n88145 , n88144 );
buf ( n88146 , n42891 );
not ( n88147 , n88146 );
or ( n88148 , n88145 , n88147 );
buf ( n88149 , n39205 );
buf ( n88150 , n41839 );
nand ( n88151 , n88149 , n88150 );
buf ( n88152 , n88151 );
buf ( n88153 , n88152 );
nand ( n88154 , n88148 , n88153 );
buf ( n88155 , n88154 );
buf ( n88156 , n88155 );
buf ( n88157 , n37452 );
and ( n88158 , n88156 , n88157 );
buf ( n88159 , n41966 );
buf ( n88160 , n87648 );
and ( n88161 , n88159 , n88160 );
buf ( n88162 , n88161 );
buf ( n88163 , n88162 );
nor ( n88164 , n88158 , n88163 );
buf ( n88165 , n88164 );
buf ( n88166 , n88165 );
not ( n88167 , n88166 );
buf ( n88168 , n88167 );
xor ( n88169 , n87627 , n88168 );
buf ( n88170 , n44670 );
buf ( n88171 , n87446 );
or ( n88172 , n88170 , n88171 );
buf ( n88173 , n44682 );
buf ( n88174 , n28306 );
buf ( n88175 , n43104 );
and ( n88176 , n88174 , n88175 );
not ( n88177 , n88174 );
buf ( n88178 , n42062 );
and ( n88179 , n88177 , n88178 );
nor ( n88180 , n88176 , n88179 );
buf ( n88181 , n88180 );
buf ( n88182 , n88181 );
or ( n88183 , n88173 , n88182 );
nand ( n88184 , n88172 , n88183 );
buf ( n88185 , n88184 );
not ( n88186 , n88185 );
xnor ( n88187 , n88169 , n88186 );
not ( n88188 , n88187 );
not ( n88189 , n39986 );
buf ( n88190 , n40010 );
not ( n88191 , n88190 );
buf ( n88192 , n38218 );
not ( n88193 , n88192 );
or ( n88194 , n88191 , n88193 );
buf ( n88195 , n47969 );
buf ( n88196 , n40009 );
nand ( n88197 , n88195 , n88196 );
buf ( n88198 , n88197 );
buf ( n88199 , n88198 );
nand ( n88200 , n88194 , n88199 );
buf ( n88201 , n88200 );
not ( n88202 , n88201 );
or ( n88203 , n88189 , n88202 );
buf ( n88204 , n87273 );
buf ( n88205 , n40002 );
nand ( n88206 , n88204 , n88205 );
buf ( n88207 , n88206 );
nand ( n88208 , n88203 , n88207 );
not ( n88209 , n88208 );
not ( n88210 , n88209 );
buf ( n88211 , n87703 );
not ( n88212 , n88211 );
buf ( n88213 , n45288 );
not ( n88214 , n88213 );
or ( n88215 , n88212 , n88214 );
not ( n88216 , n45370 );
not ( n88217 , n36500 );
or ( n88218 , n88216 , n88217 );
buf ( n88219 , n43265 );
buf ( n88220 , n42196 );
nand ( n88221 , n88219 , n88220 );
buf ( n88222 , n88221 );
nand ( n88223 , n88218 , n88222 );
nand ( n88224 , n32969 , n88223 );
buf ( n88225 , n88224 );
nand ( n88226 , n88215 , n88225 );
buf ( n88227 , n88226 );
not ( n88228 , n41862 );
not ( n88229 , n87620 );
or ( n88230 , n88228 , n88229 );
not ( n88231 , n38848 );
not ( n88232 , n41894 );
or ( n88233 , n88231 , n88232 );
nand ( n88234 , n38862 , n41895 );
nand ( n88235 , n88233 , n88234 );
buf ( n88236 , n88235 );
buf ( n88237 , n37919 );
nand ( n88238 , n88236 , n88237 );
buf ( n88239 , n88238 );
nand ( n88240 , n88230 , n88239 );
buf ( n88241 , n88240 );
xor ( n88242 , n88227 , n88241 );
buf ( n88243 , n43053 );
buf ( n88244 , n43996 );
not ( n88245 , n88244 );
buf ( n88246 , n37602 );
not ( n88247 , n88246 );
or ( n88248 , n88245 , n88247 );
buf ( n88249 , n38798 );
buf ( n88250 , n42075 );
nand ( n88251 , n88249 , n88250 );
buf ( n88252 , n88251 );
buf ( n88253 , n88252 );
nand ( n88254 , n88248 , n88253 );
buf ( n88255 , n88254 );
buf ( n88256 , n88255 );
nand ( n88257 , n88243 , n88256 );
buf ( n88258 , n88257 );
buf ( n88259 , n88258 );
nand ( n88260 , C1 , n88259 );
buf ( n88261 , n88260 );
buf ( n88262 , n88261 );
xor ( n88263 , n88242 , n88262 );
not ( n88264 , n88263 );
or ( n88265 , n88210 , n88264 );
buf ( n88266 , n88227 );
not ( n88267 , n88266 );
xnor ( n88268 , n88241 , n88262 );
not ( n88269 , n88268 );
or ( n88270 , n88267 , n88269 );
or ( n88271 , n88266 , n88268 );
nand ( n88272 , n88270 , n88271 );
or ( n88273 , n88272 , n88209 );
nand ( n88274 , n88265 , n88273 );
not ( n88275 , n88274 );
or ( n88276 , n88188 , n88275 );
and ( n88277 , n87624 , n88165 );
not ( n88278 , n87624 );
and ( n88279 , n88278 , n88168 );
nor ( n88280 , n88277 , n88279 );
not ( n88281 , n88186 );
and ( n88282 , n88280 , n88281 );
not ( n88283 , n88280 );
and ( n88284 , n88283 , n88186 );
nor ( n88285 , n88282 , n88284 );
or ( n88286 , n88285 , n88274 );
nand ( n88287 , n88276 , n88286 );
not ( n88288 , n88287 );
xnor ( n88289 , n88142 , n88288 );
buf ( n88290 , n88289 );
xor ( n88291 , n88084 , n88290 );
buf ( n88292 , n88291 );
not ( n88293 , n88292 );
not ( n88294 , n88293 );
or ( n88295 , n88048 , n88294 );
not ( n88296 , n88047 );
nand ( n88297 , n88292 , n88296 );
nand ( n88298 , n88295 , n88297 );
xor ( n88299 , n87359 , n87365 );
and ( n88300 , n88299 , n87486 );
and ( n88301 , n87359 , n87365 );
or ( n88302 , n88300 , n88301 );
buf ( n88303 , n88302 );
and ( n88304 , n88298 , n88303 );
not ( n88305 , n88298 );
not ( n88306 , n88303 );
and ( n88307 , n88305 , n88306 );
nor ( n88308 , n88304 , n88307 );
xor ( n88309 , n88042 , n88308 );
nor ( n88310 , n87787 , n88309 );
buf ( n88311 , n88235 );
not ( n88312 , n88311 );
buf ( n88313 , n37872 );
not ( n88314 , n88313 );
or ( n88315 , n88312 , n88314 );
buf ( n88316 , n44435 );
buf ( n88317 , n38830 );
and ( n88318 , n88316 , n88317 );
not ( n88319 , n88316 );
buf ( n88320 , n43470 );
and ( n88321 , n88319 , n88320 );
nor ( n88322 , n88318 , n88321 );
buf ( n88323 , n88322 );
buf ( n88324 , n88323 );
buf ( n88325 , n45617 );
nand ( n88326 , n88324 , n88325 );
buf ( n88327 , n88326 );
buf ( n88328 , n88327 );
nand ( n88329 , n88315 , n88328 );
buf ( n88330 , n88329 );
not ( n88331 , n41844 );
nand ( n88332 , n88331 , n44157 );
nand ( n88333 , n41844 , n37586 );
nand ( n88334 , n88332 , n88333 );
buf ( n88335 , n88334 );
not ( n88336 , n88335 );
buf ( n88337 , n41855 );
not ( n88338 , n88337 );
and ( n88339 , n88336 , n88338 );
buf ( n88340 , n88155 );
buf ( n88341 , n41966 );
and ( n88342 , n88340 , n88341 );
nor ( n88343 , n88339 , n88342 );
buf ( n88344 , n88343 );
buf ( n88345 , n88344 );
not ( n88346 , n88345 );
buf ( n88347 , n88346 );
xor ( n88348 , n88330 , n88347 );
not ( n88349 , n42530 );
buf ( n88350 , n41823 );
not ( n88351 , n88350 );
buf ( n88352 , n39478 );
not ( n88353 , n88352 );
or ( n88354 , n88351 , n88353 );
buf ( n88355 , n41951 );
buf ( n88356 , n51030 );
nand ( n88357 , n88355 , n88356 );
buf ( n88358 , n88357 );
buf ( n88359 , n88358 );
nand ( n88360 , n88354 , n88359 );
buf ( n88361 , n88360 );
not ( n88362 , n88361 );
or ( n88363 , n88349 , n88362 );
nand ( n88364 , n36104 , n88223 );
nand ( n88365 , n88363 , n88364 );
xnor ( n88366 , n88348 , n88365 );
not ( n88367 , n88366 );
not ( n88368 , n88367 );
buf ( n88369 , n42378 );
not ( n88370 , n88369 );
buf ( n88371 , n87813 );
not ( n88372 , n88371 );
or ( n88373 , n88370 , n88372 );
buf ( n88374 , n42339 );
not ( n88375 , n88374 );
buf ( n88376 , n88375 );
buf ( n88377 , n88376 );
not ( n88378 , n88377 );
buf ( n88379 , n42343 );
not ( n88380 , n88379 );
buf ( n88381 , n39008 );
not ( n88382 , n88381 );
or ( n88383 , n88380 , n88382 );
buf ( n88384 , n39005 );
buf ( n88385 , n42350 );
nand ( n88386 , n88384 , n88385 );
buf ( n88387 , n88386 );
buf ( n88388 , n88387 );
nand ( n88389 , n88383 , n88388 );
buf ( n88390 , n88389 );
buf ( n88391 , n88390 );
nand ( n88392 , n88378 , n88391 );
buf ( n88393 , n88392 );
buf ( n88394 , n88393 );
nand ( n88395 , n88373 , n88394 );
buf ( n88396 , n88395 );
buf ( n88397 , n88396 );
not ( n88398 , n88397 );
buf ( n88399 , n88398 );
not ( n88400 , n88399 );
or ( n88401 , n88368 , n88400 );
buf ( n88402 , n88396 );
buf ( n88403 , n88366 );
nand ( n88404 , n88402 , n88403 );
buf ( n88405 , n88404 );
nand ( n88406 , n88401 , n88405 );
buf ( n88407 , n38127 );
buf ( n88408 , n87931 );
or ( n88409 , n88407 , n88408 );
buf ( n88410 , n45141 );
buf ( n88411 , n49391 );
not ( n88412 , n88411 );
buf ( n88413 , n39672 );
not ( n88414 , n88413 );
and ( n88415 , n88412 , n88414 );
buf ( n88416 , n44004 );
buf ( n88417 , n39688 );
and ( n88418 , n88416 , n88417 );
nor ( n88419 , n88415 , n88418 );
buf ( n88420 , n88419 );
buf ( n88421 , n88420 );
or ( n88422 , n88410 , n88421 );
nand ( n88423 , n88409 , n88422 );
buf ( n88424 , n88423 );
buf ( n88425 , n87912 );
not ( n88426 , n88425 );
buf ( n88427 , n50374 );
not ( n88428 , n88427 );
or ( n88429 , n88426 , n88428 );
buf ( n88430 , n43982 );
buf ( n88431 , n41882 );
not ( n88432 , n88431 );
buf ( n88433 , n38468 );
not ( n88434 , n88433 );
or ( n88435 , n88432 , n88434 );
buf ( n88436 , n36527 );
buf ( n88437 , n41879 );
nand ( n88438 , n88436 , n88437 );
buf ( n88439 , n88438 );
buf ( n88440 , n88439 );
nand ( n88441 , n88435 , n88440 );
buf ( n88442 , n88441 );
buf ( n88443 , n88442 );
nand ( n88444 , n88430 , n88443 );
buf ( n88445 , n88444 );
buf ( n88446 , n88445 );
nand ( n88447 , n88429 , n88446 );
buf ( n88448 , n88447 );
xor ( n88449 , n88424 , n88448 );
not ( n88450 , n88181 );
not ( n88451 , n88450 );
not ( n88452 , n45158 );
or ( n88453 , n88451 , n88452 );
buf ( n88454 , n41975 );
buf ( n88455 , n49425 );
not ( n88456 , n88455 );
buf ( n88457 , n88456 );
buf ( n88458 , n88457 );
and ( n88459 , n88454 , n88458 );
not ( n88460 , n88454 );
buf ( n88461 , n39139 );
and ( n88462 , n88460 , n88461 );
nor ( n88463 , n88459 , n88462 );
buf ( n88464 , n88463 );
or ( n88465 , n36909 , n88464 );
nand ( n88466 , n88453 , n88465 );
xor ( n88467 , n88449 , n88466 );
and ( n88468 , n88406 , n88467 );
not ( n88469 , n88406 );
buf ( n88470 , n88467 );
not ( n88471 , n88470 );
buf ( n88472 , n88471 );
and ( n88473 , n88469 , n88472 );
nor ( n88474 , n88468 , n88473 );
buf ( n88475 , n87624 );
not ( n88476 , n88475 );
buf ( n88477 , n88168 );
not ( n88478 , n88477 );
or ( n88479 , n88476 , n88478 );
buf ( n88480 , n87627 );
not ( n88481 , n88480 );
buf ( n88482 , n88165 );
not ( n88483 , n88482 );
or ( n88484 , n88481 , n88483 );
buf ( n88485 , n88185 );
nand ( n88486 , n88484 , n88485 );
buf ( n88487 , n88486 );
buf ( n88488 , n88487 );
nand ( n88489 , n88479 , n88488 );
buf ( n88490 , n88489 );
buf ( n88491 , n88490 );
buf ( n88492 , n38758 );
not ( n88493 , n88492 );
and ( n88494 , n37293 , n45401 );
not ( n88495 , n37293 );
and ( n88496 , n88495 , n38413 );
or ( n88497 , n88494 , n88496 );
buf ( n88498 , n88497 );
not ( n88499 , n88498 );
or ( n88500 , n88493 , n88499 );
buf ( n88501 , n87955 );
buf ( n88502 , n38775 );
nand ( n88503 , n88501 , n88502 );
buf ( n88504 , n88503 );
buf ( n88505 , n88504 );
nand ( n88506 , n88500 , n88505 );
buf ( n88507 , n88506 );
buf ( n88508 , n88507 );
not ( n88509 , n88508 );
buf ( n88510 , n88509 );
buf ( n88511 , n88510 );
and ( n88512 , n88491 , n88511 );
not ( n88513 , n88491 );
buf ( n88514 , n88507 );
and ( n88515 , n88513 , n88514 );
nor ( n88516 , n88512 , n88515 );
buf ( n88517 , n88516 );
buf ( n88518 , n40002 );
not ( n88519 , n88518 );
buf ( n88520 , n88201 );
not ( n88521 , n88520 );
or ( n88522 , n88519 , n88521 );
buf ( n88523 , n40010 );
not ( n88524 , n88523 );
buf ( n88525 , n57073 );
not ( n88526 , n88525 );
or ( n88527 , n88524 , n88526 );
buf ( n88528 , n49804 );
buf ( n88529 , n40009 );
nand ( n88530 , n88528 , n88529 );
buf ( n88531 , n88530 );
buf ( n88532 , n88531 );
nand ( n88533 , n88527 , n88532 );
buf ( n88534 , n88533 );
buf ( n88535 , n88534 );
buf ( n88536 , n39986 );
nand ( n88537 , n88535 , n88536 );
buf ( n88538 , n88537 );
buf ( n88539 , n88538 );
nand ( n88540 , n88522 , n88539 );
buf ( n88541 , n88540 );
and ( n88542 , n88517 , n88541 );
not ( n88543 , n88517 );
buf ( n88544 , n88541 );
not ( n88545 , n88544 );
buf ( n88546 , n88545 );
and ( n88547 , n88543 , n88546 );
or ( n88548 , n88542 , n88547 );
not ( n88549 , n88548 );
xor ( n88550 , n88474 , n88549 );
xor ( n88551 , n87868 , n87893 );
and ( n88552 , n88551 , n87967 );
and ( n88553 , n87868 , n87893 );
or ( n88554 , n88552 , n88553 );
buf ( n88555 , n88554 );
not ( n88556 , n88555 );
xor ( n88557 , n88550 , n88556 );
xor ( n88558 , n87970 , n88022 );
and ( n88559 , n88558 , n88031 );
and ( n88560 , n87970 , n88022 );
or ( n88561 , n88559 , n88560 );
buf ( n88562 , n88561 );
not ( n88563 , n88562 );
xor ( n88564 , n88557 , n88563 );
not ( n88565 , n39395 );
not ( n88566 , n87831 );
or ( n88567 , n88565 , n88566 );
buf ( n88568 , n39000 );
not ( n88569 , n88568 );
buf ( n88570 , n43031 );
not ( n88571 , n88570 );
or ( n88572 , n88569 , n88571 );
nand ( n88573 , n38244 , n38997 );
buf ( n88574 , n88573 );
nand ( n88575 , n88572 , n88574 );
buf ( n88576 , n88575 );
buf ( n88577 , n88576 );
buf ( n88578 , n39374 );
nand ( n88579 , n88577 , n88578 );
buf ( n88580 , n88579 );
nand ( n88581 , n88567 , n88580 );
not ( n88582 , n88581 );
not ( n88583 , n87918 );
nand ( n88584 , n88583 , n87940 );
not ( n88585 , n88584 );
not ( n88586 , n87965 );
or ( n88587 , n88585 , n88586 );
nand ( n88588 , n87939 , n87918 );
nand ( n88589 , n88587 , n88588 );
xor ( n88590 , n88582 , n88589 );
not ( n88591 , n87882 );
not ( n88592 , n42631 );
or ( n88593 , n88591 , n88592 );
buf ( n88594 , n25160 );
not ( n88595 , n88594 );
buf ( n88596 , n37081 );
not ( n88597 , n88596 );
or ( n88598 , n88595 , n88597 );
buf ( n88599 , n39340 );
buf ( n88600 , n42581 );
nand ( n88601 , n88599 , n88600 );
buf ( n88602 , n88601 );
buf ( n88603 , n88602 );
nand ( n88604 , n88598 , n88603 );
buf ( n88605 , n88604 );
buf ( n88606 , n88605 );
buf ( n88607 , n42566 );
nand ( n88608 , n88606 , n88607 );
buf ( n88609 , n88608 );
nand ( n88610 , n88593 , n88609 );
xnor ( n88611 , n88590 , n88610 );
not ( n88612 , n88611 );
not ( n88613 , n88612 );
not ( n88614 , n88016 );
not ( n88615 , n87975 );
nand ( n88616 , n88615 , n87996 );
not ( n88617 , n88616 );
or ( n88618 , n88614 , n88617 );
not ( n88619 , n87976 );
nand ( n88620 , n88619 , n87993 );
nand ( n88621 , n88618 , n88620 );
not ( n88622 , n88621 );
not ( n88623 , n88622 );
or ( n88624 , n88613 , n88623 );
or ( n88625 , n88622 , n88612 );
nand ( n88626 , n88624 , n88625 );
not ( n88627 , n88626 );
buf ( n88628 , n88287 );
buf ( n88629 , n88127 );
buf ( n88630 , n88629 );
or ( n88631 , n88628 , n88630 );
buf ( n88632 , n88141 );
nand ( n88633 , n88631 , n88632 );
buf ( n88634 , n88633 );
buf ( n88635 , n88287 );
buf ( n88636 , n88629 );
nand ( n88637 , n88635 , n88636 );
buf ( n88638 , n88637 );
nand ( n88639 , n88634 , n88638 );
buf ( n88640 , n88639 );
not ( n88641 , n88640 );
or ( n88642 , n88627 , n88641 );
or ( n88643 , n88640 , n88626 );
nand ( n88644 , n88642 , n88643 );
xnor ( n88645 , n88564 , n88644 );
buf ( n88646 , n88645 );
xor ( n88647 , n88068 , n88083 );
and ( n88648 , n88647 , n88290 );
and ( n88649 , n88068 , n88083 );
or ( n88650 , n88648 , n88649 );
buf ( n88651 , n88650 );
buf ( n88652 , n88651 );
buf ( n88653 , n41705 );
not ( n88654 , n88653 );
buf ( n88655 , n88009 );
not ( n88656 , n88655 );
or ( n88657 , n88654 , n88656 );
buf ( n88658 , n41666 );
not ( n88659 , n88658 );
buf ( n88660 , n39582 );
not ( n88661 , n88660 );
or ( n88662 , n88659 , n88661 );
buf ( n88663 , n36611 );
buf ( n88664 , n41663 );
nand ( n88665 , n88663 , n88664 );
buf ( n88666 , n88665 );
buf ( n88667 , n88666 );
nand ( n88668 , n88662 , n88667 );
buf ( n88669 , n88668 );
buf ( n88670 , n88669 );
buf ( n88671 , n41647 );
nand ( n88672 , n88670 , n88671 );
buf ( n88673 , n88672 );
buf ( n88674 , n88673 );
nand ( n88675 , n88657 , n88674 );
buf ( n88676 , n88675 );
buf ( n88677 , n44586 );
not ( n88678 , n88677 );
buf ( n88679 , n87983 );
not ( n88680 , n88679 );
or ( n88681 , n88678 , n88680 );
and ( n88682 , n36427 , n25183 );
not ( n88683 , n36427 );
and ( n88684 , n88683 , n25184 );
or ( n88685 , n88682 , n88684 );
buf ( n88686 , n88685 );
buf ( n88687 , n43909 );
nand ( n88688 , n88686 , n88687 );
buf ( n88689 , n88688 );
buf ( n88690 , n88689 );
nand ( n88691 , n88681 , n88690 );
buf ( n88692 , n88691 );
not ( n88693 , n88692 );
xor ( n88694 , n88676 , n88693 );
xor ( n88695 , n88111 , n88116 );
and ( n88696 , n88695 , n88126 );
and ( n88697 , n88111 , n88116 );
or ( n88698 , n88696 , n88697 );
not ( n88699 , n88698 );
xor ( n88700 , n88694 , n88699 );
buf ( n88701 , n88700 );
buf ( n88702 , n38798 );
not ( n88703 , n88702 );
buf ( n88704 , n43365 );
not ( n88705 , n88704 );
and ( n88706 , n88703 , n88705 );
buf ( n88707 , n36360 );
buf ( n88708 , n43365 );
and ( n88709 , n88707 , n88708 );
nor ( n88710 , n88706 , n88709 );
buf ( n88711 , n88710 );
not ( n88712 , n88711 );
and ( n88713 , n36453 , n88712 );
nor ( n88714 , C0 , n88713 );
buf ( n88715 , n88714 );
buf ( n88716 , n37403 );
not ( n88717 , n88716 );
buf ( n88718 , n88101 );
not ( n88719 , n88718 );
or ( n88720 , n88717 , n88719 );
not ( n88721 , n88089 );
not ( n88722 , n50925 );
or ( n88723 , n88721 , n88722 );
buf ( n88724 , n43434 );
not ( n88725 , n88724 );
buf ( n88726 , n39522 );
nand ( n88727 , n88725 , n88726 );
buf ( n88728 , n88727 );
nand ( n88729 , n88723 , n88728 );
nand ( n88730 , n88729 , n38150 );
buf ( n88731 , n88730 );
nand ( n88732 , n88720 , n88731 );
buf ( n88733 , n88732 );
buf ( n88734 , n88733 );
xor ( n88735 , n88715 , n88734 );
buf ( n88736 , n88240 );
not ( n88737 , n88736 );
buf ( n88738 , n88261 );
not ( n88739 , n88738 );
or ( n88740 , n88737 , n88739 );
buf ( n88741 , n88261 );
buf ( n88742 , n88240 );
or ( n88743 , n88741 , n88742 );
buf ( n88744 , n88227 );
nand ( n88745 , n88743 , n88744 );
buf ( n88746 , n88745 );
buf ( n88747 , n88746 );
nand ( n88748 , n88740 , n88747 );
buf ( n88749 , n88748 );
buf ( n88750 , n88749 );
xor ( n88751 , n88735 , n88750 );
buf ( n88752 , n88751 );
buf ( n88753 , n87839 );
not ( n88754 , n88753 );
buf ( n88755 , n87815 );
not ( n88756 , n88755 );
or ( n88757 , n88754 , n88756 );
buf ( n88758 , n87798 );
nand ( n88759 , n88757 , n88758 );
buf ( n88760 , n88759 );
buf ( n88761 , n88760 );
buf ( n88762 , n87820 );
buf ( n88763 , n87836 );
nand ( n88764 , n88762 , n88763 );
buf ( n88765 , n88764 );
buf ( n88766 , n88765 );
nand ( n88767 , n88761 , n88766 );
buf ( n88768 , n88767 );
xor ( n88769 , n88752 , n88768 );
buf ( n88770 , n88769 );
nand ( n88771 , n88285 , n88209 );
and ( n88772 , n88771 , n88272 );
nor ( n88773 , n88285 , n88209 );
nor ( n88774 , n88772 , n88773 );
buf ( n88775 , n88774 );
xnor ( n88776 , n88770 , n88775 );
buf ( n88777 , n88776 );
buf ( n88778 , n88777 );
xor ( n88779 , n88701 , n88778 );
xor ( n88780 , n87791 , n87841 );
and ( n88781 , n88780 , n87848 );
and ( n88782 , n87791 , n87841 );
or ( n88783 , n88781 , n88782 );
buf ( n88784 , n88783 );
xor ( n88785 , n88779 , n88784 );
buf ( n88786 , n88785 );
buf ( n88787 , n88786 );
xor ( n88788 , n88652 , n88787 );
xor ( n88789 , n87850 , n87861 );
and ( n88790 , n88789 , n88034 );
and ( n88791 , n87850 , n87861 );
or ( n88792 , n88790 , n88791 );
buf ( n88793 , n88792 );
buf ( n88794 , n88793 );
xor ( n88795 , n88788 , n88794 );
buf ( n88796 , n88795 );
buf ( n88797 , n88796 );
xor ( n88798 , n88646 , n88797 );
nand ( n88799 , n88293 , n88296 );
not ( n88800 , n88799 );
not ( n88801 , n88303 );
or ( n88802 , n88800 , n88801 );
nand ( n88803 , n88292 , n88047 );
nand ( n88804 , n88802 , n88803 );
buf ( n88805 , n88804 );
xor ( n88806 , n88798 , n88805 );
buf ( n88807 , n88806 );
buf ( n88808 , n88807 );
xor ( n88809 , n88036 , n88041 );
and ( n88810 , n88809 , n88308 );
and ( n88811 , n88036 , n88041 );
or ( n88812 , n88810 , n88811 );
buf ( n88813 , n88812 );
nor ( n88814 , n88808 , n88813 );
buf ( n88815 , n88814 );
nor ( n88816 , n88310 , n88815 );
nand ( n88817 , n87779 , n88816 );
not ( n88818 , n88817 );
buf ( n88819 , n39986 );
not ( n88820 , n88819 );
buf ( n88821 , n24092 );
not ( n88822 , n88821 );
buf ( n88823 , n39861 );
not ( n88824 , n88823 );
or ( n88825 , n88822 , n88824 );
buf ( n88826 , n50876 );
buf ( n88827 , n40009 );
nand ( n88828 , n88826 , n88827 );
buf ( n88829 , n88828 );
buf ( n88830 , n88829 );
nand ( n88831 , n88825 , n88830 );
buf ( n88832 , n88831 );
buf ( n88833 , n88832 );
not ( n88834 , n88833 );
or ( n88835 , n88820 , n88834 );
buf ( n88836 , n88534 );
buf ( n88837 , n40002 );
nand ( n88838 , n88836 , n88837 );
buf ( n88839 , n88838 );
buf ( n88840 , n88839 );
nand ( n88841 , n88835 , n88840 );
buf ( n88842 , n88841 );
buf ( n88843 , n88842 );
buf ( n88844 , n42566 );
not ( n88845 , n88844 );
buf ( n88846 , n25160 );
not ( n88847 , n88846 );
buf ( n88848 , n43597 );
not ( n88849 , n88848 );
or ( n88850 , n88847 , n88849 );
buf ( n88851 , n36396 );
buf ( n88852 , n42581 );
nand ( n88853 , n88851 , n88852 );
buf ( n88854 , n88853 );
buf ( n88855 , n88854 );
nand ( n88856 , n88850 , n88855 );
buf ( n88857 , n88856 );
buf ( n88858 , n88857 );
not ( n88859 , n88858 );
or ( n88860 , n88845 , n88859 );
buf ( n88861 , n88605 );
buf ( n88862 , n42631 );
nand ( n88863 , n88861 , n88862 );
buf ( n88864 , n88863 );
buf ( n88865 , n88864 );
nand ( n88866 , n88860 , n88865 );
buf ( n88867 , n88866 );
buf ( n88868 , n88867 );
xor ( n88869 , n88843 , n88868 );
buf ( n88870 , n43719 );
buf ( n88871 , n88442 );
not ( n88872 , n88871 );
buf ( n88873 , n88872 );
buf ( n88874 , n88873 );
or ( n88875 , n88870 , n88874 );
buf ( n88876 , n39813 );
and ( n88877 , n45370 , n52246 );
not ( n88878 , n45370 );
and ( n88879 , n88878 , n38471 );
nor ( n88880 , n88877 , n88879 );
buf ( n88881 , n88880 );
or ( n88882 , n88876 , n88881 );
nand ( n88883 , n88875 , n88882 );
buf ( n88884 , n88883 );
buf ( n88885 , n88884 );
buf ( n88886 , n37452 );
not ( n88887 , n88886 );
buf ( n88888 , n88143 );
not ( n88889 , n88888 );
buf ( n88890 , n37786 );
not ( n88891 , n88890 );
or ( n88892 , n88889 , n88891 );
buf ( n88893 , n59203 );
buf ( n88894 , n37475 );
nand ( n88895 , n88893 , n88894 );
buf ( n88896 , n88895 );
buf ( n88897 , n88896 );
nand ( n88898 , n88892 , n88897 );
buf ( n88899 , n88898 );
buf ( n88900 , n88899 );
not ( n88901 , n88900 );
or ( n88902 , n88887 , n88901 );
buf ( n88903 , n88334 );
not ( n88904 , n88903 );
buf ( n88905 , n51912 );
nand ( n88906 , n88904 , n88905 );
buf ( n88907 , n88906 );
buf ( n88908 , n88907 );
nand ( n88909 , n88902 , n88908 );
buf ( n88910 , n88909 );
buf ( n88911 , n88910 );
xor ( n88912 , n88885 , n88911 );
buf ( n88913 , n38150 );
not ( n88914 , n88913 );
buf ( n88915 , n88089 );
not ( n88916 , n88915 );
buf ( n88917 , n59221 );
not ( n88918 , n88917 );
or ( n88919 , n88916 , n88918 );
buf ( n88920 , n39246 );
buf ( n88921 , n37329 );
nand ( n88922 , n88920 , n88921 );
buf ( n88923 , n88922 );
buf ( n88924 , n88923 );
nand ( n88925 , n88919 , n88924 );
buf ( n88926 , n88925 );
buf ( n88927 , n88926 );
not ( n88928 , n88927 );
or ( n88929 , n88914 , n88928 );
nand ( n88930 , n88729 , n37403 );
buf ( n88931 , n88930 );
nand ( n88932 , n88929 , n88931 );
buf ( n88933 , n88932 );
buf ( n88934 , n88933 );
xor ( n88935 , n88912 , n88934 );
buf ( n88936 , n88935 );
buf ( n88937 , n88936 );
xor ( n88938 , n88869 , n88937 );
buf ( n88939 , n88938 );
not ( n88940 , n88939 );
or ( n88941 , n88610 , n88581 );
nand ( n88942 , n88941 , n88589 );
nand ( n88943 , n88610 , n88581 );
nand ( n88944 , n88942 , n88943 );
not ( n88945 , n88944 );
nand ( n88946 , n88940 , n88945 );
not ( n88947 , n88946 );
not ( n88948 , n88676 );
not ( n88949 , n88948 );
not ( n88950 , n88693 );
or ( n88951 , n88949 , n88950 );
nand ( n88952 , n88951 , n88698 );
nand ( n88953 , n88692 , n88676 );
nand ( n88954 , n88952 , n88953 );
not ( n88955 , n88954 );
or ( n88956 , n88947 , n88955 );
nand ( n88957 , n88944 , n88939 );
nand ( n88958 , n88956 , n88957 );
buf ( n88959 , n88376 );
not ( n88960 , n88959 );
buf ( n88961 , n42375 );
not ( n88962 , n88961 );
or ( n88963 , n88960 , n88962 );
buf ( n88964 , n88390 );
nand ( n88965 , n88963 , n88964 );
buf ( n88966 , n88965 );
buf ( n88967 , n88966 );
buf ( n88968 , n38758 );
not ( n88969 , n88968 );
buf ( n88970 , n38413 );
not ( n88971 , n88970 );
buf ( n88972 , n43879 );
not ( n88973 , n88972 );
or ( n88974 , n88971 , n88973 );
buf ( n88975 , n43885 );
buf ( n88976 , n38420 );
nand ( n88977 , n88975 , n88976 );
buf ( n88978 , n88977 );
buf ( n88979 , n88978 );
nand ( n88980 , n88974 , n88979 );
buf ( n88981 , n88980 );
buf ( n88982 , n88981 );
not ( n88983 , n88982 );
or ( n88984 , n88969 , n88983 );
buf ( n88985 , n88497 );
buf ( n88986 , n38775 );
nand ( n88987 , n88985 , n88986 );
buf ( n88988 , n88987 );
buf ( n88989 , n88988 );
nand ( n88990 , n88984 , n88989 );
buf ( n88991 , n88990 );
buf ( n88992 , n88991 );
xor ( n88993 , n88967 , n88992 );
xor ( n88994 , n88715 , n88734 );
and ( n88995 , n88994 , n88750 );
and ( n88996 , n88715 , n88734 );
or ( n88997 , n88995 , n88996 );
buf ( n88998 , n88997 );
buf ( n88999 , n88998 );
and ( n89000 , n88993 , n88999 );
and ( n89001 , n88967 , n88992 );
or ( n89002 , n89000 , n89001 );
buf ( n89003 , n89002 );
not ( n89004 , n39986 );
not ( n89005 , n24092 );
not ( n89006 , n37081 );
or ( n89007 , n89005 , n89006 );
not ( n89008 , n24092 );
nand ( n89009 , n89008 , n40089 );
nand ( n89010 , n89007 , n89009 );
not ( n89011 , n89010 );
or ( n89012 , n89004 , n89011 );
buf ( n89013 , n88832 );
buf ( n89014 , n40002 );
nand ( n89015 , n89013 , n89014 );
buf ( n89016 , n89015 );
nand ( n89017 , n89012 , n89016 );
not ( n89018 , n89017 );
not ( n89019 , n44586 );
buf ( n89020 , n25184 );
not ( n89021 , n89020 );
buf ( n89022 , n39927 );
not ( n89023 , n89022 );
or ( n89024 , n89021 , n89023 );
buf ( n89025 , n36562 );
buf ( n89026 , n25183 );
nand ( n89027 , n89025 , n89026 );
buf ( n89028 , n89027 );
buf ( n89029 , n89028 );
nand ( n89030 , n89024 , n89029 );
buf ( n89031 , n89030 );
not ( n89032 , n89031 );
or ( n89033 , n89019 , n89032 );
buf ( n89034 , n25184 );
not ( n89035 , n89034 );
buf ( n89036 , n36614 );
not ( n89037 , n89036 );
or ( n89038 , n89035 , n89037 );
buf ( n89039 , n36617 );
buf ( n89040 , n25183 );
nand ( n89041 , n89039 , n89040 );
buf ( n89042 , n89041 );
buf ( n89043 , n89042 );
nand ( n89044 , n89038 , n89043 );
buf ( n89045 , n89044 );
nand ( n89046 , n43909 , n89045 );
nand ( n89047 , n89033 , n89046 );
not ( n89048 , n89047 );
not ( n89049 , n43053 );
buf ( n89050 , n41882 );
not ( n89051 , n89050 );
buf ( n89052 , n37602 );
not ( n89053 , n89052 );
or ( n89054 , n89051 , n89053 );
buf ( n89055 , n36360 );
buf ( n89056 , n41879 );
nand ( n89057 , n89055 , n89056 );
buf ( n89058 , n89057 );
buf ( n89059 , n89058 );
nand ( n89060 , n89054 , n89059 );
buf ( n89061 , n89060 );
not ( n89062 , n89061 );
or ( n89063 , n89049 , n89062 );
and ( n89064 , n38798 , n42152 );
not ( n89065 , n38798 );
and ( n89066 , n89065 , n42160 );
nor ( n89067 , n89064 , n89066 );
nand ( n89068 , n89063 , C1 );
buf ( n89069 , n89068 );
buf ( n89070 , n38865 );
not ( n89071 , n89070 );
buf ( n89072 , n47898 );
not ( n89073 , n89072 );
or ( n89074 , n89071 , n89073 );
buf ( n89075 , n44983 );
buf ( n89076 , n49391 );
nand ( n89077 , n89075 , n89076 );
buf ( n89078 , n89077 );
buf ( n89079 , n89078 );
nand ( n89080 , n89074 , n89079 );
buf ( n89081 , n89080 );
buf ( n89082 , n89081 );
not ( n89083 , n89082 );
buf ( n89084 , n43991 );
not ( n89085 , n89084 );
or ( n89086 , n89083 , n89085 );
buf ( n89087 , n38830 );
not ( n89088 , n89087 );
buf ( n89089 , n38068 );
not ( n89090 , n89089 );
or ( n89091 , n89088 , n89090 );
buf ( n89092 , n49391 );
buf ( n89093 , n39742 );
nand ( n89094 , n89092 , n89093 );
buf ( n89095 , n89094 );
buf ( n89096 , n89095 );
nand ( n89097 , n89091 , n89096 );
buf ( n89098 , n89097 );
buf ( n89099 , n89098 );
buf ( n89100 , n38060 );
nand ( n89101 , n89099 , n89100 );
buf ( n89102 , n89101 );
buf ( n89103 , n89102 );
nand ( n89104 , n89086 , n89103 );
buf ( n89105 , n89104 );
buf ( n89106 , n89105 );
xor ( n89107 , n89069 , n89106 );
buf ( n89108 , n43719 );
buf ( n89109 , n88880 );
or ( n89110 , n89108 , n89109 );
buf ( n89111 , n39813 );
buf ( n89112 , n41951 );
buf ( n89113 , n36527 );
and ( n89114 , n89112 , n89113 );
not ( n89115 , n89112 );
buf ( n89116 , n39726 );
and ( n89117 , n89115 , n89116 );
nor ( n89118 , n89114 , n89117 );
buf ( n89119 , n89118 );
buf ( n89120 , n89119 );
or ( n89121 , n89111 , n89120 );
nand ( n89122 , n89110 , n89121 );
buf ( n89123 , n89122 );
buf ( n89124 , n89123 );
xor ( n89125 , n89107 , n89124 );
buf ( n89126 , n89125 );
buf ( n89127 , n89126 );
not ( n89128 , n89127 );
buf ( n89129 , n89128 );
and ( n89130 , n89048 , n89129 );
not ( n89131 , n89048 );
and ( n89132 , n89131 , n89126 );
nor ( n89133 , n89130 , n89132 );
not ( n89134 , n89133 );
or ( n89135 , n89018 , n89134 );
not ( n89136 , n89129 );
nand ( n89137 , n89136 , n89048 );
not ( n89138 , n89126 );
nand ( n89139 , n89138 , n89047 );
not ( n89140 , n89017 );
nand ( n89141 , n89137 , n89139 , n89140 );
nand ( n89142 , n89135 , n89141 );
xor ( n89143 , n89003 , n89142 );
xor ( n89144 , n88843 , n88868 );
and ( n89145 , n89144 , n88937 );
and ( n89146 , n88843 , n88868 );
or ( n89147 , n89145 , n89146 );
buf ( n89148 , n89147 );
xnor ( n89149 , n89143 , n89148 );
not ( n89150 , n88714 );
not ( n89151 , n89150 );
not ( n89152 , n43991 );
not ( n89153 , n44004 );
not ( n89154 , n39688 );
or ( n89155 , n89153 , n89154 );
or ( n89156 , n49391 , n39672 );
nand ( n89157 , n89155 , n89156 );
not ( n89158 , n89157 );
or ( n89159 , n89152 , n89158 );
buf ( n89160 , n89081 );
buf ( n89161 , n43414 );
nand ( n89162 , n89160 , n89161 );
buf ( n89163 , n89162 );
nand ( n89164 , n89159 , n89163 );
not ( n89165 , n89164 );
or ( n89166 , n89151 , n89165 );
not ( n89167 , n88714 );
buf ( n89168 , n89164 );
not ( n89169 , n89168 );
buf ( n89170 , n89169 );
not ( n89171 , n89170 );
or ( n89172 , n89167 , n89171 );
buf ( n89173 , n45426 );
buf ( n89174 , n88464 );
or ( n89175 , n89173 , n89174 );
buf ( n89176 , n36909 );
buf ( n89177 , n39656 );
buf ( n89178 , n43095 );
and ( n89179 , n89177 , n89178 );
not ( n89180 , n89177 );
buf ( n89181 , n44689 );
and ( n89182 , n89180 , n89181 );
nor ( n89183 , n89179 , n89182 );
buf ( n89184 , n89183 );
buf ( n89185 , n89184 );
or ( n89186 , n89176 , n89185 );
nand ( n89187 , n89175 , n89186 );
buf ( n89188 , n89187 );
nand ( n89189 , n89172 , n89188 );
nand ( n89190 , n89166 , n89189 );
not ( n89191 , n89190 );
not ( n89192 , n89191 );
buf ( n89193 , n41647 );
not ( n89194 , n89193 );
buf ( n89195 , n41666 );
not ( n89196 , n89195 );
buf ( n89197 , n35971 );
not ( n89198 , n89197 );
or ( n89199 , n89196 , n89198 );
buf ( n89200 , n53159 );
buf ( n89201 , n41663 );
nand ( n89202 , n89200 , n89201 );
buf ( n89203 , n89202 );
buf ( n89204 , n89203 );
nand ( n89205 , n89199 , n89204 );
buf ( n89206 , n89205 );
buf ( n89207 , n89206 );
not ( n89208 , n89207 );
or ( n89209 , n89194 , n89208 );
buf ( n89210 , n41666 );
not ( n89211 , n89210 );
buf ( n89212 , n36054 );
not ( n89213 , n89212 );
or ( n89214 , n89211 , n89213 );
buf ( n89215 , n44718 );
buf ( n89216 , n41663 );
nand ( n89217 , n89215 , n89216 );
buf ( n89218 , n89217 );
buf ( n89219 , n89218 );
nand ( n89220 , n89214 , n89219 );
buf ( n89221 , n89220 );
buf ( n89222 , n89221 );
buf ( n89223 , n41705 );
nand ( n89224 , n89222 , n89223 );
buf ( n89225 , n89224 );
buf ( n89226 , n89225 );
nand ( n89227 , n89209 , n89226 );
buf ( n89228 , n89227 );
not ( n89229 , n89228 );
or ( n89230 , n89192 , n89229 );
not ( n89231 , n89228 );
nand ( n89232 , n89231 , n89190 );
nand ( n89233 , n89230 , n89232 );
not ( n89234 , n39395 );
buf ( n89235 , n39000 );
not ( n89236 , n89235 );
buf ( n89237 , n39407 );
not ( n89238 , n89237 );
or ( n89239 , n89236 , n89238 );
buf ( n89240 , n42941 );
buf ( n89241 , n38997 );
nand ( n89242 , n89240 , n89241 );
buf ( n89243 , n89242 );
buf ( n89244 , n89243 );
nand ( n89245 , n89239 , n89244 );
buf ( n89246 , n89245 );
not ( n89247 , n89246 );
or ( n89248 , n89234 , n89247 );
buf ( n89249 , n39000 );
not ( n89250 , n89249 );
buf ( n89251 , n39280 );
not ( n89252 , n89251 );
or ( n89253 , n89250 , n89252 );
buf ( n89254 , n39277 );
buf ( n89255 , n38997 );
nand ( n89256 , n89254 , n89255 );
buf ( n89257 , n89256 );
buf ( n89258 , n89257 );
nand ( n89259 , n89253 , n89258 );
buf ( n89260 , n89259 );
buf ( n89261 , n89260 );
buf ( n89262 , n39374 );
nand ( n89263 , n89261 , n89262 );
buf ( n89264 , n89263 );
nand ( n89265 , n89248 , n89264 );
not ( n89266 , n89265 );
and ( n89267 , n89233 , n89266 );
not ( n89268 , n89233 );
and ( n89269 , n89268 , n89265 );
nor ( n89270 , n89267 , n89269 );
buf ( n89271 , n41647 );
not ( n89272 , n89271 );
buf ( n89273 , n89221 );
not ( n89274 , n89273 );
or ( n89275 , n89272 , n89274 );
buf ( n89276 , n41705 );
buf ( n89277 , n88669 );
nand ( n89278 , n89276 , n89277 );
buf ( n89279 , n89278 );
buf ( n89280 , n89279 );
nand ( n89281 , n89275 , n89280 );
buf ( n89282 , n89281 );
buf ( n89283 , n89282 );
xor ( n89284 , n88424 , n88448 );
and ( n89285 , n89284 , n88466 );
and ( n89286 , n88424 , n88448 );
or ( n89287 , n89285 , n89286 );
buf ( n89288 , n89287 );
xor ( n89289 , n89283 , n89288 );
buf ( n89290 , n89164 );
buf ( n89291 , n88714 );
xor ( n89292 , n89290 , n89291 );
buf ( n89293 , n89188 );
not ( n89294 , n89293 );
xor ( n89295 , n89292 , n89294 );
buf ( n89296 , n89295 );
buf ( n89297 , n89296 );
and ( n89298 , n89289 , n89297 );
and ( n89299 , n89283 , n89288 );
or ( n89300 , n89298 , n89299 );
buf ( n89301 , n89300 );
and ( n89302 , n89270 , n89301 );
not ( n89303 , n89270 );
not ( n89304 , n89301 );
and ( n89305 , n89303 , n89304 );
nor ( n89306 , n89302 , n89305 );
xor ( n89307 , n88885 , n88911 );
and ( n89308 , n89307 , n88934 );
and ( n89309 , n88885 , n88911 );
or ( n89310 , n89308 , n89309 );
buf ( n89311 , n89310 );
not ( n89312 , n89311 );
not ( n89313 , n89312 );
buf ( n89314 , n38775 );
not ( n89315 , n89314 );
buf ( n89316 , n88981 );
not ( n89317 , n89316 );
or ( n89318 , n89315 , n89317 );
buf ( n89319 , n38413 );
not ( n89320 , n89319 );
buf ( n89321 , n43031 );
not ( n89322 , n89321 );
or ( n89323 , n89320 , n89322 );
buf ( n89324 , n38247 );
buf ( n89325 , n38420 );
nand ( n89326 , n89324 , n89325 );
buf ( n89327 , n89326 );
buf ( n89328 , n89327 );
nand ( n89329 , n89323 , n89328 );
buf ( n89330 , n89329 );
buf ( n89331 , n89330 );
buf ( n89332 , n38758 );
nand ( n89333 , n89331 , n89332 );
buf ( n89334 , n89333 );
buf ( n89335 , n89334 );
nand ( n89336 , n89318 , n89335 );
buf ( n89337 , n89336 );
not ( n89338 , n89337 );
not ( n89339 , n89338 );
buf ( n89340 , n43806 );
not ( n89341 , n89340 );
buf ( n89342 , n39478 );
not ( n89343 , n89342 );
or ( n89344 , n89341 , n89343 );
buf ( n89345 , n33077 );
buf ( n89346 , n75045 );
nand ( n89347 , n89345 , n89346 );
buf ( n89348 , n89347 );
buf ( n89349 , n89348 );
nand ( n89350 , n89344 , n89349 );
buf ( n89351 , n89350 );
buf ( n89352 , n89351 );
not ( n89353 , n89352 );
buf ( n89354 , n51937 );
not ( n89355 , n89354 );
or ( n89356 , n89353 , n89355 );
buf ( n89357 , n32969 );
buf ( n89358 , n28723 );
not ( n89359 , n89358 );
buf ( n89360 , n39493 );
not ( n89361 , n89360 );
or ( n89362 , n89359 , n89361 );
buf ( n89363 , n51030 );
buf ( n89364 , n41975 );
nand ( n89365 , n89363 , n89364 );
buf ( n89366 , n89365 );
buf ( n89367 , n89366 );
nand ( n89368 , n89362 , n89367 );
buf ( n89369 , n89368 );
buf ( n89370 , n89369 );
nand ( n89371 , n89357 , n89370 );
buf ( n89372 , n89371 );
buf ( n89373 , n89372 );
nand ( n89374 , n89356 , n89373 );
buf ( n89375 , n89374 );
buf ( n89376 , n89375 );
not ( n89377 , n89376 );
buf ( n89378 , n37919 );
not ( n89379 , n89378 );
buf ( n89380 , n41947 );
not ( n89381 , n89380 );
buf ( n89382 , n37589 );
not ( n89383 , n89382 );
or ( n89384 , n89381 , n89383 );
buf ( n89385 , n39489 );
buf ( n89386 , n41925 );
nand ( n89387 , n89385 , n89386 );
buf ( n89388 , n89387 );
buf ( n89389 , n89388 );
nand ( n89390 , n89384 , n89389 );
buf ( n89391 , n89390 );
buf ( n89392 , n89391 );
not ( n89393 , n89392 );
or ( n89394 , n89379 , n89393 );
buf ( n89395 , n37872 );
and ( n89396 , n42891 , n41925 );
not ( n89397 , n42891 );
and ( n89398 , n89397 , n37879 );
nor ( n89399 , n89396 , n89398 );
buf ( n89400 , n89399 );
nand ( n89401 , n89395 , n89400 );
buf ( n89402 , n89401 );
buf ( n89403 , n89402 );
nand ( n89404 , n89394 , n89403 );
buf ( n89405 , n89404 );
buf ( n89406 , n89405 );
not ( n89407 , n89406 );
buf ( n89408 , n89407 );
buf ( n89409 , n89408 );
not ( n89410 , n89409 );
or ( n89411 , n89377 , n89410 );
buf ( n89412 , n89405 );
buf ( n89413 , n89375 );
not ( n89414 , n89413 );
buf ( n89415 , n89414 );
buf ( n89416 , n89415 );
nand ( n89417 , n89412 , n89416 );
buf ( n89418 , n89417 );
buf ( n89419 , n89418 );
nand ( n89420 , n89411 , n89419 );
buf ( n89421 , n89420 );
not ( n89422 , n44679 );
buf ( n89423 , n39688 );
not ( n89424 , n89423 );
buf ( n89425 , n89424 );
buf ( n89426 , n89425 );
not ( n89427 , n89426 );
buf ( n89428 , n36932 );
not ( n89429 , n89428 );
or ( n89430 , n89427 , n89429 );
buf ( n89431 , n42062 );
buf ( n89432 , n39688 );
nand ( n89433 , n89431 , n89432 );
buf ( n89434 , n89433 );
buf ( n89435 , n89434 );
nand ( n89436 , n89430 , n89435 );
buf ( n89437 , n89436 );
not ( n89438 , n89437 );
or ( n89439 , n89422 , n89438 );
not ( n89440 , n89184 );
nand ( n89441 , n89440 , n45158 );
nand ( n89442 , n89439 , n89441 );
buf ( n89443 , n89442 );
not ( n89444 , n89443 );
buf ( n89445 , n89444 );
and ( n89446 , n89421 , n89445 );
not ( n89447 , n89421 );
and ( n89448 , n89447 , n89442 );
nor ( n89449 , n89446 , n89448 );
not ( n89450 , n89449 );
not ( n89451 , n89450 );
or ( n89452 , n89339 , n89451 );
or ( n89453 , n89450 , n89338 );
nand ( n89454 , n89452 , n89453 );
not ( n89455 , n89454 );
or ( n89456 , n89313 , n89455 );
or ( n89457 , n89454 , n89312 );
nand ( n89458 , n89456 , n89457 );
xor ( n89459 , n89306 , n89458 );
not ( n89460 , n89459 );
nor ( n89461 , n88958 , n89149 , n89460 );
not ( n89462 , n89461 );
not ( n89463 , n89149 );
nand ( n89464 , n88958 , n89463 , n89460 );
not ( n89465 , n88958 );
buf ( n89466 , n89149 );
nand ( n89467 , n89465 , n89466 , n89460 );
nand ( n89468 , n89466 , n88958 , n89459 );
nand ( n89469 , n89462 , n89464 , n89467 , n89468 );
not ( n89470 , n89469 );
not ( n89471 , n88330 );
nand ( n89472 , n89471 , n88344 );
not ( n89473 , n89472 );
not ( n89474 , n88365 );
or ( n89475 , n89473 , n89474 );
buf ( n89476 , n88347 );
buf ( n89477 , n88330 );
nand ( n89478 , n89476 , n89477 );
buf ( n89479 , n89478 );
nand ( n89480 , n89475 , n89479 );
buf ( n89481 , n89480 );
buf ( n89482 , n88361 );
not ( n89483 , n89482 );
buf ( n89484 , n42521 );
not ( n89485 , n89484 );
or ( n89486 , n89483 , n89485 );
buf ( n89487 , n42530 );
buf ( n89488 , n89351 );
nand ( n89489 , n89487 , n89488 );
buf ( n89490 , n89489 );
buf ( n89491 , n89490 );
nand ( n89492 , n89486 , n89491 );
buf ( n89493 , n89492 );
buf ( n89494 , n89493 );
not ( n89495 , n89399 );
not ( n89496 , n41905 );
or ( n89497 , n89495 , n89496 );
buf ( n89498 , n37872 );
buf ( n89499 , n88323 );
nand ( n89500 , n89498 , n89499 );
buf ( n89501 , n89500 );
nand ( n89502 , n89497 , n89501 );
buf ( n89503 , n89502 );
xor ( n89504 , n89494 , n89503 );
not ( n89505 , n42004 );
nand ( n89506 , n89505 , n89067 );
nand ( n89507 , C1 , n89506 );
buf ( n89508 , n89507 );
xor ( n89509 , n89504 , n89508 );
buf ( n89510 , n89509 );
buf ( n89511 , n89510 );
xor ( n89512 , n89481 , n89511 );
buf ( n89513 , n39374 );
not ( n89514 , n89513 );
buf ( n89515 , n89246 );
not ( n89516 , n89515 );
or ( n89517 , n89514 , n89516 );
buf ( n89518 , n88576 );
buf ( n89519 , n39395 );
nand ( n89520 , n89518 , n89519 );
buf ( n89521 , n89520 );
buf ( n89522 , n89521 );
nand ( n89523 , n89517 , n89522 );
buf ( n89524 , n89523 );
buf ( n89525 , n89524 );
xor ( n89526 , n89512 , n89525 );
buf ( n89527 , n89526 );
buf ( n89528 , n89527 );
xor ( n89529 , n88967 , n88992 );
xor ( n89530 , n89529 , n88999 );
buf ( n89531 , n89530 );
buf ( n89532 , n89531 );
xor ( n89533 , n89528 , n89532 );
xor ( n89534 , n89283 , n89288 );
xor ( n89535 , n89534 , n89297 );
buf ( n89536 , n89535 );
buf ( n89537 , n89536 );
xor ( n89538 , n89533 , n89537 );
buf ( n89539 , n89538 );
buf ( n89540 , n89539 );
buf ( n89541 , n88612 );
not ( n89542 , n89541 );
buf ( n89543 , n88622 );
not ( n89544 , n89543 );
or ( n89545 , n89542 , n89544 );
buf ( n89546 , n88639 );
nand ( n89547 , n89545 , n89546 );
buf ( n89548 , n89547 );
buf ( n89549 , n89548 );
buf ( n89550 , n88621 );
buf ( n89551 , n88611 );
nand ( n89552 , n89550 , n89551 );
buf ( n89553 , n89552 );
buf ( n89554 , n89553 );
nand ( n89555 , n89549 , n89554 );
buf ( n89556 , n89555 );
buf ( n89557 , n89556 );
xor ( n89558 , n89540 , n89557 );
nand ( n89559 , n88940 , n88944 );
nand ( n89560 , n88939 , n88945 );
nand ( n89561 , n89559 , n89560 );
xor ( n89562 , n89561 , n88954 );
buf ( n89563 , n89562 );
and ( n89564 , n89558 , n89563 );
and ( n89565 , n89540 , n89557 );
or ( n89566 , n89564 , n89565 );
buf ( n89567 , n89566 );
buf ( n89568 , n89567 );
buf ( n89569 , n88768 );
buf ( n89570 , n88752 );
nor ( n89571 , n89569 , n89570 );
buf ( n89572 , n89571 );
buf ( n89573 , n89572 );
buf ( n89574 , n88774 );
or ( n89575 , n89573 , n89574 );
buf ( n89576 , n88768 );
buf ( n89577 , n88752 );
nand ( n89578 , n89576 , n89577 );
buf ( n89579 , n89578 );
buf ( n89580 , n89579 );
nand ( n89581 , n89575 , n89580 );
buf ( n89582 , n89581 );
buf ( n89583 , n89582 );
not ( n89584 , n88396 );
nand ( n89585 , n89584 , n88366 );
not ( n89586 , n89585 );
not ( n89587 , n88467 );
or ( n89588 , n89586 , n89587 );
not ( n89589 , n88366 );
nand ( n89590 , n89589 , n88396 );
nand ( n89591 , n89588 , n89590 );
buf ( n89592 , n88546 );
buf ( n89593 , n88510 );
nand ( n89594 , n89592 , n89593 );
buf ( n89595 , n89594 );
buf ( n89596 , n89595 );
buf ( n89597 , n88490 );
and ( n89598 , n89596 , n89597 );
buf ( n89599 , n88541 );
buf ( n89600 , n88507 );
and ( n89601 , n89599 , n89600 );
buf ( n89602 , n89601 );
buf ( n89603 , n89602 );
nor ( n89604 , n89598 , n89603 );
buf ( n89605 , n89604 );
buf ( n89606 , n89605 );
not ( n89607 , n89606 );
buf ( n89608 , n89607 );
buf ( n89609 , n89608 );
not ( n89610 , n89609 );
buf ( n89611 , n88685 );
buf ( n89612 , n44586 );
and ( n89613 , n89611 , n89612 );
buf ( n89614 , n89031 );
not ( n89615 , n89614 );
buf ( n89616 , n43906 );
nor ( n89617 , n89615 , n89616 );
buf ( n89618 , n89617 );
buf ( n89619 , n89618 );
nor ( n89620 , n89613 , n89619 );
buf ( n89621 , n89620 );
buf ( n89622 , n89621 );
not ( n89623 , n89622 );
or ( n89624 , n89610 , n89623 );
buf ( n89625 , n89621 );
not ( n89626 , n89625 );
buf ( n89627 , n89626 );
buf ( n89628 , n89627 );
buf ( n89629 , n89605 );
nand ( n89630 , n89628 , n89629 );
buf ( n89631 , n89630 );
buf ( n89632 , n89631 );
nand ( n89633 , n89624 , n89632 );
buf ( n89634 , n89633 );
xor ( n89635 , n89591 , n89634 );
buf ( n89636 , n89635 );
xor ( n89637 , n89583 , n89636 );
not ( n89638 , n88555 );
not ( n89639 , n88474 );
buf ( n89640 , n89639 );
buf ( n89641 , n88549 );
nand ( n89642 , n89640 , n89641 );
buf ( n89643 , n89642 );
not ( n89644 , n89643 );
or ( n89645 , n89638 , n89644 );
not ( n89646 , n89639 );
nand ( n89647 , n89646 , n88548 );
nand ( n89648 , n89645 , n89647 );
buf ( n89649 , n89648 );
and ( n89650 , n89637 , n89649 );
and ( n89651 , n89583 , n89636 );
or ( n89652 , n89650 , n89651 );
buf ( n89653 , n89652 );
buf ( n89654 , n89653 );
not ( n89655 , n89608 );
not ( n89656 , n89627 );
or ( n89657 , n89655 , n89656 );
not ( n89658 , n89605 );
not ( n89659 , n89621 );
or ( n89660 , n89658 , n89659 );
nand ( n89661 , n89660 , n89591 );
nand ( n89662 , n89657 , n89661 );
buf ( n89663 , n42566 );
not ( n89664 , n89663 );
buf ( n89665 , n25160 );
not ( n89666 , n89665 );
buf ( n89667 , n40067 );
not ( n89668 , n89667 );
or ( n89669 , n89666 , n89668 );
buf ( n89670 , n36427 );
buf ( n89671 , n42581 );
nand ( n89672 , n89670 , n89671 );
buf ( n89673 , n89672 );
buf ( n89674 , n89673 );
nand ( n89675 , n89669 , n89674 );
buf ( n89676 , n89675 );
buf ( n89677 , n89676 );
not ( n89678 , n89677 );
or ( n89679 , n89664 , n89678 );
buf ( n89680 , n88857 );
buf ( n89681 , n42631 );
nand ( n89682 , n89680 , n89681 );
buf ( n89683 , n89682 );
buf ( n89684 , n89683 );
nand ( n89685 , n89679 , n89684 );
buf ( n89686 , n89685 );
buf ( n89687 , n51912 );
not ( n89688 , n89687 );
buf ( n89689 , n88899 );
not ( n89690 , n89689 );
or ( n89691 , n89688 , n89690 );
buf ( n89692 , n88143 );
not ( n89693 , n89692 );
buf ( n89694 , n44316 );
not ( n89695 , n89694 );
or ( n89696 , n89693 , n89695 );
buf ( n89697 , n39522 );
buf ( n89698 , n37475 );
nand ( n89699 , n89697 , n89698 );
buf ( n89700 , n89699 );
buf ( n89701 , n89700 );
nand ( n89702 , n89696 , n89701 );
buf ( n89703 , n89702 );
buf ( n89704 , n89703 );
buf ( n89705 , n37452 );
nand ( n89706 , n89704 , n89705 );
buf ( n89707 , n89706 );
buf ( n89708 , n89707 );
nand ( n89709 , n89691 , n89708 );
buf ( n89710 , n89709 );
buf ( n89711 , n89710 );
buf ( n89712 , n37403 );
not ( n89713 , n89712 );
buf ( n89714 , n88926 );
not ( n89715 , n89714 );
or ( n89716 , n89713 , n89715 );
buf ( n89717 , n88089 );
not ( n89718 , n89717 );
buf ( n89719 , n37295 );
not ( n89720 , n89719 );
or ( n89721 , n89718 , n89720 );
buf ( n89722 , n49179 );
buf ( n89723 , n37329 );
nand ( n89724 , n89722 , n89723 );
buf ( n89725 , n89724 );
buf ( n89726 , n89725 );
nand ( n89727 , n89721 , n89726 );
buf ( n89728 , n89727 );
buf ( n89729 , n89728 );
buf ( n89730 , n38150 );
nand ( n89731 , n89729 , n89730 );
buf ( n89732 , n89731 );
buf ( n89733 , n89732 );
nand ( n89734 , n89716 , n89733 );
buf ( n89735 , n89734 );
buf ( n89736 , n89735 );
xor ( n89737 , n89711 , n89736 );
xor ( n89738 , n89494 , n89503 );
and ( n89739 , n89738 , n89508 );
and ( n89740 , n89494 , n89503 );
or ( n89741 , n89739 , n89740 );
buf ( n89742 , n89741 );
buf ( n89743 , n89742 );
xor ( n89744 , n89737 , n89743 );
buf ( n89745 , n89744 );
xor ( n89746 , n89686 , n89745 );
xor ( n89747 , n89481 , n89511 );
and ( n89748 , n89747 , n89525 );
and ( n89749 , n89481 , n89511 );
or ( n89750 , n89748 , n89749 );
buf ( n89751 , n89750 );
xor ( n89752 , n89746 , n89751 );
xor ( n89753 , n89662 , n89752 );
xor ( n89754 , n89528 , n89532 );
and ( n89755 , n89754 , n89537 );
and ( n89756 , n89528 , n89532 );
or ( n89757 , n89755 , n89756 );
buf ( n89758 , n89757 );
xor ( n89759 , n89753 , n89758 );
buf ( n89760 , n89759 );
not ( n89761 , n89760 );
buf ( n89762 , n89761 );
buf ( n89763 , n89762 );
and ( n89764 , n89654 , n89763 );
not ( n89765 , n89654 );
buf ( n89766 , n89759 );
and ( n89767 , n89765 , n89766 );
nor ( n89768 , n89764 , n89767 );
buf ( n89769 , n89768 );
buf ( n89770 , n89769 );
and ( n89771 , n89568 , n89770 );
not ( n89772 , n89568 );
buf ( n89773 , n89769 );
not ( n89774 , n89773 );
buf ( n89775 , n89774 );
buf ( n89776 , n89775 );
and ( n89777 , n89772 , n89776 );
nor ( n89778 , n89771 , n89777 );
buf ( n89779 , n89778 );
not ( n89780 , n89779 );
not ( n89781 , n89780 );
or ( n89782 , n89470 , n89781 );
not ( n89783 , n89469 );
nand ( n89784 , n89779 , n89783 );
nand ( n89785 , n89782 , n89784 );
xor ( n89786 , n89583 , n89636 );
xor ( n89787 , n89786 , n89649 );
buf ( n89788 , n89787 );
not ( n89789 , n89788 );
xor ( n89790 , n88701 , n88778 );
and ( n89791 , n89790 , n88784 );
and ( n89792 , n88701 , n88778 );
or ( n89793 , n89791 , n89792 );
buf ( n89794 , n89793 );
not ( n89795 , n89794 );
nand ( n89796 , n89789 , n89795 );
not ( n89797 , n89796 );
not ( n89798 , n88644 );
not ( n89799 , n88557 );
nand ( n89800 , n88563 , n89799 );
not ( n89801 , n89800 );
or ( n89802 , n89798 , n89801 );
nand ( n89803 , n88562 , n88557 );
nand ( n89804 , n89802 , n89803 );
not ( n89805 , n89804 );
or ( n89806 , n89797 , n89805 );
nand ( n89807 , n89788 , n89794 );
nand ( n89808 , n89806 , n89807 );
buf ( n89809 , n89808 );
not ( n89810 , n89809 );
buf ( n89811 , n89810 );
and ( n89812 , n89785 , n89811 );
not ( n89813 , n89785 );
and ( n89814 , n89813 , n89808 );
nor ( n89815 , n89812 , n89814 );
xor ( n89816 , n89540 , n89557 );
xor ( n89817 , n89816 , n89563 );
buf ( n89818 , n89817 );
buf ( n89819 , n89818 );
xor ( n89820 , n88652 , n88787 );
and ( n89821 , n89820 , n88794 );
and ( n89822 , n88652 , n88787 );
or ( n89823 , n89821 , n89822 );
buf ( n89824 , n89823 );
buf ( n89825 , n89824 );
xor ( n89826 , n89819 , n89825 );
not ( n89827 , n89794 );
not ( n89828 , n89788 );
not ( n89829 , n89828 );
or ( n89830 , n89827 , n89829 );
nand ( n89831 , n89795 , n89788 );
nand ( n89832 , n89830 , n89831 );
and ( n89833 , n89832 , n89804 );
not ( n89834 , n89832 );
not ( n89835 , n89804 );
and ( n89836 , n89834 , n89835 );
nor ( n89837 , n89833 , n89836 );
buf ( n89838 , n89837 );
and ( n89839 , n89826 , n89838 );
and ( n89840 , n89819 , n89825 );
or ( n89841 , n89839 , n89840 );
buf ( n89842 , n89841 );
nor ( n89843 , n89815 , n89842 );
buf ( n89844 , n89843 );
not ( n89845 , n89844 );
buf ( n89846 , n89845 );
xor ( n89847 , n89819 , n89825 );
xor ( n89848 , n89847 , n89838 );
buf ( n89849 , n89848 );
xor ( n89850 , n88646 , n88797 );
and ( n89851 , n89850 , n88805 );
and ( n89852 , n88646 , n88797 );
or ( n89853 , n89851 , n89852 );
buf ( n89854 , n89853 );
or ( n89855 , n89849 , n89854 );
nand ( n89856 , n89846 , n89855 );
not ( n89857 , n41644 );
not ( n89858 , n41704 );
or ( n89859 , n89857 , n89858 );
nand ( n89860 , n89859 , n89206 );
not ( n89861 , n89728 );
not ( n89862 , n37403 );
or ( n89863 , n89861 , n89862 );
not ( n89864 , n37416 );
not ( n89865 , n43143 );
not ( n89866 , n37330 );
or ( n89867 , n89865 , n89866 );
buf ( n89868 , n37271 );
buf ( n89869 , n37329 );
nand ( n89870 , n89868 , n89869 );
buf ( n89871 , n89870 );
nand ( n89872 , n89867 , n89871 );
nand ( n89873 , n89864 , n89872 );
nand ( n89874 , n89863 , n89873 );
xor ( n89875 , n89860 , n89874 );
buf ( n89876 , n89068 );
not ( n89877 , n89876 );
buf ( n89878 , n89123 );
not ( n89879 , n89878 );
buf ( n89880 , n89879 );
buf ( n89881 , n89880 );
not ( n89882 , n89881 );
or ( n89883 , n89877 , n89882 );
buf ( n89884 , n89105 );
nand ( n89885 , n89883 , n89884 );
buf ( n89886 , n89885 );
not ( n89887 , n89068 );
nand ( n89888 , n89123 , n89887 );
nand ( n89889 , n89886 , n89888 );
and ( n89890 , n89875 , n89889 );
and ( n89891 , n89860 , n89874 );
or ( n89892 , n89890 , n89891 );
buf ( n89893 , n89375 );
not ( n89894 , n89893 );
buf ( n89895 , n89405 );
not ( n89896 , n89895 );
or ( n89897 , n89894 , n89896 );
buf ( n89898 , n89442 );
buf ( n89899 , n89408 );
buf ( n89900 , n89415 );
nand ( n89901 , n89899 , n89900 );
buf ( n89902 , n89901 );
buf ( n89903 , n89902 );
nand ( n89904 , n89898 , n89903 );
buf ( n89905 , n89904 );
buf ( n89906 , n89905 );
nand ( n89907 , n89897 , n89906 );
buf ( n89908 , n89907 );
not ( n89909 , n89908 );
buf ( n89910 , n43909 );
not ( n89911 , n89910 );
buf ( n89912 , n25184 );
not ( n89913 , n89912 );
buf ( n89914 , n36054 );
not ( n89915 , n89914 );
or ( n89916 , n89913 , n89915 );
buf ( n89917 , n43851 );
buf ( n89918 , n25183 );
nand ( n89919 , n89917 , n89918 );
buf ( n89920 , n89919 );
buf ( n89921 , n89920 );
nand ( n89922 , n89916 , n89921 );
buf ( n89923 , n89922 );
buf ( n89924 , n89923 );
not ( n89925 , n89924 );
or ( n89926 , n89911 , n89925 );
buf ( n89927 , n89045 );
buf ( n89928 , n44586 );
nand ( n89929 , n89927 , n89928 );
buf ( n89930 , n89929 );
buf ( n89931 , n89930 );
nand ( n89932 , n89926 , n89931 );
buf ( n89933 , n89932 );
not ( n89934 , n89933 );
or ( n89935 , n89909 , n89934 );
not ( n89936 , n89908 );
not ( n89937 , n89936 );
not ( n89938 , n89933 );
not ( n89939 , n89938 );
or ( n89940 , n89937 , n89939 );
buf ( n89941 , n42854 );
buf ( n89942 , n42196 );
buf ( n89943 , n36363 );
and ( n89944 , n89942 , n89943 );
not ( n89945 , n89942 );
buf ( n89946 , n38837 );
and ( n89947 , n89945 , n89946 );
nor ( n89948 , n89944 , n89947 );
buf ( n89949 , n89948 );
buf ( n89950 , n89949 );
or ( n89951 , n89941 , n89950 );
nand ( n89952 , C1 , n89951 );
buf ( n89953 , n89952 );
buf ( n89954 , n89953 );
buf ( n89955 , n89369 );
not ( n89956 , n89955 );
buf ( n89957 , n36104 );
not ( n89958 , n89957 );
or ( n89959 , n89956 , n89958 );
buf ( n89960 , n29290 );
buf ( n89961 , n33077 );
and ( n89962 , n89960 , n89961 );
not ( n89963 , n89960 );
buf ( n89964 , n39478 );
and ( n89965 , n89963 , n89964 );
or ( n89966 , n89962 , n89965 );
buf ( n89967 , n89966 );
buf ( n89968 , n89967 );
not ( n89969 , n89968 );
buf ( n89970 , n32972 );
nand ( n89971 , n89969 , n89970 );
buf ( n89972 , n89971 );
buf ( n89973 , n89972 );
nand ( n89974 , n89959 , n89973 );
buf ( n89975 , n89974 );
buf ( n89976 , n89975 );
xor ( n89977 , n89954 , n89976 );
buf ( n89978 , n36985 );
buf ( n89979 , n89437 );
not ( n89980 , n89979 );
buf ( n89981 , n89980 );
buf ( n89982 , n89981 );
or ( n89983 , n89978 , n89982 );
buf ( n89984 , n37005 );
buf ( n89985 , n38851 );
buf ( n89986 , n39235 );
and ( n89987 , n89985 , n89986 );
not ( n89988 , n89985 );
buf ( n89989 , n36932 );
and ( n89990 , n89988 , n89989 );
nor ( n89991 , n89987 , n89990 );
buf ( n89992 , n89991 );
buf ( n89993 , n89992 );
or ( n89994 , n89984 , n89993 );
nand ( n89995 , n89983 , n89994 );
buf ( n89996 , n89995 );
buf ( n89997 , n89996 );
xor ( n89998 , n89977 , n89997 );
buf ( n89999 , n89998 );
nand ( n90000 , n89940 , n89999 );
nand ( n90001 , n89935 , n90000 );
xor ( n90002 , n89892 , n90001 );
buf ( n90003 , n37875 );
not ( n90004 , n90003 );
buf ( n90005 , n37892 );
not ( n90006 , n90005 );
buf ( n90007 , n37786 );
not ( n90008 , n90007 );
or ( n90009 , n90006 , n90008 );
buf ( n90010 , n37792 );
buf ( n90011 , n41890 );
nand ( n90012 , n90010 , n90011 );
buf ( n90013 , n90012 );
buf ( n90014 , n90013 );
nand ( n90015 , n90009 , n90014 );
buf ( n90016 , n90015 );
buf ( n90017 , n90016 );
not ( n90018 , n90017 );
or ( n90019 , n90004 , n90018 );
buf ( n90020 , n37892 );
not ( n90021 , n90020 );
buf ( n90022 , n42597 );
not ( n90023 , n90022 );
or ( n90024 , n90021 , n90023 );
buf ( n90025 , n50925 );
not ( n90026 , n90025 );
buf ( n90027 , n41890 );
nand ( n90028 , n90026 , n90027 );
buf ( n90029 , n90028 );
buf ( n90030 , n90029 );
nand ( n90031 , n90024 , n90030 );
buf ( n90032 , n90031 );
buf ( n90033 , n90032 );
buf ( n90034 , n37922 );
nand ( n90035 , n90033 , n90034 );
buf ( n90036 , n90035 );
buf ( n90037 , n90036 );
nand ( n90038 , n90019 , n90037 );
buf ( n90039 , n90038 );
buf ( n90040 , n90039 );
buf ( n90041 , n38775 );
not ( n90042 , n90041 );
buf ( n90043 , n38413 );
not ( n90044 , n90043 );
buf ( n90045 , n38221 );
not ( n90046 , n90045 );
or ( n90047 , n90044 , n90046 );
buf ( n90048 , n42941 );
buf ( n90049 , n38420 );
nand ( n90050 , n90048 , n90049 );
buf ( n90051 , n90050 );
buf ( n90052 , n90051 );
nand ( n90053 , n90047 , n90052 );
buf ( n90054 , n90053 );
buf ( n90055 , n90054 );
not ( n90056 , n90055 );
or ( n90057 , n90042 , n90056 );
not ( n90058 , n38413 );
not ( n90059 , n37970 );
or ( n90060 , n90058 , n90059 );
nand ( n90061 , n42929 , n38420 );
nand ( n90062 , n90060 , n90061 );
nand ( n90063 , n90062 , n38758 );
buf ( n90064 , n90063 );
nand ( n90065 , n90057 , n90064 );
buf ( n90066 , n90065 );
buf ( n90067 , n90066 );
xor ( n90068 , n90040 , n90067 );
xor ( n90069 , n89954 , n89976 );
and ( n90070 , n90069 , n89997 );
and ( n90071 , n89954 , n89976 );
or ( n90072 , n90070 , n90071 );
buf ( n90073 , n90072 );
buf ( n90074 , n90073 );
xor ( n90075 , n90068 , n90074 );
buf ( n90076 , n90075 );
xor ( n90077 , n90002 , n90076 );
buf ( n90078 , n90077 );
buf ( n90079 , n89017 );
buf ( n90080 , n89047 );
or ( n90081 , n90079 , n90080 );
buf ( n90082 , n89129 );
nand ( n90083 , n90081 , n90082 );
buf ( n90084 , n90083 );
buf ( n90085 , n90084 );
buf ( n90086 , n89017 );
buf ( n90087 , n89047 );
nand ( n90088 , n90086 , n90087 );
buf ( n90089 , n90088 );
buf ( n90090 , n90089 );
and ( n90091 , n90085 , n90090 );
buf ( n90092 , n90091 );
buf ( n90093 , n90092 );
not ( n90094 , n90093 );
buf ( n90095 , n90094 );
buf ( n90096 , n90095 );
not ( n90097 , n90096 );
xor ( n90098 , n89860 , n89874 );
xor ( n90099 , n90098 , n89889 );
buf ( n90100 , n90099 );
not ( n90101 , n90100 );
or ( n90102 , n90097 , n90101 );
buf ( n90103 , n39374 );
not ( n90104 , n90103 );
buf ( n90105 , n39000 );
not ( n90106 , n90105 );
buf ( n90107 , n42360 );
not ( n90108 , n90107 );
or ( n90109 , n90106 , n90108 );
buf ( n90110 , n50876 );
buf ( n90111 , n38997 );
nand ( n90112 , n90110 , n90111 );
buf ( n90113 , n90112 );
buf ( n90114 , n90113 );
nand ( n90115 , n90109 , n90114 );
buf ( n90116 , n90115 );
buf ( n90117 , n90116 );
not ( n90118 , n90117 );
or ( n90119 , n90104 , n90118 );
buf ( n90120 , n89260 );
buf ( n90121 , n39395 );
nand ( n90122 , n90120 , n90121 );
buf ( n90123 , n90122 );
buf ( n90124 , n90123 );
nand ( n90125 , n90119 , n90124 );
buf ( n90126 , n90125 );
buf ( n90127 , n89068 );
buf ( n90128 , n89098 );
not ( n90129 , n90128 );
buf ( n90130 , n43389 );
not ( n90131 , n90130 );
or ( n90132 , n90129 , n90131 );
buf ( n90133 , n43400 );
not ( n90134 , n90133 );
buf ( n90135 , n45394 );
not ( n90136 , n90135 );
or ( n90137 , n90134 , n90136 );
buf ( n90138 , n39205 );
buf ( n90139 , n43371 );
nand ( n90140 , n90138 , n90139 );
buf ( n90141 , n90140 );
buf ( n90142 , n90141 );
nand ( n90143 , n90137 , n90142 );
buf ( n90144 , n90143 );
buf ( n90145 , n90144 );
buf ( n90146 , n43414 );
nand ( n90147 , n90145 , n90146 );
buf ( n90148 , n90147 );
buf ( n90149 , n90148 );
nand ( n90150 , n90132 , n90149 );
buf ( n90151 , n90150 );
buf ( n90152 , n90151 );
xor ( n90153 , n90127 , n90152 );
and ( n90154 , n28306 , n60583 );
not ( n90155 , n28306 );
and ( n90156 , n90155 , n36533 );
or ( n90157 , n90154 , n90156 );
not ( n90158 , n90157 );
not ( n90159 , n39816 );
or ( n90160 , n90158 , n90159 );
not ( n90161 , n89119 );
nand ( n90162 , n90161 , n39806 );
nand ( n90163 , n90160 , n90162 );
buf ( n90164 , n90163 );
not ( n90165 , n90164 );
buf ( n90166 , n90165 );
buf ( n90167 , n90166 );
xor ( n90168 , n90153 , n90167 );
buf ( n90169 , n90168 );
xor ( n90170 , n90126 , n90169 );
xor ( n90171 , n89711 , n89736 );
and ( n90172 , n90171 , n89743 );
and ( n90173 , n89711 , n89736 );
or ( n90174 , n90172 , n90173 );
buf ( n90175 , n90174 );
xnor ( n90176 , n90170 , n90175 );
buf ( n90177 , n90176 );
buf ( n90178 , n90099 );
not ( n90179 , n90178 );
buf ( n90180 , n90092 );
nand ( n90181 , n90179 , n90180 );
buf ( n90182 , n90181 );
buf ( n90183 , n90182 );
nand ( n90184 , n90177 , n90183 );
buf ( n90185 , n90184 );
buf ( n90186 , n90185 );
nand ( n90187 , n90102 , n90186 );
buf ( n90188 , n90187 );
buf ( n90189 , n90188 );
xor ( n90190 , n90078 , n90189 );
buf ( n90191 , n37403 );
not ( n90192 , n90191 );
buf ( n90193 , n89872 );
not ( n90194 , n90193 );
or ( n90195 , n90192 , n90194 );
buf ( n90196 , n37330 );
not ( n90197 , n90196 );
buf ( n90198 , n53044 );
not ( n90199 , n90198 );
or ( n90200 , n90197 , n90199 );
buf ( n90201 , n38247 );
buf ( n90202 , n37329 );
nand ( n90203 , n90201 , n90202 );
buf ( n90204 , n90203 );
buf ( n90205 , n90204 );
nand ( n90206 , n90200 , n90205 );
buf ( n90207 , n90206 );
buf ( n90208 , n90207 );
buf ( n90209 , n38150 );
nand ( n90210 , n90208 , n90209 );
buf ( n90211 , n90210 );
buf ( n90212 , n90211 );
nand ( n90213 , n90195 , n90212 );
buf ( n90214 , n90213 );
buf ( n90215 , n39395 );
not ( n90216 , n90215 );
buf ( n90217 , n90116 );
not ( n90218 , n90217 );
or ( n90219 , n90216 , n90218 );
buf ( n90220 , n39000 );
not ( n90221 , n90220 );
buf ( n90222 , n38098 );
not ( n90223 , n90222 );
or ( n90224 , n90221 , n90223 );
buf ( n90225 , n39340 );
buf ( n90226 , n38997 );
nand ( n90227 , n90225 , n90226 );
buf ( n90228 , n90227 );
buf ( n90229 , n90228 );
nand ( n90230 , n90224 , n90229 );
buf ( n90231 , n90230 );
buf ( n90232 , n90231 );
buf ( n90233 , n39374 );
nand ( n90234 , n90232 , n90233 );
buf ( n90235 , n90234 );
buf ( n90236 , n90235 );
nand ( n90237 , n90219 , n90236 );
buf ( n90238 , n90237 );
not ( n90239 , n90238 );
xor ( n90240 , n90214 , n90239 );
buf ( n90241 , n43283 );
buf ( n90242 , n38798 );
not ( n90243 , n90242 );
buf ( n90244 , n41951 );
not ( n90245 , n90244 );
and ( n90246 , n90243 , n90245 );
buf ( n90247 , n38834 );
buf ( n90248 , n41951 );
and ( n90249 , n90247 , n90248 );
nor ( n90250 , n90246 , n90249 );
buf ( n90251 , n90250 );
buf ( n90252 , n90251 );
or ( n90253 , n90241 , n90252 );
nand ( n90254 , C1 , n90253 );
buf ( n90255 , n90254 );
not ( n90256 , n90255 );
buf ( n90257 , n90256 );
buf ( n90258 , n90157 );
not ( n90259 , n90258 );
buf ( n90260 , n39806 );
not ( n90261 , n90260 );
or ( n90262 , n90259 , n90261 );
buf ( n90263 , n39816 );
buf ( n90264 , n28723 );
not ( n90265 , n90264 );
buf ( n90266 , n60583 );
not ( n90267 , n90266 );
or ( n90268 , n90265 , n90267 );
buf ( n90269 , n39729 );
not ( n90270 , n28723 );
buf ( n90271 , n90270 );
nand ( n90272 , n90269 , n90271 );
buf ( n90273 , n90272 );
buf ( n90274 , n90273 );
nand ( n90275 , n90268 , n90274 );
buf ( n90276 , n90275 );
buf ( n90277 , n90276 );
nand ( n90278 , n90263 , n90277 );
buf ( n90279 , n90278 );
buf ( n90280 , n90279 );
nand ( n90281 , n90262 , n90280 );
buf ( n90282 , n90281 );
buf ( n90283 , n90282 );
xor ( n90284 , n90257 , n90283 );
not ( n90285 , n51912 );
buf ( n90286 , n88143 );
buf ( n90287 , n37692 );
and ( n90288 , n90286 , n90287 );
not ( n90289 , n90286 );
buf ( n90290 , n37717 );
and ( n90291 , n90289 , n90290 );
nor ( n90292 , n90288 , n90291 );
buf ( n90293 , n90292 );
not ( n90294 , n90293 );
or ( n90295 , n90285 , n90294 );
buf ( n90296 , n37476 );
not ( n90297 , n90296 );
buf ( n90298 , n49178 );
not ( n90299 , n90298 );
or ( n90300 , n90297 , n90299 );
buf ( n90301 , n38287 );
buf ( n90302 , n37475 );
nand ( n90303 , n90301 , n90302 );
buf ( n90304 , n90303 );
buf ( n90305 , n90304 );
nand ( n90306 , n90300 , n90305 );
buf ( n90307 , n90306 );
nand ( n90308 , n37452 , n90307 );
nand ( n90309 , n90295 , n90308 );
buf ( n90310 , n90309 );
xor ( n90311 , n90284 , n90310 );
buf ( n90312 , n90311 );
xnor ( n90313 , n90240 , n90312 );
not ( n90314 , n43909 );
buf ( n90315 , n25184 );
buf ( n90316 , n39005 );
and ( n90317 , n90315 , n90316 );
not ( n90318 , n90315 );
buf ( n90319 , n35971 );
and ( n90320 , n90318 , n90319 );
nor ( n90321 , n90317 , n90320 );
buf ( n90322 , n90321 );
not ( n90323 , n90322 );
or ( n90324 , n90314 , n90323 );
buf ( n90325 , n89923 );
buf ( n90326 , n44586 );
nand ( n90327 , n90325 , n90326 );
buf ( n90328 , n90327 );
nand ( n90329 , n90324 , n90328 );
not ( n90330 , n89887 );
not ( n90331 , n90166 );
or ( n90332 , n90330 , n90331 );
nand ( n90333 , n90332 , n90151 );
buf ( n90334 , n90163 );
buf ( n90335 , n89068 );
nand ( n90336 , n90334 , n90335 );
buf ( n90337 , n90336 );
nand ( n90338 , n90333 , n90337 );
xor ( n90339 , n90329 , n90338 );
buf ( n90340 , n36985 );
buf ( n90341 , n89992 );
or ( n90342 , n90340 , n90341 );
buf ( n90343 , n37005 );
buf ( n90344 , n42062 );
buf ( n90345 , n39742 );
and ( n90346 , n90344 , n90345 );
not ( n90347 , n90344 );
buf ( n90348 , n38824 );
not ( n90349 , n90348 );
buf ( n90350 , n90349 );
buf ( n90351 , n90350 );
and ( n90352 , n90347 , n90351 );
nor ( n90353 , n90346 , n90352 );
buf ( n90354 , n90353 );
buf ( n90355 , n90354 );
or ( n90356 , n90343 , n90355 );
nand ( n90357 , n90342 , n90356 );
buf ( n90358 , n90357 );
buf ( n90359 , n90144 );
not ( n90360 , n90359 );
buf ( n90361 , n43389 );
not ( n90362 , n90361 );
or ( n90363 , n90360 , n90362 );
buf ( n90364 , n43400 );
not ( n90365 , n90364 );
buf ( n90366 , n37589 );
not ( n90367 , n90366 );
or ( n90368 , n90365 , n90367 );
buf ( n90369 , n39489 );
buf ( n90370 , n44635 );
nand ( n90371 , n90369 , n90370 );
buf ( n90372 , n90371 );
buf ( n90373 , n90372 );
nand ( n90374 , n90368 , n90373 );
buf ( n90375 , n90374 );
buf ( n90376 , n90375 );
buf ( n90377 , n38060 );
nand ( n90378 , n90376 , n90377 );
buf ( n90379 , n90378 );
buf ( n90380 , n90379 );
nand ( n90381 , n90363 , n90380 );
buf ( n90382 , n90381 );
buf ( n90383 , n90382 );
buf ( n90384 , n36104 );
not ( n90385 , n90384 );
buf ( n90386 , n90385 );
buf ( n90387 , n90386 );
buf ( n90388 , n89967 );
or ( n90389 , n90387 , n90388 );
buf ( n90390 , n32966 );
buf ( n90391 , n90390 );
buf ( n90392 , n39688 );
not ( n90393 , n90392 );
buf ( n90394 , n33077 );
not ( n90395 , n90394 );
and ( n90396 , n90393 , n90395 );
buf ( n90397 , n43503 );
buf ( n90398 , n39688 );
and ( n90399 , n90397 , n90398 );
nor ( n90400 , n90396 , n90399 );
buf ( n90401 , n90400 );
buf ( n90402 , n90401 );
or ( n90403 , n90391 , n90402 );
nand ( n90404 , n90389 , n90403 );
buf ( n90405 , n90404 );
buf ( n90406 , n90405 );
and ( n90407 , n90383 , n90406 );
not ( n90408 , n90383 );
buf ( n90409 , n90405 );
not ( n90410 , n90409 );
buf ( n90411 , n90410 );
buf ( n90412 , n90411 );
and ( n90413 , n90408 , n90412 );
nor ( n90414 , n90407 , n90413 );
buf ( n90415 , n90414 );
xor ( n90416 , n90358 , n90415 );
xor ( n90417 , n90339 , n90416 );
xor ( n90418 , n90313 , n90417 );
buf ( n90419 , n37922 );
not ( n90420 , n90419 );
buf ( n90421 , n90016 );
not ( n90422 , n90421 );
or ( n90423 , n90420 , n90422 );
buf ( n90424 , n89391 );
buf ( n90425 , n37875 );
nand ( n90426 , n90424 , n90425 );
buf ( n90427 , n90426 );
buf ( n90428 , n90427 );
nand ( n90429 , n90423 , n90428 );
buf ( n90430 , n90429 );
not ( n90431 , n90430 );
not ( n90432 , n37452 );
not ( n90433 , n90293 );
or ( n90434 , n90432 , n90433 );
nand ( n90435 , n89703 , n37517 );
nand ( n90436 , n90434 , n90435 );
not ( n90437 , n90436 );
not ( n90438 , n90437 );
or ( n90439 , n90431 , n90438 );
not ( n90440 , n90430 );
nand ( n90441 , n90440 , n90436 );
nand ( n90442 , n90439 , n90441 );
not ( n90443 , n38382 );
not ( n90444 , n90054 );
or ( n90445 , n90443 , n90444 );
buf ( n90446 , n89330 );
buf ( n90447 , n38775 );
nand ( n90448 , n90446 , n90447 );
buf ( n90449 , n90448 );
nand ( n90450 , n90445 , n90449 );
and ( n90451 , n90442 , n90450 );
not ( n90452 , n90442 );
not ( n90453 , n90450 );
and ( n90454 , n90452 , n90453 );
nor ( n90455 , n90451 , n90454 );
not ( n90456 , n90455 );
buf ( n90457 , n39986 );
not ( n90458 , n90457 );
buf ( n90459 , n24092 );
not ( n90460 , n90459 );
buf ( n90461 , n39897 );
not ( n90462 , n90461 );
or ( n90463 , n90460 , n90462 );
buf ( n90464 , n55813 );
buf ( n90465 , n40009 );
nand ( n90466 , n90464 , n90465 );
buf ( n90467 , n90466 );
buf ( n90468 , n90467 );
nand ( n90469 , n90463 , n90468 );
buf ( n90470 , n90469 );
buf ( n90471 , n90470 );
not ( n90472 , n90471 );
or ( n90473 , n90458 , n90472 );
buf ( n90474 , n89010 );
buf ( n90475 , n40002 );
nand ( n90476 , n90474 , n90475 );
buf ( n90477 , n90476 );
buf ( n90478 , n90477 );
nand ( n90479 , n90473 , n90478 );
buf ( n90480 , n90479 );
buf ( n90481 , n90480 );
buf ( n90482 , n42631 );
not ( n90483 , n90482 );
buf ( n90484 , n89676 );
not ( n90485 , n90484 );
or ( n90486 , n90483 , n90485 );
buf ( n90487 , n25160 );
not ( n90488 , n90487 );
buf ( n90489 , n42277 );
not ( n90490 , n90489 );
or ( n90491 , n90488 , n90490 );
buf ( n90492 , n42280 );
buf ( n90493 , n42581 );
nand ( n90494 , n90492 , n90493 );
buf ( n90495 , n90494 );
buf ( n90496 , n90495 );
nand ( n90497 , n90491 , n90496 );
buf ( n90498 , n90497 );
buf ( n90499 , n90498 );
buf ( n90500 , n42566 );
nand ( n90501 , n90499 , n90500 );
buf ( n90502 , n90501 );
buf ( n90503 , n90502 );
nand ( n90504 , n90486 , n90503 );
buf ( n90505 , n90504 );
buf ( n90506 , n90505 );
or ( n90507 , n90481 , n90506 );
buf ( n90508 , n90507 );
not ( n90509 , n90508 );
or ( n90510 , n90456 , n90509 );
buf ( n90511 , n90505 );
buf ( n90512 , n90480 );
and ( n90513 , n90511 , n90512 );
buf ( n90514 , n90513 );
not ( n90515 , n90514 );
nand ( n90516 , n90510 , n90515 );
xor ( n90517 , n90418 , n90516 );
buf ( n90518 , n90517 );
xor ( n90519 , n90190 , n90518 );
buf ( n90520 , n90519 );
buf ( n90521 , n90520 );
not ( n90522 , n89463 );
not ( n90523 , n89460 );
or ( n90524 , n90522 , n90523 );
not ( n90525 , n89459 );
not ( n90526 , n89149 );
or ( n90527 , n90525 , n90526 );
nand ( n90528 , n90527 , n88958 );
nand ( n90529 , n90524 , n90528 );
buf ( n90530 , n90529 );
not ( n90531 , n90530 );
xor ( n90532 , n89662 , n89752 );
and ( n90533 , n90532 , n89758 );
and ( n90534 , n89662 , n89752 );
or ( n90535 , n90533 , n90534 );
buf ( n90536 , n90535 );
not ( n90537 , n90536 );
buf ( n90538 , n90537 );
xor ( n90539 , n90511 , n90512 );
buf ( n90540 , n90539 );
not ( n90541 , n90455 );
and ( n90542 , n90540 , n90541 );
not ( n90543 , n90540 );
and ( n90544 , n90543 , n90455 );
nor ( n90545 , n90542 , n90544 );
xor ( n90546 , n89686 , n89745 );
and ( n90547 , n90546 , n89751 );
and ( n90548 , n89686 , n89745 );
or ( n90549 , n90547 , n90548 );
and ( n90550 , n90545 , n90549 );
not ( n90551 , n90545 );
not ( n90552 , n90549 );
and ( n90553 , n90551 , n90552 );
or ( n90554 , n90550 , n90553 );
not ( n90555 , n89458 );
nand ( n90556 , n89270 , n89304 );
not ( n90557 , n90556 );
or ( n90558 , n90555 , n90557 );
not ( n90559 , n89270 );
nand ( n90560 , n90559 , n89301 );
nand ( n90561 , n90558 , n90560 );
not ( n90562 , n90561 );
and ( n90563 , n90554 , n90562 );
not ( n90564 , n90554 );
and ( n90565 , n90564 , n90561 );
nor ( n90566 , n90563 , n90565 );
nand ( n90567 , n90538 , n90566 );
buf ( n90568 , n90567 );
not ( n90569 , n90568 );
or ( n90570 , n90531 , n90569 );
not ( n90571 , n90566 );
buf ( n90572 , n90571 );
buf ( n90573 , n90535 );
nand ( n90574 , n90572 , n90573 );
buf ( n90575 , n90574 );
buf ( n90576 , n90575 );
nand ( n90577 , n90570 , n90576 );
buf ( n90578 , n90577 );
buf ( n90579 , n90578 );
xor ( n90580 , n90521 , n90579 );
buf ( n90581 , n90175 );
buf ( n90582 , n90126 );
or ( n90583 , n90581 , n90582 );
buf ( n90584 , n90169 );
not ( n90585 , n90584 );
buf ( n90586 , n90585 );
buf ( n90587 , n90586 );
nand ( n90588 , n90583 , n90587 );
buf ( n90589 , n90588 );
buf ( n90590 , n90589 );
buf ( n90591 , n90175 );
buf ( n90592 , n90126 );
nand ( n90593 , n90591 , n90592 );
buf ( n90594 , n90593 );
buf ( n90595 , n90594 );
and ( n90596 , n90590 , n90595 );
buf ( n90597 , n90596 );
buf ( n90598 , n90597 );
not ( n90599 , n90450 );
nand ( n90600 , n90437 , n90440 );
not ( n90601 , n90600 );
or ( n90602 , n90599 , n90601 );
nand ( n90603 , n90430 , n90436 );
nand ( n90604 , n90602 , n90603 );
not ( n90605 , n40002 );
not ( n90606 , n90470 );
or ( n90607 , n90605 , n90606 );
buf ( n90608 , n40010 );
not ( n90609 , n90608 );
buf ( n90610 , n40067 );
not ( n90611 , n90610 );
or ( n90612 , n90609 , n90611 );
buf ( n90613 , n36427 );
buf ( n90614 , n40009 );
nand ( n90615 , n90613 , n90614 );
buf ( n90616 , n90615 );
buf ( n90617 , n90616 );
nand ( n90618 , n90612 , n90617 );
buf ( n90619 , n90618 );
buf ( n90620 , n90619 );
buf ( n90621 , n39986 );
nand ( n90622 , n90620 , n90621 );
buf ( n90623 , n90622 );
nand ( n90624 , n90607 , n90623 );
not ( n90625 , n90624 );
not ( n90626 , n42631 );
not ( n90627 , n90498 );
or ( n90628 , n90626 , n90627 );
buf ( n90629 , n25160 );
not ( n90630 , n90629 );
buf ( n90631 , n39582 );
not ( n90632 , n90631 );
or ( n90633 , n90630 , n90632 );
buf ( n90634 , n36611 );
buf ( n90635 , n42581 );
nand ( n90636 , n90634 , n90635 );
buf ( n90637 , n90636 );
buf ( n90638 , n90637 );
nand ( n90639 , n90633 , n90638 );
buf ( n90640 , n90639 );
buf ( n90641 , n90640 );
buf ( n90642 , n42566 );
nand ( n90643 , n90641 , n90642 );
buf ( n90644 , n90643 );
nand ( n90645 , n90628 , n90644 );
and ( n90646 , n90604 , n90625 , n90645 );
not ( n90647 , n90646 );
not ( n90648 , n90645 );
and ( n90649 , n90604 , n90624 , n90648 );
not ( n90650 , n90604 );
nor ( n90651 , n90624 , n90645 );
and ( n90652 , n90650 , n90651 );
nor ( n90653 , n90649 , n90652 );
nand ( n90654 , n90624 , n90645 , n90650 );
nand ( n90655 , n90647 , n90653 , n90654 );
buf ( n90656 , n90655 );
xor ( n90657 , n90598 , n90656 );
not ( n90658 , n89450 );
not ( n90659 , n89337 );
or ( n90660 , n90658 , n90659 );
not ( n90661 , n89338 );
not ( n90662 , n89449 );
or ( n90663 , n90661 , n90662 );
nand ( n90664 , n90663 , n89311 );
nand ( n90665 , n90660 , n90664 );
not ( n90666 , n90665 );
not ( n90667 , n90666 );
not ( n90668 , n89190 );
not ( n90669 , n89228 );
or ( n90670 , n90668 , n90669 );
not ( n90671 , n89191 );
not ( n90672 , n89231 );
or ( n90673 , n90671 , n90672 );
nand ( n90674 , n90673 , n89265 );
nand ( n90675 , n90670 , n90674 );
buf ( n90676 , n90675 );
not ( n90677 , n90676 );
buf ( n90678 , n90677 );
not ( n90679 , n90678 );
and ( n90680 , n90667 , n90679 );
not ( n90681 , n89999 );
and ( n90682 , n89908 , n89933 );
not ( n90683 , n89908 );
and ( n90684 , n90683 , n89938 );
nor ( n90685 , n90682 , n90684 );
not ( n90686 , n90685 );
not ( n90687 , n90686 );
or ( n90688 , n90681 , n90687 );
not ( n90689 , n89999 );
nand ( n90690 , n90689 , n90685 );
nand ( n90691 , n90688 , n90690 );
or ( n90692 , n90665 , n90675 );
and ( n90693 , n90691 , n90692 );
nor ( n90694 , n90680 , n90693 );
buf ( n90695 , n90694 );
xor ( n90696 , n90657 , n90695 );
buf ( n90697 , n90696 );
buf ( n90698 , n90697 );
not ( n90699 , n90552 );
not ( n90700 , n90545 );
and ( n90701 , n90699 , n90700 );
nand ( n90702 , n90552 , n90545 );
and ( n90703 , n90561 , n90702 );
nor ( n90704 , n90701 , n90703 );
buf ( n90705 , n90704 );
and ( n90706 , n90698 , n90705 );
not ( n90707 , n90698 );
buf ( n90708 , n90704 );
not ( n90709 , n90708 );
buf ( n90710 , n90709 );
buf ( n90711 , n90710 );
and ( n90712 , n90707 , n90711 );
nor ( n90713 , n90706 , n90712 );
buf ( n90714 , n90713 );
buf ( n90715 , n90714 );
buf ( n90716 , n90675 );
not ( n90717 , n90716 );
buf ( n90718 , n90666 );
not ( n90719 , n90718 );
or ( n90720 , n90717 , n90719 );
buf ( n90721 , n90665 );
buf ( n90722 , n90678 );
nand ( n90723 , n90721 , n90722 );
buf ( n90724 , n90723 );
buf ( n90725 , n90724 );
nand ( n90726 , n90720 , n90725 );
buf ( n90727 , n90726 );
not ( n90728 , n90691 );
and ( n90729 , n90727 , n90728 );
not ( n90730 , n90727 );
and ( n90731 , n90730 , n90691 );
nor ( n90732 , n90729 , n90731 );
buf ( n90733 , n90732 );
not ( n90734 , n90733 );
xor ( n90735 , n90099 , n90092 );
xor ( n90736 , n90735 , n90176 );
buf ( n90737 , n90736 );
not ( n90738 , n90737 );
or ( n90739 , n90734 , n90738 );
not ( n90740 , n89003 );
buf ( n90741 , n89142 );
not ( n90742 , n90741 );
or ( n90743 , n90740 , n90742 );
or ( n90744 , n90741 , n89003 );
nand ( n90745 , n90744 , n89148 );
nand ( n90746 , n90743 , n90745 );
buf ( n90747 , n90746 );
nand ( n90748 , n90739 , n90747 );
buf ( n90749 , n90748 );
buf ( n90750 , n90749 );
buf ( n90751 , n90732 );
not ( n90752 , n90751 );
buf ( n90753 , n90736 );
not ( n90754 , n90753 );
buf ( n90755 , n90754 );
buf ( n90756 , n90755 );
nand ( n90757 , n90752 , n90756 );
buf ( n90758 , n90757 );
buf ( n90759 , n90758 );
nand ( n90760 , n90750 , n90759 );
buf ( n90761 , n90760 );
buf ( n90762 , n90761 );
xor ( n90763 , n90715 , n90762 );
buf ( n90764 , n90763 );
buf ( n90765 , n90764 );
xor ( n90766 , n90580 , n90765 );
buf ( n90767 , n90766 );
not ( n90768 , n90767 );
not ( n90769 , n90746 );
and ( n90770 , n90732 , n90769 );
not ( n90771 , n90732 );
and ( n90772 , n90771 , n90746 );
nor ( n90773 , n90770 , n90772 );
and ( n90774 , n90773 , n90736 );
not ( n90775 , n90773 );
and ( n90776 , n90775 , n90755 );
nor ( n90777 , n90774 , n90776 );
not ( n90778 , n90535 );
not ( n90779 , n90566 );
or ( n90780 , n90778 , n90779 );
buf ( n90781 , n90571 );
buf ( n90782 , n90538 );
nand ( n90783 , n90781 , n90782 );
buf ( n90784 , n90783 );
nand ( n90785 , n90780 , n90784 );
not ( n90786 , n90529 );
and ( n90787 , n90785 , n90786 );
not ( n90788 , n90785 );
and ( n90789 , n90788 , n90529 );
nor ( n90790 , n90787 , n90789 );
xor ( n90791 , n90777 , n90790 );
buf ( n90792 , n89567 );
buf ( n90793 , n89653 );
not ( n90794 , n90793 );
buf ( n90795 , n89762 );
nand ( n90796 , n90794 , n90795 );
buf ( n90797 , n90796 );
buf ( n90798 , n90797 );
and ( n90799 , n90792 , n90798 );
buf ( n90800 , n89653 );
not ( n90801 , n90800 );
buf ( n90802 , n89762 );
nor ( n90803 , n90801 , n90802 );
buf ( n90804 , n90803 );
buf ( n90805 , n90804 );
nor ( n90806 , n90799 , n90805 );
buf ( n90807 , n90806 );
and ( n90808 , n90791 , n90807 );
and ( n90809 , n90777 , n90790 );
or ( n90810 , n90808 , n90809 );
nand ( n90811 , n90768 , n90810 );
not ( n90812 , n90811 );
not ( n90813 , n89811 );
buf ( n90814 , n89469 );
not ( n90815 , n90814 );
buf ( n90816 , n90815 );
not ( n90817 , n90816 );
and ( n90818 , n90813 , n90817 );
buf ( n90819 , n89811 );
buf ( n90820 , n90816 );
nand ( n90821 , n90819 , n90820 );
buf ( n90822 , n90821 );
buf ( n90823 , n89779 );
not ( n90824 , n90823 );
buf ( n90825 , n90824 );
and ( n90826 , n90822 , n90825 );
nor ( n90827 , n90818 , n90826 );
xor ( n90828 , n90777 , n90790 );
xor ( n90829 , n90828 , n90807 );
nand ( n90830 , n90827 , n90829 );
not ( n90831 , n90830 );
nor ( n90832 , n89856 , n90812 , n90831 );
xor ( n90833 , n90521 , n90579 );
and ( n90834 , n90833 , n90765 );
and ( n90835 , n90521 , n90579 );
or ( n90836 , n90834 , n90835 );
buf ( n90837 , n90836 );
not ( n90838 , n90837 );
xor ( n90839 , n90040 , n90067 );
and ( n90840 , n90839 , n90074 );
and ( n90841 , n90040 , n90067 );
or ( n90842 , n90840 , n90841 );
buf ( n90843 , n90842 );
buf ( n90844 , n90843 );
not ( n90845 , n90844 );
buf ( n90846 , n90845 );
buf ( n90847 , n90846 );
not ( n90848 , n90847 );
buf ( n90849 , n38063 );
not ( n90850 , n90849 );
buf ( n90851 , n43371 );
buf ( n90852 , n43678 );
and ( n90853 , n90851 , n90852 );
not ( n90854 , n90851 );
buf ( n90855 , n51833 );
and ( n90856 , n90854 , n90855 );
nor ( n90857 , n90853 , n90856 );
buf ( n90858 , n90857 );
buf ( n90859 , n90858 );
not ( n90860 , n90859 );
or ( n90861 , n90850 , n90860 );
buf ( n90862 , n38133 );
buf ( n90863 , n90375 );
nand ( n90864 , n90862 , n90863 );
buf ( n90865 , n90864 );
buf ( n90866 , n90865 );
nand ( n90867 , n90861 , n90866 );
buf ( n90868 , n90867 );
not ( n90869 , n37403 );
not ( n90870 , n90207 );
or ( n90871 , n90869 , n90870 );
buf ( n90872 , n37330 );
not ( n90873 , n90872 );
buf ( n90874 , n39407 );
not ( n90875 , n90874 );
or ( n90876 , n90873 , n90875 );
buf ( n90877 , n52072 );
buf ( n90878 , n37329 );
nand ( n90879 , n90877 , n90878 );
buf ( n90880 , n90879 );
buf ( n90881 , n90880 );
nand ( n90882 , n90876 , n90881 );
buf ( n90883 , n90882 );
nand ( n90884 , n90883 , n38150 );
nand ( n90885 , n90871 , n90884 );
xor ( n90886 , n90868 , n90885 );
buf ( n90887 , n90405 );
not ( n90888 , n90887 );
buf ( n90889 , n90382 );
not ( n90890 , n90889 );
or ( n90891 , n90888 , n90890 );
buf ( n90892 , n90411 );
not ( n90893 , n90892 );
buf ( n90894 , n90382 );
not ( n90895 , n90894 );
buf ( n90896 , n90895 );
buf ( n90897 , n90896 );
not ( n90898 , n90897 );
or ( n90899 , n90893 , n90898 );
buf ( n90900 , n90358 );
nand ( n90901 , n90899 , n90900 );
buf ( n90902 , n90901 );
buf ( n90903 , n90902 );
nand ( n90904 , n90891 , n90903 );
buf ( n90905 , n90904 );
xnor ( n90906 , n90886 , n90905 );
buf ( n90907 , n90906 );
not ( n90908 , n90907 );
buf ( n90909 , n90908 );
buf ( n90910 , n90909 );
not ( n90911 , n90910 );
or ( n90912 , n90848 , n90911 );
buf ( n90913 , n90906 );
buf ( n90914 , n90843 );
nand ( n90915 , n90913 , n90914 );
buf ( n90916 , n90915 );
buf ( n90917 , n90916 );
nand ( n90918 , n90912 , n90917 );
buf ( n90919 , n90918 );
xor ( n90920 , n90329 , n90338 );
and ( n90921 , n90920 , n90416 );
and ( n90922 , n90329 , n90338 );
or ( n90923 , n90921 , n90922 );
and ( n90924 , n90919 , n90923 );
not ( n90925 , n90919 );
not ( n90926 , n90923 );
and ( n90927 , n90925 , n90926 );
nor ( n90928 , n90924 , n90927 );
buf ( n90929 , n90928 );
buf ( n90930 , n42566 );
not ( n90931 , n90930 );
buf ( n90932 , n25160 );
not ( n90933 , n90932 );
buf ( n90934 , n43857 );
not ( n90935 , n90934 );
or ( n90936 , n90933 , n90935 );
buf ( n90937 , n36038 );
buf ( n90938 , n42581 );
nand ( n90939 , n90937 , n90938 );
buf ( n90940 , n90939 );
buf ( n90941 , n90940 );
nand ( n90942 , n90936 , n90941 );
buf ( n90943 , n90942 );
buf ( n90944 , n90943 );
not ( n90945 , n90944 );
or ( n90946 , n90931 , n90945 );
buf ( n90947 , n90640 );
buf ( n90948 , n42631 );
nand ( n90949 , n90947 , n90948 );
buf ( n90950 , n90949 );
buf ( n90951 , n90950 );
nand ( n90952 , n90946 , n90951 );
buf ( n90953 , n90952 );
buf ( n90954 , n90953 );
buf ( n90955 , n37452 );
not ( n90956 , n90955 );
buf ( n90957 , n88143 );
not ( n90958 , n90957 );
buf ( n90959 , n37268 );
not ( n90960 , n90959 );
or ( n90961 , n90958 , n90960 );
buf ( n90962 , n43142 );
buf ( n90963 , n37475 );
nand ( n90964 , n90962 , n90963 );
buf ( n90965 , n90964 );
buf ( n90966 , n90965 );
nand ( n90967 , n90961 , n90966 );
buf ( n90968 , n90967 );
buf ( n90969 , n90968 );
not ( n90970 , n90969 );
or ( n90971 , n90956 , n90970 );
buf ( n90972 , n90307 );
buf ( n90973 , n37517 );
nand ( n90974 , n90972 , n90973 );
buf ( n90975 , n90974 );
buf ( n90976 , n90975 );
nand ( n90977 , n90971 , n90976 );
buf ( n90978 , n90977 );
buf ( n90979 , n90978 );
xor ( n90980 , n90954 , n90979 );
buf ( n90981 , n43053 );
buf ( n90982 , n43806 );
not ( n90983 , n90982 );
buf ( n90984 , n37649 );
not ( n90985 , n90984 );
or ( n90986 , n90983 , n90985 );
buf ( n90987 , n38798 );
buf ( n90988 , n75045 );
nand ( n90989 , n90987 , n90988 );
buf ( n90990 , n90989 );
buf ( n90991 , n90990 );
nand ( n90992 , n90986 , n90991 );
buf ( n90993 , n90992 );
buf ( n90994 , n90993 );
nand ( n90995 , n90981 , n90994 );
buf ( n90996 , n90995 );
buf ( n90997 , n90996 );
nand ( n90998 , C1 , n90997 );
buf ( n90999 , n90998 );
buf ( n91000 , n90999 );
not ( n91001 , n42530 );
buf ( n91002 , n33077 );
not ( n91003 , n91002 );
buf ( n91004 , n38851 );
not ( n91005 , n91004 );
or ( n91006 , n91003 , n91005 );
buf ( n91007 , n38865 );
buf ( n91008 , n39478 );
nand ( n91009 , n91007 , n91008 );
buf ( n91010 , n91009 );
buf ( n91011 , n91010 );
nand ( n91012 , n91006 , n91011 );
buf ( n91013 , n91012 );
not ( n91014 , n91013 );
or ( n91015 , n91001 , n91014 );
not ( n91016 , n90401 );
nand ( n91017 , n91016 , n36104 );
nand ( n91018 , n91015 , n91017 );
buf ( n91019 , n91018 );
xor ( n91020 , n91000 , n91019 );
buf ( n91021 , n45426 );
buf ( n91022 , n90354 );
or ( n91023 , n91021 , n91022 );
and ( n91024 , n39209 , n88457 );
not ( n91025 , n39209 );
and ( n91026 , n91025 , n42082 );
nor ( n91027 , n91024 , n91026 );
buf ( n91028 , n91027 );
buf ( n91029 , n44682 );
or ( n91030 , n91028 , n91029 );
nand ( n91031 , n91023 , n91030 );
buf ( n91032 , n91031 );
buf ( n91033 , n91032 );
xor ( n91034 , n91020 , n91033 );
buf ( n91035 , n91034 );
buf ( n91036 , n91035 );
xor ( n91037 , n90980 , n91036 );
buf ( n91038 , n91037 );
buf ( n91039 , n91038 );
not ( n91040 , n90312 );
not ( n91041 , n90214 );
nand ( n91042 , n91041 , n90239 );
not ( n91043 , n91042 );
or ( n91044 , n91040 , n91043 );
nand ( n91045 , n90238 , n90214 );
nand ( n91046 , n91044 , n91045 );
buf ( n91047 , n91046 );
and ( n91048 , n91039 , n91047 );
not ( n91049 , n91039 );
buf ( n91050 , n91046 );
not ( n91051 , n91050 );
buf ( n91052 , n91051 );
buf ( n91053 , n91052 );
and ( n91054 , n91049 , n91053 );
nor ( n91055 , n91048 , n91054 );
buf ( n91056 , n91055 );
buf ( n91057 , n91056 );
buf ( n91058 , n43906 );
not ( n91059 , n91058 );
buf ( n91060 , n43941 );
not ( n91061 , n91060 );
or ( n91062 , n91059 , n91061 );
buf ( n91063 , n90322 );
nand ( n91064 , n91062 , n91063 );
buf ( n91065 , n91064 );
xor ( n91066 , n90257 , n90283 );
and ( n91067 , n91066 , n90310 );
and ( n91068 , n90257 , n90283 );
or ( n91069 , n91067 , n91068 );
buf ( n91070 , n91069 );
xor ( n91071 , n91065 , n91070 );
buf ( n91072 , n90276 );
not ( n91073 , n91072 );
buf ( n91074 , n50374 );
not ( n91075 , n91074 );
or ( n91076 , n91073 , n91075 );
buf ( n91077 , n39816 );
and ( n91078 , n43777 , n39729 );
not ( n91079 , n43777 );
and ( n91080 , n91079 , n52246 );
or ( n91081 , n91078 , n91080 );
buf ( n91082 , n91081 );
nand ( n91083 , n91077 , n91082 );
buf ( n91084 , n91083 );
buf ( n91085 , n91084 );
nand ( n91086 , n91076 , n91085 );
buf ( n91087 , n91086 );
xor ( n91088 , n91087 , n90256 );
buf ( n91089 , n37892 );
buf ( n91090 , n37717 );
and ( n91091 , n91089 , n91090 );
not ( n91092 , n91089 );
buf ( n91093 , n39246 );
and ( n91094 , n91092 , n91093 );
nor ( n91095 , n91091 , n91094 );
buf ( n91096 , n91095 );
buf ( n91097 , n91096 );
buf ( n91098 , n40276 );
or ( n91099 , n91097 , n91098 );
buf ( n91100 , n90032 );
buf ( n91101 , n37875 );
nand ( n91102 , n91100 , n91101 );
buf ( n91103 , n91102 );
buf ( n91104 , n91103 );
nand ( n91105 , n91099 , n91104 );
buf ( n91106 , n91105 );
xnor ( n91107 , n91088 , n91106 );
xor ( n91108 , n91071 , n91107 );
buf ( n91109 , n91108 );
not ( n91110 , n91109 );
buf ( n91111 , n91110 );
buf ( n91112 , n91111 );
and ( n91113 , n91057 , n91112 );
not ( n91114 , n91057 );
buf ( n91115 , n91108 );
and ( n91116 , n91114 , n91115 );
nor ( n91117 , n91113 , n91116 );
buf ( n91118 , n91117 );
buf ( n91119 , n91118 );
xor ( n91120 , n90929 , n91119 );
not ( n91121 , n90313 );
not ( n91122 , n90417 );
nor ( n91123 , n91121 , n91122 );
or ( n91124 , n91123 , n90516 );
not ( n91125 , n90417 );
nand ( n91126 , n91125 , n91121 );
nand ( n91127 , n91124 , n91126 );
buf ( n91128 , n91127 );
xnor ( n91129 , n91120 , n91128 );
buf ( n91130 , n91129 );
buf ( n91131 , n91130 );
buf ( n91132 , n90704 );
not ( n91133 , n91132 );
buf ( n91134 , n90697 );
not ( n91135 , n91134 );
or ( n91136 , n91133 , n91135 );
buf ( n91137 , n90761 );
nand ( n91138 , n91136 , n91137 );
buf ( n91139 , n91138 );
buf ( n91140 , n91139 );
buf ( n91141 , n90697 );
not ( n91142 , n91141 );
buf ( n91143 , n90710 );
nand ( n91144 , n91142 , n91143 );
buf ( n91145 , n91144 );
buf ( n91146 , n91145 );
and ( n91147 , n91140 , n91146 );
buf ( n91148 , n91147 );
buf ( n91149 , n91148 );
xor ( n91150 , n91131 , n91149 );
buf ( n91151 , n38382 );
not ( n91152 , n91151 );
buf ( n91153 , n38413 );
not ( n91154 , n91153 );
buf ( n91155 , n42360 );
not ( n91156 , n91155 );
or ( n91157 , n91154 , n91156 );
nand ( n91158 , n38436 , n38420 );
buf ( n91159 , n91158 );
nand ( n91160 , n91157 , n91159 );
buf ( n91161 , n91160 );
buf ( n91162 , n91161 );
not ( n91163 , n91162 );
or ( n91164 , n91152 , n91163 );
buf ( n91165 , n90062 );
buf ( n91166 , n38775 );
nand ( n91167 , n91165 , n91166 );
buf ( n91168 , n91167 );
buf ( n91169 , n91168 );
nand ( n91170 , n91164 , n91169 );
buf ( n91171 , n91170 );
buf ( n91172 , n91171 );
buf ( n91173 , n39374 );
not ( n91174 , n91173 );
buf ( n91175 , n39000 );
not ( n91176 , n91175 );
buf ( n91177 , n39891 );
not ( n91178 , n91177 );
or ( n91179 , n91176 , n91178 );
buf ( n91180 , n36396 );
buf ( n91181 , n38997 );
nand ( n91182 , n91180 , n91181 );
buf ( n91183 , n91182 );
buf ( n91184 , n91183 );
nand ( n91185 , n91179 , n91184 );
buf ( n91186 , n91185 );
buf ( n91187 , n91186 );
not ( n91188 , n91187 );
or ( n91189 , n91174 , n91188 );
buf ( n91190 , n90231 );
buf ( n91191 , n39395 );
nand ( n91192 , n91190 , n91191 );
buf ( n91193 , n91192 );
buf ( n91194 , n91193 );
nand ( n91195 , n91189 , n91194 );
buf ( n91196 , n91195 );
buf ( n91197 , n91196 );
xor ( n91198 , n91172 , n91197 );
buf ( n91199 , n90619 );
buf ( n91200 , n40002 );
and ( n91201 , n91199 , n91200 );
buf ( n91202 , n24092 );
not ( n91203 , n91202 );
buf ( n91204 , n39927 );
not ( n91205 , n91204 );
or ( n91206 , n91203 , n91205 );
buf ( n91207 , n39924 );
buf ( n91208 , n40009 );
nand ( n91209 , n91207 , n91208 );
buf ( n91210 , n91209 );
buf ( n91211 , n91210 );
nand ( n91212 , n91206 , n91211 );
buf ( n91213 , n91212 );
buf ( n91214 , n91213 );
not ( n91215 , n91214 );
buf ( n91216 , n39989 );
nor ( n91217 , n91215 , n91216 );
buf ( n91218 , n91217 );
buf ( n91219 , n91218 );
nor ( n91220 , n91201 , n91219 );
buf ( n91221 , n91220 );
buf ( n91222 , n91221 );
not ( n91223 , n91222 );
buf ( n91224 , n91223 );
buf ( n91225 , n91224 );
xnor ( n91226 , n91198 , n91225 );
buf ( n91227 , n91226 );
buf ( n91228 , n91227 );
not ( n91229 , n91228 );
buf ( n91230 , n91229 );
buf ( n91231 , n91230 );
not ( n91232 , n91231 );
or ( n91233 , n90650 , n90651 );
nand ( n91234 , n90624 , n90645 );
nand ( n91235 , n91233 , n91234 );
buf ( n91236 , n91235 );
not ( n91237 , n91236 );
buf ( n91238 , n91237 );
buf ( n91239 , n91238 );
not ( n91240 , n91239 );
or ( n91241 , n91232 , n91240 );
buf ( n91242 , n91227 );
buf ( n91243 , n91235 );
nand ( n91244 , n91242 , n91243 );
buf ( n91245 , n91244 );
buf ( n91246 , n91245 );
nand ( n91247 , n91241 , n91246 );
buf ( n91248 , n91247 );
buf ( n91249 , n91248 );
xor ( n91250 , n89892 , n90001 );
and ( n91251 , n91250 , n90076 );
and ( n91252 , n89892 , n90001 );
or ( n91253 , n91251 , n91252 );
buf ( n91254 , n91253 );
and ( n91255 , n91249 , n91254 );
not ( n91256 , n91249 );
buf ( n91257 , n91253 );
not ( n91258 , n91257 );
buf ( n91259 , n91258 );
buf ( n91260 , n91259 );
and ( n91261 , n91256 , n91260 );
nor ( n91262 , n91255 , n91261 );
buf ( n91263 , n91262 );
xor ( n91264 , n90598 , n90656 );
and ( n91265 , n91264 , n90695 );
and ( n91266 , n90598 , n90656 );
or ( n91267 , n91265 , n91266 );
buf ( n91268 , n91267 );
xor ( n91269 , n91263 , n91268 );
xor ( n91270 , n90078 , n90189 );
and ( n91271 , n91270 , n90518 );
and ( n91272 , n90078 , n90189 );
or ( n91273 , n91271 , n91272 );
buf ( n91274 , n91273 );
xor ( n91275 , n91269 , n91274 );
buf ( n91276 , n91275 );
xor ( n91277 , n91150 , n91276 );
buf ( n91278 , n91277 );
nand ( n91279 , n90838 , n91278 );
buf ( n91280 , n39000 );
buf ( n91281 , n40067 );
and ( n91282 , n91280 , n91281 );
not ( n91283 , n91280 );
buf ( n91284 , n36427 );
and ( n91285 , n91283 , n91284 );
nor ( n91286 , n91282 , n91285 );
buf ( n91287 , n91286 );
buf ( n91288 , n91287 );
not ( n91289 , n91288 );
buf ( n91290 , n38974 );
not ( n91291 , n91290 );
and ( n91292 , n91289 , n91291 );
buf ( n91293 , n91186 );
buf ( n91294 , n39395 );
and ( n91295 , n91293 , n91294 );
nor ( n91296 , n91292 , n91295 );
buf ( n91297 , n91296 );
not ( n91298 , n90868 );
not ( n91299 , n91298 );
not ( n91300 , n90885 );
not ( n91301 , n91300 );
or ( n91302 , n91299 , n91301 );
nand ( n91303 , n91302 , n90905 );
nand ( n91304 , n90868 , n90885 );
nand ( n91305 , n91303 , n91304 );
xor ( n91306 , n91297 , n91305 );
xor ( n91307 , n90954 , n90979 );
and ( n91308 , n91307 , n91036 );
and ( n91309 , n90954 , n90979 );
or ( n91310 , n91308 , n91309 );
buf ( n91311 , n91310 );
xnor ( n91312 , n91306 , n91311 );
buf ( n91313 , n91038 );
not ( n91314 , n91313 );
buf ( n91315 , n91046 );
not ( n91316 , n91315 );
or ( n91317 , n91314 , n91316 );
buf ( n91318 , n91046 );
buf ( n91319 , n91038 );
or ( n91320 , n91318 , n91319 );
buf ( n91321 , n91108 );
nand ( n91322 , n91320 , n91321 );
buf ( n91323 , n91322 );
buf ( n91324 , n91323 );
nand ( n91325 , n91317 , n91324 );
buf ( n91326 , n91325 );
xor ( n91327 , n91312 , n91326 );
xor ( n91328 , n91000 , n91019 );
and ( n91329 , n91328 , n91033 );
and ( n91330 , n91000 , n91019 );
or ( n91331 , n91329 , n91330 );
buf ( n91332 , n91331 );
buf ( n91333 , n91332 );
buf ( n91334 , n42631 );
not ( n91335 , n91334 );
buf ( n91336 , n90943 );
not ( n91337 , n91336 );
or ( n91338 , n91335 , n91337 );
buf ( n91339 , n25160 );
not ( n91340 , n91339 );
buf ( n91341 , n39008 );
not ( n91342 , n91341 );
or ( n91343 , n91340 , n91342 );
buf ( n91344 , n41619 );
not ( n91345 , n91344 );
buf ( n91346 , n42581 );
nand ( n91347 , n91345 , n91346 );
buf ( n91348 , n91347 );
buf ( n91349 , n91348 );
nand ( n91350 , n91343 , n91349 );
buf ( n91351 , n91350 );
buf ( n91352 , n91351 );
buf ( n91353 , n42566 );
nand ( n91354 , n91352 , n91353 );
buf ( n91355 , n91354 );
buf ( n91356 , n91355 );
nand ( n91357 , n91338 , n91356 );
buf ( n91358 , n91357 );
buf ( n91359 , n91358 );
xor ( n91360 , n91333 , n91359 );
buf ( n91361 , n37403 );
not ( n91362 , n91361 );
buf ( n91363 , n90883 );
not ( n91364 , n91363 );
or ( n91365 , n91362 , n91364 );
buf ( n91366 , n37330 );
not ( n91367 , n91366 );
buf ( n91368 , n37971 );
not ( n91369 , n91368 );
or ( n91370 , n91367 , n91369 );
buf ( n91371 , n39277 );
buf ( n91372 , n37329 );
nand ( n91373 , n91371 , n91372 );
buf ( n91374 , n91373 );
buf ( n91375 , n91374 );
nand ( n91376 , n91370 , n91375 );
buf ( n91377 , n91376 );
buf ( n91378 , n91377 );
buf ( n91379 , n38150 );
nand ( n91380 , n91378 , n91379 );
buf ( n91381 , n91380 );
buf ( n91382 , n91381 );
nand ( n91383 , n91365 , n91382 );
buf ( n91384 , n91383 );
buf ( n91385 , n91384 );
xor ( n91386 , n91360 , n91385 );
buf ( n91387 , n91386 );
buf ( n91388 , n91387 );
buf ( n91389 , n37517 );
not ( n91390 , n91389 );
buf ( n91391 , n90968 );
not ( n91392 , n91391 );
or ( n91393 , n91390 , n91392 );
buf ( n91394 , n88143 );
not ( n91395 , n91394 );
buf ( n91396 , n43031 );
not ( n91397 , n91396 );
or ( n91398 , n91395 , n91397 );
buf ( n91399 , n38247 );
buf ( n91400 , n37475 );
nand ( n91401 , n91399 , n91400 );
buf ( n91402 , n91401 );
buf ( n91403 , n91402 );
nand ( n91404 , n91398 , n91403 );
buf ( n91405 , n91404 );
buf ( n91406 , n91405 );
buf ( n91407 , n37452 );
nand ( n91408 , n91406 , n91407 );
buf ( n91409 , n91408 );
buf ( n91410 , n91409 );
nand ( n91411 , n91393 , n91410 );
buf ( n91412 , n91411 );
buf ( n91413 , n91412 );
buf ( n91414 , n40002 );
not ( n91415 , n91414 );
buf ( n91416 , n91213 );
not ( n91417 , n91416 );
or ( n91418 , n91415 , n91417 );
buf ( n91419 , n40010 );
not ( n91420 , n91419 );
buf ( n91421 , n39582 );
not ( n91422 , n91421 );
or ( n91423 , n91420 , n91422 );
buf ( n91424 , n36617 );
buf ( n91425 , n40009 );
nand ( n91426 , n91424 , n91425 );
buf ( n91427 , n91426 );
buf ( n91428 , n91427 );
nand ( n91429 , n91423 , n91428 );
buf ( n91430 , n91429 );
buf ( n91431 , n91430 );
buf ( n91432 , n39986 );
nand ( n91433 , n91431 , n91432 );
buf ( n91434 , n91433 );
buf ( n91435 , n91434 );
nand ( n91436 , n91418 , n91435 );
buf ( n91437 , n91436 );
buf ( n91438 , n91437 );
xor ( n91439 , n91413 , n91438 );
buf ( n91440 , n91013 );
not ( n91441 , n91440 );
buf ( n91442 , n36104 );
not ( n91443 , n91442 );
or ( n91444 , n91441 , n91443 );
buf ( n91445 , n39481 );
buf ( n91446 , n39742 );
and ( n91447 , n91445 , n91446 );
not ( n91448 , n91445 );
buf ( n91449 , n38830 );
and ( n91450 , n91448 , n91449 );
nor ( n91451 , n91447 , n91450 );
buf ( n91452 , n91451 );
buf ( n91453 , n91452 );
not ( n91454 , n91453 );
buf ( n91455 , n32972 );
nand ( n91456 , n91454 , n91455 );
buf ( n91457 , n91456 );
buf ( n91458 , n91457 );
nand ( n91459 , n91444 , n91458 );
buf ( n91460 , n91459 );
buf ( n91461 , n91460 );
not ( n91462 , n60583 );
not ( n91463 , n89425 );
or ( n91464 , n91462 , n91463 );
buf ( n91465 , n38471 );
buf ( n91466 , n39688 );
nand ( n91467 , n91465 , n91466 );
buf ( n91468 , n91467 );
nand ( n91469 , n91464 , n91468 );
not ( n91470 , n91469 );
not ( n91471 , n39816 );
or ( n91472 , n91470 , n91471 );
nand ( n91473 , n39806 , n91081 );
nand ( n91474 , n91472 , n91473 );
buf ( n91475 , n91474 );
xor ( n91476 , n91461 , n91475 );
buf ( n91477 , n36985 );
buf ( n91478 , n91027 );
or ( n91479 , n91477 , n91478 );
buf ( n91480 , n36932 );
buf ( n91481 , n37598 );
and ( n91482 , n91480 , n91481 );
not ( n91483 , n91480 );
buf ( n91484 , n42991 );
and ( n91485 , n91483 , n91484 );
nor ( n91486 , n91482 , n91485 );
buf ( n91487 , n91486 );
buf ( n91488 , n91487 );
buf ( n91489 , n36909 );
or ( n91490 , n91488 , n91489 );
nand ( n91491 , n91479 , n91490 );
buf ( n91492 , n91491 );
buf ( n91493 , n91492 );
xor ( n91494 , n91476 , n91493 );
buf ( n91495 , n91494 );
buf ( n91496 , n91495 );
xor ( n91497 , n91439 , n91496 );
buf ( n91498 , n91497 );
buf ( n91499 , n91498 );
xor ( n91500 , n91388 , n91499 );
xor ( n91501 , n91065 , n91070 );
and ( n91502 , n91501 , n91107 );
and ( n91503 , n91065 , n91070 );
or ( n91504 , n91502 , n91503 );
buf ( n91505 , n91504 );
xor ( n91506 , n91500 , n91505 );
buf ( n91507 , n91506 );
xnor ( n91508 , n91327 , n91507 );
buf ( n91509 , n91508 );
not ( n91510 , n91230 );
not ( n91511 , n91235 );
or ( n91512 , n91510 , n91511 );
not ( n91513 , n91227 );
not ( n91514 , n91238 );
or ( n91515 , n91513 , n91514 );
nand ( n91516 , n91515 , n91253 );
nand ( n91517 , n91512 , n91516 );
not ( n91518 , n91087 );
nand ( n91519 , n90256 , n91518 );
and ( n91520 , n91106 , n91519 );
nor ( n91521 , n90256 , n91518 );
nor ( n91522 , n91520 , n91521 );
not ( n91523 , n91522 );
buf ( n91524 , n38775 );
not ( n91525 , n91524 );
buf ( n91526 , n91161 );
not ( n91527 , n91526 );
or ( n91528 , n91525 , n91527 );
buf ( n91529 , n38413 );
not ( n91530 , n91529 );
buf ( n91531 , n38098 );
not ( n91532 , n91531 );
or ( n91533 , n91530 , n91532 );
buf ( n91534 , n39340 );
buf ( n91535 , n38420 );
nand ( n91536 , n91534 , n91535 );
buf ( n91537 , n91536 );
buf ( n91538 , n91537 );
nand ( n91539 , n91533 , n91538 );
buf ( n91540 , n91539 );
buf ( n91541 , n91540 );
buf ( n91542 , n38758 );
nand ( n91543 , n91541 , n91542 );
buf ( n91544 , n91543 );
buf ( n91545 , n91544 );
nand ( n91546 , n91528 , n91545 );
buf ( n91547 , n91546 );
and ( n91548 , n91523 , n91547 );
not ( n91549 , n91523 );
not ( n91550 , n91547 );
and ( n91551 , n91549 , n91550 );
nor ( n91552 , n91548 , n91551 );
not ( n91553 , n36450 );
buf ( n91554 , n36363 );
not ( n91555 , n91554 );
buf ( n91556 , n90270 );
not ( n91557 , n91556 );
and ( n91558 , n91555 , n91557 );
buf ( n91559 , n36360 );
buf ( n91560 , n41975 );
and ( n91561 , n91559 , n91560 );
nor ( n91562 , n91558 , n91561 );
buf ( n91563 , n91562 );
not ( n91564 , n91563 );
and ( n91565 , n91553 , n91564 );
nor ( n91566 , n91565 , C0 );
buf ( n91567 , n38133 );
not ( n91568 , n91567 );
buf ( n91569 , n90858 );
not ( n91570 , n91569 );
or ( n91571 , n91568 , n91570 );
buf ( n91572 , n38074 );
not ( n91573 , n91572 );
buf ( n91574 , n39518 );
not ( n91575 , n91574 );
or ( n91576 , n91573 , n91575 );
buf ( n91577 , n42596 );
buf ( n91578 , n43371 );
nand ( n91579 , n91577 , n91578 );
buf ( n91580 , n91579 );
buf ( n91581 , n91580 );
nand ( n91582 , n91576 , n91581 );
buf ( n91583 , n91582 );
buf ( n91584 , n91583 );
buf ( n91585 , n38063 );
nand ( n91586 , n91584 , n91585 );
buf ( n91587 , n91586 );
buf ( n91588 , n91587 );
nand ( n91589 , n91571 , n91588 );
buf ( n91590 , n91589 );
xor ( n91591 , n91566 , n91590 );
buf ( n91592 , n37922 );
not ( n91593 , n91592 );
buf ( n91594 , n37892 );
not ( n91595 , n91594 );
buf ( n91596 , n49178 );
not ( n91597 , n91596 );
or ( n91598 , n91595 , n91597 );
buf ( n91599 , n49179 );
buf ( n91600 , n41890 );
nand ( n91601 , n91599 , n91600 );
buf ( n91602 , n91601 );
buf ( n91603 , n91602 );
nand ( n91604 , n91598 , n91603 );
buf ( n91605 , n91604 );
buf ( n91606 , n91605 );
not ( n91607 , n91606 );
or ( n91608 , n91593 , n91607 );
buf ( n91609 , n91096 );
not ( n91610 , n91609 );
buf ( n91611 , n37875 );
nand ( n91612 , n91610 , n91611 );
buf ( n91613 , n91612 );
buf ( n91614 , n91613 );
nand ( n91615 , n91608 , n91614 );
buf ( n91616 , n91615 );
xor ( n91617 , n91591 , n91616 );
not ( n91618 , n91617 );
and ( n91619 , n91552 , n91618 );
not ( n91620 , n91552 );
and ( n91621 , n91620 , n91617 );
nor ( n91622 , n91619 , n91621 );
not ( n91623 , n91224 );
not ( n91624 , n91171 );
or ( n91625 , n91623 , n91624 );
buf ( n91626 , n91171 );
not ( n91627 , n91626 );
buf ( n91628 , n91627 );
not ( n91629 , n91628 );
not ( n91630 , n91221 );
or ( n91631 , n91629 , n91630 );
nand ( n91632 , n91631 , n91196 );
nand ( n91633 , n91625 , n91632 );
and ( n91634 , n91622 , n91633 );
not ( n91635 , n91622 );
buf ( n91636 , n91633 );
not ( n91637 , n91636 );
buf ( n91638 , n91637 );
and ( n91639 , n91635 , n91638 );
nor ( n91640 , n91634 , n91639 );
buf ( n91641 , n90843 );
not ( n91642 , n91641 );
buf ( n91643 , n90909 );
not ( n91644 , n91643 );
or ( n91645 , n91642 , n91644 );
not ( n91646 , n90846 );
not ( n91647 , n90906 );
or ( n91648 , n91646 , n91647 );
nand ( n91649 , n91648 , n90923 );
buf ( n91650 , n91649 );
nand ( n91651 , n91645 , n91650 );
buf ( n91652 , n91651 );
xor ( n91653 , n91640 , n91652 );
xor ( n91654 , n91517 , n91653 );
not ( n91655 , n91118 );
not ( n91656 , n91127 );
and ( n91657 , n91655 , n91656 );
nand ( n91658 , n91118 , n91127 );
buf ( n91659 , n90919 );
and ( n91660 , n91659 , n90923 );
not ( n91661 , n91659 );
and ( n91662 , n91661 , n90926 );
nor ( n91663 , n91660 , n91662 );
and ( n91664 , n91658 , n91663 );
nor ( n91665 , n91657 , n91664 );
xnor ( n91666 , n91654 , n91665 );
buf ( n91667 , n91666 );
xor ( n91668 , n91509 , n91667 );
buf ( n91669 , n91274 );
buf ( n91670 , n91263 );
not ( n91671 , n91670 );
buf ( n91672 , n91268 );
nand ( n91673 , n91671 , n91672 );
buf ( n91674 , n91673 );
buf ( n91675 , n91674 );
nand ( n91676 , n91669 , n91675 );
buf ( n91677 , n91676 );
buf ( n91678 , n91677 );
buf ( n91679 , n91268 );
not ( n91680 , n91679 );
buf ( n91681 , n91263 );
nand ( n91682 , n91680 , n91681 );
buf ( n91683 , n91682 );
buf ( n91684 , n91683 );
and ( n91685 , n91678 , n91684 );
buf ( n91686 , n91685 );
buf ( n91687 , n91686 );
xor ( n91688 , n91668 , n91687 );
buf ( n91689 , n91688 );
xor ( n91690 , n91131 , n91149 );
and ( n91691 , n91690 , n91276 );
and ( n91692 , n91131 , n91149 );
or ( n91693 , n91691 , n91692 );
buf ( n91694 , n91693 );
nand ( n91695 , n91689 , n91694 );
nand ( n91696 , n91279 , n91695 );
not ( n91697 , n91696 );
xor ( n91698 , n91388 , n91499 );
and ( n91699 , n91698 , n91505 );
and ( n91700 , n91388 , n91499 );
or ( n91701 , n91699 , n91700 );
buf ( n91702 , n91701 );
buf ( n91703 , n91702 );
buf ( n91704 , n38997 );
buf ( n91705 , n42280 );
and ( n91706 , n91704 , n91705 );
not ( n91707 , n91704 );
buf ( n91708 , n42277 );
and ( n91709 , n91707 , n91708 );
nor ( n91710 , n91706 , n91709 );
buf ( n91711 , n91710 );
not ( n91712 , n91711 );
not ( n91713 , n38974 );
and ( n91714 , n91712 , n91713 );
buf ( n91715 , n91287 );
not ( n91716 , n91715 );
buf ( n91717 , n91716 );
and ( n91718 , n91717 , n39395 );
nor ( n91719 , n91714 , n91718 );
buf ( n91720 , n91719 );
buf ( n91721 , n38420 );
not ( n91722 , n91721 );
buf ( n91723 , n36399 );
not ( n91724 , n91723 );
or ( n91725 , n91722 , n91724 );
buf ( n91726 , n55813 );
not ( n91727 , n91726 );
buf ( n91728 , n38413 );
nand ( n91729 , n91727 , n91728 );
buf ( n91730 , n91729 );
buf ( n91731 , n91730 );
nand ( n91732 , n91725 , n91731 );
buf ( n91733 , n91732 );
buf ( n91734 , n91733 );
buf ( n91735 , n38758 );
and ( n91736 , n91734 , n91735 );
buf ( n91737 , n91540 );
not ( n91738 , n91737 );
buf ( n91739 , n38407 );
nor ( n91740 , n91738 , n91739 );
buf ( n91741 , n91740 );
buf ( n91742 , n91741 );
nor ( n91743 , n91736 , n91742 );
buf ( n91744 , n91743 );
buf ( n91745 , n91744 );
xor ( n91746 , n91720 , n91745 );
buf ( n91747 , n91746 );
buf ( n91748 , n91747 );
xor ( n91749 , n91333 , n91359 );
and ( n91750 , n91749 , n91385 );
and ( n91751 , n91333 , n91359 );
or ( n91752 , n91750 , n91751 );
buf ( n91753 , n91752 );
buf ( n91754 , n91753 );
xnor ( n91755 , n91748 , n91754 );
buf ( n91756 , n91755 );
buf ( n91757 , n91756 );
not ( n91758 , n91757 );
buf ( n91759 , n91758 );
buf ( n91760 , n91759 );
and ( n91761 , n91703 , n91760 );
not ( n91762 , n91703 );
buf ( n91763 , n91756 );
and ( n91764 , n91762 , n91763 );
nor ( n91765 , n91761 , n91764 );
buf ( n91766 , n91765 );
buf ( n91767 , n91766 );
xor ( n91768 , n91413 , n91438 );
and ( n91769 , n91768 , n91496 );
and ( n91770 , n91413 , n91438 );
or ( n91771 , n91769 , n91770 );
buf ( n91772 , n91771 );
buf ( n91773 , n37922 );
not ( n91774 , n91773 );
not ( n91775 , n37892 );
not ( n91776 , n47319 );
or ( n91777 , n91775 , n91776 );
nand ( n91778 , n37271 , n38660 );
nand ( n91779 , n91777 , n91778 );
buf ( n91780 , n91779 );
not ( n91781 , n91780 );
or ( n91782 , n91774 , n91781 );
buf ( n91783 , n91605 );
buf ( n91784 , n37875 );
nand ( n91785 , n91783 , n91784 );
buf ( n91786 , n91785 );
buf ( n91787 , n91786 );
nand ( n91788 , n91782 , n91787 );
buf ( n91789 , n91788 );
buf ( n91790 , n91789 );
buf ( n91791 , n42565 );
not ( n91792 , n91791 );
buf ( n91793 , n42631 );
not ( n91794 , n91793 );
buf ( n91795 , n91794 );
buf ( n91796 , n91795 );
not ( n91797 , n91796 );
or ( n91798 , n91792 , n91797 );
buf ( n91799 , n91351 );
nand ( n91800 , n91798 , n91799 );
buf ( n91801 , n91800 );
buf ( n91802 , n91801 );
not ( n91803 , n91802 );
buf ( n91804 , n91803 );
buf ( n91805 , n91804 );
and ( n91806 , n91790 , n91805 );
not ( n91807 , n91790 );
buf ( n91808 , n91801 );
and ( n91809 , n91807 , n91808 );
nor ( n91810 , n91806 , n91809 );
buf ( n91811 , n91810 );
xor ( n91812 , n91461 , n91475 );
and ( n91813 , n91812 , n91493 );
and ( n91814 , n91461 , n91475 );
or ( n91815 , n91813 , n91814 );
buf ( n91816 , n91815 );
xor ( n91817 , n91811 , n91816 );
and ( n91818 , n91772 , n91817 );
not ( n91819 , n91772 );
buf ( n91820 , n91817 );
not ( n91821 , n91820 );
buf ( n91822 , n91821 );
and ( n91823 , n91819 , n91822 );
or ( n91824 , n91818 , n91823 );
buf ( n91825 , n91824 );
buf ( n91826 , n37452 );
not ( n91827 , n91826 );
buf ( n91828 , n37476 );
not ( n91829 , n91828 );
buf ( n91830 , n39407 );
not ( n91831 , n91830 );
or ( n91832 , n91829 , n91831 );
buf ( n91833 , n42941 );
buf ( n91834 , n37475 );
nand ( n91835 , n91833 , n91834 );
buf ( n91836 , n91835 );
buf ( n91837 , n91836 );
nand ( n91838 , n91832 , n91837 );
buf ( n91839 , n91838 );
buf ( n91840 , n91839 );
not ( n91841 , n91840 );
or ( n91842 , n91827 , n91841 );
buf ( n91843 , n91405 );
buf ( n91844 , n37517 );
nand ( n91845 , n91843 , n91844 );
buf ( n91846 , n91845 );
buf ( n91847 , n91846 );
nand ( n91848 , n91842 , n91847 );
buf ( n91849 , n91848 );
buf ( n91850 , n91849 );
buf ( n91851 , n39986 );
not ( n91852 , n91851 );
buf ( n91853 , n40010 );
not ( n91854 , n91853 );
buf ( n91855 , n36041 );
not ( n91856 , n91855 );
or ( n91857 , n91854 , n91856 );
buf ( n91858 , n36038 );
buf ( n91859 , n40009 );
nand ( n91860 , n91858 , n91859 );
buf ( n91861 , n91860 );
buf ( n91862 , n91861 );
nand ( n91863 , n91857 , n91862 );
buf ( n91864 , n91863 );
buf ( n91865 , n91864 );
not ( n91866 , n91865 );
or ( n91867 , n91852 , n91866 );
buf ( n91868 , n91430 );
buf ( n91869 , n40002 );
nand ( n91870 , n91868 , n91869 );
buf ( n91871 , n91870 );
buf ( n91872 , n91871 );
nand ( n91873 , n91867 , n91872 );
buf ( n91874 , n91873 );
buf ( n91875 , n91874 );
xor ( n91876 , n91850 , n91875 );
buf ( n91877 , n87681 );
not ( n91878 , n91877 );
buf ( n91879 , n91452 );
not ( n91880 , n91879 );
and ( n91881 , n91878 , n91880 );
buf ( n91882 , n39708 );
buf ( n91883 , n42530 );
and ( n91884 , n91882 , n91883 );
nor ( n91885 , n91881 , n91884 );
buf ( n91886 , n91885 );
not ( n91887 , n91886 );
not ( n91888 , n91887 );
buf ( n91889 , n43283 );
buf ( n91890 , n39664 );
nor ( n91891 , n91889 , n91890 );
buf ( n91892 , n91891 );
buf ( n91893 , n91892 );
nor ( n91894 , C0 , n91893 );
buf ( n91895 , n91894 );
not ( n91896 , n91895 );
or ( n91897 , n91888 , n91896 );
buf ( n91898 , n91895 );
not ( n91899 , n91898 );
buf ( n91900 , n91899 );
nand ( n91901 , n91900 , n91886 );
nand ( n91902 , n91897 , n91901 );
buf ( n91903 , n91566 );
not ( n91904 , n91903 );
buf ( n91905 , n91904 );
buf ( n91906 , n91905 );
not ( n91907 , n91906 );
buf ( n91908 , n91907 );
xnor ( n91909 , n91902 , n91908 );
buf ( n91910 , n91909 );
xor ( n91911 , n91876 , n91910 );
buf ( n91912 , n91911 );
buf ( n91913 , n91912 );
not ( n91914 , n91913 );
buf ( n91915 , n91914 );
buf ( n91916 , n91915 );
and ( n91917 , n91825 , n91916 );
not ( n91918 , n91825 );
buf ( n91919 , n91912 );
and ( n91920 , n91918 , n91919 );
nor ( n91921 , n91917 , n91920 );
buf ( n91922 , n91921 );
buf ( n91923 , n91922 );
buf ( n91924 , n91923 );
buf ( n91925 , n91924 );
buf ( n91926 , n91925 );
xor ( n91927 , n91767 , n91926 );
buf ( n91928 , n91927 );
buf ( n91929 , n91928 );
not ( n91930 , n91929 );
buf ( n91931 , n91930 );
buf ( n91932 , n91931 );
not ( n91933 , n91932 );
not ( n91934 , n91523 );
not ( n91935 , n91547 );
or ( n91936 , n91934 , n91935 );
and ( n91937 , n91106 , n91519 );
nor ( n91938 , n91937 , n91521 );
not ( n91939 , n91938 );
not ( n91940 , n91550 );
or ( n91941 , n91939 , n91940 );
nand ( n91942 , n91941 , n91617 );
nand ( n91943 , n91936 , n91942 );
buf ( n91944 , n91943 );
buf ( n91945 , n38150 );
not ( n91946 , n91945 );
buf ( n91947 , n37330 );
not ( n91948 , n91947 );
buf ( n91949 , n39861 );
not ( n91950 , n91949 );
or ( n91951 , n91948 , n91950 );
buf ( n91952 , n37148 );
buf ( n91953 , n37329 );
nand ( n91954 , n91952 , n91953 );
buf ( n91955 , n91954 );
buf ( n91956 , n91955 );
nand ( n91957 , n91951 , n91956 );
buf ( n91958 , n91957 );
buf ( n91959 , n91958 );
not ( n91960 , n91959 );
or ( n91961 , n91946 , n91960 );
buf ( n91962 , n91377 );
buf ( n91963 , n37403 );
nand ( n91964 , n91962 , n91963 );
buf ( n91965 , n91964 );
buf ( n91966 , n91965 );
nand ( n91967 , n91961 , n91966 );
buf ( n91968 , n91967 );
buf ( n91969 , n91968 );
buf ( n91970 , n91908 );
not ( n91971 , n91970 );
buf ( n91972 , n91616 );
not ( n91973 , n91972 );
or ( n91974 , n91971 , n91973 );
buf ( n91975 , n91616 );
buf ( n91976 , n91908 );
or ( n91977 , n91975 , n91976 );
buf ( n91978 , n91590 );
nand ( n91979 , n91977 , n91978 );
buf ( n91980 , n91979 );
buf ( n91981 , n91980 );
nand ( n91982 , n91974 , n91981 );
buf ( n91983 , n91982 );
buf ( n91984 , n91983 );
xor ( n91985 , n91969 , n91984 );
buf ( n91986 , n91469 );
not ( n91987 , n91986 );
buf ( n91988 , n39806 );
not ( n91989 , n91988 );
or ( n91990 , n91987 , n91989 );
buf ( n91991 , n39737 );
not ( n91992 , n91991 );
buf ( n91993 , n39816 );
nand ( n91994 , n91992 , n91993 );
buf ( n91995 , n91994 );
buf ( n91996 , n91995 );
nand ( n91997 , n91990 , n91996 );
buf ( n91998 , n91997 );
buf ( n91999 , n91998 );
buf ( n92000 , n36915 );
not ( n92001 , n92000 );
buf ( n92002 , n39235 );
not ( n92003 , n92002 );
buf ( n92004 , n37786 );
not ( n92005 , n92004 );
or ( n92006 , n92003 , n92005 );
buf ( n92007 , n38480 );
buf ( n92008 , n39139 );
nand ( n92009 , n92007 , n92008 );
buf ( n92010 , n92009 );
buf ( n92011 , n92010 );
nand ( n92012 , n92006 , n92011 );
buf ( n92013 , n92012 );
buf ( n92014 , n92013 );
not ( n92015 , n92014 );
or ( n92016 , n92001 , n92015 );
buf ( n92017 , n91487 );
not ( n92018 , n92017 );
buf ( n92019 , n39257 );
nand ( n92020 , n92018 , n92019 );
buf ( n92021 , n92020 );
buf ( n92022 , n92021 );
nand ( n92023 , n92016 , n92022 );
buf ( n92024 , n92023 );
buf ( n92025 , n92024 );
xor ( n92026 , n91999 , n92025 );
buf ( n92027 , n38063 );
not ( n92028 , n92027 );
buf ( n92029 , n38074 );
not ( n92030 , n92029 );
buf ( n92031 , n37717 );
not ( n92032 , n92031 );
or ( n92033 , n92030 , n92032 );
buf ( n92034 , n37695 );
buf ( n92035 , n38071 );
nand ( n92036 , n92034 , n92035 );
buf ( n92037 , n92036 );
buf ( n92038 , n92037 );
nand ( n92039 , n92033 , n92038 );
buf ( n92040 , n92039 );
buf ( n92041 , n92040 );
not ( n92042 , n92041 );
or ( n92043 , n92028 , n92042 );
buf ( n92044 , n38133 );
buf ( n92045 , n91583 );
nand ( n92046 , n92044 , n92045 );
buf ( n92047 , n92046 );
buf ( n92048 , n92047 );
nand ( n92049 , n92043 , n92048 );
buf ( n92050 , n92049 );
buf ( n92051 , n92050 );
xor ( n92052 , n92026 , n92051 );
buf ( n92053 , n92052 );
buf ( n92054 , n92053 );
xor ( n92055 , n91985 , n92054 );
buf ( n92056 , n92055 );
buf ( n92057 , n92056 );
xor ( n92058 , n91944 , n92057 );
buf ( n92059 , n92058 );
buf ( n92060 , n92059 );
not ( n92061 , n91305 );
buf ( n92062 , n91297 );
not ( n92063 , n92062 );
buf ( n92064 , n92063 );
not ( n92065 , n92064 );
or ( n92066 , n92061 , n92065 );
not ( n92067 , n91305 );
buf ( n92068 , n92067 );
not ( n92069 , n92068 );
buf ( n92070 , n91297 );
not ( n92071 , n92070 );
or ( n92072 , n92069 , n92071 );
buf ( n92073 , n91311 );
nand ( n92074 , n92072 , n92073 );
buf ( n92075 , n92074 );
nand ( n92076 , n92066 , n92075 );
buf ( n92077 , n92076 );
and ( n92078 , n92060 , n92077 );
not ( n92079 , n92060 );
buf ( n92080 , n92076 );
not ( n92081 , n92080 );
buf ( n92082 , n92081 );
buf ( n92083 , n92082 );
and ( n92084 , n92079 , n92083 );
nor ( n92085 , n92078 , n92084 );
buf ( n92086 , n92085 );
buf ( n92087 , n92086 );
buf ( n92088 , n91622 );
not ( n92089 , n92088 );
buf ( n92090 , n91638 );
not ( n92091 , n92090 );
or ( n92092 , n92089 , n92091 );
buf ( n92093 , n91652 );
nand ( n92094 , n92092 , n92093 );
buf ( n92095 , n92094 );
buf ( n92096 , n92095 );
not ( n92097 , n91622 );
nand ( n92098 , n92097 , n91633 );
buf ( n92099 , n92098 );
nand ( n92100 , n92096 , n92099 );
buf ( n92101 , n92100 );
buf ( n92102 , n92101 );
xor ( n92103 , n92087 , n92102 );
buf ( n92104 , n92103 );
buf ( n92105 , n91312 );
not ( n92106 , n92105 );
buf ( n92107 , n91507 );
not ( n92108 , n92107 );
or ( n92109 , n92106 , n92108 );
buf ( n92110 , n91507 );
buf ( n92111 , n91312 );
or ( n92112 , n92110 , n92111 );
buf ( n92113 , n91326 );
nand ( n92114 , n92112 , n92113 );
buf ( n92115 , n92114 );
buf ( n92116 , n92115 );
nand ( n92117 , n92109 , n92116 );
buf ( n92118 , n92117 );
and ( n92119 , n92104 , n92118 );
not ( n92120 , n92104 );
buf ( n92121 , n92118 );
not ( n92122 , n92121 );
buf ( n92123 , n92122 );
and ( n92124 , n92120 , n92123 );
nor ( n92125 , n92119 , n92124 );
not ( n92126 , n92125 );
buf ( n92127 , n92126 );
not ( n92128 , n92127 );
or ( n92129 , n91933 , n92128 );
nand ( n92130 , n91928 , n92125 );
buf ( n92131 , n92130 );
nand ( n92132 , n92129 , n92131 );
buf ( n92133 , n92132 );
buf ( n92134 , n92133 );
buf ( n92135 , n91517 );
not ( n92136 , n92135 );
buf ( n92137 , n91653 );
nand ( n92138 , n92136 , n92137 );
buf ( n92139 , n92138 );
buf ( n92140 , n92139 );
not ( n92141 , n92140 );
buf ( n92142 , n91665 );
not ( n92143 , n92142 );
buf ( n92144 , n92143 );
buf ( n92145 , n92144 );
not ( n92146 , n92145 );
or ( n92147 , n92141 , n92146 );
buf ( n92148 , n91653 );
not ( n92149 , n92148 );
buf ( n92150 , n91517 );
nand ( n92151 , n92149 , n92150 );
buf ( n92152 , n92151 );
buf ( n92153 , n92152 );
nand ( n92154 , n92147 , n92153 );
buf ( n92155 , n92154 );
buf ( n92156 , n92155 );
xnor ( n92157 , n92134 , n92156 );
buf ( n92158 , n92157 );
xor ( n92159 , n91509 , n91667 );
and ( n92160 , n92159 , n91687 );
and ( n92161 , n91509 , n91667 );
or ( n92162 , n92160 , n92161 );
buf ( n92163 , n92162 );
nand ( n92164 , n92158 , n92163 );
not ( n92165 , n91931 );
not ( n92166 , n92125 );
or ( n92167 , n92165 , n92166 );
buf ( n92168 , n91928 );
not ( n92169 , n92168 );
buf ( n92170 , n92126 );
not ( n92171 , n92170 );
or ( n92172 , n92169 , n92171 );
buf ( n92173 , n92155 );
nand ( n92174 , n92172 , n92173 );
buf ( n92175 , n92174 );
nand ( n92176 , n92167 , n92175 );
not ( n92177 , n92176 );
xor ( n92178 , n91850 , n91875 );
and ( n92179 , n92178 , n91910 );
and ( n92180 , n91850 , n91875 );
or ( n92181 , n92179 , n92180 );
buf ( n92182 , n92181 );
buf ( n92183 , n92182 );
buf ( n92184 , n91804 );
not ( n92185 , n92184 );
buf ( n92186 , n91789 );
not ( n92187 , n92186 );
buf ( n92188 , n92187 );
buf ( n92189 , n92188 );
not ( n92190 , n92189 );
or ( n92191 , n92185 , n92190 );
buf ( n92192 , n91816 );
nand ( n92193 , n92191 , n92192 );
buf ( n92194 , n92193 );
buf ( n92195 , n92194 );
buf ( n92196 , n91804 );
not ( n92197 , n92196 );
buf ( n92198 , n91789 );
nand ( n92199 , n92197 , n92198 );
buf ( n92200 , n92199 );
buf ( n92201 , n92200 );
nand ( n92202 , n92195 , n92201 );
buf ( n92203 , n92202 );
buf ( n92204 , n92203 );
xor ( n92205 , n92183 , n92204 );
buf ( n92206 , n91900 );
not ( n92207 , n92206 );
buf ( n92208 , n91887 );
not ( n92209 , n92208 );
or ( n92210 , n92207 , n92209 );
buf ( n92211 , n91895 );
not ( n92212 , n92211 );
buf ( n92213 , n91886 );
not ( n92214 , n92213 );
or ( n92215 , n92212 , n92214 );
buf ( n92216 , n91905 );
nand ( n92217 , n92215 , n92216 );
buf ( n92218 , n92217 );
buf ( n92219 , n92218 );
nand ( n92220 , n92210 , n92219 );
buf ( n92221 , n92220 );
buf ( n92222 , n92221 );
buf ( n92223 , n37875 );
not ( n92224 , n92223 );
buf ( n92225 , n91779 );
not ( n92226 , n92225 );
or ( n92227 , n92224 , n92226 );
buf ( n92228 , n39551 );
buf ( n92229 , n37922 );
nand ( n92230 , n92228 , n92229 );
buf ( n92231 , n92230 );
buf ( n92232 , n92231 );
nand ( n92233 , n92227 , n92232 );
buf ( n92234 , n92233 );
buf ( n92235 , n92234 );
xor ( n92236 , n92222 , n92235 );
buf ( n92237 , n39986 );
not ( n92238 , n92237 );
buf ( n92239 , n40022 );
not ( n92240 , n92239 );
or ( n92241 , n92238 , n92240 );
buf ( n92242 , n91864 );
buf ( n92243 , n40002 );
nand ( n92244 , n92242 , n92243 );
buf ( n92245 , n92244 );
buf ( n92246 , n92245 );
nand ( n92247 , n92241 , n92246 );
buf ( n92248 , n92247 );
buf ( n92249 , n92248 );
xor ( n92250 , n92236 , n92249 );
buf ( n92251 , n92250 );
buf ( n92252 , n92251 );
xor ( n92253 , n92205 , n92252 );
buf ( n92254 , n92253 );
buf ( n92255 , n92254 );
buf ( n92256 , n91822 );
not ( n92257 , n92256 );
buf ( n92258 , n91772 );
not ( n92259 , n92258 );
or ( n92260 , n92257 , n92259 );
buf ( n92261 , n91822 );
buf ( n92262 , n91772 );
or ( n92263 , n92261 , n92262 );
buf ( n92264 , n91912 );
nand ( n92265 , n92263 , n92264 );
buf ( n92266 , n92265 );
buf ( n92267 , n92266 );
nand ( n92268 , n92260 , n92267 );
buf ( n92269 , n92268 );
buf ( n92270 , n92269 );
xor ( n92271 , n91999 , n92025 );
and ( n92272 , n92271 , n92051 );
and ( n92273 , n91999 , n92025 );
or ( n92274 , n92272 , n92273 );
buf ( n92275 , n92274 );
buf ( n92276 , n92275 );
buf ( n92277 , n38775 );
not ( n92278 , n92277 );
buf ( n92279 , n91733 );
not ( n92280 , n92279 );
or ( n92281 , n92278 , n92280 );
buf ( n92282 , n40071 );
buf ( n92283 , n38758 );
nand ( n92284 , n92282 , n92283 );
buf ( n92285 , n92284 );
buf ( n92286 , n92285 );
nand ( n92287 , n92281 , n92286 );
buf ( n92288 , n92287 );
buf ( n92289 , n92288 );
xor ( n92290 , n92276 , n92289 );
buf ( n92291 , n38133 );
not ( n92292 , n92291 );
buf ( n92293 , n92040 );
not ( n92294 , n92293 );
or ( n92295 , n92292 , n92294 );
buf ( n92296 , n39628 );
buf ( n92297 , n38063 );
nand ( n92298 , n92296 , n92297 );
buf ( n92299 , n92298 );
buf ( n92300 , n92299 );
nand ( n92301 , n92295 , n92300 );
buf ( n92302 , n92301 );
buf ( n92303 , n92302 );
buf ( n92304 , n36988 );
not ( n92305 , n92304 );
buf ( n92306 , n92013 );
not ( n92307 , n92306 );
or ( n92308 , n92305 , n92307 );
buf ( n92309 , n39529 );
buf ( n92310 , n36915 );
nand ( n92311 , n92309 , n92310 );
buf ( n92312 , n92311 );
buf ( n92313 , n92312 );
nand ( n92314 , n92308 , n92313 );
buf ( n92315 , n92314 );
buf ( n92316 , n92315 );
xor ( n92317 , n92303 , n92316 );
buf ( n92318 , n37517 );
not ( n92319 , n92318 );
buf ( n92320 , n91839 );
not ( n92321 , n92320 );
or ( n92322 , n92319 , n92321 );
buf ( n92323 , n37449 );
not ( n92324 , n92323 );
buf ( n92325 , n40044 );
nand ( n92326 , n92324 , n92325 );
buf ( n92327 , n92326 );
buf ( n92328 , n92327 );
nand ( n92329 , n92322 , n92328 );
buf ( n92330 , n92329 );
buf ( n92331 , n92330 );
xor ( n92332 , n92317 , n92331 );
buf ( n92333 , n92332 );
buf ( n92334 , n92333 );
xor ( n92335 , n92290 , n92334 );
buf ( n92336 , n92335 );
buf ( n92337 , n92336 );
xor ( n92338 , n92270 , n92337 );
buf ( n92339 , n92338 );
buf ( n92340 , n92339 );
not ( n92341 , n92340 );
xor ( n92342 , n92255 , n92341 );
buf ( n92343 , n92342 );
buf ( n92344 , n92343 );
buf ( n92345 , n92086 );
buf ( n92346 , n92101 );
or ( n92347 , n92345 , n92346 );
buf ( n92348 , n92347 );
buf ( n92349 , n92348 );
buf ( n92350 , n92118 );
and ( n92351 , n92349 , n92350 );
and ( n92352 , n92087 , n92102 );
buf ( n92353 , n92352 );
buf ( n92354 , n92353 );
nor ( n92355 , n92351 , n92354 );
buf ( n92356 , n92355 );
buf ( n92357 , n92356 );
xor ( n92358 , n92344 , n92357 );
or ( n92359 , n91943 , n92056 );
buf ( n92360 , n92359 );
buf ( n92361 , n92076 );
and ( n92362 , n92360 , n92361 );
and ( n92363 , n91944 , n92057 );
buf ( n92364 , n92363 );
buf ( n92365 , n92364 );
nor ( n92366 , n92362 , n92365 );
buf ( n92367 , n92366 );
buf ( n92368 , n92367 );
xor ( n92369 , n91969 , n91984 );
and ( n92370 , n92369 , n92054 );
and ( n92371 , n91969 , n91984 );
or ( n92372 , n92370 , n92371 );
buf ( n92373 , n92372 );
xor ( n92374 , n39699 , n39723 );
xor ( n92375 , n92374 , n39756 );
buf ( n92376 , n92375 );
buf ( n92377 , n92376 );
buf ( n92378 , n37403 );
not ( n92379 , n92378 );
buf ( n92380 , n91958 );
not ( n92381 , n92380 );
or ( n92382 , n92379 , n92381 );
nand ( n92383 , n40093 , n38150 );
buf ( n92384 , n92383 );
nand ( n92385 , n92382 , n92384 );
buf ( n92386 , n92385 );
buf ( n92387 , n92386 );
xor ( n92388 , n92377 , n92387 );
buf ( n92389 , n39395 );
not ( n92390 , n92389 );
buf ( n92391 , n91711 );
not ( n92392 , n92391 );
buf ( n92393 , n92392 );
buf ( n92394 , n92393 );
not ( n92395 , n92394 );
or ( n92396 , n92390 , n92395 );
buf ( n92397 , n39592 );
buf ( n92398 , n39374 );
nand ( n92399 , n92397 , n92398 );
buf ( n92400 , n92399 );
buf ( n92401 , n92400 );
nand ( n92402 , n92396 , n92401 );
buf ( n92403 , n92402 );
buf ( n92404 , n92403 );
xor ( n92405 , n92388 , n92404 );
buf ( n92406 , n92405 );
buf ( n92407 , n92406 );
not ( n92408 , n92407 );
buf ( n92409 , n92408 );
and ( n92410 , n92373 , n92409 );
not ( n92411 , n92373 );
and ( n92412 , n92411 , n92406 );
nor ( n92413 , n92410 , n92412 );
buf ( n92414 , n91753 );
buf ( n92415 , n91719 );
buf ( n92416 , n91744 );
nand ( n92417 , n92415 , n92416 );
buf ( n92418 , n92417 );
buf ( n92419 , n92418 );
and ( n92420 , n92414 , n92419 );
buf ( n92421 , n91744 );
buf ( n92422 , n91719 );
nor ( n92423 , n92421 , n92422 );
buf ( n92424 , n92423 );
buf ( n92425 , n92424 );
nor ( n92426 , n92420 , n92425 );
buf ( n92427 , n92426 );
buf ( n92428 , n92427 );
not ( n92429 , n92428 );
buf ( n92430 , n92429 );
and ( n92431 , n92413 , n92430 );
not ( n92432 , n92413 );
and ( n92433 , n92432 , n92427 );
nor ( n92434 , n92431 , n92433 );
buf ( n92435 , n92434 );
xor ( n92436 , n92368 , n92435 );
buf ( n92437 , n91922 );
buf ( n92438 , n91756 );
nand ( n92439 , n92437 , n92438 );
buf ( n92440 , n92439 );
buf ( n92441 , n92440 );
buf ( n92442 , n91702 );
and ( n92443 , n92441 , n92442 );
buf ( n92444 , n91922 );
buf ( n92445 , n91756 );
nor ( n92446 , n92444 , n92445 );
buf ( n92447 , n92446 );
buf ( n92448 , n92447 );
nor ( n92449 , n92443 , n92448 );
buf ( n92450 , n92449 );
buf ( n92451 , n92450 );
xor ( n92452 , n92436 , n92451 );
buf ( n92453 , n92452 );
buf ( n92454 , n92453 );
xor ( n92455 , n92358 , n92454 );
buf ( n92456 , n92455 );
nand ( n92457 , n92177 , n92456 );
nand ( n92458 , n91697 , n92164 , n92457 );
buf ( n92459 , n92458 );
not ( n92460 , n92459 );
buf ( n92461 , n92460 );
buf ( n92462 , n39949 );
not ( n92463 , n92462 );
buf ( n92464 , n39878 );
not ( n92465 , n92464 );
or ( n92466 , n92463 , n92465 );
buf ( n92467 , n39878 );
buf ( n92468 , n39949 );
or ( n92469 , n92467 , n92468 );
nand ( n92470 , n92466 , n92469 );
buf ( n92471 , n92470 );
buf ( n92472 , n92471 );
buf ( n92473 , n39913 );
and ( n92474 , n92472 , n92473 );
not ( n92475 , n92472 );
buf ( n92476 , n39959 );
and ( n92477 , n92475 , n92476 );
nor ( n92478 , n92474 , n92477 );
buf ( n92479 , n92478 );
buf ( n92480 , n92479 );
buf ( n92481 , n39563 );
buf ( n92482 , n39568 );
xor ( n92483 , n92481 , n92482 );
buf ( n92484 , n39766 );
xnor ( n92485 , n92483 , n92484 );
buf ( n92486 , n92485 );
buf ( n92487 , n92486 );
xor ( n92488 , n92480 , n92487 );
xor ( n92489 , n92303 , n92316 );
and ( n92490 , n92489 , n92331 );
and ( n92491 , n92303 , n92316 );
or ( n92492 , n92490 , n92491 );
buf ( n92493 , n92492 );
buf ( n92494 , n92493 );
not ( n92495 , n92494 );
xor ( n92496 , n39599 , n39639 );
xor ( n92497 , n92496 , n39760 );
buf ( n92498 , n92497 );
nand ( n92499 , n92495 , n92498 );
buf ( n92500 , n92499 );
buf ( n92501 , n92500 );
xor ( n92502 , n92222 , n92235 );
and ( n92503 , n92502 , n92249 );
and ( n92504 , n92222 , n92235 );
or ( n92505 , n92503 , n92504 );
buf ( n92506 , n92505 );
buf ( n92507 , n92506 );
and ( n92508 , n92501 , n92507 );
buf ( n92509 , n92493 );
not ( n92510 , n92509 );
buf ( n92511 , n92497 );
nor ( n92512 , n92510 , n92511 );
buf ( n92513 , n92512 );
buf ( n92514 , n92513 );
nor ( n92515 , n92508 , n92514 );
buf ( n92516 , n92515 );
buf ( n92517 , n92516 );
and ( n92518 , n92488 , n92517 );
and ( n92519 , n92480 , n92487 );
or ( n92520 , n92518 , n92519 );
buf ( n92521 , n92520 );
not ( n92522 , n92521 );
buf ( n92523 , n39969 );
buf ( n92524 , n40121 );
and ( n92525 , n92523 , n92524 );
not ( n92526 , n92523 );
buf ( n92527 , n40124 );
and ( n92528 , n92526 , n92527 );
nor ( n92529 , n92525 , n92528 );
buf ( n92530 , n92529 );
buf ( n92531 , n92530 );
buf ( n92532 , n39780 );
and ( n92533 , n92531 , n92532 );
not ( n92534 , n92531 );
buf ( n92535 , n39780 );
not ( n92536 , n92535 );
buf ( n92537 , n92536 );
buf ( n92538 , n92537 );
and ( n92539 , n92534 , n92538 );
or ( n92540 , n92533 , n92539 );
buf ( n92541 , n92540 );
xor ( n92542 , n92522 , n92541 );
xor ( n92543 , n40057 , n40061 );
xor ( n92544 , n92543 , n40117 );
buf ( n92545 , n92544 );
buf ( n92546 , n92545 );
not ( n92547 , n92546 );
buf ( n92548 , n92547 );
buf ( n92549 , n92548 );
not ( n92550 , n92549 );
xor ( n92551 , n92493 , n92506 );
buf ( n92552 , n92551 );
buf ( n92553 , n92497 );
not ( n92554 , n92553 );
buf ( n92555 , n92554 );
buf ( n92556 , n92555 );
and ( n92557 , n92552 , n92556 );
not ( n92558 , n92552 );
buf ( n92559 , n92497 );
and ( n92560 , n92558 , n92559 );
nor ( n92561 , n92557 , n92560 );
buf ( n92562 , n92561 );
buf ( n92563 , n92562 );
not ( n92564 , n92563 );
buf ( n92565 , n40104 );
buf ( n92566 , n40081 );
and ( n92567 , n92565 , n92566 );
not ( n92568 , n92565 );
buf ( n92569 , n40084 );
and ( n92570 , n92568 , n92569 );
nor ( n92571 , n92567 , n92570 );
buf ( n92572 , n92571 );
buf ( n92573 , n92572 );
not ( n92574 , n92573 );
buf ( n92575 , n40098 );
buf ( n92576 , n92575 );
not ( n92577 , n92576 );
or ( n92578 , n92574 , n92577 );
buf ( n92579 , n92572 );
not ( n92580 , n92579 );
buf ( n92581 , n92580 );
buf ( n92582 , n92581 );
not ( n92583 , n92575 );
buf ( n92584 , n92583 );
nand ( n92585 , n92582 , n92584 );
buf ( n92586 , n92585 );
buf ( n92587 , n92586 );
nand ( n92588 , n92578 , n92587 );
buf ( n92589 , n92588 );
buf ( n92590 , n92589 );
not ( n92591 , n92590 );
or ( n92592 , n92564 , n92591 );
buf ( n92593 , n92562 );
buf ( n92594 , n92589 );
or ( n92595 , n92593 , n92594 );
xor ( n92596 , n92183 , n92204 );
and ( n92597 , n92596 , n92252 );
and ( n92598 , n92183 , n92204 );
or ( n92599 , n92597 , n92598 );
buf ( n92600 , n92599 );
buf ( n92601 , n92600 );
nand ( n92602 , n92595 , n92601 );
buf ( n92603 , n92602 );
buf ( n92604 , n92603 );
nand ( n92605 , n92592 , n92604 );
buf ( n92606 , n92605 );
buf ( n92607 , n92606 );
not ( n92608 , n92607 );
buf ( n92609 , n92608 );
buf ( n92610 , n92609 );
not ( n92611 , n92610 );
or ( n92612 , n92550 , n92611 );
xor ( n92613 , n40026 , n40030 );
xor ( n92614 , n92613 , n40052 );
buf ( n92615 , n92614 );
buf ( n92616 , n92615 );
xor ( n92617 , n92377 , n92387 );
and ( n92618 , n92617 , n92404 );
and ( n92619 , n92377 , n92387 );
or ( n92620 , n92618 , n92619 );
buf ( n92621 , n92620 );
buf ( n92622 , n92621 );
or ( n92623 , n92616 , n92622 );
xor ( n92624 , n92276 , n92289 );
and ( n92625 , n92624 , n92334 );
and ( n92626 , n92276 , n92289 );
or ( n92627 , n92625 , n92626 );
buf ( n92628 , n92627 );
buf ( n92629 , n92628 );
nand ( n92630 , n92623 , n92629 );
buf ( n92631 , n92630 );
buf ( n92632 , n92631 );
buf ( n92633 , n92621 );
buf ( n92634 , n92615 );
nand ( n92635 , n92633 , n92634 );
buf ( n92636 , n92635 );
buf ( n92637 , n92636 );
nand ( n92638 , n92632 , n92637 );
buf ( n92639 , n92638 );
buf ( n92640 , n92639 );
nand ( n92641 , n92612 , n92640 );
buf ( n92642 , n92641 );
buf ( n92643 , n92642 );
buf ( n92644 , n92606 );
buf ( n92645 , n92545 );
nand ( n92646 , n92644 , n92645 );
buf ( n92647 , n92646 );
buf ( n92648 , n92647 );
and ( n92649 , n92643 , n92648 );
buf ( n92650 , n92649 );
xnor ( n92651 , n92542 , n92650 );
xor ( n92652 , n92480 , n92487 );
xor ( n92653 , n92652 , n92517 );
buf ( n92654 , n92653 );
not ( n92655 , n92430 );
not ( n92656 , n92406 );
or ( n92657 , n92655 , n92656 );
not ( n92658 , n92427 );
not ( n92659 , n92409 );
or ( n92660 , n92658 , n92659 );
nand ( n92661 , n92660 , n92373 );
nand ( n92662 , n92657 , n92661 );
buf ( n92663 , n92662 );
not ( n92664 , n92663 );
buf ( n92665 , n92621 );
buf ( n92666 , n92615 );
xor ( n92667 , n92665 , n92666 );
buf ( n92668 , n92628 );
xnor ( n92669 , n92667 , n92668 );
buf ( n92670 , n92669 );
buf ( n92671 , n92670 );
not ( n92672 , n92671 );
buf ( n92673 , n92672 );
buf ( n92674 , n92673 );
not ( n92675 , n92674 );
or ( n92676 , n92664 , n92675 );
buf ( n92677 , n92662 );
not ( n92678 , n92677 );
buf ( n92679 , n92678 );
buf ( n92680 , n92679 );
not ( n92681 , n92680 );
buf ( n92682 , n92670 );
not ( n92683 , n92682 );
or ( n92684 , n92681 , n92683 );
buf ( n92685 , n92254 );
buf ( n92686 , n92336 );
or ( n92687 , n92685 , n92686 );
buf ( n92688 , n92269 );
nand ( n92689 , n92687 , n92688 );
buf ( n92690 , n92689 );
buf ( n92691 , n92690 );
buf ( n92692 , n92254 );
buf ( n92693 , n92336 );
nand ( n92694 , n92692 , n92693 );
buf ( n92695 , n92694 );
buf ( n92696 , n92695 );
nand ( n92697 , n92691 , n92696 );
buf ( n92698 , n92697 );
buf ( n92699 , n92698 );
nand ( n92700 , n92684 , n92699 );
buf ( n92701 , n92700 );
buf ( n92702 , n92701 );
nand ( n92703 , n92676 , n92702 );
buf ( n92704 , n92703 );
buf ( n92705 , n92704 );
not ( n92706 , n92705 );
buf ( n92707 , n92706 );
xor ( n92708 , n92654 , n92707 );
buf ( n92709 , n92545 );
buf ( n92710 , n92639 );
xor ( n92711 , n92709 , n92710 );
buf ( n92712 , n92711 );
buf ( n92713 , n92712 );
buf ( n92714 , n92609 );
and ( n92715 , n92713 , n92714 );
not ( n92716 , n92713 );
buf ( n92717 , n92606 );
and ( n92718 , n92716 , n92717 );
nor ( n92719 , n92715 , n92718 );
buf ( n92720 , n92719 );
and ( n92721 , n92708 , n92720 );
and ( n92722 , n92654 , n92707 );
or ( n92723 , n92721 , n92722 );
nand ( n92724 , n92651 , n92723 );
buf ( n92725 , n92589 );
buf ( n92726 , n92600 );
xor ( n92727 , n92725 , n92726 );
buf ( n92728 , n92562 );
xnor ( n92729 , n92727 , n92728 );
buf ( n92730 , n92729 );
buf ( n92731 , n92730 );
xor ( n92732 , n92368 , n92435 );
and ( n92733 , n92732 , n92451 );
and ( n92734 , n92368 , n92435 );
or ( n92735 , n92733 , n92734 );
buf ( n92736 , n92735 );
buf ( n92737 , n92736 );
xor ( n92738 , n92731 , n92737 );
buf ( n92739 , n92670 );
buf ( n92740 , n92679 );
and ( n92741 , n92739 , n92740 );
not ( n92742 , n92739 );
buf ( n92743 , n92662 );
and ( n92744 , n92742 , n92743 );
nor ( n92745 , n92741 , n92744 );
buf ( n92746 , n92745 );
buf ( n92747 , n92746 );
buf ( n92748 , n92698 );
not ( n92749 , n92748 );
buf ( n92750 , n92749 );
buf ( n92751 , n92750 );
and ( n92752 , n92747 , n92751 );
not ( n92753 , n92747 );
buf ( n92754 , n92698 );
and ( n92755 , n92753 , n92754 );
nor ( n92756 , n92752 , n92755 );
buf ( n92757 , n92756 );
buf ( n92758 , n92757 );
and ( n92759 , n92738 , n92758 );
and ( n92760 , n92731 , n92737 );
or ( n92761 , n92759 , n92760 );
buf ( n92762 , n92761 );
xor ( n92763 , n92654 , n92707 );
xor ( n92764 , n92763 , n92720 );
nand ( n92765 , n92762 , n92764 );
xor ( n92766 , n92731 , n92737 );
xor ( n92767 , n92766 , n92758 );
buf ( n92768 , n92767 );
xor ( n92769 , n92344 , n92357 );
and ( n92770 , n92769 , n92454 );
and ( n92771 , n92344 , n92357 );
or ( n92772 , n92770 , n92771 );
buf ( n92773 , n92772 );
nand ( n92774 , n92768 , n92773 );
nand ( n92775 , n92724 , n92765 , n92774 );
buf ( n92776 , n92775 );
buf ( n92777 , n92530 );
buf ( n92778 , n39780 );
and ( n92779 , n92777 , n92778 );
not ( n92780 , n92777 );
buf ( n92781 , n92537 );
and ( n92782 , n92780 , n92781 );
or ( n92783 , n92779 , n92782 );
buf ( n92784 , n92783 );
or ( n92785 , n92784 , n92521 );
and ( n92786 , n92785 , n92650 );
and ( n92787 , n92784 , n92521 );
nor ( n92788 , n92786 , n92787 );
not ( n92789 , n92788 );
not ( n92790 , n40162 );
not ( n92791 , n40137 );
not ( n92792 , n92791 );
or ( n92793 , n92790 , n92792 );
nand ( n92794 , n40137 , n40161 );
nand ( n92795 , n92793 , n92794 );
and ( n92796 , n92795 , n40155 );
not ( n92797 , n92795 );
and ( n92798 , n92797 , n40156 );
nor ( n92799 , n92796 , n92798 );
nand ( n92800 , n92789 , n92799 );
buf ( n92801 , n92800 );
not ( n92802 , n92801 );
buf ( n92803 , n92802 );
buf ( n92804 , n92803 );
nor ( n92805 , n92776 , n92804 );
buf ( n92806 , n92805 );
and ( n92807 , n88818 , n90832 , n92461 , n92806 );
nand ( n92808 , n86691 , n92807 );
buf ( n92809 , n90811 );
not ( n92810 , n92809 );
not ( n92811 , n90830 );
buf ( n92812 , n89849 );
buf ( n92813 , n89854 );
nand ( n92814 , n92812 , n92813 );
buf ( n92815 , n92814 );
or ( n92816 , n89843 , n92815 );
buf ( n92817 , n89815 );
buf ( n92818 , n89842 );
nand ( n92819 , n92817 , n92818 );
buf ( n92820 , n92819 );
nand ( n92821 , n92816 , n92820 );
not ( n92822 , n92821 );
or ( n92823 , n92811 , n92822 );
not ( n92824 , n90827 );
not ( n92825 , n90829 );
nand ( n92826 , n92824 , n92825 );
nand ( n92827 , n92823 , n92826 );
not ( n92828 , n92827 );
or ( n92829 , n92810 , n92828 );
nor ( n92830 , n92768 , n92773 );
not ( n92831 , n92830 );
not ( n92832 , n92765 );
or ( n92833 , n92831 , n92832 );
buf ( n92834 , n92764 );
not ( n92835 , n92834 );
buf ( n92836 , n92835 );
buf ( n92837 , n92762 );
not ( n92838 , n92837 );
buf ( n92839 , n92838 );
nand ( n92840 , n92836 , n92839 );
nand ( n92841 , n92833 , n92840 );
nand ( n92842 , n92841 , n92800 , n92724 );
nor ( n92843 , n92723 , n92651 );
and ( n92844 , n92843 , n92800 );
not ( n92845 , n92788 );
nor ( n92846 , n92845 , n92799 );
nor ( n92847 , n92844 , n92846 );
nand ( n92848 , n92842 , n92847 );
not ( n92849 , n90810 );
nand ( n92850 , n92849 , n90767 );
not ( n92851 , n92850 );
nor ( n92852 , n92848 , n92851 );
nand ( n92853 , n92829 , n92852 );
not ( n92854 , n92457 );
buf ( n92855 , n92164 );
not ( n92856 , n92855 );
not ( n92857 , n91695 );
not ( n92858 , n90837 );
nor ( n92859 , n92858 , n91278 );
not ( n92860 , n92859 );
or ( n92861 , n92857 , n92860 );
buf ( n92862 , n91689 );
not ( n92863 , n92862 );
buf ( n92864 , n92863 );
buf ( n92865 , n91694 );
not ( n92866 , n92865 );
buf ( n92867 , n92866 );
nand ( n92868 , n92864 , n92867 );
nand ( n92869 , n92861 , n92868 );
buf ( n92870 , n92869 );
not ( n92871 , n92870 );
or ( n92872 , n92856 , n92871 );
buf ( n92873 , n92158 );
buf ( n92874 , n92163 );
or ( n92875 , n92873 , n92874 );
buf ( n92876 , n92875 );
buf ( n92877 , n92876 );
nand ( n92878 , n92872 , n92877 );
buf ( n92879 , n92878 );
not ( n92880 , n92879 );
or ( n92881 , n92854 , n92880 );
not ( n92882 , n92456 );
nand ( n92883 , n92882 , n92176 );
nand ( n92884 , n92881 , n92883 );
nor ( n92885 , n92853 , n92884 );
not ( n92886 , n92885 );
not ( n92887 , n87768 );
buf ( n92888 , n87775 );
not ( n92889 , n92888 );
buf ( n92890 , n92889 );
nand ( n92891 , n92887 , n92890 );
nand ( n92892 , n87246 , n86705 );
nand ( n92893 , n92891 , n92892 );
not ( n92894 , n87776 );
nor ( n92895 , n88310 , n92894 );
not ( n92896 , n88815 );
nand ( n92897 , n92893 , n92895 , n92896 );
buf ( n92898 , n88807 );
buf ( n92899 , n88812 );
nand ( n92900 , n92898 , n92899 );
buf ( n92901 , n92900 );
not ( n92902 , n92901 );
nand ( n92903 , n88309 , n87787 );
not ( n92904 , n92903 );
or ( n92905 , n92902 , n92904 );
nand ( n92906 , n92905 , n92896 );
nand ( n92907 , n92897 , n92906 );
nand ( n92908 , n92907 , n90832 );
not ( n92909 , n92908 );
or ( n92910 , n92886 , n92909 );
not ( n92911 , n92457 );
not ( n92912 , n92879 );
or ( n92913 , n92911 , n92912 );
nand ( n92914 , n92913 , n92883 );
not ( n92915 , n92914 );
not ( n92916 , n92848 );
buf ( n92917 , n92916 );
buf ( n92918 , n92458 );
nand ( n92919 , n92917 , n92918 );
buf ( n92920 , n92919 );
not ( n92921 , n92920 );
and ( n92922 , n92915 , n92921 );
buf ( n92923 , n92806 );
buf ( n92924 , n92848 );
nor ( n92925 , n92923 , n92924 );
buf ( n92926 , n92925 );
nor ( n92927 , n92922 , n92926 );
nand ( n92928 , n92910 , n92927 );
not ( n92929 , n49693 );
nor ( n92930 , n53388 , n53376 );
nand ( n92931 , n52859 , n92930 );
not ( n92932 , n92931 );
not ( n92933 , n52858 );
not ( n92934 , n92933 );
not ( n92935 , n51584 );
not ( n92936 , n92935 );
or ( n92937 , n92934 , n92936 );
buf ( n92938 , n53427 );
not ( n92939 , n92938 );
buf ( n92940 , n92939 );
not ( n92941 , n53431 );
nand ( n92942 , n92940 , n92941 );
nand ( n92943 , n92937 , n92942 );
or ( n92944 , n92932 , n92943 );
nand ( n92945 , n53435 , n53440 );
and ( n92946 , n92945 , n53432 );
nand ( n92947 , n92944 , n92946 );
buf ( n92948 , n92947 );
or ( n92949 , n53435 , n53440 );
buf ( n92950 , n92949 );
nand ( n92951 , n92948 , n92950 );
buf ( n92952 , n92951 );
not ( n92953 , n92952 );
or ( n92954 , n92929 , n92953 );
buf ( n92955 , n47221 );
buf ( n92956 , n46538 );
nor ( n92957 , n92955 , n92956 );
buf ( n92958 , n92957 );
buf ( n92959 , n92958 );
buf ( n92960 , n48099 );
buf ( n92961 , n47228 );
nor ( n92962 , n92960 , n92961 );
buf ( n92963 , n92962 );
buf ( n92964 , n92963 );
nor ( n92965 , n92959 , n92964 );
buf ( n92966 , n92965 );
nor ( n92967 , n48105 , n49128 );
nand ( n92968 , n92967 , n48102 );
nand ( n92969 , n92966 , n92968 );
buf ( n92970 , n47224 );
buf ( n92971 , n49690 );
buf ( n92972 , n92971 );
buf ( n92973 , n92972 );
and ( n92974 , n92969 , n92970 , n92973 );
buf ( n92975 , n49136 );
not ( n92976 , n92975 );
buf ( n92977 , n49687 );
buf ( n92978 , n92977 );
nor ( n92979 , n92976 , n92978 );
buf ( n92980 , n92979 );
nor ( n92981 , n92974 , n92980 );
nand ( n92982 , n92954 , n92981 );
not ( n92983 , n92982 );
not ( n92984 , n92983 );
buf ( n92985 , n53391 );
buf ( n92986 , n53442 );
and ( n92987 , n92985 , n92986 );
buf ( n92988 , n92987 );
and ( n92989 , n92988 , n49693 );
nand ( n92990 , n63510 , n63519 );
not ( n92991 , n92990 );
nor ( n92992 , n59126 , n92991 );
not ( n92993 , n92992 );
buf ( n92994 , n61208 );
buf ( n92995 , n62044 );
nand ( n92996 , n92994 , n92995 );
buf ( n92997 , n92996 );
nand ( n92998 , n62052 , n63471 );
nand ( n92999 , n92997 , n92998 );
nand ( n93000 , n92999 , n63502 , n62048 );
buf ( n93001 , n63507 );
buf ( n93002 , n63516 );
nand ( n93003 , n93001 , n93002 );
buf ( n93004 , n93003 );
nand ( n93005 , n63491 , n63498 );
buf ( n93006 , n93005 );
nand ( n93007 , n93000 , n93004 , n93006 );
not ( n93008 , n93007 );
or ( n93009 , n92993 , n93008 );
buf ( n93010 , n55500 );
not ( n93011 , n93010 );
buf ( n93012 , n93011 );
nand ( n93013 , n57034 , n57038 );
buf ( n93014 , n57028 );
not ( n93015 , n93014 );
buf ( n93016 , n93015 );
nand ( n93017 , n93012 , n93013 , n93016 );
not ( n93018 , n57034 );
not ( n93019 , n57038 );
nand ( n93020 , n93018 , n93019 );
nand ( n93021 , n93017 , n93020 );
nor ( n93022 , n57951 , n59122 );
not ( n93023 , n93022 );
nand ( n93024 , n57946 , n57942 );
not ( n93025 , n93024 );
or ( n93026 , n93023 , n93025 );
buf ( n93027 , n57946 );
not ( n93028 , n93027 );
buf ( n93029 , n93028 );
buf ( n93030 , n57942 );
not ( n93031 , n93030 );
buf ( n93032 , n93031 );
nand ( n93033 , n93029 , n93032 );
nand ( n93034 , n93026 , n93033 );
nor ( n93035 , n93021 , n93034 );
nand ( n93036 , n93009 , n93035 );
not ( n93037 , n93020 );
buf ( n93038 , n57029 );
not ( n93039 , n93038 );
buf ( n93040 , n93039 );
not ( n93041 , n93040 );
or ( n93042 , n93037 , n93041 );
not ( n93043 , n57039 );
not ( n93044 , n93043 );
nand ( n93045 , n93042 , n93044 );
not ( n93046 , n93045 );
nand ( n93047 , n92989 , n93036 , n93046 );
not ( n93048 , n93047 );
or ( n93049 , n92984 , n93048 );
nand ( n93050 , n93049 , n92807 );
nand ( n93051 , n92808 , n92928 , n93050 );
not ( n93052 , n93051 );
or ( n93053 , n41567 , n93052 );
not ( n93054 , n41562 );
not ( n93055 , n41322 );
buf ( n93056 , n40495 );
not ( n93057 , n93056 );
buf ( n93058 , n39463 );
not ( n93059 , n93058 );
buf ( n93060 , n40184 );
buf ( n93061 , n40170 );
nand ( n93062 , n93060 , n93061 );
buf ( n93063 , n93062 );
or ( n93064 , n93063 , n40201 );
buf ( n93065 , n40190 );
buf ( n93066 , n40200 );
nand ( n93067 , n93065 , n93066 );
buf ( n93068 , n93067 );
nand ( n93069 , n93064 , n93068 );
buf ( n93070 , n93069 );
not ( n93071 , n93070 );
or ( n93072 , n93059 , n93071 );
buf ( n93073 , n39109 );
buf ( n93074 , n39460 );
or ( n93075 , n93073 , n93074 );
buf ( n93076 , n93075 );
buf ( n93077 , n93076 );
nand ( n93078 , n93072 , n93077 );
buf ( n93079 , n93078 );
buf ( n93080 , n93079 );
not ( n93081 , n93080 );
or ( n93082 , n93057 , n93081 );
buf ( n93083 , n40492 );
buf ( n93084 , n40486 );
or ( n93085 , n93083 , n93084 );
buf ( n93086 , n93085 );
buf ( n93087 , n93086 );
nand ( n93088 , n93082 , n93087 );
buf ( n93089 , n93088 );
not ( n93090 , n93089 );
or ( n93091 , n93055 , n93090 );
buf ( n93092 , n41259 );
not ( n93093 , n93092 );
not ( n93094 , n41052 );
buf ( n93095 , n41301 );
buf ( n93096 , n41317 );
buf ( n93097 , n41314 );
nand ( n93098 , n93096 , n93097 );
buf ( n93099 , n93098 );
buf ( n93100 , n93099 );
or ( n93101 , n93095 , n93100 );
buf ( n93102 , n41265 );
buf ( n93103 , n41298 );
nand ( n93104 , n93102 , n93103 );
buf ( n93105 , n93104 );
buf ( n93106 , n93105 );
nand ( n93107 , n93101 , n93106 );
buf ( n93108 , n93107 );
not ( n93109 , n93108 );
or ( n93110 , n93094 , n93109 );
buf ( n93111 , n40998 );
buf ( n93112 , n41051 );
or ( n93113 , n93111 , n93112 );
buf ( n93114 , n93113 );
nand ( n93115 , n93110 , n93114 );
buf ( n93116 , n93115 );
not ( n93117 , n93116 );
or ( n93118 , n93093 , n93117 );
buf ( n93119 , n41250 );
buf ( n93120 , n41256 );
or ( n93121 , n93119 , n93120 );
buf ( n93122 , n93121 );
buf ( n93123 , n93122 );
nand ( n93124 , n93118 , n93123 );
buf ( n93125 , n93124 );
buf ( n93126 , n93125 );
not ( n93127 , n93126 );
buf ( n93128 , n93127 );
nand ( n93129 , n93091 , n93128 );
not ( n93130 , n93129 );
or ( n93131 , n93054 , n93130 );
buf ( n93132 , n41544 );
not ( n93133 , n93132 );
nand ( n93134 , n41434 , n41341 );
or ( n93135 , n93134 , n41486 );
buf ( n93136 , n41477 );
buf ( n93137 , n41483 );
nand ( n93138 , n93136 , n93137 );
buf ( n93139 , n93138 );
nand ( n93140 , n93135 , n93139 );
buf ( n93141 , n93140 );
not ( n93142 , n93141 );
or ( n93143 , n93133 , n93142 );
buf ( n93144 , n41541 );
not ( n93145 , n93144 );
buf ( n93146 , n41497 );
nand ( n93147 , n93145 , n93146 );
buf ( n93148 , n93147 );
buf ( n93149 , n93148 );
nand ( n93150 , n93143 , n93149 );
buf ( n93151 , n93150 );
and ( n93152 , n93151 , n41558 );
buf ( n93153 , n41548 );
not ( n93154 , n93153 );
buf ( n93155 , n41555 );
nor ( n93156 , n93154 , n93155 );
buf ( n93157 , n93156 );
nor ( n93158 , n93152 , n93157 );
nand ( n93159 , n93131 , n93158 );
not ( n93160 , n93159 );
nand ( n93161 , n93053 , n93160 );
not ( n93162 , n93161 );
or ( n93163 , n37244 , n93162 );
not ( n93164 , n37242 );
and ( n93165 , n93164 , n37221 );
not ( n93166 , n93165 );
nand ( n93167 , n93163 , n93166 );
buf ( n93168 , n93167 );
and ( n93169 , n93168 , n36842 );
not ( n93170 , n93168 );
and ( n93171 , n93170 , n36838 );
nor ( n93172 , n93169 , n93171 );
buf ( n93173 , n93172 );
buf ( n93174 , n93157 );
not ( n93175 , n93174 );
buf ( n93176 , n41558 );
nand ( n93177 , n93175 , n93176 );
buf ( n93178 , n93177 );
buf ( n93179 , n93178 );
buf ( n93180 , n93178 );
not ( n93181 , n93180 );
buf ( n93182 , n93181 );
buf ( n93183 , n93182 );
buf ( n93184 , n41544 );
not ( n93185 , n93184 );
not ( n93186 , n41325 );
nor ( n93187 , n93186 , n41492 );
not ( n93188 , n93187 );
not ( n93189 , n93051 );
or ( n93190 , n93188 , n93189 );
not ( n93191 , n41492 );
nand ( n93192 , n93191 , n93129 );
nand ( n93193 , n93190 , n93192 );
buf ( n93194 , n93193 );
not ( n93195 , n93194 );
or ( n93196 , n93185 , n93195 );
buf ( n93197 , n93151 );
not ( n93198 , n93197 );
buf ( n93199 , n93198 );
buf ( n93200 , n93199 );
nand ( n93201 , n93196 , n93200 );
buf ( n93202 , n93201 );
buf ( n93203 , n93202 );
and ( n93204 , n93203 , n93183 );
not ( n93205 , n93203 );
and ( n93206 , n93205 , n93179 );
nor ( n93207 , n93204 , n93206 );
buf ( n93208 , n93207 );
buf ( n93209 , n93139 );
buf ( n93210 , n41489 );
nand ( n93211 , n93209 , n93210 );
buf ( n93212 , n93211 );
buf ( n93213 , n93212 );
buf ( n93214 , n93212 );
not ( n93215 , n93214 );
buf ( n93216 , n93215 );
buf ( n93217 , n93216 );
not ( n93218 , n41437 );
not ( n93219 , n41325 );
nand ( n93220 , n92808 , n93050 , n92928 );
not ( n93221 , n93220 );
or ( n93222 , n93219 , n93221 );
not ( n93223 , n93129 );
nand ( n93224 , n93222 , n93223 );
not ( n93225 , n93224 );
or ( n93226 , n93218 , n93225 );
buf ( n93227 , n93134 );
nand ( n93228 , n93226 , n93227 );
buf ( n93229 , n93228 );
and ( n93230 , n93229 , n93217 );
not ( n93231 , n93229 );
and ( n93232 , n93231 , n93213 );
nor ( n93233 , n93230 , n93232 );
buf ( n93234 , n93233 );
not ( n93235 , n41301 );
nand ( n93236 , n93235 , n93105 );
buf ( n93237 , n93236 );
buf ( n93238 , n93236 );
not ( n93239 , n93238 );
buf ( n93240 , n93239 );
buf ( n93241 , n93240 );
buf ( n93242 , n41318 );
not ( n93243 , n93242 );
not ( n93244 , n40498 );
not ( n93245 , n93220 );
or ( n93246 , n93244 , n93245 );
buf ( n93247 , n93089 );
not ( n93248 , n93247 );
buf ( n93249 , n93248 );
nand ( n93250 , n93246 , n93249 );
buf ( n93251 , n93250 );
not ( n93252 , n93251 );
or ( n93253 , n93243 , n93252 );
buf ( n93254 , n93099 );
buf ( n93255 , n93254 );
buf ( n93256 , n93255 );
buf ( n93257 , n93256 );
nand ( n93258 , n93253 , n93257 );
buf ( n93259 , n93258 );
buf ( n93260 , n93259 );
and ( n93261 , n93260 , n93241 );
not ( n93262 , n93260 );
and ( n93263 , n93262 , n93237 );
nor ( n93264 , n93261 , n93263 );
buf ( n93265 , n93264 );
buf ( n93266 , n41544 );
buf ( n93267 , n93148 );
nand ( n93268 , n93266 , n93267 );
buf ( n93269 , n93268 );
buf ( n93270 , n93269 );
not ( n93271 , n93270 );
buf ( n93272 , n93271 );
buf ( n93273 , n93272 );
buf ( n93274 , n93269 );
buf ( n93275 , n93193 );
buf ( n93276 , n93140 );
nor ( n93277 , n93275 , n93276 );
buf ( n93278 , n93277 );
buf ( n93279 , n93278 );
and ( n93280 , n93279 , n93274 );
not ( n93281 , n93279 );
and ( n93282 , n93281 , n93273 );
nor ( n93283 , n93280 , n93282 );
buf ( n93284 , n93283 );
buf ( n93285 , n41052 );
buf ( n93286 , n93114 );
nand ( n93287 , n93285 , n93286 );
buf ( n93288 , n93287 );
buf ( n93289 , n93288 );
not ( n93290 , n93289 );
buf ( n93291 , n93290 );
buf ( n93292 , n93291 );
buf ( n93293 , n93288 );
not ( n93294 , n40498 );
nor ( n93295 , n93294 , n41319 );
not ( n93296 , n93295 );
not ( n93297 , n93220 );
or ( n93298 , n93296 , n93297 );
not ( n93299 , n41319 );
nand ( n93300 , n93299 , n93089 );
nand ( n93301 , n93298 , n93300 );
buf ( n93302 , n93108 );
nor ( n93303 , n93301 , n93302 );
buf ( n93304 , n93303 );
and ( n93305 , n93304 , n93293 );
not ( n93306 , n93304 );
and ( n93307 , n93306 , n93292 );
nor ( n93308 , n93305 , n93307 );
buf ( n93309 , n93308 );
not ( n93310 , n92843 );
buf ( n93311 , n92724 );
nand ( n93312 , n93310 , n93311 );
buf ( n93313 , n93312 );
not ( n93314 , n93313 );
buf ( n93315 , n93314 );
buf ( n93316 , n93315 );
buf ( n93317 , n93312 );
nor ( n93318 , n89856 , n90831 , n90812 );
not ( n93319 , n93318 );
not ( n93320 , n92458 );
buf ( n93321 , n88818 );
buf ( n93322 , n93321 );
buf ( n93323 , n93322 );
nand ( n93324 , n93320 , n93323 );
nor ( n93325 , n93319 , n93324 );
not ( n93326 , n93325 );
nand ( n93327 , n92989 , n93036 , n93046 );
and ( n93328 , n86690 , n92983 , n93327 );
not ( n93329 , n93328 );
not ( n93330 , n93329 );
or ( n93331 , n93326 , n93330 );
and ( n93332 , n92827 , n92809 );
nor ( n93333 , n93332 , n92851 );
nand ( n93334 , n93333 , n92908 );
not ( n93335 , n92164 );
nor ( n93336 , n93335 , n91696 );
and ( n93337 , n93336 , n92457 );
and ( n93338 , n93334 , n93337 );
buf ( n93339 , n92914 );
nor ( n93340 , n93338 , n93339 );
nand ( n93341 , n93331 , n93340 );
and ( n93342 , n92774 , n92765 );
and ( n93343 , n93341 , n93342 );
buf ( n93344 , n92765 );
not ( n93345 , n93344 );
nor ( n93346 , n92768 , n92773 );
buf ( n93347 , n93346 );
not ( n93348 , n93347 );
or ( n93349 , n93345 , n93348 );
buf ( n93350 , n92840 );
nand ( n93351 , n93349 , n93350 );
buf ( n93352 , n93351 );
nor ( n93353 , n93343 , n93352 );
buf ( n93354 , n93353 );
and ( n93355 , n93354 , n93317 );
not ( n93356 , n93354 );
and ( n93357 , n93356 , n93316 );
nor ( n93358 , n93355 , n93357 );
buf ( n93359 , n93358 );
nand ( n93360 , n93068 , n40202 );
buf ( n93361 , n93360 );
buf ( n93362 , n93360 );
not ( n93363 , n93362 );
buf ( n93364 , n93363 );
buf ( n93365 , n93364 );
buf ( n93366 , n40186 );
not ( n93367 , n93366 );
buf ( n93368 , n93051 );
buf ( n93369 , n93368 );
not ( n93370 , n93369 );
or ( n93371 , n93367 , n93370 );
buf ( n93372 , n93063 );
buf ( n93373 , n93372 );
nand ( n93374 , n93371 , n93373 );
buf ( n93375 , n93374 );
buf ( n93376 , n93375 );
and ( n93377 , n93376 , n93365 );
not ( n93378 , n93376 );
and ( n93379 , n93378 , n93361 );
nor ( n93380 , n93377 , n93379 );
buf ( n93381 , n93380 );
nand ( n93382 , n41437 , n93227 );
buf ( n93383 , n93382 );
buf ( n93384 , n93382 );
not ( n93385 , n93384 );
buf ( n93386 , n93385 );
buf ( n93387 , n93386 );
buf ( n93388 , n93224 );
and ( n93389 , n93388 , n93387 );
not ( n93390 , n93388 );
and ( n93391 , n93390 , n93383 );
nor ( n93392 , n93389 , n93391 );
buf ( n93393 , n93392 );
buf ( n93394 , n93256 );
buf ( n93395 , n41318 );
nand ( n93396 , n93394 , n93395 );
buf ( n93397 , n93396 );
buf ( n93398 , n93397 );
buf ( n93399 , n93397 );
not ( n93400 , n93399 );
buf ( n93401 , n93400 );
buf ( n93402 , n93401 );
buf ( n93403 , n93250 );
and ( n93404 , n93403 , n93402 );
not ( n93405 , n93403 );
and ( n93406 , n93405 , n93398 );
nor ( n93407 , n93404 , n93406 );
buf ( n93408 , n93407 );
buf ( n93409 , n93086 );
buf ( n93410 , n40495 );
nand ( n93411 , n93409 , n93410 );
buf ( n93412 , n93411 );
buf ( n93413 , n93412 );
buf ( n93414 , n93412 );
not ( n93415 , n93414 );
buf ( n93416 , n93415 );
buf ( n93417 , n93416 );
buf ( n93418 , n40206 );
not ( n93419 , n93418 );
buf ( n93420 , n93368 );
not ( n93421 , n93420 );
or ( n93422 , n93419 , n93421 );
buf ( n93423 , n93079 );
not ( n93424 , n93423 );
buf ( n93425 , n93424 );
buf ( n93426 , n93425 );
nand ( n93427 , n93422 , n93426 );
buf ( n93428 , n93427 );
buf ( n93429 , n93428 );
and ( n93430 , n93429 , n93417 );
not ( n93431 , n93429 );
and ( n93432 , n93431 , n93413 );
nor ( n93433 , n93430 , n93432 );
buf ( n93434 , n93433 );
buf ( n93435 , n93076 );
buf ( n93436 , n39463 );
nand ( n93437 , n93435 , n93436 );
buf ( n93438 , n93437 );
buf ( n93439 , n93438 );
buf ( n93440 , n93438 );
not ( n93441 , n93440 );
buf ( n93442 , n93441 );
buf ( n93443 , n93442 );
buf ( n93444 , n40203 );
not ( n93445 , n93444 );
buf ( n93446 , n93445 );
buf ( n93447 , n93446 );
not ( n93448 , n93447 );
buf ( n93449 , n93368 );
not ( n93450 , n93449 );
or ( n93451 , n93448 , n93450 );
buf ( n93452 , n93069 );
buf ( n93453 , n93452 );
not ( n93454 , n93453 );
buf ( n93455 , n93454 );
buf ( n93456 , n93455 );
nand ( n93457 , n93451 , n93456 );
buf ( n93458 , n93457 );
buf ( n93459 , n93458 );
and ( n93460 , n93459 , n93443 );
not ( n93461 , n93459 );
and ( n93462 , n93461 , n93439 );
nor ( n93463 , n93460 , n93462 );
buf ( n93464 , n93463 );
not ( n93465 , n92846 );
nand ( n93466 , n93465 , n92800 );
buf ( n93467 , n93466 );
buf ( n93468 , n93466 );
not ( n93469 , n93468 );
buf ( n93470 , n93469 );
buf ( n93471 , n93470 );
buf ( n93472 , n92775 );
not ( n93473 , n93472 );
buf ( n93474 , n93473 );
buf ( n93475 , n93474 );
not ( n93476 , n93475 );
buf ( n93477 , n93341 );
not ( n93478 , n93477 );
or ( n93479 , n93476 , n93478 );
not ( n93480 , n93311 );
not ( n93481 , n92841 );
or ( n93482 , n93480 , n93481 );
nand ( n93483 , n93482 , n93310 );
buf ( n93484 , n93483 );
not ( n93485 , n93484 );
buf ( n93486 , n93485 );
buf ( n93487 , n93486 );
nand ( n93488 , n93479 , n93487 );
buf ( n93489 , n93488 );
buf ( n93490 , n93489 );
and ( n93491 , n93490 , n93471 );
not ( n93492 , n93490 );
and ( n93493 , n93492 , n93467 );
nor ( n93494 , n93491 , n93493 );
buf ( n93495 , n93494 );
buf ( n93496 , n92840 );
buf ( n93497 , n92765 );
nand ( n93498 , n93496 , n93497 );
buf ( n93499 , n93498 );
buf ( n93500 , n93499 );
buf ( n93501 , n93499 );
not ( n93502 , n93501 );
buf ( n93503 , n93502 );
buf ( n93504 , n93503 );
buf ( n93505 , n92774 );
not ( n93506 , n93505 );
buf ( n93507 , n93341 );
not ( n93508 , n93507 );
or ( n93509 , n93506 , n93508 );
buf ( n93510 , n93346 );
not ( n93511 , n93510 );
buf ( n93512 , n93511 );
buf ( n93513 , n93512 );
nand ( n93514 , n93509 , n93513 );
buf ( n93515 , n93514 );
buf ( n93516 , n93515 );
and ( n93517 , n93516 , n93504 );
not ( n93518 , n93516 );
and ( n93519 , n93518 , n93500 );
nor ( n93520 , n93517 , n93519 );
buf ( n93521 , n93520 );
buf ( n93522 , n93512 );
buf ( n93523 , n92774 );
nand ( n93524 , n93522 , n93523 );
buf ( n93525 , n93524 );
buf ( n93526 , n93525 );
buf ( n93527 , n93525 );
not ( n93528 , n93527 );
buf ( n93529 , n93528 );
buf ( n93530 , n93529 );
buf ( n93531 , n92461 );
not ( n93532 , n93531 );
and ( n93533 , n93318 , n93323 );
not ( n93534 , n93533 );
not ( n93535 , n93329 );
or ( n93536 , n93534 , n93535 );
not ( n93537 , n93334 );
nand ( n93538 , n93536 , n93537 );
buf ( n93539 , n93538 );
not ( n93540 , n93539 );
or ( n93541 , n93532 , n93540 );
not ( n93542 , n93339 );
buf ( n93543 , n93542 );
nand ( n93544 , n93541 , n93543 );
buf ( n93545 , n93544 );
buf ( n93546 , n93545 );
and ( n93547 , n93546 , n93530 );
not ( n93548 , n93546 );
and ( n93549 , n93548 , n93526 );
nor ( n93550 , n93547 , n93549 );
buf ( n93551 , n93550 );
buf ( n93552 , n92883 );
buf ( n93553 , n92457 );
nand ( n93554 , n93552 , n93553 );
buf ( n93555 , n93554 );
buf ( n93556 , n93555 );
buf ( n93557 , n93555 );
not ( n93558 , n93557 );
buf ( n93559 , n93558 );
buf ( n93560 , n93559 );
buf ( n93561 , n93336 );
not ( n93562 , n93561 );
buf ( n93563 , n93538 );
not ( n93564 , n93563 );
or ( n93565 , n93562 , n93564 );
buf ( n93566 , n92879 );
not ( n93567 , n93566 );
buf ( n93568 , n93567 );
buf ( n93569 , n93568 );
nand ( n93570 , n93565 , n93569 );
buf ( n93571 , n93570 );
buf ( n93572 , n93571 );
and ( n93573 , n93572 , n93560 );
not ( n93574 , n93572 );
and ( n93575 , n93574 , n93556 );
nor ( n93576 , n93573 , n93575 );
buf ( n93577 , n93576 );
nand ( n93578 , n92809 , n92850 );
buf ( n93579 , n93578 );
buf ( n93580 , n93578 );
not ( n93581 , n93580 );
buf ( n93582 , n93581 );
buf ( n93583 , n93582 );
nor ( n93584 , n89856 , n90831 );
not ( n93585 , n93584 );
not ( n93586 , n93323 );
not ( n93587 , n93329 );
or ( n93588 , n93586 , n93587 );
buf ( n93589 , n92907 );
buf ( n93590 , n93589 );
not ( n93591 , n93590 );
buf ( n93592 , n93591 );
nand ( n93593 , n93588 , n93592 );
not ( n93594 , n93593 );
or ( n93595 , n93585 , n93594 );
buf ( n93596 , n92827 );
not ( n93597 , n93596 );
buf ( n93598 , n93597 );
nand ( n93599 , n93595 , n93598 );
buf ( n93600 , n93599 );
and ( n93601 , n93600 , n93583 );
not ( n93602 , n93600 );
and ( n93603 , n93602 , n93579 );
nor ( n93604 , n93601 , n93603 );
buf ( n93605 , n93604 );
buf ( n93606 , n90830 );
buf ( n93607 , n92826 );
nand ( n93608 , n93606 , n93607 );
buf ( n93609 , n93608 );
buf ( n93610 , n93609 );
buf ( n93611 , n93609 );
not ( n93612 , n93611 );
buf ( n93613 , n93612 );
buf ( n93614 , n93613 );
not ( n93615 , n89856 );
not ( n93616 , n93615 );
not ( n93617 , n93593 );
or ( n93618 , n93616 , n93617 );
buf ( n93619 , n92821 );
not ( n93620 , n93619 );
nand ( n93621 , n93618 , n93620 );
buf ( n93622 , n93621 );
and ( n93623 , n93622 , n93614 );
not ( n93624 , n93622 );
and ( n93625 , n93624 , n93610 );
nor ( n93626 , n93623 , n93625 );
buf ( n93627 , n93626 );
buf ( n93628 , n92820 );
buf ( n93629 , n93628 );
buf ( n93630 , n89846 );
nand ( n93631 , n93629 , n93630 );
buf ( n93632 , n93631 );
buf ( n93633 , n93632 );
buf ( n93634 , n93632 );
not ( n93635 , n93634 );
buf ( n93636 , n93635 );
buf ( n93637 , n93636 );
buf ( n93638 , n89855 );
not ( n93639 , n93638 );
buf ( n93640 , n93593 );
not ( n93641 , n93640 );
or ( n93642 , n93639 , n93641 );
buf ( n93643 , n92815 );
buf ( n93644 , n93643 );
buf ( n93645 , n93644 );
buf ( n93646 , n93645 );
nand ( n93647 , n93642 , n93646 );
buf ( n93648 , n93647 );
buf ( n93649 , n93648 );
and ( n93650 , n93649 , n93637 );
not ( n93651 , n93649 );
and ( n93652 , n93651 , n93633 );
nor ( n93653 , n93650 , n93652 );
buf ( n93654 , n93653 );
buf ( n93655 , n92980 );
not ( n93656 , n93655 );
buf ( n93657 , n92973 );
nand ( n93658 , n93656 , n93657 );
buf ( n93659 , n93658 );
buf ( n93660 , n93659 );
buf ( n93661 , n93659 );
not ( n93662 , n93661 );
buf ( n93663 , n93662 );
buf ( n93664 , n93663 );
buf ( n93665 , n47224 );
buf ( n93666 , n48102 );
buf ( n93667 , n93666 );
buf ( n93668 , n49129 );
buf ( n93669 , n93668 );
and ( n93670 , n93665 , n93667 , n93669 );
buf ( n93671 , n93670 );
not ( n93672 , n93671 );
buf ( n93673 , n53445 );
buf ( n93674 , n93673 );
buf ( n93675 , n93674 );
buf ( n93676 , n93675 );
not ( n93677 , n93676 );
buf ( n93678 , n86689 );
buf ( n93679 , n63523 );
buf ( n93680 , n59133 );
nand ( n93681 , n93678 , n93679 , n93680 );
buf ( n93682 , n93034 );
buf ( n93683 , n93682 );
buf ( n93684 , n93683 );
buf ( n93685 , n57042 );
and ( n93686 , n93684 , n93685 );
buf ( n93687 , n93021 );
nor ( n93688 , n93686 , n93687 );
buf ( n93689 , n63522 );
not ( n93690 , n93689 );
nand ( n93691 , n93006 , n93000 );
buf ( n93692 , n93691 );
not ( n93693 , n93692 );
or ( n93694 , n93690 , n93693 );
buf ( n93695 , n93004 );
buf ( n93696 , n93695 );
nand ( n93697 , n93694 , n93696 );
buf ( n93698 , n93697 );
nand ( n93699 , n93680 , n93698 );
nand ( n93700 , n93681 , n93688 , n93699 );
buf ( n93701 , n93700 );
not ( n93702 , n93701 );
or ( n93703 , n93677 , n93702 );
buf ( n93704 , n92952 );
buf ( n93705 , n93704 );
buf ( n93706 , n93705 );
buf ( n93707 , n93706 );
not ( n93708 , n93707 );
buf ( n93709 , n93708 );
buf ( n93710 , n93709 );
nand ( n93711 , n93703 , n93710 );
buf ( n93712 , n93711 );
not ( n93713 , n93712 );
or ( n93714 , n93672 , n93713 );
nand ( n93715 , n92969 , n92970 );
nand ( n93716 , n93714 , n93715 );
buf ( n93717 , n93716 );
and ( n93718 , n93717 , n93664 );
not ( n93719 , n93717 );
and ( n93720 , n93719 , n93660 );
nor ( n93721 , n93718 , n93720 );
buf ( n93722 , n93721 );
buf ( n93723 , n92958 );
not ( n93724 , n93723 );
buf ( n93725 , n47224 );
buf ( n93726 , n93725 );
nand ( n93727 , n93724 , n93726 );
buf ( n93728 , n93727 );
buf ( n93729 , n93728 );
buf ( n93730 , n93728 );
not ( n93731 , n93730 );
buf ( n93732 , n93731 );
buf ( n93733 , n93732 );
not ( n93734 , n93666 );
buf ( n93735 , n93675 );
not ( n93736 , n93735 );
buf ( n93737 , n93668 );
not ( n93738 , n93737 );
buf ( n93739 , n93738 );
buf ( n93740 , n93739 );
nor ( n93741 , n93736 , n93740 );
buf ( n93742 , n93741 );
buf ( n93743 , n93742 );
not ( n93744 , n93743 );
nand ( n93745 , n93681 , n93699 );
buf ( n93746 , n93745 );
not ( n93747 , n93746 );
or ( n93748 , n93744 , n93747 );
buf ( n93749 , n93709 );
not ( n93750 , n93749 );
buf ( n93751 , n93739 );
not ( n93752 , n93751 );
and ( n93753 , n93750 , n93752 );
buf ( n93754 , n93688 );
not ( n93755 , n93754 );
buf ( n93756 , n93755 );
buf ( n93757 , n93756 );
buf ( n93758 , n93742 );
and ( n93759 , n93757 , n93758 );
nor ( n93760 , n93753 , n93759 );
buf ( n93761 , n93760 );
buf ( n93762 , n93761 );
nand ( n93763 , n93748 , n93762 );
buf ( n93764 , n93763 );
not ( n93765 , n93764 );
or ( n93766 , n93734 , n93765 );
not ( n93767 , n92968 );
buf ( n93768 , n92963 );
buf ( n93769 , n93768 );
nor ( n93770 , n93767 , n93769 );
nand ( n93771 , n93766 , n93770 );
buf ( n93772 , n93771 );
and ( n93773 , n93772 , n93733 );
not ( n93774 , n93772 );
and ( n93775 , n93774 , n93729 );
nor ( n93776 , n93773 , n93775 );
buf ( n93777 , n93776 );
buf ( n93778 , n93768 );
not ( n93779 , n93778 );
buf ( n93780 , n93666 );
nand ( n93781 , n93779 , n93780 );
buf ( n93782 , n93781 );
buf ( n93783 , n93782 );
not ( n93784 , n93783 );
buf ( n93785 , n93784 );
buf ( n93786 , n93785 );
buf ( n93787 , n93782 );
nor ( n93788 , n49128 , n48105 );
nor ( n93789 , n93764 , n93788 );
buf ( n93790 , n93789 );
and ( n93791 , n93790 , n93787 );
not ( n93792 , n93790 );
and ( n93793 , n93792 , n93786 );
nor ( n93794 , n93791 , n93793 );
buf ( n93795 , n93794 );
buf ( n93796 , n92891 );
not ( n93797 , n92894 );
buf ( n93798 , n93797 );
nand ( n93799 , n93796 , n93798 );
buf ( n93800 , n93799 );
buf ( n93801 , n93800 );
buf ( n93802 , n93800 );
not ( n93803 , n93802 );
buf ( n93804 , n93803 );
buf ( n93805 , n93804 );
buf ( n93806 , n87252 );
not ( n93807 , n93806 );
buf ( n93808 , n93329 );
not ( n93809 , n93808 );
or ( n93810 , n93807 , n93809 );
buf ( n93811 , n92892 );
buf ( n93812 , n93811 );
nand ( n93813 , n93810 , n93812 );
buf ( n93814 , n93813 );
buf ( n93815 , n93814 );
and ( n93816 , n93815 , n93805 );
not ( n93817 , n93815 );
and ( n93818 , n93817 , n93801 );
nor ( n93819 , n93816 , n93818 );
buf ( n93820 , n93819 );
buf ( n93821 , n93024 );
buf ( n93822 , n93033 );
nand ( n93823 , n93821 , n93822 );
buf ( n93824 , n93823 );
buf ( n93825 , n93823 );
not ( n93826 , n93825 );
buf ( n93827 , n93826 );
buf ( n93828 , n93827 );
nand ( n93829 , n67885 , n67890 );
not ( n93830 , n93829 );
nand ( n93831 , n63476 , n63522 , n63505 );
nor ( n93832 , n93830 , n93831 );
not ( n93833 , n93832 );
not ( n93834 , n67879 );
not ( n93835 , n67869 );
or ( n93836 , n93834 , n93835 );
nand ( n93837 , n86684 , n86677 );
nand ( n93838 , n93836 , n93837 );
not ( n93839 , n93838 );
or ( n93840 , n93833 , n93839 );
not ( n93841 , n86688 );
not ( n93842 , n93831 );
and ( n93843 , n93841 , n93842 );
nor ( n93844 , n93843 , n93698 );
nand ( n93845 , n93840 , n93844 );
buf ( n93846 , n93845 );
not ( n93847 , n93846 );
buf ( n93848 , n93847 );
buf ( n93849 , n93848 );
buf ( n93850 , n59125 );
not ( n93851 , n93850 );
buf ( n93852 , n93851 );
or ( n93853 , n93849 , n93852 );
buf ( n93854 , n93022 );
not ( n93855 , n93854 );
buf ( n93856 , n93855 );
buf ( n93857 , n93856 );
nand ( n93858 , n93853 , n93857 );
buf ( n93859 , n93858 );
buf ( n93860 , n93859 );
and ( n93861 , n93860 , n93828 );
not ( n93862 , n93860 );
and ( n93863 , n93862 , n93824 );
nor ( n93864 , n93861 , n93863 );
buf ( n93865 , n93864 );
buf ( n93866 , n57029 );
nand ( n93867 , n93012 , n93016 );
buf ( n93868 , n93867 );
nand ( n93869 , n93866 , n93868 );
buf ( n93870 , n93869 );
buf ( n93871 , n93870 );
buf ( n93872 , n93870 );
not ( n93873 , n93872 );
buf ( n93874 , n93873 );
buf ( n93875 , n93874 );
not ( n93876 , n59127 );
not ( n93877 , n93845 );
or ( n93878 , n93876 , n93877 );
buf ( n93879 , n93684 );
not ( n93880 , n93879 );
buf ( n93881 , n93880 );
nand ( n93882 , n93878 , n93881 );
buf ( n93883 , n93882 );
and ( n93884 , n93883 , n93875 );
not ( n93885 , n93883 );
and ( n93886 , n93885 , n93871 );
nor ( n93887 , n93884 , n93886 );
buf ( n93888 , n93887 );
nand ( n93889 , n92949 , n92945 );
buf ( n93890 , n93889 );
buf ( n93891 , n93889 );
not ( n93892 , n93891 );
buf ( n93893 , n93892 );
buf ( n93894 , n93893 );
buf ( n93895 , n53391 );
buf ( n93896 , n93895 );
buf ( n93897 , n93896 );
buf ( n93898 , n93897 );
buf ( n93899 , n53432 );
buf ( n93900 , n93899 );
and ( n93901 , n93898 , n93900 );
buf ( n93902 , n93901 );
buf ( n93903 , n93902 );
not ( n93904 , n93903 );
buf ( n93905 , n93745 );
not ( n93906 , n93905 );
or ( n93907 , n93904 , n93906 );
and ( n93908 , n93902 , n93756 );
not ( n93909 , n93899 );
buf ( n93910 , n92931 );
buf ( n93911 , n93910 );
nand ( n93912 , n92935 , n92933 );
buf ( n93913 , n93912 );
nand ( n93914 , n93911 , n93913 );
buf ( n93915 , n93914 );
not ( n93916 , n93915 );
or ( n93917 , n93909 , n93916 );
nand ( n93918 , n93917 , n92942 );
nor ( n93919 , n93908 , n93918 );
buf ( n93920 , n93919 );
nand ( n93921 , n93907 , n93920 );
buf ( n93922 , n93921 );
buf ( n93923 , n93922 );
and ( n93924 , n93923 , n93894 );
not ( n93925 , n93923 );
and ( n93926 , n93925 , n93890 );
nor ( n93927 , n93924 , n93926 );
buf ( n93928 , n93927 );
buf ( n93929 , n52859 );
nand ( n93930 , n93912 , n93929 );
buf ( n93931 , n93930 );
buf ( n93932 , n93930 );
not ( n93933 , n93932 );
buf ( n93934 , n93933 );
buf ( n93935 , n93934 );
buf ( n93936 , n53389 );
buf ( n93937 , n93936 );
buf ( n93938 , n93937 );
not ( n93939 , n93938 );
buf ( n93940 , n93700 );
not ( n93941 , n93940 );
or ( n93942 , n93939 , n93941 );
buf ( n93943 , n92930 );
buf ( n93944 , n93943 );
not ( n93945 , n93944 );
nand ( n93946 , n93942 , n93945 );
buf ( n93947 , n93946 );
and ( n93948 , n93947 , n93935 );
not ( n93949 , n93947 );
and ( n93950 , n93949 , n93931 );
nor ( n93951 , n93948 , n93950 );
buf ( n93952 , n93951 );
buf ( n93953 , n40186 );
buf ( n93954 , n93372 );
and ( n93955 , n93953 , n93954 );
buf ( n93956 , n93955 );
buf ( n93957 , n93956 );
buf ( n93958 , n93368 );
not ( n93959 , n93958 );
buf ( n93960 , n93959 );
buf ( n93961 , n93960 );
buf ( n93962 , n93956 );
buf ( n93963 , n93960 );
not ( n93964 , n93957 );
not ( n93965 , n93961 );
or ( n93966 , n93964 , n93965 );
or ( n93967 , n93962 , n93963 );
nand ( n93968 , n93966 , n93967 );
buf ( n93969 , n93968 );
buf ( n93970 , n91279 );
buf ( n93971 , n93970 );
not ( n93972 , n92859 );
buf ( n93973 , n93972 );
nand ( n93974 , n93971 , n93973 );
buf ( n93975 , n93974 );
buf ( n93976 , n93975 );
buf ( n93977 , n93538 );
buf ( n93978 , n93977 );
buf ( n93979 , n93975 );
buf ( n93980 , n93977 );
not ( n93981 , n93976 );
not ( n93982 , n93978 );
or ( n93983 , n93981 , n93982 );
or ( n93984 , n93979 , n93980 );
nand ( n93985 , n93983 , n93984 );
buf ( n93986 , n93985 );
buf ( n93987 , n93645 );
buf ( n93988 , n89855 );
nand ( n93989 , n93987 , n93988 );
buf ( n93990 , n93989 );
buf ( n93991 , n93990 );
buf ( n93992 , n93990 );
not ( n93993 , n93992 );
buf ( n93994 , n93993 );
buf ( n93995 , n93994 );
buf ( n93996 , n93593 );
and ( n93997 , n93996 , n93995 );
not ( n93998 , n93996 );
and ( n93999 , n93998 , n93991 );
nor ( n94000 , n93997 , n93999 );
buf ( n94001 , n94000 );
buf ( n94002 , n92942 );
buf ( n94003 , n93899 );
nand ( n94004 , n94002 , n94003 );
buf ( n94005 , n94004 );
buf ( n94006 , n94005 );
buf ( n94007 , n94005 );
not ( n94008 , n94007 );
buf ( n94009 , n94008 );
buf ( n94010 , n94009 );
buf ( n94011 , n93897 );
not ( n94012 , n94011 );
buf ( n94013 , n93940 );
not ( n94014 , n94013 );
or ( n94015 , n94012 , n94014 );
buf ( n94016 , n93915 );
not ( n94017 , n94016 );
buf ( n94018 , n94017 );
buf ( n94019 , n94018 );
nand ( n94020 , n94015 , n94019 );
buf ( n94021 , n94020 );
buf ( n94022 , n94021 );
and ( n94023 , n94022 , n94010 );
not ( n94024 , n94022 );
and ( n94025 , n94024 , n94006 );
nor ( n94026 , n94023 , n94025 );
buf ( n94027 , n94026 );
not ( n94028 , n93788 );
nand ( n94029 , n94028 , n93668 );
buf ( n94030 , n94029 );
buf ( n94031 , n94029 );
not ( n94032 , n94031 );
buf ( n94033 , n94032 );
buf ( n94034 , n94033 );
buf ( n94035 , n93712 );
and ( n94036 , n94035 , n94034 );
not ( n94037 , n94035 );
and ( n94038 , n94037 , n94030 );
nor ( n94039 , n94036 , n94038 );
buf ( n94040 , n94039 );
buf ( n94041 , n66130 );
buf ( n94042 , n67876 );
nand ( n94043 , n94041 , n94042 );
buf ( n94044 , n94043 );
buf ( n94045 , n94044 );
buf ( n94046 , n94044 );
not ( n94047 , n94046 );
buf ( n94048 , n94047 );
buf ( n94049 , n94048 );
buf ( n94050 , n67867 );
not ( n94051 , n86681 );
and ( n94052 , n94050 , n94051 );
buf ( n94053 , n67871 );
not ( n94054 , n71014 );
not ( n94055 , n86653 );
or ( n94056 , n94054 , n94055 );
nand ( n94057 , n94056 , n86676 );
nand ( n94058 , n94052 , n94053 , n94057 );
not ( n94059 , n67866 );
not ( n94060 , n94050 );
or ( n94061 , n94059 , n94060 );
buf ( n94062 , n66005 );
nand ( n94063 , n94062 , n65910 );
nand ( n94064 , n94061 , n94063 );
and ( n94065 , n94064 , n94053 );
nand ( n94066 , n66088 , n66093 );
not ( n94067 , n94066 );
nor ( n94068 , n94065 , n94067 );
nand ( n94069 , n94058 , n94068 );
buf ( n94070 , n94069 );
and ( n94071 , n94070 , n94049 );
not ( n94072 , n94070 );
and ( n94073 , n94072 , n94045 );
nor ( n94074 , n94071 , n94073 );
buf ( n94075 , n94074 );
buf ( n94076 , n93856 );
buf ( n94077 , n93850 );
nand ( n94078 , n94076 , n94077 );
buf ( n94079 , n94078 );
buf ( n94080 , n94079 );
not ( n94081 , n94080 );
buf ( n94082 , n94081 );
buf ( n94083 , n94082 );
buf ( n94084 , n94079 );
buf ( n94085 , n93848 );
and ( n94086 , n94085 , n94084 );
not ( n94087 , n94085 );
and ( n94088 , n94087 , n94083 );
nor ( n94089 , n94086 , n94088 );
buf ( n94090 , n94089 );
not ( n94091 , n93944 );
nand ( n94092 , n94091 , n93938 );
buf ( n94093 , n94092 );
buf ( n94094 , n93940 );
buf ( n94095 , n94092 );
buf ( n94096 , n93940 );
not ( n94097 , n94093 );
not ( n94098 , n94094 );
or ( n94099 , n94097 , n94098 );
or ( n94100 , n94095 , n94096 );
nand ( n94101 , n94099 , n94100 );
buf ( n94102 , n94101 );
buf ( n94103 , n63505 );
not ( n94104 , n94103 );
buf ( n94105 , n94104 );
not ( n94106 , n94105 );
nand ( n94107 , n94106 , n93006 );
buf ( n94108 , n94107 );
buf ( n94109 , n94107 );
not ( n94110 , n94109 );
buf ( n94111 , n94110 );
buf ( n94112 , n94111 );
buf ( n94113 , n63476 );
not ( n94114 , n94113 );
buf ( n94115 , n93678 );
not ( n94116 , n94115 );
or ( n94117 , n94114 , n94116 );
nand ( n94118 , n62047 , n61209 );
buf ( n94119 , n94118 );
buf ( n94120 , n92999 );
nand ( n94121 , n94119 , n94120 );
buf ( n94122 , n94121 );
nand ( n94123 , n94117 , n94122 );
buf ( n94124 , n94123 );
and ( n94125 , n94124 , n94112 );
not ( n94126 , n94124 );
and ( n94127 , n94126 , n94108 );
nor ( n94128 , n94125 , n94127 );
buf ( n94129 , n94128 );
buf ( n94130 , n93695 );
buf ( n94131 , n92990 );
nand ( n94132 , n94130 , n94131 );
buf ( n94133 , n94132 );
buf ( n94134 , n94133 );
buf ( n94135 , n94133 );
not ( n94136 , n94135 );
buf ( n94137 , n94136 );
buf ( n94138 , n94137 );
buf ( n94139 , n94113 );
not ( n94140 , n94139 );
buf ( n94141 , n94105 );
nor ( n94142 , n94140 , n94141 );
buf ( n94143 , n94142 );
not ( n94144 , n94143 );
not ( n94145 , n94115 );
or ( n94146 , n94144 , n94145 );
buf ( n94147 , n93691 );
not ( n94148 , n94147 );
buf ( n94149 , n94148 );
nand ( n94150 , n94146 , n94149 );
buf ( n94151 , n94150 );
and ( n94152 , n94151 , n94138 );
not ( n94153 , n94151 );
and ( n94154 , n94153 , n94134 );
nor ( n94155 , n94152 , n94154 );
buf ( n94156 , n94155 );
buf ( n94157 , n93329 );
buf ( n94158 , n94157 );
buf ( n94159 , n94158 );
buf ( n94160 , n86675 );
not ( n94161 , n94160 );
buf ( n94162 , n67907 );
buf ( n94163 , n94162 );
buf ( n94164 , n69269 );
nand ( n94165 , n94163 , n94164 );
buf ( n94166 , n94165 );
buf ( n94167 , n94166 );
nand ( n94168 , n94161 , n94167 );
buf ( n94169 , n94168 );
buf ( n94170 , n94169 );
buf ( n94171 , n94169 );
not ( n94172 , n94171 );
buf ( n94173 , n94172 );
buf ( n94174 , n94173 );
buf ( n94175 , n71011 );
buf ( n94176 , n86337 );
buf ( n94177 , n94176 );
buf ( n94178 , n86355 );
buf ( n94179 , n86360 );
nand ( n94180 , n94177 , n94178 , n94179 );
buf ( n94181 , n94180 );
buf ( n94182 , n94181 );
buf ( n94183 , n86521 );
buf ( n94184 , n86608 );
nand ( n94185 , n94182 , n94183 , n94184 );
buf ( n94186 , n94185 );
buf ( n94187 , n94186 );
buf ( n94188 , n86650 );
buf ( n94189 , n94188 );
buf ( n94190 , n94189 );
nand ( n94191 , n94187 , n94190 );
buf ( n94192 , n94191 );
buf ( n94193 , n94192 );
nand ( n94194 , n94175 , n94193 );
buf ( n94195 , n94194 );
buf ( n94196 , n69350 );
buf ( n94197 , n94196 );
buf ( n94198 , n94197 );
buf ( n94199 , n94198 );
not ( n94200 , n94199 );
buf ( n94201 , n94200 );
or ( n94202 , n94195 , n94201 );
not ( n94203 , n86673 );
nand ( n94204 , n94202 , n94203 );
buf ( n94205 , n94204 );
and ( n94206 , n94205 , n94174 );
not ( n94207 , n94205 );
and ( n94208 , n94207 , n94170 );
nor ( n94209 , n94206 , n94208 );
buf ( n94210 , n94209 );
buf ( n94211 , n86672 );
buf ( n94212 , n94198 );
nand ( n94213 , n94211 , n94212 );
buf ( n94214 , n94213 );
buf ( n94215 , n94214 );
buf ( n94216 , n94214 );
not ( n94217 , n94216 );
buf ( n94218 , n94217 );
buf ( n94219 , n94218 );
buf ( n94220 , n94195 );
buf ( n94221 , n86660 );
buf ( n94222 , n94221 );
not ( n94223 , n94222 );
buf ( n94224 , n94223 );
buf ( n94225 , n94224 );
nand ( n94226 , n94220 , n94225 );
buf ( n94227 , n94226 );
buf ( n94228 , n94227 );
and ( n94229 , n94228 , n94219 );
not ( n94230 , n94228 );
and ( n94231 , n94230 , n94215 );
nor ( n94232 , n94229 , n94231 );
buf ( n94233 , n94232 );
buf ( n94234 , n86649 );
buf ( n94235 , n86637 );
nand ( n94236 , n94234 , n94235 );
buf ( n94237 , n94236 );
buf ( n94238 , n94237 );
buf ( n94239 , n94237 );
not ( n94240 , n94239 );
buf ( n94241 , n94240 );
buf ( n94242 , n94241 );
buf ( n94243 , n86494 );
not ( n94244 , n94243 );
buf ( n94245 , n86631 );
not ( n94246 , n94245 );
buf ( n94247 , n86608 );
buf ( n94248 , n94176 );
buf ( n94249 , n86355 );
buf ( n94250 , n86360 );
nand ( n94251 , n94248 , n94249 , n94250 );
buf ( n94252 , n94251 );
buf ( n94253 , n94252 );
nand ( n94254 , n94247 , n94253 );
buf ( n94255 , n94254 );
buf ( n94256 , n94255 );
nand ( n94257 , n94246 , n94256 );
buf ( n94258 , n94257 );
buf ( n94259 , n94258 );
not ( n94260 , n94259 );
or ( n94261 , n94244 , n94260 );
buf ( n94262 , n86424 );
buf ( n94263 , n86488 );
nand ( n94264 , n94262 , n94263 );
buf ( n94265 , n94264 );
buf ( n94266 , n94265 );
nand ( n94267 , n94261 , n94266 );
buf ( n94268 , n94267 );
buf ( n94269 , n94268 );
and ( n94270 , n94269 , n94242 );
not ( n94271 , n94269 );
and ( n94272 , n94271 , n94238 );
nor ( n94273 , n94270 , n94272 );
buf ( n94274 , n94273 );
buf ( n94275 , n94265 );
buf ( n94276 , n86494 );
nand ( n94277 , n94275 , n94276 );
buf ( n94278 , n94277 );
buf ( n94279 , n94278 );
buf ( n94280 , n94278 );
not ( n94281 , n94280 );
buf ( n94282 , n94281 );
buf ( n94283 , n94282 );
buf ( n94284 , n94258 );
and ( n94285 , n94284 , n94283 );
not ( n94286 , n94284 );
and ( n94287 , n94286 , n94279 );
nor ( n94288 , n94285 , n94287 );
buf ( n94289 , n94288 );
buf ( n94290 , n86630 );
buf ( n94291 , n86605 );
nand ( n94292 , n94290 , n94291 );
buf ( n94293 , n94292 );
buf ( n94294 , n94293 );
buf ( n94295 , n94293 );
not ( n94296 , n94295 );
buf ( n94297 , n94296 );
buf ( n94298 , n94297 );
buf ( n94299 , n86581 );
not ( n94300 , n94299 );
buf ( n94301 , n94252 );
not ( n94302 , n94301 );
or ( n94303 , n94300 , n94302 );
buf ( n94304 , n86618 );
not ( n94305 , n94304 );
buf ( n94306 , n94305 );
buf ( n94307 , n94306 );
nand ( n94308 , n94303 , n94307 );
buf ( n94309 , n94308 );
buf ( n94310 , n94309 );
and ( n94311 , n94310 , n94298 );
not ( n94312 , n94310 );
and ( n94313 , n94312 , n94294 );
nor ( n94314 , n94311 , n94313 );
buf ( n94315 , n94314 );
buf ( n94316 , n86350 );
buf ( n94317 , n86312 );
nand ( n94318 , n94316 , n94317 );
buf ( n94319 , n94318 );
buf ( n94320 , n94319 );
buf ( n94321 , n94319 );
not ( n94322 , n94321 );
buf ( n94323 , n94322 );
buf ( n94324 , n94323 );
not ( n94325 , n86331 );
buf ( n94326 , n94325 );
not ( n94327 , n94326 );
not ( n94328 , n84435 );
not ( n94329 , n85673 );
or ( n94330 , n94328 , n94329 );
nand ( n94331 , n94330 , n85696 );
buf ( n94332 , n94331 );
not ( n94333 , n94332 );
or ( n94334 , n94327 , n94333 );
buf ( n94335 , n86343 );
not ( n94336 , n94335 );
buf ( n94337 , n94336 );
buf ( n94338 , n94337 );
nand ( n94339 , n94334 , n94338 );
buf ( n94340 , n94339 );
buf ( n94341 , n94340 );
and ( n94342 , n94341 , n94324 );
not ( n94343 , n94341 );
and ( n94344 , n94343 , n94320 );
nor ( n94345 , n94342 , n94344 );
buf ( n94346 , n94345 );
buf ( n94347 , n85684 );
buf ( n94348 , n85363 );
nand ( n94349 , n94347 , n94348 );
buf ( n94350 , n94349 );
buf ( n94351 , n94350 );
buf ( n94352 , n94350 );
not ( n94353 , n94352 );
buf ( n94354 , n94353 );
buf ( n94355 , n94354 );
buf ( n94356 , n85380 );
not ( n94357 , n94356 );
buf ( n94358 , n94357 );
not ( n94359 , n94358 );
buf ( n94360 , n84435 );
buf ( n94361 , n94360 );
buf ( n94362 , n94361 );
not ( n94363 , n94362 );
or ( n94364 , n94359 , n94363 );
not ( n94365 , n85678 );
nand ( n94366 , n94364 , n94365 );
buf ( n94367 , n94366 );
and ( n94368 , n94367 , n94355 );
not ( n94369 , n94367 );
and ( n94370 , n94369 , n94351 );
nor ( n94371 , n94368 , n94370 );
buf ( n94372 , n94371 );
buf ( n94373 , n94362 );
buf ( n94374 , n85363 );
buf ( n94375 , n94358 );
buf ( n94376 , n85685 );
and ( n94377 , n94373 , n94374 , n94375 );
nor ( n94378 , n94377 , n94376 );
buf ( n94379 , n94378 );
buf ( n94380 , n84340 );
buf ( n94381 , n80146 );
nand ( n94382 , n94380 , n94381 );
buf ( n94383 , n94382 );
buf ( n94384 , n94383 );
buf ( n94385 , n94383 );
not ( n94386 , n94385 );
buf ( n94387 , n94386 );
buf ( n94388 , n94387 );
buf ( n94389 , n79236 );
buf ( n94390 , n94389 );
buf ( n94391 , n94390 );
buf ( n94392 , n94391 );
not ( n94393 , n94392 );
buf ( n94394 , n80057 );
not ( n94395 , n94394 );
buf ( n94396 , n80150 );
not ( n94397 , n94396 );
buf ( n94398 , n94397 );
buf ( n94399 , n94398 );
not ( n94400 , n94399 );
buf ( n94401 , n84338 );
not ( n94402 , n94401 );
or ( n94403 , n94400 , n94402 );
buf ( n94404 , n80051 );
nand ( n94405 , n94403 , n94404 );
buf ( n94406 , n94405 );
buf ( n94407 , n94406 );
not ( n94408 , n94407 );
or ( n94409 , n94395 , n94408 );
buf ( n94410 , n79324 );
nand ( n94411 , n94409 , n94410 );
buf ( n94412 , n94411 );
buf ( n94413 , n94412 );
not ( n94414 , n94413 );
or ( n94415 , n94393 , n94414 );
buf ( n94416 , n80075 );
nand ( n94417 , n94415 , n94416 );
buf ( n94418 , n94417 );
buf ( n94419 , n94418 );
and ( n94420 , n94419 , n94388 );
not ( n94421 , n94419 );
and ( n94422 , n94421 , n94384 );
nor ( n94423 , n94420 , n94422 );
buf ( n94424 , n94423 );
buf ( n94425 , n80075 );
buf ( n94426 , n94391 );
nand ( n94427 , n94425 , n94426 );
buf ( n94428 , n94427 );
buf ( n94429 , n94428 );
buf ( n94430 , n94428 );
not ( n94431 , n94430 );
buf ( n94432 , n94431 );
buf ( n94433 , n94432 );
buf ( n94434 , n94412 );
and ( n94435 , n94434 , n94433 );
not ( n94436 , n94434 );
and ( n94437 , n94436 , n94429 );
nor ( n94438 , n94435 , n94437 );
buf ( n94439 , n94438 );
buf ( n94440 , n84390 );
buf ( n94441 , n84420 );
not ( n94442 , n94441 );
buf ( n94443 , n94442 );
buf ( n94444 , n94443 );
nand ( n94445 , n94440 , n94444 );
buf ( n94446 , n94445 );
buf ( n94447 , n79324 );
buf ( n94448 , n80057 );
nand ( n94449 , n94447 , n94448 );
buf ( n94450 , n94449 );
buf ( n94451 , n94450 );
buf ( n94452 , n94450 );
not ( n94453 , n94452 );
buf ( n94454 , n94453 );
buf ( n94455 , n94454 );
buf ( n94456 , n94406 );
and ( n94457 , n94456 , n94455 );
not ( n94458 , n94456 );
and ( n94459 , n94458 , n94451 );
nor ( n94460 , n94457 , n94459 );
buf ( n94461 , n94460 );
xor ( n94462 , n81116 , n81120 );
xor ( n94463 , n94462 , n84324 );
buf ( n94464 , n94463 );
buf ( n94465 , n85670 );
buf ( n94466 , n85692 );
nand ( n94467 , n94465 , n94466 );
buf ( n94468 , n94467 );
buf ( n94469 , n94337 );
buf ( n94470 , n94325 );
nand ( n94471 , n94469 , n94470 );
buf ( n94472 , n94471 );
buf ( n94473 , n94472 );
not ( n94474 , n94473 );
buf ( n94475 , n94474 );
xor ( n94476 , n81434 , n81438 );
xor ( n94477 , n94476 , n84319 );
buf ( n94478 , n94477 );
buf ( n94479 , n94306 );
buf ( n94480 , n86581 );
nand ( n94481 , n94479 , n94480 );
buf ( n94482 , n94481 );
buf ( n94483 , n94482 );
not ( n94484 , n94483 );
buf ( n94485 , n94484 );
buf ( n94486 , n94224 );
buf ( n94487 , n71011 );
nand ( n94488 , n94486 , n94487 );
buf ( n94489 , n94488 );
xor ( n94490 , n81557 , n81561 );
xor ( n94491 , n94490 , n84314 );
buf ( n94492 , n94491 );
buf ( n94493 , n94050 );
buf ( n94494 , n94063 );
nand ( n94495 , n94493 , n94494 );
buf ( n94496 , n94495 );
buf ( n94497 , n94496 );
not ( n94498 , n94497 );
buf ( n94499 , n94498 );
nand ( n94500 , n94066 , n94053 );
buf ( n94501 , n94500 );
not ( n94502 , n94501 );
buf ( n94503 , n94502 );
buf ( n94504 , n94398 );
buf ( n94505 , n80051 );
nand ( n94506 , n94504 , n94505 );
buf ( n94507 , n94506 );
xor ( n94508 , n81986 , n81990 );
xor ( n94509 , n94508 , n84309 );
buf ( n94510 , n94509 );
not ( n94511 , n93830 );
nand ( n94512 , n94511 , n86688 );
buf ( n94513 , n94512 );
not ( n94514 , n94513 );
buf ( n94515 , n94514 );
buf ( n94516 , n82434 );
buf ( n94517 , n84307 );
nand ( n94518 , n94516 , n94517 );
buf ( n94519 , n94518 );
buf ( n94520 , n84292 );
buf ( n94521 , n82594 );
not ( n94522 , n94520 );
nor ( n94523 , n94522 , n94521 );
buf ( n94524 , n94523 );
buf ( n94525 , n84260 );
buf ( n94526 , n84253 );
nand ( n94527 , n94525 , n94526 );
buf ( n94528 , n94527 );
buf ( n94529 , n94528 );
buf ( n94530 , n84200 );
buf ( n94531 , n84200 );
buf ( n94532 , n94528 );
not ( n94533 , n94529 );
not ( n94534 , n94530 );
or ( n94535 , n94533 , n94534 );
or ( n94536 , n94531 , n94532 );
nand ( n94537 , n94535 , n94536 );
buf ( n94538 , n94537 );
buf ( n94539 , n83180 );
buf ( n94540 , n84199 );
nand ( n94541 , n94539 , n94540 );
buf ( n94542 , n94541 );
buf ( n94543 , n84168 );
buf ( n94544 , n84171 );
buf ( n94545 , n84183 );
not ( n94546 , n94545 );
buf ( n94547 , n84189 );
nand ( n94548 , n94546 , n94547 );
buf ( n94549 , n94548 );
buf ( n94550 , n94549 );
and ( n94551 , n94550 , n94544 );
not ( n94552 , n94550 );
and ( n94553 , n94552 , n94543 );
nor ( n94554 , n94551 , n94553 );
buf ( n94555 , n94554 );
xor ( n94556 , n83475 , n84149 );
xor ( n94557 , n94556 , n84164 );
buf ( n94558 , n94557 );
buf ( n94559 , n84135 );
buf ( n94560 , n84147 );
nand ( n94561 , n94559 , n94560 );
buf ( n94562 , n94561 );
buf ( n94563 , n94562 );
buf ( n94564 , n84096 );
buf ( n94565 , n84096 );
buf ( n94566 , n94562 );
not ( n94567 , n94563 );
not ( n94568 , n94564 );
or ( n94569 , n94567 , n94568 );
or ( n94570 , n94565 , n94566 );
nand ( n94571 , n94569 , n94570 );
buf ( n94572 , n94571 );
buf ( n94573 , n93811 );
buf ( n94574 , n87252 );
and ( n94575 , n94573 , n94574 );
buf ( n94576 , n94575 );
buf ( n94577 , n83771 );
buf ( n94578 , n84048 );
nand ( n94579 , n94577 , n94578 );
buf ( n94580 , n94579 );
buf ( n94581 , n94580 );
buf ( n94582 , n84043 );
buf ( n94583 , n84043 );
buf ( n94584 , n94580 );
not ( n94585 , n94581 );
not ( n94586 , n94582 );
or ( n94587 , n94585 , n94586 );
or ( n94588 , n94583 , n94584 );
nand ( n94589 , n94587 , n94588 );
buf ( n94590 , n94589 );
buf ( n94591 , n88815 );
not ( n94592 , n94591 );
buf ( n94593 , n92901 );
nand ( n94594 , n94592 , n94593 );
buf ( n94595 , n94594 );
buf ( n94596 , n94595 );
not ( n94597 , n94596 );
buf ( n94598 , n94597 );
buf ( n94599 , n84042 );
buf ( n94600 , n84036 );
nand ( n94601 , n94599 , n94600 );
buf ( n94602 , n94601 );
buf ( n94603 , n94602 );
buf ( n94604 , n84015 );
buf ( n94605 , n84015 );
buf ( n94606 , n94602 );
not ( n94607 , n94603 );
not ( n94608 , n94604 );
or ( n94609 , n94607 , n94608 );
or ( n94610 , n94605 , n94606 );
nand ( n94611 , n94609 , n94610 );
buf ( n94612 , n94611 );
xor ( n94613 , n83960 , n84004 );
xor ( n94614 , n94613 , n84012 );
buf ( n94615 , n94614 );
xor ( n94616 , C0 , n84002 );
buf ( n94617 , n94616 );
xor ( n94618 , C0 , n83998 );
buf ( n94619 , n94618 );
buf ( n94620 , n83993 );
not ( n94621 , n94620 );
buf ( n94622 , n83994 );
nand ( n94623 , n94621 , n94622 );
buf ( n94624 , n94623 );
buf ( n94625 , n83985 );
buf ( n94626 , n94624 );
or ( n94627 , n94625 , n94626 );
nand ( n94628 , C1 , n94627 );
buf ( n94629 , n94628 );
xor ( n94630 , n83964 , n83982 );
xor ( n94631 , n94630 , n83984 );
buf ( n94632 , n94631 );
buf ( n94633 , n37243 );
buf ( n94634 , n93166 );
nand ( n94635 , n94633 , n94634 );
buf ( n94636 , n94635 );
buf ( n94637 , n94636 );
not ( n94638 , n94637 );
buf ( n94639 , n94638 );
xor ( n94640 , n83968 , n83978 );
xor ( n94641 , n94640 , n83980 );
buf ( n94642 , n94641 );
xor ( n94643 , n36713 , n36733 );
and ( n94644 , n94643 , n36791 );
and ( n94645 , n36713 , n36733 );
or ( n94646 , n94644 , n94645 );
buf ( n94647 , n94646 );
buf ( n94648 , n36712 );
not ( n94649 , n94648 );
buf ( n94650 , n36688 );
buf ( n94651 , n36706 );
nand ( n94652 , n94650 , n94651 );
buf ( n94653 , n94652 );
buf ( n94654 , n94653 );
not ( n94655 , n94654 );
buf ( n94656 , n36702 );
nor ( n94657 , n94655 , n94656 );
buf ( n94658 , n94657 );
buf ( n94659 , n36363 );
buf ( n94660 , n36044 );
and ( n94661 , n94659 , n94660 );
not ( n94662 , n94659 );
buf ( n94663 , n36057 );
and ( n94664 , n94662 , n94663 );
nor ( n94665 , n94661 , n94664 );
buf ( n94666 , n94665 );
buf ( n94667 , n94666 );
not ( n94668 , n94667 );
buf ( n94669 , n36456 );
nand ( n94670 , n94668 , n94669 );
buf ( n94671 , n94670 );
buf ( n94672 , n94671 );
nand ( n94673 , C1 , n94672 );
buf ( n94674 , n94673 );
buf ( n94675 , n94674 );
buf ( n94676 , n94658 );
or ( n94677 , n94675 , n94676 );
nand ( n94678 , C1 , n94677 );
buf ( n94679 , n94678 );
buf ( n94680 , n94679 );
not ( n94681 , n94680 );
or ( n94682 , n94649 , n94681 );
buf ( n94683 , n94679 );
buf ( n94684 , n36712 );
or ( n94685 , n94683 , n94684 );
nand ( n94686 , n94682 , n94685 );
buf ( n94687 , n94686 );
buf ( n94688 , C0 );
buf ( n94689 , C1 );
xor ( n94690 , n83970 , n83974 );
xor ( n94691 , n94690 , n83976 );
buf ( n94692 , n94691 );
buf ( n94693 , n83870 );
buf ( n94694 , n83882 );
xor ( n94695 , n94693 , n94694 );
buf ( n94696 , n94695 );
buf ( n94697 , n94647 );
buf ( n94698 , n94687 );
and ( n94699 , n94697 , n94698 );
buf ( n94700 , n94699 );
buf ( n94701 , n94576 );
buf ( n94702 , n94159 );
xor ( n94703 , n94701 , n94702 );
buf ( n94704 , n94703 );
buf ( n94705 , n94362 );
nand ( n94706 , n94358 , n94365 );
buf ( n94707 , n94706 );
xnor ( n94708 , n94705 , n94707 );
buf ( n94709 , n94708 );
buf ( n94710 , n94446 );
buf ( n94711 , n84415 );
buf ( n94712 , n84424 );
or ( n94713 , n94711 , n94712 );
buf ( n94714 , n94713 );
buf ( n94715 , n94714 );
xnor ( n94716 , n94710 , n94715 );
buf ( n94717 , n94716 );
buf ( n94718 , n94379 );
buf ( n94719 , n94468 );
xor ( n94720 , n94718 , n94719 );
buf ( n94721 , n94720 );
buf ( n94722 , n84388 );
buf ( n94723 , n94443 );
not ( n94724 , n94722 );
nand ( n94725 , n94724 , n94723 );
buf ( n94726 , n94725 );
buf ( n94727 , n82503 );
buf ( n94728 , n84299 );
not ( n94729 , n94727 );
nand ( n94730 , n94729 , n94728 );
buf ( n94731 , n94730 );
buf ( n94732 , n92998 );
buf ( n94733 , n94732 );
buf ( n94734 , n63473 );
nand ( n94735 , n94733 , n94734 );
buf ( n94736 , n94735 );
nand ( n94737 , n67865 , n94051 );
xnor ( n94738 , n94057 , n94737 );
buf ( n94739 , n94192 );
buf ( n94740 , n94489 );
xnor ( n94741 , n94739 , n94740 );
buf ( n94742 , n94741 );
buf ( n94743 , n84300 );
buf ( n94744 , n94519 );
xnor ( n94745 , n94743 , n94744 );
buf ( n94746 , n94745 );
buf ( n94747 , n92807 );
buf ( n94748 , n93329 );
buf ( n94749 , n92928 );
buf ( n94750 , n94749 );
not ( n94751 , n94747 );
not ( n94752 , n94748 );
or ( n94753 , n94751 , n94752 );
nand ( n94754 , n94753 , n94750 );
buf ( n94755 , n94754 );
buf ( n94756 , n84192 );
buf ( n94757 , n94542 );
buf ( n94758 , n84171 );
buf ( n94759 , n84183 );
or ( n94760 , n94758 , n94759 );
buf ( n94761 , n84189 );
nand ( n94762 , n94760 , n94761 );
buf ( n94763 , n94762 );
buf ( n94764 , n94763 );
buf ( n94765 , n94542 );
not ( n94766 , n94756 );
not ( n94767 , n94757 );
or ( n94768 , n94766 , n94767 );
or ( n94769 , n94764 , n94765 );
nand ( n94770 , n94768 , n94769 );
buf ( n94771 , n94770 );
nand ( n94772 , n93160 , n94639 );
or ( n94773 , n94755 , n94772 );
not ( n94774 , n41566 );
nor ( n94775 , n94774 , n94639 );
nand ( n94776 , n94775 , n94755 );
nor ( n94777 , n94772 , n41566 );
and ( n94778 , n93159 , n94636 );
nor ( n94779 , n94777 , n94778 );
nand ( n94780 , n94773 , n94776 , n94779 );
not ( n94781 , n87779 );
not ( n94782 , n93329 );
or ( n94783 , n94781 , n94782 );
nand ( n94784 , n92893 , n93797 );
nand ( n94785 , n94783 , n94784 );
not ( n94786 , n94785 );
not ( n94787 , n92903 );
nor ( n94788 , n94595 , n94787 );
nand ( n94789 , n94786 , n94788 );
not ( n94790 , n88310 );
not ( n94791 , n94790 );
nor ( n94792 , n94791 , n94598 );
nand ( n94793 , n94785 , n94792 );
not ( n94794 , n94598 );
not ( n94795 , n92903 );
and ( n94796 , n94794 , n94795 );
nor ( n94797 , n94595 , n94790 , n94787 );
nor ( n94798 , n94796 , n94797 );
nand ( n94799 , n94789 , n94793 , n94798 );
and ( n94800 , n93838 , n94515 );
not ( n94801 , n93838 );
and ( n94802 , n94801 , n94512 );
nor ( n94803 , n94800 , n94802 );
nand ( n94804 , n94118 , n92997 );
not ( n94805 , n94804 );
not ( n94806 , n63473 );
not ( n94807 , n94115 );
or ( n94808 , n94806 , n94807 );
nand ( n94809 , n94808 , n94732 );
not ( n94810 , n94809 );
or ( n94811 , n94805 , n94810 );
or ( n94812 , n94804 , n94809 );
nand ( n94813 , n94811 , n94812 );
nand ( n94814 , n92808 , n93050 , n92928 );
not ( n94815 , n36827 );
nand ( n94816 , n94815 , n37243 );
nor ( n94817 , n94816 , n94688 );
not ( n94818 , n94817 );
not ( n94819 , n94818 );
nand ( n94820 , n94819 , C1 );
nor ( n94821 , n41563 , n94820 );
nand ( n94822 , n94814 , n94821 );
not ( n94823 , n94815 );
not ( n94824 , n93165 );
or ( n94825 , n94823 , n94824 );
nand ( n94826 , n94825 , n36834 );
and ( n94827 , n94826 , n94689 );
nor ( n94828 , n94827 , n94700 );
and ( n94829 , n94828 , C1 );
not ( n94830 , n94829 );
not ( n94831 , n93160 );
or ( n94832 , n94830 , n94831 );
nand ( n94833 , n94832 , C1 );
nand ( n94834 , n94822 , n94833 );
and ( n94835 , n94834 , C1 );
not ( n94836 , n94834 );
and ( n94837 , n94836 , C0 );
nor ( n94838 , n94835 , n94837 );
not ( n94839 , n93115 );
nand ( n94840 , n93122 , n41259 );
not ( n94841 , n94840 );
nor ( n94842 , n41563 , n94818 );
not ( n94843 , n94842 );
not ( n94844 , n93368 );
or ( n94845 , n94843 , n94844 );
not ( n94846 , n94828 );
and ( n94847 , n93159 , n94817 );
nor ( n94848 , n94846 , n94847 );
nand ( n94849 , n94845 , n94848 );
and ( n94850 , n94849 , C1 );
not ( n94851 , n94849 );
and ( n94852 , n94851 , C0 );
nor ( n94853 , n94850 , n94852 );
not ( n94854 , n93970 );
not ( n94855 , n93538 );
or ( n94856 , n94854 , n94855 );
buf ( n94857 , n93972 );
nand ( n94858 , n94856 , n94857 );
buf ( n94859 , n91695 );
nand ( n94860 , n92868 , n94859 );
not ( n94861 , n94860 );
and ( n94862 , n94858 , n94861 );
not ( n94863 , n94858 );
and ( n94864 , n94863 , n94860 );
nor ( n94865 , n94862 , n94864 );
not ( n94866 , n91696 );
not ( n94867 , n94866 );
not ( n94868 , n93538 );
or ( n94869 , n94867 , n94868 );
not ( n94870 , n92869 );
nand ( n94871 , n94869 , n94870 );
buf ( n94872 , n92876 );
nand ( n94873 , n94872 , n92164 );
not ( n94874 , n94873 );
and ( n94875 , n94871 , n94874 );
not ( n94876 , n94871 );
and ( n94877 , n94876 , n94873 );
nor ( n94878 , n94875 , n94877 );
buf ( n94879 , n84333 );
or ( n94880 , n80732 , n80717 );
or ( n94881 , n94879 , n94880 );
nand ( n94882 , n80717 , n80732 );
or ( n94883 , n94882 , n94879 );
not ( n94884 , n84337 );
not ( n94885 , n80733 );
or ( n94886 , n94884 , n94885 );
nand ( n94887 , n94886 , n94879 );
nand ( n94888 , n94881 , n94883 , n94887 );
not ( n94889 , n57029 );
not ( n94890 , n93882 );
or ( n94891 , n94889 , n94890 );
nand ( n94892 , n94891 , n93867 );
not ( n94893 , n93043 );
nand ( n94894 , n94893 , n93020 );
not ( n94895 , n94894 );
and ( n94896 , n94892 , n94895 );
not ( n94897 , n94892 );
and ( n94898 , n94897 , n94894 );
nor ( n94899 , n94896 , n94898 );
nand ( n94900 , n94822 , n94833 , C1 );
nand ( n94901 , n94900 , C1 );
buf ( n94902 , n94901 );
and ( n94903 , n94057 , n94052 );
nor ( n94904 , n94903 , n94064 );
and ( n94905 , n94904 , n94500 );
not ( n94906 , n94904 );
and ( n94907 , n94906 , n94503 );
nor ( n94908 , n94905 , n94907 );
not ( n94909 , n94051 );
not ( n94910 , n94057 );
or ( n94911 , n94909 , n94910 );
nand ( n94912 , n94911 , n67865 );
and ( n94913 , n94912 , n94499 );
not ( n94914 , n94912 );
and ( n94915 , n94914 , n94496 );
nor ( n94916 , n94913 , n94915 );
not ( n94917 , n84284 );
and ( n94918 , n94731 , n84294 );
not ( n94919 , n94731 );
and ( n94920 , n94919 , n84293 );
nor ( n94921 , n94918 , n94920 );
not ( n94922 , n84287 );
not ( n94923 , n94524 );
or ( n94924 , n94922 , n94923 );
or ( n94925 , n94524 , n84287 );
nand ( n94926 , n94924 , n94925 );
not ( n94927 , n41052 );
nor ( n94928 , n94927 , n94841 );
not ( n94929 , n94839 );
nor ( n94930 , n94840 , n94929 , n41052 );
not ( n94931 , n94726 );
buf ( n94932 , n84341 );
not ( n94933 , n94932 );
or ( n94934 , n94931 , n94933 );
or ( n94935 , n94932 , n94726 );
nand ( n94936 , n94934 , n94935 );
not ( n94937 , n94736 );
not ( n94938 , n94115 );
or ( n94939 , n94937 , n94938 );
or ( n94940 , n94736 , n94115 );
nand ( n94941 , n94939 , n94940 );
buf ( n94942 , n94482 );
buf ( n94943 , n94485 );
buf ( n94944 , n94252 );
and ( n94945 , n94944 , n94943 );
not ( n94946 , n94944 );
and ( n94947 , n94946 , n94942 );
nor ( n94948 , n94945 , n94947 );
buf ( n94949 , n94948 );
xor ( n94950 , n76413 , n76905 );
xor ( n94951 , n94950 , n84431 );
buf ( n94952 , n94951 );
buf ( n94953 , n94472 );
buf ( n94954 , n94475 );
buf ( n94955 , n94331 );
and ( n94956 , n94955 , n94954 );
not ( n94957 , n94955 );
and ( n94958 , n94957 , n94953 );
nor ( n94959 , n94956 , n94958 );
buf ( n94960 , n94959 );
and ( n94961 , n84278 , n84283 );
not ( n94962 , n84278 );
and ( n94963 , n94962 , n84282 );
nor ( n94964 , n94961 , n94963 );
not ( n94965 , n94840 );
nand ( n94966 , n94965 , n94839 );
or ( n94967 , n94966 , n93301 );
nand ( n94968 , n93301 , n94928 );
not ( n94969 , n94841 );
not ( n94970 , n94839 );
and ( n94971 , n94969 , n94970 );
nor ( n94972 , n94971 , n94930 );
nand ( n94973 , n94967 , n94968 , n94972 );
buf ( n94974 , n86268 );
buf ( n94975 , n86360 );
nand ( n94976 , n94974 , n94975 );
buf ( n94977 , n94976 );
buf ( n94978 , n94977 );
buf ( n94979 , n94977 );
not ( n94980 , n94979 );
buf ( n94981 , n94980 );
buf ( n94982 , n94981 );
and ( n94983 , n94331 , n94325 , n86312 );
nor ( n94984 , n94983 , n86351 );
not ( n94985 , n94984 );
buf ( n94986 , n94985 );
and ( n94987 , n94986 , n94982 );
not ( n94988 , n94986 );
and ( n94989 , n94988 , n94978 );
nor ( n94990 , n94987 , n94989 );
buf ( n94991 , n94990 );
nand ( n94992 , n94790 , n92903 );
not ( n94993 , n94992 );
and ( n94994 , n94785 , n94993 );
not ( n94995 , n94785 );
and ( n94996 , n94995 , n94992 );
nor ( n94997 , n94994 , n94996 );
xor ( n94998 , n80953 , n80956 );
xor ( n94999 , n94998 , n84329 );
buf ( n95000 , n94999 );
buf ( n95001 , n84338 );
buf ( n95002 , n94507 );
xnor ( n95003 , n95001 , n95002 );
buf ( n95004 , n95003 );
nand ( n95005 , n84093 , n84087 );
not ( n95006 , n95005 );
nand ( n95007 , n84051 , n83771 );
not ( n95008 , n95007 );
or ( n95009 , n95006 , n95008 );
or ( n95010 , n95007 , n95005 );
nand ( n95011 , n95009 , n95010 );
not ( n95012 , n29666 );
xnor ( n95013 , n29538 , n26042 );
not ( n95014 , n95013 );
or ( n95015 , n95012 , n95014 );
or ( n95016 , n95013 , n29666 );
nand ( n95017 , n95015 , n95016 );
xor ( n95018 , n29570 , n29571 );
xor ( n95019 , n95018 , n29573 );
buf ( n95020 , n95019 );
not ( n95021 , n94917 );
not ( n95022 , n84261 );
or ( n95023 , n95021 , n95022 );
not ( n95024 , n84261 );
not ( n95025 , n94964 );
and ( n95026 , n95024 , n95025 );
and ( n95027 , n84261 , n84286 );
nor ( n95028 , n95026 , n95027 );
nand ( n95029 , n95023 , n95028 );
xor ( n95030 , n29366 , n29838 );
xor ( n95031 , n95030 , n29842 );
buf ( n95032 , n95031 );
xor ( n95033 , n29384 , n29388 );
xor ( n95034 , n95033 , n29833 );
buf ( n95035 , n95034 );
xor ( n95036 , n25866 , n25530 );
xor ( n95037 , n24718 , n24698 );
xor ( n95038 , n95037 , n25491 );
not ( n95039 , n94816 );
not ( n95040 , n95039 );
not ( n95041 , n93161 );
or ( n95042 , n95040 , n95041 );
not ( n95043 , n94826 );
nand ( n95044 , n95042 , n95043 );
nor ( n95045 , n94700 , n94688 );
and ( n95046 , n95044 , n95045 );
not ( n95047 , n95044 );
not ( n95048 , n95045 );
and ( n95049 , n95047 , n95048 );
nor ( n95050 , n95046 , n95049 );
xor ( n95051 , n25862 , n25527 );
xor ( n95052 , n24693 , n24670 );
not ( n95053 , n25487 );
xor ( n95054 , n95052 , n95053 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
