module mul_21_11_21(a, b, c);
  input [20:0] a;
  input [10:0] b;
  output [20:0] c;
  assign c = a * b;
endmodule
