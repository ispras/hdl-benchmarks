module OptKuznechikEncoder(
  input wire clk,
  input wire [127:0] _block,
  input wire [255:0] key,
  output wire [127:0] out
);
  wire [7:0] arr[256] = '{8'hfc, 8'hee, 8'hdd, 8'h11, 8'hcf, 8'h6e, 8'h31, 8'h16, 8'hfb, 8'hc4, 8'hfa, 8'hda, 8'h23, 8'hc5, 8'h04, 8'h4d, 8'he9, 8'h77, 8'hf0, 8'hdb, 8'h93, 8'h2e, 8'h99, 8'hba, 8'h17, 8'h36, 8'hf1, 8'hbb, 8'h14, 8'hcd, 8'h5f, 8'hc1, 8'hf9, 8'h18, 8'h65, 8'h5a, 8'he2, 8'h5c, 8'hef, 8'h21, 8'h81, 8'h1c, 8'h3c, 8'h42, 8'h8b, 8'h01, 8'h8e, 8'h4f, 8'h05, 8'h84, 8'h02, 8'hae, 8'he3, 8'h6a, 8'h8f, 8'ha0, 8'h06, 8'h0b, 8'hed, 8'h98, 8'h7f, 8'hd4, 8'hd3, 8'h1f, 8'heb, 8'h34, 8'h2c, 8'h51, 8'hea, 8'hc8, 8'h48, 8'hab, 8'hf2, 8'h2a, 8'h68, 8'ha2, 8'hfd, 8'h3a, 8'hce, 8'hcc, 8'hb5, 8'h70, 8'h0e, 8'h56, 8'h08, 8'h0c, 8'h76, 8'h12, 8'hbf, 8'h72, 8'h13, 8'h47, 8'h9c, 8'hb7, 8'h5d, 8'h87, 8'h15, 8'ha1, 8'h96, 8'h29, 8'h10, 8'h7b, 8'h9a, 8'hc7, 8'hf3, 8'h91, 8'h78, 8'h6f, 8'h9d, 8'h9e, 8'hb2, 8'hb1, 8'h32, 8'h75, 8'h19, 8'h3d, 8'hff, 8'h35, 8'h8a, 8'h7e, 8'h6d, 8'h54, 8'hc6, 8'h80, 8'hc3, 8'hbd, 8'h0d, 8'h57, 8'hdf, 8'hf5, 8'h24, 8'ha9, 8'h3e, 8'ha8, 8'h43, 8'hc9, 8'hd7, 8'h79, 8'hd6, 8'hf6, 8'h7c, 8'h22, 8'hb9, 8'h03, 8'he0, 8'h0f, 8'hec, 8'hde, 8'h7a, 8'h94, 8'hb0, 8'hbc, 8'hdc, 8'he8, 8'h28, 8'h50, 8'h4e, 8'h33, 8'h0a, 8'h4a, 8'ha7, 8'h97, 8'h60, 8'h73, 8'h1e, 8'h00, 8'h62, 8'h44, 8'h1a, 8'hb8, 8'h38, 8'h82, 8'h64, 8'h9f, 8'h26, 8'h41, 8'had, 8'h45, 8'h46, 8'h92, 8'h27, 8'h5e, 8'h55, 8'h2f, 8'h8c, 8'ha3, 8'ha5, 8'h7d, 8'h69, 8'hd5, 8'h95, 8'h3b, 8'h07, 8'h58, 8'hb3, 8'h40, 8'h86, 8'hac, 8'h1d, 8'hf7, 8'h30, 8'h37, 8'h6b, 8'he4, 8'h88, 8'hd9, 8'he7, 8'h89, 8'he1, 8'h1b, 8'h83, 8'h49, 8'h4c, 8'h3f, 8'hf8, 8'hfe, 8'h8d, 8'h53, 8'haa, 8'h90, 8'hca, 8'hd8, 8'h85, 8'h61, 8'h20, 8'h71, 8'h67, 8'ha4, 8'h2d, 8'h2b, 8'h09, 8'h5b, 8'hcb, 8'h9b, 8'h25, 8'hd0, 8'hbe, 8'he5, 8'h6c, 8'h52, 8'h59, 8'ha6, 8'h74, 8'hd2, 8'he6, 8'hf4, 8'hb4, 8'hc0, 8'hd1, 8'h66, 8'haf, 8'hc2, 8'h39, 8'h4b, 8'h63, 8'hb6};
  wire [7:0] literal_1076345[256] = '{8'h00, 8'h94, 8'heb, 8'h7f, 8'h15, 8'h81, 8'hfe, 8'h6a, 8'h2a, 8'hbe, 8'hc1, 8'h55, 8'h3f, 8'hab, 8'hd4, 8'h40, 8'h54, 8'hc0, 8'hbf, 8'h2b, 8'h41, 8'hd5, 8'haa, 8'h3e, 8'h7e, 8'hea, 8'h95, 8'h01, 8'h6b, 8'hff, 8'h80, 8'h14, 8'ha8, 8'h3c, 8'h43, 8'hd7, 8'hbd, 8'h29, 8'h56, 8'hc2, 8'h82, 8'h16, 8'h69, 8'hfd, 8'h97, 8'h03, 8'h7c, 8'he8, 8'hfc, 8'h68, 8'h17, 8'h83, 8'he9, 8'h7d, 8'h02, 8'h96, 8'hd6, 8'h42, 8'h3d, 8'ha9, 8'hc3, 8'h57, 8'h28, 8'hbc, 8'h93, 8'h07, 8'h78, 8'hec, 8'h86, 8'h12, 8'h6d, 8'hf9, 8'hb9, 8'h2d, 8'h52, 8'hc6, 8'hac, 8'h38, 8'h47, 8'hd3, 8'hc7, 8'h53, 8'h2c, 8'hb8, 8'hd2, 8'h46, 8'h39, 8'had, 8'hed, 8'h79, 8'h06, 8'h92, 8'hf8, 8'h6c, 8'h13, 8'h87, 8'h3b, 8'haf, 8'hd0, 8'h44, 8'h2e, 8'hba, 8'hc5, 8'h51, 8'h11, 8'h85, 8'hfa, 8'h6e, 8'h04, 8'h90, 8'hef, 8'h7b, 8'h6f, 8'hfb, 8'h84, 8'h10, 8'h7a, 8'hee, 8'h91, 8'h05, 8'h45, 8'hd1, 8'hae, 8'h3a, 8'h50, 8'hc4, 8'hbb, 8'h2f, 8'he5, 8'h71, 8'h0e, 8'h9a, 8'hf0, 8'h64, 8'h1b, 8'h8f, 8'hcf, 8'h5b, 8'h24, 8'hb0, 8'hda, 8'h4e, 8'h31, 8'ha5, 8'hb1, 8'h25, 8'h5a, 8'hce, 8'ha4, 8'h30, 8'h4f, 8'hdb, 8'h9b, 8'h0f, 8'h70, 8'he4, 8'h8e, 8'h1a, 8'h65, 8'hf1, 8'h4d, 8'hd9, 8'ha6, 8'h32, 8'h58, 8'hcc, 8'hb3, 8'h27, 8'h67, 8'hf3, 8'h8c, 8'h18, 8'h72, 8'he6, 8'h99, 8'h0d, 8'h19, 8'h8d, 8'hf2, 8'h66, 8'h0c, 8'h98, 8'he7, 8'h73, 8'h33, 8'ha7, 8'hd8, 8'h4c, 8'h26, 8'hb2, 8'hcd, 8'h59, 8'h76, 8'he2, 8'h9d, 8'h09, 8'h63, 8'hf7, 8'h88, 8'h1c, 8'h5c, 8'hc8, 8'hb7, 8'h23, 8'h49, 8'hdd, 8'ha2, 8'h36, 8'h22, 8'hb6, 8'hc9, 8'h5d, 8'h37, 8'ha3, 8'hdc, 8'h48, 8'h08, 8'h9c, 8'he3, 8'h77, 8'h1d, 8'h89, 8'hf6, 8'h62, 8'hde, 8'h4a, 8'h35, 8'ha1, 8'hcb, 8'h5f, 8'h20, 8'hb4, 8'hf4, 8'h60, 8'h1f, 8'h8b, 8'he1, 8'h75, 8'h0a, 8'h9e, 8'h8a, 8'h1e, 8'h61, 8'hf5, 8'h9f, 8'h0b, 8'h74, 8'he0, 8'ha0, 8'h34, 8'h4b, 8'hdf, 8'hb5, 8'h21, 8'h5e, 8'hca};
  wire [7:0] literal_1076347[256] = '{8'h00, 8'h20, 8'h40, 8'h60, 8'h80, 8'ha0, 8'hc0, 8'he0, 8'hc3, 8'he3, 8'h83, 8'ha3, 8'h43, 8'h63, 8'h03, 8'h23, 8'h45, 8'h65, 8'h05, 8'h25, 8'hc5, 8'he5, 8'h85, 8'ha5, 8'h86, 8'ha6, 8'hc6, 8'he6, 8'h06, 8'h26, 8'h46, 8'h66, 8'h8a, 8'haa, 8'hca, 8'hea, 8'h0a, 8'h2a, 8'h4a, 8'h6a, 8'h49, 8'h69, 8'h09, 8'h29, 8'hc9, 8'he9, 8'h89, 8'ha9, 8'hcf, 8'hef, 8'h8f, 8'haf, 8'h4f, 8'h6f, 8'h0f, 8'h2f, 8'h0c, 8'h2c, 8'h4c, 8'h6c, 8'h8c, 8'hac, 8'hcc, 8'hec, 8'hd7, 8'hf7, 8'h97, 8'hb7, 8'h57, 8'h77, 8'h17, 8'h37, 8'h14, 8'h34, 8'h54, 8'h74, 8'h94, 8'hb4, 8'hd4, 8'hf4, 8'h92, 8'hb2, 8'hd2, 8'hf2, 8'h12, 8'h32, 8'h52, 8'h72, 8'h51, 8'h71, 8'h11, 8'h31, 8'hd1, 8'hf1, 8'h91, 8'hb1, 8'h5d, 8'h7d, 8'h1d, 8'h3d, 8'hdd, 8'hfd, 8'h9d, 8'hbd, 8'h9e, 8'hbe, 8'hde, 8'hfe, 8'h1e, 8'h3e, 8'h5e, 8'h7e, 8'h18, 8'h38, 8'h58, 8'h78, 8'h98, 8'hb8, 8'hd8, 8'hf8, 8'hdb, 8'hfb, 8'h9b, 8'hbb, 8'h5b, 8'h7b, 8'h1b, 8'h3b, 8'h6d, 8'h4d, 8'h2d, 8'h0d, 8'hed, 8'hcd, 8'had, 8'h8d, 8'hae, 8'h8e, 8'hee, 8'hce, 8'h2e, 8'h0e, 8'h6e, 8'h4e, 8'h28, 8'h08, 8'h68, 8'h48, 8'ha8, 8'h88, 8'he8, 8'hc8, 8'heb, 8'hcb, 8'hab, 8'h8b, 8'h6b, 8'h4b, 8'h2b, 8'h0b, 8'he7, 8'hc7, 8'ha7, 8'h87, 8'h67, 8'h47, 8'h27, 8'h07, 8'h24, 8'h04, 8'h64, 8'h44, 8'ha4, 8'h84, 8'he4, 8'hc4, 8'ha2, 8'h82, 8'he2, 8'hc2, 8'h22, 8'h02, 8'h62, 8'h42, 8'h61, 8'h41, 8'h21, 8'h01, 8'he1, 8'hc1, 8'ha1, 8'h81, 8'hba, 8'h9a, 8'hfa, 8'hda, 8'h3a, 8'h1a, 8'h7a, 8'h5a, 8'h79, 8'h59, 8'h39, 8'h19, 8'hf9, 8'hd9, 8'hb9, 8'h99, 8'hff, 8'hdf, 8'hbf, 8'h9f, 8'h7f, 8'h5f, 8'h3f, 8'h1f, 8'h3c, 8'h1c, 8'h7c, 8'h5c, 8'hbc, 8'h9c, 8'hfc, 8'hdc, 8'h30, 8'h10, 8'h70, 8'h50, 8'hb0, 8'h90, 8'hf0, 8'hd0, 8'hf3, 8'hd3, 8'hb3, 8'h93, 8'h73, 8'h53, 8'h33, 8'h13, 8'h75, 8'h55, 8'h35, 8'h15, 8'hf5, 8'hd5, 8'hb5, 8'h95, 8'hb6, 8'h96, 8'hf6, 8'hd6, 8'h36, 8'h16, 8'h76, 8'h56};
  wire [7:0] literal_1076349[256] = '{8'h00, 8'h85, 8'hc9, 8'h4c, 8'h51, 8'hd4, 8'h98, 8'h1d, 8'ha2, 8'h27, 8'h6b, 8'hee, 8'hf3, 8'h76, 8'h3a, 8'hbf, 8'h87, 8'h02, 8'h4e, 8'hcb, 8'hd6, 8'h53, 8'h1f, 8'h9a, 8'h25, 8'ha0, 8'hec, 8'h69, 8'h74, 8'hf1, 8'hbd, 8'h38, 8'hcd, 8'h48, 8'h04, 8'h81, 8'h9c, 8'h19, 8'h55, 8'hd0, 8'h6f, 8'hea, 8'ha6, 8'h23, 8'h3e, 8'hbb, 8'hf7, 8'h72, 8'h4a, 8'hcf, 8'h83, 8'h06, 8'h1b, 8'h9e, 8'hd2, 8'h57, 8'he8, 8'h6d, 8'h21, 8'ha4, 8'hb9, 8'h3c, 8'h70, 8'hf5, 8'h59, 8'hdc, 8'h90, 8'h15, 8'h08, 8'h8d, 8'hc1, 8'h44, 8'hfb, 8'h7e, 8'h32, 8'hb7, 8'haa, 8'h2f, 8'h63, 8'he6, 8'hde, 8'h5b, 8'h17, 8'h92, 8'h8f, 8'h0a, 8'h46, 8'hc3, 8'h7c, 8'hf9, 8'hb5, 8'h30, 8'h2d, 8'ha8, 8'he4, 8'h61, 8'h94, 8'h11, 8'h5d, 8'hd8, 8'hc5, 8'h40, 8'h0c, 8'h89, 8'h36, 8'hb3, 8'hff, 8'h7a, 8'h67, 8'he2, 8'hae, 8'h2b, 8'h13, 8'h96, 8'hda, 8'h5f, 8'h42, 8'hc7, 8'h8b, 8'h0e, 8'hb1, 8'h34, 8'h78, 8'hfd, 8'he0, 8'h65, 8'h29, 8'hac, 8'hb2, 8'h37, 8'h7b, 8'hfe, 8'he3, 8'h66, 8'h2a, 8'haf, 8'h10, 8'h95, 8'hd9, 8'h5c, 8'h41, 8'hc4, 8'h88, 8'h0d, 8'h35, 8'hb0, 8'hfc, 8'h79, 8'h64, 8'he1, 8'had, 8'h28, 8'h97, 8'h12, 8'h5e, 8'hdb, 8'hc6, 8'h43, 8'h0f, 8'h8a, 8'h7f, 8'hfa, 8'hb6, 8'h33, 8'h2e, 8'hab, 8'he7, 8'h62, 8'hdd, 8'h58, 8'h14, 8'h91, 8'h8c, 8'h09, 8'h45, 8'hc0, 8'hf8, 8'h7d, 8'h31, 8'hb4, 8'ha9, 8'h2c, 8'h60, 8'he5, 8'h5a, 8'hdf, 8'h93, 8'h16, 8'h0b, 8'h8e, 8'hc2, 8'h47, 8'heb, 8'h6e, 8'h22, 8'ha7, 8'hba, 8'h3f, 8'h73, 8'hf6, 8'h49, 8'hcc, 8'h80, 8'h05, 8'h18, 8'h9d, 8'hd1, 8'h54, 8'h6c, 8'he9, 8'ha5, 8'h20, 8'h3d, 8'hb8, 8'hf4, 8'h71, 8'hce, 8'h4b, 8'h07, 8'h82, 8'h9f, 8'h1a, 8'h56, 8'hd3, 8'h26, 8'ha3, 8'hef, 8'h6a, 8'h77, 8'hf2, 8'hbe, 8'h3b, 8'h84, 8'h01, 8'h4d, 8'hc8, 8'hd5, 8'h50, 8'h1c, 8'h99, 8'ha1, 8'h24, 8'h68, 8'hed, 8'hf0, 8'h75, 8'h39, 8'hbc, 8'h03, 8'h86, 8'hca, 8'h4f, 8'h52, 8'hd7, 8'h9b, 8'h1e};
  wire [7:0] literal_1076351[256] = '{8'h00, 8'h10, 8'h20, 8'h30, 8'h40, 8'h50, 8'h60, 8'h70, 8'h80, 8'h90, 8'ha0, 8'hb0, 8'hc0, 8'hd0, 8'he0, 8'hf0, 8'hc3, 8'hd3, 8'he3, 8'hf3, 8'h83, 8'h93, 8'ha3, 8'hb3, 8'h43, 8'h53, 8'h63, 8'h73, 8'h03, 8'h13, 8'h23, 8'h33, 8'h45, 8'h55, 8'h65, 8'h75, 8'h05, 8'h15, 8'h25, 8'h35, 8'hc5, 8'hd5, 8'he5, 8'hf5, 8'h85, 8'h95, 8'ha5, 8'hb5, 8'h86, 8'h96, 8'ha6, 8'hb6, 8'hc6, 8'hd6, 8'he6, 8'hf6, 8'h06, 8'h16, 8'h26, 8'h36, 8'h46, 8'h56, 8'h66, 8'h76, 8'h8a, 8'h9a, 8'haa, 8'hba, 8'hca, 8'hda, 8'hea, 8'hfa, 8'h0a, 8'h1a, 8'h2a, 8'h3a, 8'h4a, 8'h5a, 8'h6a, 8'h7a, 8'h49, 8'h59, 8'h69, 8'h79, 8'h09, 8'h19, 8'h29, 8'h39, 8'hc9, 8'hd9, 8'he9, 8'hf9, 8'h89, 8'h99, 8'ha9, 8'hb9, 8'hcf, 8'hdf, 8'hef, 8'hff, 8'h8f, 8'h9f, 8'haf, 8'hbf, 8'h4f, 8'h5f, 8'h6f, 8'h7f, 8'h0f, 8'h1f, 8'h2f, 8'h3f, 8'h0c, 8'h1c, 8'h2c, 8'h3c, 8'h4c, 8'h5c, 8'h6c, 8'h7c, 8'h8c, 8'h9c, 8'hac, 8'hbc, 8'hcc, 8'hdc, 8'hec, 8'hfc, 8'hd7, 8'hc7, 8'hf7, 8'he7, 8'h97, 8'h87, 8'hb7, 8'ha7, 8'h57, 8'h47, 8'h77, 8'h67, 8'h17, 8'h07, 8'h37, 8'h27, 8'h14, 8'h04, 8'h34, 8'h24, 8'h54, 8'h44, 8'h74, 8'h64, 8'h94, 8'h84, 8'hb4, 8'ha4, 8'hd4, 8'hc4, 8'hf4, 8'he4, 8'h92, 8'h82, 8'hb2, 8'ha2, 8'hd2, 8'hc2, 8'hf2, 8'he2, 8'h12, 8'h02, 8'h32, 8'h22, 8'h52, 8'h42, 8'h72, 8'h62, 8'h51, 8'h41, 8'h71, 8'h61, 8'h11, 8'h01, 8'h31, 8'h21, 8'hd1, 8'hc1, 8'hf1, 8'he1, 8'h91, 8'h81, 8'hb1, 8'ha1, 8'h5d, 8'h4d, 8'h7d, 8'h6d, 8'h1d, 8'h0d, 8'h3d, 8'h2d, 8'hdd, 8'hcd, 8'hfd, 8'hed, 8'h9d, 8'h8d, 8'hbd, 8'had, 8'h9e, 8'h8e, 8'hbe, 8'hae, 8'hde, 8'hce, 8'hfe, 8'hee, 8'h1e, 8'h0e, 8'h3e, 8'h2e, 8'h5e, 8'h4e, 8'h7e, 8'h6e, 8'h18, 8'h08, 8'h38, 8'h28, 8'h58, 8'h48, 8'h78, 8'h68, 8'h98, 8'h88, 8'hb8, 8'ha8, 8'hd8, 8'hc8, 8'hf8, 8'he8, 8'hdb, 8'hcb, 8'hfb, 8'heb, 8'h9b, 8'h8b, 8'hbb, 8'hab, 8'h5b, 8'h4b, 8'h7b, 8'h6b, 8'h1b, 8'h0b, 8'h3b, 8'h2b};
  wire [7:0] literal_1076353[256] = '{8'h00, 8'hc2, 8'h47, 8'h85, 8'h8e, 8'h4c, 8'hc9, 8'h0b, 8'hdf, 8'h1d, 8'h98, 8'h5a, 8'h51, 8'h93, 8'h16, 8'hd4, 8'h7d, 8'hbf, 8'h3a, 8'hf8, 8'hf3, 8'h31, 8'hb4, 8'h76, 8'ha2, 8'h60, 8'he5, 8'h27, 8'h2c, 8'hee, 8'h6b, 8'ha9, 8'hfa, 8'h38, 8'hbd, 8'h7f, 8'h74, 8'hb6, 8'h33, 8'hf1, 8'h25, 8'he7, 8'h62, 8'ha0, 8'hab, 8'h69, 8'hec, 8'h2e, 8'h87, 8'h45, 8'hc0, 8'h02, 8'h09, 8'hcb, 8'h4e, 8'h8c, 8'h58, 8'h9a, 8'h1f, 8'hdd, 8'hd6, 8'h14, 8'h91, 8'h53, 8'h37, 8'hf5, 8'h70, 8'hb2, 8'hb9, 8'h7b, 8'hfe, 8'h3c, 8'he8, 8'h2a, 8'haf, 8'h6d, 8'h66, 8'ha4, 8'h21, 8'he3, 8'h4a, 8'h88, 8'h0d, 8'hcf, 8'hc4, 8'h06, 8'h83, 8'h41, 8'h95, 8'h57, 8'hd2, 8'h10, 8'h1b, 8'hd9, 8'h5c, 8'h9e, 8'hcd, 8'h0f, 8'h8a, 8'h48, 8'h43, 8'h81, 8'h04, 8'hc6, 8'h12, 8'hd0, 8'h55, 8'h97, 8'h9c, 8'h5e, 8'hdb, 8'h19, 8'hb0, 8'h72, 8'hf7, 8'h35, 8'h3e, 8'hfc, 8'h79, 8'hbb, 8'h6f, 8'had, 8'h28, 8'hea, 8'he1, 8'h23, 8'ha6, 8'h64, 8'h6e, 8'hac, 8'h29, 8'heb, 8'he0, 8'h22, 8'ha7, 8'h65, 8'hb1, 8'h73, 8'hf6, 8'h34, 8'h3f, 8'hfd, 8'h78, 8'hba, 8'h13, 8'hd1, 8'h54, 8'h96, 8'h9d, 8'h5f, 8'hda, 8'h18, 8'hcc, 8'h0e, 8'h8b, 8'h49, 8'h42, 8'h80, 8'h05, 8'hc7, 8'h94, 8'h56, 8'hd3, 8'h11, 8'h1a, 8'hd8, 8'h5d, 8'h9f, 8'h4b, 8'h89, 8'h0c, 8'hce, 8'hc5, 8'h07, 8'h82, 8'h40, 8'he9, 8'h2b, 8'hae, 8'h6c, 8'h67, 8'ha5, 8'h20, 8'he2, 8'h36, 8'hf4, 8'h71, 8'hb3, 8'hb8, 8'h7a, 8'hff, 8'h3d, 8'h59, 8'h9b, 8'h1e, 8'hdc, 8'hd7, 8'h15, 8'h90, 8'h52, 8'h86, 8'h44, 8'hc1, 8'h03, 8'h08, 8'hca, 8'h4f, 8'h8d, 8'h24, 8'he6, 8'h63, 8'ha1, 8'haa, 8'h68, 8'hed, 8'h2f, 8'hfb, 8'h39, 8'hbc, 8'h7e, 8'h75, 8'hb7, 8'h32, 8'hf0, 8'ha3, 8'h61, 8'he4, 8'h26, 8'h2d, 8'hef, 8'h6a, 8'ha8, 8'h7c, 8'hbe, 8'h3b, 8'hf9, 8'hf2, 8'h30, 8'hb5, 8'h77, 8'hde, 8'h1c, 8'h99, 8'h5b, 8'h50, 8'h92, 8'h17, 8'hd5, 8'h01, 8'hc3, 8'h46, 8'h84, 8'h8f, 8'h4d, 8'hc8, 8'h0a};
  wire [7:0] literal_1076355[256] = '{8'h00, 8'hc0, 8'h43, 8'h83, 8'h86, 8'h46, 8'hc5, 8'h05, 8'hcf, 8'h0f, 8'h8c, 8'h4c, 8'h49, 8'h89, 8'h0a, 8'hca, 8'h5d, 8'h9d, 8'h1e, 8'hde, 8'hdb, 8'h1b, 8'h98, 8'h58, 8'h92, 8'h52, 8'hd1, 8'h11, 8'h14, 8'hd4, 8'h57, 8'h97, 8'hba, 8'h7a, 8'hf9, 8'h39, 8'h3c, 8'hfc, 8'h7f, 8'hbf, 8'h75, 8'hb5, 8'h36, 8'hf6, 8'hf3, 8'h33, 8'hb0, 8'h70, 8'he7, 8'h27, 8'ha4, 8'h64, 8'h61, 8'ha1, 8'h22, 8'he2, 8'h28, 8'he8, 8'h6b, 8'hab, 8'hae, 8'h6e, 8'hed, 8'h2d, 8'hb7, 8'h77, 8'hf4, 8'h34, 8'h31, 8'hf1, 8'h72, 8'hb2, 8'h78, 8'hb8, 8'h3b, 8'hfb, 8'hfe, 8'h3e, 8'hbd, 8'h7d, 8'hea, 8'h2a, 8'ha9, 8'h69, 8'h6c, 8'hac, 8'h2f, 8'hef, 8'h25, 8'he5, 8'h66, 8'ha6, 8'ha3, 8'h63, 8'he0, 8'h20, 8'h0d, 8'hcd, 8'h4e, 8'h8e, 8'h8b, 8'h4b, 8'hc8, 8'h08, 8'hc2, 8'h02, 8'h81, 8'h41, 8'h44, 8'h84, 8'h07, 8'hc7, 8'h50, 8'h90, 8'h13, 8'hd3, 8'hd6, 8'h16, 8'h95, 8'h55, 8'h9f, 8'h5f, 8'hdc, 8'h1c, 8'h19, 8'hd9, 8'h5a, 8'h9a, 8'had, 8'h6d, 8'hee, 8'h2e, 8'h2b, 8'heb, 8'h68, 8'ha8, 8'h62, 8'ha2, 8'h21, 8'he1, 8'he4, 8'h24, 8'ha7, 8'h67, 8'hf0, 8'h30, 8'hb3, 8'h73, 8'h76, 8'hb6, 8'h35, 8'hf5, 8'h3f, 8'hff, 8'h7c, 8'hbc, 8'hb9, 8'h79, 8'hfa, 8'h3a, 8'h17, 8'hd7, 8'h54, 8'h94, 8'h91, 8'h51, 8'hd2, 8'h12, 8'hd8, 8'h18, 8'h9b, 8'h5b, 8'h5e, 8'h9e, 8'h1d, 8'hdd, 8'h4a, 8'h8a, 8'h09, 8'hc9, 8'hcc, 8'h0c, 8'h8f, 8'h4f, 8'h85, 8'h45, 8'hc6, 8'h06, 8'h03, 8'hc3, 8'h40, 8'h80, 8'h1a, 8'hda, 8'h59, 8'h99, 8'h9c, 8'h5c, 8'hdf, 8'h1f, 8'hd5, 8'h15, 8'h96, 8'h56, 8'h53, 8'h93, 8'h10, 8'hd0, 8'h47, 8'h87, 8'h04, 8'hc4, 8'hc1, 8'h01, 8'h82, 8'h42, 8'h88, 8'h48, 8'hcb, 8'h0b, 8'h0e, 8'hce, 8'h4d, 8'h8d, 8'ha0, 8'h60, 8'he3, 8'h23, 8'h26, 8'he6, 8'h65, 8'ha5, 8'h6f, 8'haf, 8'h2c, 8'hec, 8'he9, 8'h29, 8'haa, 8'h6a, 8'hfd, 8'h3d, 8'hbe, 8'h7e, 8'h7b, 8'hbb, 8'h38, 8'hf8, 8'h32, 8'hf2, 8'h71, 8'hb1, 8'hb4, 8'h74, 8'hf7, 8'h37};
  wire [7:0] literal_1076358[256] = '{8'h00, 8'hfb, 8'h35, 8'hce, 8'h6a, 8'h91, 8'h5f, 8'ha4, 8'hd4, 8'h2f, 8'he1, 8'h1a, 8'hbe, 8'h45, 8'h8b, 8'h70, 8'h6b, 8'h90, 8'h5e, 8'ha5, 8'h01, 8'hfa, 8'h34, 8'hcf, 8'hbf, 8'h44, 8'h8a, 8'h71, 8'hd5, 8'h2e, 8'he0, 8'h1b, 8'hd6, 8'h2d, 8'he3, 8'h18, 8'hbc, 8'h47, 8'h89, 8'h72, 8'h02, 8'hf9, 8'h37, 8'hcc, 8'h68, 8'h93, 8'h5d, 8'ha6, 8'hbd, 8'h46, 8'h88, 8'h73, 8'hd7, 8'h2c, 8'he2, 8'h19, 8'h69, 8'h92, 8'h5c, 8'ha7, 8'h03, 8'hf8, 8'h36, 8'hcd, 8'h6f, 8'h94, 8'h5a, 8'ha1, 8'h05, 8'hfe, 8'h30, 8'hcb, 8'hbb, 8'h40, 8'h8e, 8'h75, 8'hd1, 8'h2a, 8'he4, 8'h1f, 8'h04, 8'hff, 8'h31, 8'hca, 8'h6e, 8'h95, 8'h5b, 8'ha0, 8'hd0, 8'h2b, 8'he5, 8'h1e, 8'hba, 8'h41, 8'h8f, 8'h74, 8'hb9, 8'h42, 8'h8c, 8'h77, 8'hd3, 8'h28, 8'he6, 8'h1d, 8'h6d, 8'h96, 8'h58, 8'ha3, 8'h07, 8'hfc, 8'h32, 8'hc9, 8'hd2, 8'h29, 8'he7, 8'h1c, 8'hb8, 8'h43, 8'h8d, 8'h76, 8'h06, 8'hfd, 8'h33, 8'hc8, 8'h6c, 8'h97, 8'h59, 8'ha2, 8'hde, 8'h25, 8'heb, 8'h10, 8'hb4, 8'h4f, 8'h81, 8'h7a, 8'h0a, 8'hf1, 8'h3f, 8'hc4, 8'h60, 8'h9b, 8'h55, 8'hae, 8'hb5, 8'h4e, 8'h80, 8'h7b, 8'hdf, 8'h24, 8'hea, 8'h11, 8'h61, 8'h9a, 8'h54, 8'haf, 8'h0b, 8'hf0, 8'h3e, 8'hc5, 8'h08, 8'hf3, 8'h3d, 8'hc6, 8'h62, 8'h99, 8'h57, 8'hac, 8'hdc, 8'h27, 8'he9, 8'h12, 8'hb6, 8'h4d, 8'h83, 8'h78, 8'h63, 8'h98, 8'h56, 8'had, 8'h09, 8'hf2, 8'h3c, 8'hc7, 8'hb7, 8'h4c, 8'h82, 8'h79, 8'hdd, 8'h26, 8'he8, 8'h13, 8'hb1, 8'h4a, 8'h84, 8'h7f, 8'hdb, 8'h20, 8'hee, 8'h15, 8'h65, 8'h9e, 8'h50, 8'hab, 8'h0f, 8'hf4, 8'h3a, 8'hc1, 8'hda, 8'h21, 8'hef, 8'h14, 8'hb0, 8'h4b, 8'h85, 8'h7e, 8'h0e, 8'hf5, 8'h3b, 8'hc0, 8'h64, 8'h9f, 8'h51, 8'haa, 8'h67, 8'h9c, 8'h52, 8'ha9, 8'h0d, 8'hf6, 8'h38, 8'hc3, 8'hb3, 8'h48, 8'h86, 8'h7d, 8'hd9, 8'h22, 8'hec, 8'h17, 8'h0c, 8'hf7, 8'h39, 8'hc2, 8'h66, 8'h9d, 8'h53, 8'ha8, 8'hd8, 8'h23, 8'hed, 8'h16, 8'hb2, 8'h49, 8'h87, 8'h7c};

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [127:0] p0__block;
  reg [255:0] p0_key;
  reg [7:0] p1_arr[256];
  reg [7:0] p1_literal_1076345[256];
  reg [7:0] p1_literal_1076347[256];
  reg [7:0] p1_literal_1076349[256];
  reg [7:0] p1_literal_1076351[256];
  reg [7:0] p1_literal_1076353[256];
  reg [7:0] p1_literal_1076355[256];
  reg [7:0] p1_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p0__block <= _block;
    p0_key <= key;
    p1_arr <= arr;
    p1_literal_1076345 <= literal_1076345;
    p1_literal_1076347 <= literal_1076347;
    p1_literal_1076349 <= literal_1076349;
    p1_literal_1076351 <= literal_1076351;
    p1_literal_1076353 <= literal_1076353;
    p1_literal_1076355 <= literal_1076355;
    p1_literal_1076358 <= literal_1076358;
  end

  // ===== Pipe stage 1:
  wire [127:0] p1_bit_slice_1076328_comb;
  wire [127:0] p1_addedKey__41_comb;
  wire [127:0] p1_addedKey__32_comb;
  wire [7:0] p1_array_index_1076346_comb;
  wire [7:0] p1_array_index_1076348_comb;
  wire [7:0] p1_array_index_1076350_comb;
  wire [7:0] p1_array_index_1076352_comb;
  wire [7:0] p1_array_index_1076354_comb;
  wire [7:0] p1_array_index_1076356_comb;
  wire [7:0] p1_array_index_1076359_comb;
  wire [7:0] p1_array_index_1076361_comb;
  wire [7:0] p1_array_index_1076362_comb;
  wire [7:0] p1_array_index_1076363_comb;
  wire [7:0] p1_array_index_1076364_comb;
  wire [7:0] p1_array_index_1076365_comb;
  wire [7:0] p1_array_index_1076366_comb;
  wire [7:0] p1_array_index_1076455_comb;
  wire [7:0] p1_array_index_1076456_comb;
  wire [7:0] p1_array_index_1076457_comb;
  wire [7:0] p1_array_index_1076458_comb;
  wire [7:0] p1_array_index_1076459_comb;
  wire [7:0] p1_array_index_1076460_comb;
  wire [7:0] p1_array_index_1076462_comb;
  wire [7:0] p1_array_index_1076464_comb;
  wire [7:0] p1_array_index_1076465_comb;
  wire [7:0] p1_array_index_1076466_comb;
  wire [7:0] p1_array_index_1076467_comb;
  wire [7:0] p1_array_index_1076468_comb;
  wire [7:0] p1_array_index_1076469_comb;
  wire [7:0] p1_array_index_1076368_comb;
  wire [7:0] p1_array_index_1076369_comb;
  wire [7:0] p1_array_index_1076370_comb;
  wire [7:0] p1_array_index_1076371_comb;
  wire [7:0] p1_array_index_1076372_comb;
  wire [7:0] p1_array_index_1076373_comb;
  wire [7:0] p1_array_index_1076374_comb;
  wire [7:0] p1_array_index_1076376_comb;
  wire [7:0] p1_array_index_1076471_comb;
  wire [7:0] p1_array_index_1076472_comb;
  wire [7:0] p1_array_index_1076473_comb;
  wire [7:0] p1_array_index_1076474_comb;
  wire [7:0] p1_array_index_1076475_comb;
  wire [7:0] p1_array_index_1076476_comb;
  wire [7:0] p1_array_index_1076477_comb;
  wire [7:0] p1_array_index_1076479_comb;
  wire [7:0] p1_res7_comb;
  wire [7:0] p1_res7__512_comb;
  wire [7:0] p1_array_index_1076385_comb;
  wire [7:0] p1_array_index_1076386_comb;
  wire [7:0] p1_array_index_1076387_comb;
  wire [7:0] p1_array_index_1076388_comb;
  wire [7:0] p1_array_index_1076389_comb;
  wire [7:0] p1_array_index_1076390_comb;
  wire [7:0] p1_array_index_1076488_comb;
  wire [7:0] p1_array_index_1076489_comb;
  wire [7:0] p1_array_index_1076490_comb;
  wire [7:0] p1_array_index_1076491_comb;
  wire [7:0] p1_array_index_1076492_comb;
  wire [7:0] p1_array_index_1076493_comb;
  wire [7:0] p1_res7__1_comb;
  wire [7:0] p1_res7__513_comb;
  wire [7:0] p1_array_index_1076400_comb;
  wire [7:0] p1_array_index_1076401_comb;
  wire [7:0] p1_array_index_1076402_comb;
  wire [7:0] p1_array_index_1076403_comb;
  wire [7:0] p1_array_index_1076404_comb;
  wire [7:0] p1_array_index_1076503_comb;
  wire [7:0] p1_array_index_1076504_comb;
  wire [7:0] p1_array_index_1076505_comb;
  wire [7:0] p1_array_index_1076506_comb;
  wire [7:0] p1_array_index_1076507_comb;
  wire [7:0] p1_res7__2_comb;
  wire [7:0] p1_res7__514_comb;
  wire [7:0] p1_array_index_1076414_comb;
  wire [7:0] p1_array_index_1076415_comb;
  wire [7:0] p1_array_index_1076416_comb;
  wire [7:0] p1_array_index_1076417_comb;
  wire [7:0] p1_array_index_1076418_comb;
  wire [7:0] p1_array_index_1076517_comb;
  wire [7:0] p1_array_index_1076518_comb;
  wire [7:0] p1_array_index_1076519_comb;
  wire [7:0] p1_array_index_1076520_comb;
  wire [7:0] p1_array_index_1076521_comb;
  wire [7:0] p1_res7__3_comb;
  wire [7:0] p1_res7__515_comb;
  wire [7:0] p1_array_index_1076429_comb;
  wire [7:0] p1_array_index_1076430_comb;
  wire [7:0] p1_array_index_1076431_comb;
  wire [7:0] p1_array_index_1076432_comb;
  wire [7:0] p1_array_index_1076532_comb;
  wire [7:0] p1_array_index_1076533_comb;
  wire [7:0] p1_array_index_1076534_comb;
  wire [7:0] p1_array_index_1076535_comb;
  wire [7:0] p1_res7__4_comb;
  wire [127:0] p1_bit_slice_1076440_comb;
  wire [7:0] p1_res7__516_comb;
  assign p1_bit_slice_1076328_comb = p0_key[255:128];
  assign p1_addedKey__41_comb = p1_bit_slice_1076328_comb ^ 128'h6ea2_7672_6c48_7ab8_5d27_bd10_dd84_9401;
  assign p1_addedKey__32_comb = p1_bit_slice_1076328_comb ^ p0__block;
  assign p1_array_index_1076346_comb = arr[p1_addedKey__41_comb[127:120]];
  assign p1_array_index_1076348_comb = arr[p1_addedKey__41_comb[119:112]];
  assign p1_array_index_1076350_comb = arr[p1_addedKey__41_comb[111:104]];
  assign p1_array_index_1076352_comb = arr[p1_addedKey__41_comb[103:96]];
  assign p1_array_index_1076354_comb = arr[p1_addedKey__41_comb[95:88]];
  assign p1_array_index_1076356_comb = arr[p1_addedKey__41_comb[87:80]];
  assign p1_array_index_1076359_comb = arr[p1_addedKey__41_comb[71:64]];
  assign p1_array_index_1076361_comb = arr[p1_addedKey__41_comb[55:48]];
  assign p1_array_index_1076362_comb = arr[p1_addedKey__41_comb[47:40]];
  assign p1_array_index_1076363_comb = arr[p1_addedKey__41_comb[39:32]];
  assign p1_array_index_1076364_comb = arr[p1_addedKey__41_comb[31:24]];
  assign p1_array_index_1076365_comb = arr[p1_addedKey__41_comb[23:16]];
  assign p1_array_index_1076366_comb = arr[p1_addedKey__41_comb[15:8]];
  assign p1_array_index_1076455_comb = arr[p1_addedKey__32_comb[127:120]];
  assign p1_array_index_1076456_comb = arr[p1_addedKey__32_comb[119:112]];
  assign p1_array_index_1076457_comb = arr[p1_addedKey__32_comb[111:104]];
  assign p1_array_index_1076458_comb = arr[p1_addedKey__32_comb[103:96]];
  assign p1_array_index_1076459_comb = arr[p1_addedKey__32_comb[95:88]];
  assign p1_array_index_1076460_comb = arr[p1_addedKey__32_comb[87:80]];
  assign p1_array_index_1076462_comb = arr[p1_addedKey__32_comb[71:64]];
  assign p1_array_index_1076464_comb = arr[p1_addedKey__32_comb[55:48]];
  assign p1_array_index_1076465_comb = arr[p1_addedKey__32_comb[47:40]];
  assign p1_array_index_1076466_comb = arr[p1_addedKey__32_comb[39:32]];
  assign p1_array_index_1076467_comb = arr[p1_addedKey__32_comb[31:24]];
  assign p1_array_index_1076468_comb = arr[p1_addedKey__32_comb[23:16]];
  assign p1_array_index_1076469_comb = arr[p1_addedKey__32_comb[15:8]];
  assign p1_array_index_1076368_comb = literal_1076345[p1_array_index_1076346_comb];
  assign p1_array_index_1076369_comb = literal_1076347[p1_array_index_1076348_comb];
  assign p1_array_index_1076370_comb = literal_1076349[p1_array_index_1076350_comb];
  assign p1_array_index_1076371_comb = literal_1076351[p1_array_index_1076352_comb];
  assign p1_array_index_1076372_comb = literal_1076353[p1_array_index_1076354_comb];
  assign p1_array_index_1076373_comb = literal_1076355[p1_array_index_1076356_comb];
  assign p1_array_index_1076374_comb = arr[p1_addedKey__41_comb[79:72]];
  assign p1_array_index_1076376_comb = arr[p1_addedKey__41_comb[63:56]];
  assign p1_array_index_1076471_comb = literal_1076345[p1_array_index_1076455_comb];
  assign p1_array_index_1076472_comb = literal_1076347[p1_array_index_1076456_comb];
  assign p1_array_index_1076473_comb = literal_1076349[p1_array_index_1076457_comb];
  assign p1_array_index_1076474_comb = literal_1076351[p1_array_index_1076458_comb];
  assign p1_array_index_1076475_comb = literal_1076353[p1_array_index_1076459_comb];
  assign p1_array_index_1076476_comb = literal_1076355[p1_array_index_1076460_comb];
  assign p1_array_index_1076477_comb = arr[p1_addedKey__32_comb[79:72]];
  assign p1_array_index_1076479_comb = arr[p1_addedKey__32_comb[63:56]];
  assign p1_res7_comb = p1_array_index_1076368_comb ^ p1_array_index_1076369_comb ^ p1_array_index_1076370_comb ^ p1_array_index_1076371_comb ^ p1_array_index_1076372_comb ^ p1_array_index_1076373_comb ^ p1_array_index_1076374_comb ^ literal_1076358[p1_array_index_1076359_comb] ^ p1_array_index_1076376_comb ^ literal_1076355[p1_array_index_1076361_comb] ^ literal_1076353[p1_array_index_1076362_comb] ^ literal_1076351[p1_array_index_1076363_comb] ^ literal_1076349[p1_array_index_1076364_comb] ^ literal_1076347[p1_array_index_1076365_comb] ^ literal_1076345[p1_array_index_1076366_comb] ^ arr[p1_addedKey__41_comb[7:0]];
  assign p1_res7__512_comb = p1_array_index_1076471_comb ^ p1_array_index_1076472_comb ^ p1_array_index_1076473_comb ^ p1_array_index_1076474_comb ^ p1_array_index_1076475_comb ^ p1_array_index_1076476_comb ^ p1_array_index_1076477_comb ^ literal_1076358[p1_array_index_1076462_comb] ^ p1_array_index_1076479_comb ^ literal_1076355[p1_array_index_1076464_comb] ^ literal_1076353[p1_array_index_1076465_comb] ^ literal_1076351[p1_array_index_1076466_comb] ^ literal_1076349[p1_array_index_1076467_comb] ^ literal_1076347[p1_array_index_1076468_comb] ^ literal_1076345[p1_array_index_1076469_comb] ^ arr[p1_addedKey__32_comb[7:0]];
  assign p1_array_index_1076385_comb = literal_1076345[p1_res7_comb];
  assign p1_array_index_1076386_comb = literal_1076347[p1_array_index_1076346_comb];
  assign p1_array_index_1076387_comb = literal_1076349[p1_array_index_1076348_comb];
  assign p1_array_index_1076388_comb = literal_1076351[p1_array_index_1076350_comb];
  assign p1_array_index_1076389_comb = literal_1076353[p1_array_index_1076352_comb];
  assign p1_array_index_1076390_comb = literal_1076355[p1_array_index_1076354_comb];
  assign p1_array_index_1076488_comb = literal_1076345[p1_res7__512_comb];
  assign p1_array_index_1076489_comb = literal_1076347[p1_array_index_1076455_comb];
  assign p1_array_index_1076490_comb = literal_1076349[p1_array_index_1076456_comb];
  assign p1_array_index_1076491_comb = literal_1076351[p1_array_index_1076457_comb];
  assign p1_array_index_1076492_comb = literal_1076353[p1_array_index_1076458_comb];
  assign p1_array_index_1076493_comb = literal_1076355[p1_array_index_1076459_comb];
  assign p1_res7__1_comb = p1_array_index_1076385_comb ^ p1_array_index_1076386_comb ^ p1_array_index_1076387_comb ^ p1_array_index_1076388_comb ^ p1_array_index_1076389_comb ^ p1_array_index_1076390_comb ^ p1_array_index_1076356_comb ^ literal_1076358[p1_array_index_1076374_comb] ^ p1_array_index_1076359_comb ^ literal_1076355[p1_array_index_1076376_comb] ^ literal_1076353[p1_array_index_1076361_comb] ^ literal_1076351[p1_array_index_1076362_comb] ^ literal_1076349[p1_array_index_1076363_comb] ^ literal_1076347[p1_array_index_1076364_comb] ^ literal_1076345[p1_array_index_1076365_comb] ^ p1_array_index_1076366_comb;
  assign p1_res7__513_comb = p1_array_index_1076488_comb ^ p1_array_index_1076489_comb ^ p1_array_index_1076490_comb ^ p1_array_index_1076491_comb ^ p1_array_index_1076492_comb ^ p1_array_index_1076493_comb ^ p1_array_index_1076460_comb ^ literal_1076358[p1_array_index_1076477_comb] ^ p1_array_index_1076462_comb ^ literal_1076355[p1_array_index_1076479_comb] ^ literal_1076353[p1_array_index_1076464_comb] ^ literal_1076351[p1_array_index_1076465_comb] ^ literal_1076349[p1_array_index_1076466_comb] ^ literal_1076347[p1_array_index_1076467_comb] ^ literal_1076345[p1_array_index_1076468_comb] ^ p1_array_index_1076469_comb;
  assign p1_array_index_1076400_comb = literal_1076347[p1_res7_comb];
  assign p1_array_index_1076401_comb = literal_1076349[p1_array_index_1076346_comb];
  assign p1_array_index_1076402_comb = literal_1076351[p1_array_index_1076348_comb];
  assign p1_array_index_1076403_comb = literal_1076353[p1_array_index_1076350_comb];
  assign p1_array_index_1076404_comb = literal_1076355[p1_array_index_1076352_comb];
  assign p1_array_index_1076503_comb = literal_1076347[p1_res7__512_comb];
  assign p1_array_index_1076504_comb = literal_1076349[p1_array_index_1076455_comb];
  assign p1_array_index_1076505_comb = literal_1076351[p1_array_index_1076456_comb];
  assign p1_array_index_1076506_comb = literal_1076353[p1_array_index_1076457_comb];
  assign p1_array_index_1076507_comb = literal_1076355[p1_array_index_1076458_comb];
  assign p1_res7__2_comb = literal_1076345[p1_res7__1_comb] ^ p1_array_index_1076400_comb ^ p1_array_index_1076401_comb ^ p1_array_index_1076402_comb ^ p1_array_index_1076403_comb ^ p1_array_index_1076404_comb ^ p1_array_index_1076354_comb ^ literal_1076358[p1_array_index_1076356_comb] ^ p1_array_index_1076374_comb ^ literal_1076355[p1_array_index_1076359_comb] ^ literal_1076353[p1_array_index_1076376_comb] ^ literal_1076351[p1_array_index_1076361_comb] ^ literal_1076349[p1_array_index_1076362_comb] ^ literal_1076347[p1_array_index_1076363_comb] ^ literal_1076345[p1_array_index_1076364_comb] ^ p1_array_index_1076365_comb;
  assign p1_res7__514_comb = literal_1076345[p1_res7__513_comb] ^ p1_array_index_1076503_comb ^ p1_array_index_1076504_comb ^ p1_array_index_1076505_comb ^ p1_array_index_1076506_comb ^ p1_array_index_1076507_comb ^ p1_array_index_1076459_comb ^ literal_1076358[p1_array_index_1076460_comb] ^ p1_array_index_1076477_comb ^ literal_1076355[p1_array_index_1076462_comb] ^ literal_1076353[p1_array_index_1076479_comb] ^ literal_1076351[p1_array_index_1076464_comb] ^ literal_1076349[p1_array_index_1076465_comb] ^ literal_1076347[p1_array_index_1076466_comb] ^ literal_1076345[p1_array_index_1076467_comb] ^ p1_array_index_1076468_comb;
  assign p1_array_index_1076414_comb = literal_1076347[p1_res7__1_comb];
  assign p1_array_index_1076415_comb = literal_1076349[p1_res7_comb];
  assign p1_array_index_1076416_comb = literal_1076351[p1_array_index_1076346_comb];
  assign p1_array_index_1076417_comb = literal_1076353[p1_array_index_1076348_comb];
  assign p1_array_index_1076418_comb = literal_1076355[p1_array_index_1076350_comb];
  assign p1_array_index_1076517_comb = literal_1076347[p1_res7__513_comb];
  assign p1_array_index_1076518_comb = literal_1076349[p1_res7__512_comb];
  assign p1_array_index_1076519_comb = literal_1076351[p1_array_index_1076455_comb];
  assign p1_array_index_1076520_comb = literal_1076353[p1_array_index_1076456_comb];
  assign p1_array_index_1076521_comb = literal_1076355[p1_array_index_1076457_comb];
  assign p1_res7__3_comb = literal_1076345[p1_res7__2_comb] ^ p1_array_index_1076414_comb ^ p1_array_index_1076415_comb ^ p1_array_index_1076416_comb ^ p1_array_index_1076417_comb ^ p1_array_index_1076418_comb ^ p1_array_index_1076352_comb ^ literal_1076358[p1_array_index_1076354_comb] ^ p1_array_index_1076356_comb ^ literal_1076355[p1_array_index_1076374_comb] ^ literal_1076353[p1_array_index_1076359_comb] ^ literal_1076351[p1_array_index_1076376_comb] ^ literal_1076349[p1_array_index_1076361_comb] ^ literal_1076347[p1_array_index_1076362_comb] ^ literal_1076345[p1_array_index_1076363_comb] ^ p1_array_index_1076364_comb;
  assign p1_res7__515_comb = literal_1076345[p1_res7__514_comb] ^ p1_array_index_1076517_comb ^ p1_array_index_1076518_comb ^ p1_array_index_1076519_comb ^ p1_array_index_1076520_comb ^ p1_array_index_1076521_comb ^ p1_array_index_1076458_comb ^ literal_1076358[p1_array_index_1076459_comb] ^ p1_array_index_1076460_comb ^ literal_1076355[p1_array_index_1076477_comb] ^ literal_1076353[p1_array_index_1076462_comb] ^ literal_1076351[p1_array_index_1076479_comb] ^ literal_1076349[p1_array_index_1076464_comb] ^ literal_1076347[p1_array_index_1076465_comb] ^ literal_1076345[p1_array_index_1076466_comb] ^ p1_array_index_1076467_comb;
  assign p1_array_index_1076429_comb = literal_1076349[p1_res7__1_comb];
  assign p1_array_index_1076430_comb = literal_1076351[p1_res7_comb];
  assign p1_array_index_1076431_comb = literal_1076353[p1_array_index_1076346_comb];
  assign p1_array_index_1076432_comb = literal_1076355[p1_array_index_1076348_comb];
  assign p1_array_index_1076532_comb = literal_1076349[p1_res7__513_comb];
  assign p1_array_index_1076533_comb = literal_1076351[p1_res7__512_comb];
  assign p1_array_index_1076534_comb = literal_1076353[p1_array_index_1076455_comb];
  assign p1_array_index_1076535_comb = literal_1076355[p1_array_index_1076456_comb];
  assign p1_res7__4_comb = literal_1076345[p1_res7__3_comb] ^ literal_1076347[p1_res7__2_comb] ^ p1_array_index_1076429_comb ^ p1_array_index_1076430_comb ^ p1_array_index_1076431_comb ^ p1_array_index_1076432_comb ^ p1_array_index_1076350_comb ^ literal_1076358[p1_array_index_1076352_comb] ^ p1_array_index_1076354_comb ^ p1_array_index_1076373_comb ^ literal_1076353[p1_array_index_1076374_comb] ^ literal_1076351[p1_array_index_1076359_comb] ^ literal_1076349[p1_array_index_1076376_comb] ^ literal_1076347[p1_array_index_1076361_comb] ^ literal_1076345[p1_array_index_1076362_comb] ^ p1_array_index_1076363_comb;
  assign p1_bit_slice_1076440_comb = p0_key[127:0];
  assign p1_res7__516_comb = literal_1076345[p1_res7__515_comb] ^ literal_1076347[p1_res7__514_comb] ^ p1_array_index_1076532_comb ^ p1_array_index_1076533_comb ^ p1_array_index_1076534_comb ^ p1_array_index_1076535_comb ^ p1_array_index_1076457_comb ^ literal_1076358[p1_array_index_1076458_comb] ^ p1_array_index_1076459_comb ^ p1_array_index_1076476_comb ^ literal_1076353[p1_array_index_1076477_comb] ^ literal_1076351[p1_array_index_1076462_comb] ^ literal_1076349[p1_array_index_1076479_comb] ^ literal_1076347[p1_array_index_1076464_comb] ^ literal_1076345[p1_array_index_1076465_comb] ^ p1_array_index_1076466_comb;

  // Registers for pipe stage 1:
  reg [127:0] p1_bit_slice_1076328;
  reg [7:0] p1_array_index_1076346;
  reg [7:0] p1_array_index_1076348;
  reg [7:0] p1_array_index_1076350;
  reg [7:0] p1_array_index_1076352;
  reg [7:0] p1_array_index_1076354;
  reg [7:0] p1_array_index_1076356;
  reg [7:0] p1_array_index_1076359;
  reg [7:0] p1_array_index_1076361;
  reg [7:0] p1_array_index_1076362;
  reg [7:0] p1_array_index_1076368;
  reg [7:0] p1_array_index_1076369;
  reg [7:0] p1_array_index_1076370;
  reg [7:0] p1_array_index_1076371;
  reg [7:0] p1_array_index_1076372;
  reg [7:0] p1_array_index_1076374;
  reg [7:0] p1_array_index_1076376;
  reg [7:0] p1_res7;
  reg [7:0] p1_array_index_1076385;
  reg [7:0] p1_array_index_1076386;
  reg [7:0] p1_array_index_1076387;
  reg [7:0] p1_array_index_1076388;
  reg [7:0] p1_array_index_1076389;
  reg [7:0] p1_array_index_1076390;
  reg [7:0] p1_res7__1;
  reg [7:0] p1_array_index_1076400;
  reg [7:0] p1_array_index_1076401;
  reg [7:0] p1_array_index_1076402;
  reg [7:0] p1_array_index_1076403;
  reg [7:0] p1_array_index_1076404;
  reg [7:0] p1_res7__2;
  reg [7:0] p1_array_index_1076414;
  reg [7:0] p1_array_index_1076415;
  reg [7:0] p1_array_index_1076416;
  reg [7:0] p1_array_index_1076417;
  reg [7:0] p1_array_index_1076418;
  reg [7:0] p1_res7__3;
  reg [7:0] p1_array_index_1076429;
  reg [7:0] p1_array_index_1076430;
  reg [7:0] p1_array_index_1076431;
  reg [7:0] p1_array_index_1076432;
  reg [7:0] p1_res7__4;
  reg [127:0] p1_bit_slice_1076440;
  reg [7:0] p1_array_index_1076455;
  reg [7:0] p1_array_index_1076456;
  reg [7:0] p1_array_index_1076457;
  reg [7:0] p1_array_index_1076458;
  reg [7:0] p1_array_index_1076459;
  reg [7:0] p1_array_index_1076460;
  reg [7:0] p1_array_index_1076462;
  reg [7:0] p1_array_index_1076464;
  reg [7:0] p1_array_index_1076465;
  reg [7:0] p1_array_index_1076471;
  reg [7:0] p1_array_index_1076472;
  reg [7:0] p1_array_index_1076473;
  reg [7:0] p1_array_index_1076474;
  reg [7:0] p1_array_index_1076475;
  reg [7:0] p1_array_index_1076477;
  reg [7:0] p1_array_index_1076479;
  reg [7:0] p1_res7__512;
  reg [7:0] p1_array_index_1076488;
  reg [7:0] p1_array_index_1076489;
  reg [7:0] p1_array_index_1076490;
  reg [7:0] p1_array_index_1076491;
  reg [7:0] p1_array_index_1076492;
  reg [7:0] p1_array_index_1076493;
  reg [7:0] p1_res7__513;
  reg [7:0] p1_array_index_1076503;
  reg [7:0] p1_array_index_1076504;
  reg [7:0] p1_array_index_1076505;
  reg [7:0] p1_array_index_1076506;
  reg [7:0] p1_array_index_1076507;
  reg [7:0] p1_res7__514;
  reg [7:0] p1_array_index_1076517;
  reg [7:0] p1_array_index_1076518;
  reg [7:0] p1_array_index_1076519;
  reg [7:0] p1_array_index_1076520;
  reg [7:0] p1_array_index_1076521;
  reg [7:0] p1_res7__515;
  reg [7:0] p1_array_index_1076532;
  reg [7:0] p1_array_index_1076533;
  reg [7:0] p1_array_index_1076534;
  reg [7:0] p1_array_index_1076535;
  reg [7:0] p1_res7__516;
  reg [7:0] p2_arr[256];
  reg [7:0] p2_literal_1076345[256];
  reg [7:0] p2_literal_1076347[256];
  reg [7:0] p2_literal_1076349[256];
  reg [7:0] p2_literal_1076351[256];
  reg [7:0] p2_literal_1076353[256];
  reg [7:0] p2_literal_1076355[256];
  reg [7:0] p2_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p1_bit_slice_1076328 <= p1_bit_slice_1076328_comb;
    p1_array_index_1076346 <= p1_array_index_1076346_comb;
    p1_array_index_1076348 <= p1_array_index_1076348_comb;
    p1_array_index_1076350 <= p1_array_index_1076350_comb;
    p1_array_index_1076352 <= p1_array_index_1076352_comb;
    p1_array_index_1076354 <= p1_array_index_1076354_comb;
    p1_array_index_1076356 <= p1_array_index_1076356_comb;
    p1_array_index_1076359 <= p1_array_index_1076359_comb;
    p1_array_index_1076361 <= p1_array_index_1076361_comb;
    p1_array_index_1076362 <= p1_array_index_1076362_comb;
    p1_array_index_1076368 <= p1_array_index_1076368_comb;
    p1_array_index_1076369 <= p1_array_index_1076369_comb;
    p1_array_index_1076370 <= p1_array_index_1076370_comb;
    p1_array_index_1076371 <= p1_array_index_1076371_comb;
    p1_array_index_1076372 <= p1_array_index_1076372_comb;
    p1_array_index_1076374 <= p1_array_index_1076374_comb;
    p1_array_index_1076376 <= p1_array_index_1076376_comb;
    p1_res7 <= p1_res7_comb;
    p1_array_index_1076385 <= p1_array_index_1076385_comb;
    p1_array_index_1076386 <= p1_array_index_1076386_comb;
    p1_array_index_1076387 <= p1_array_index_1076387_comb;
    p1_array_index_1076388 <= p1_array_index_1076388_comb;
    p1_array_index_1076389 <= p1_array_index_1076389_comb;
    p1_array_index_1076390 <= p1_array_index_1076390_comb;
    p1_res7__1 <= p1_res7__1_comb;
    p1_array_index_1076400 <= p1_array_index_1076400_comb;
    p1_array_index_1076401 <= p1_array_index_1076401_comb;
    p1_array_index_1076402 <= p1_array_index_1076402_comb;
    p1_array_index_1076403 <= p1_array_index_1076403_comb;
    p1_array_index_1076404 <= p1_array_index_1076404_comb;
    p1_res7__2 <= p1_res7__2_comb;
    p1_array_index_1076414 <= p1_array_index_1076414_comb;
    p1_array_index_1076415 <= p1_array_index_1076415_comb;
    p1_array_index_1076416 <= p1_array_index_1076416_comb;
    p1_array_index_1076417 <= p1_array_index_1076417_comb;
    p1_array_index_1076418 <= p1_array_index_1076418_comb;
    p1_res7__3 <= p1_res7__3_comb;
    p1_array_index_1076429 <= p1_array_index_1076429_comb;
    p1_array_index_1076430 <= p1_array_index_1076430_comb;
    p1_array_index_1076431 <= p1_array_index_1076431_comb;
    p1_array_index_1076432 <= p1_array_index_1076432_comb;
    p1_res7__4 <= p1_res7__4_comb;
    p1_bit_slice_1076440 <= p1_bit_slice_1076440_comb;
    p1_array_index_1076455 <= p1_array_index_1076455_comb;
    p1_array_index_1076456 <= p1_array_index_1076456_comb;
    p1_array_index_1076457 <= p1_array_index_1076457_comb;
    p1_array_index_1076458 <= p1_array_index_1076458_comb;
    p1_array_index_1076459 <= p1_array_index_1076459_comb;
    p1_array_index_1076460 <= p1_array_index_1076460_comb;
    p1_array_index_1076462 <= p1_array_index_1076462_comb;
    p1_array_index_1076464 <= p1_array_index_1076464_comb;
    p1_array_index_1076465 <= p1_array_index_1076465_comb;
    p1_array_index_1076471 <= p1_array_index_1076471_comb;
    p1_array_index_1076472 <= p1_array_index_1076472_comb;
    p1_array_index_1076473 <= p1_array_index_1076473_comb;
    p1_array_index_1076474 <= p1_array_index_1076474_comb;
    p1_array_index_1076475 <= p1_array_index_1076475_comb;
    p1_array_index_1076477 <= p1_array_index_1076477_comb;
    p1_array_index_1076479 <= p1_array_index_1076479_comb;
    p1_res7__512 <= p1_res7__512_comb;
    p1_array_index_1076488 <= p1_array_index_1076488_comb;
    p1_array_index_1076489 <= p1_array_index_1076489_comb;
    p1_array_index_1076490 <= p1_array_index_1076490_comb;
    p1_array_index_1076491 <= p1_array_index_1076491_comb;
    p1_array_index_1076492 <= p1_array_index_1076492_comb;
    p1_array_index_1076493 <= p1_array_index_1076493_comb;
    p1_res7__513 <= p1_res7__513_comb;
    p1_array_index_1076503 <= p1_array_index_1076503_comb;
    p1_array_index_1076504 <= p1_array_index_1076504_comb;
    p1_array_index_1076505 <= p1_array_index_1076505_comb;
    p1_array_index_1076506 <= p1_array_index_1076506_comb;
    p1_array_index_1076507 <= p1_array_index_1076507_comb;
    p1_res7__514 <= p1_res7__514_comb;
    p1_array_index_1076517 <= p1_array_index_1076517_comb;
    p1_array_index_1076518 <= p1_array_index_1076518_comb;
    p1_array_index_1076519 <= p1_array_index_1076519_comb;
    p1_array_index_1076520 <= p1_array_index_1076520_comb;
    p1_array_index_1076521 <= p1_array_index_1076521_comb;
    p1_res7__515 <= p1_res7__515_comb;
    p1_array_index_1076532 <= p1_array_index_1076532_comb;
    p1_array_index_1076533 <= p1_array_index_1076533_comb;
    p1_array_index_1076534 <= p1_array_index_1076534_comb;
    p1_array_index_1076535 <= p1_array_index_1076535_comb;
    p1_res7__516 <= p1_res7__516_comb;
    p2_arr <= p1_arr;
    p2_literal_1076345 <= p1_literal_1076345;
    p2_literal_1076347 <= p1_literal_1076347;
    p2_literal_1076349 <= p1_literal_1076349;
    p2_literal_1076351 <= p1_literal_1076351;
    p2_literal_1076353 <= p1_literal_1076353;
    p2_literal_1076355 <= p1_literal_1076355;
    p2_literal_1076358 <= p1_literal_1076358;
  end

  // ===== Pipe stage 2:
  wire [7:0] p2_array_index_1076729_comb;
  wire [7:0] p2_array_index_1076730_comb;
  wire [7:0] p2_array_index_1076731_comb;
  wire [7:0] p2_array_index_1076732_comb;
  wire [7:0] p2_array_index_1076797_comb;
  wire [7:0] p2_array_index_1076798_comb;
  wire [7:0] p2_array_index_1076799_comb;
  wire [7:0] p2_array_index_1076800_comb;
  wire [7:0] p2_res7__5_comb;
  wire [7:0] p2_res7__517_comb;
  wire [7:0] p2_array_index_1076743_comb;
  wire [7:0] p2_array_index_1076744_comb;
  wire [7:0] p2_array_index_1076745_comb;
  wire [7:0] p2_array_index_1076811_comb;
  wire [7:0] p2_array_index_1076812_comb;
  wire [7:0] p2_array_index_1076813_comb;
  wire [7:0] p2_res7__6_comb;
  wire [7:0] p2_res7__518_comb;
  wire [7:0] p2_array_index_1076755_comb;
  wire [7:0] p2_array_index_1076756_comb;
  wire [7:0] p2_array_index_1076757_comb;
  wire [7:0] p2_array_index_1076823_comb;
  wire [7:0] p2_array_index_1076824_comb;
  wire [7:0] p2_array_index_1076825_comb;
  wire [7:0] p2_res7__7_comb;
  wire [7:0] p2_res7__519_comb;
  wire [7:0] p2_array_index_1076768_comb;
  wire [7:0] p2_array_index_1076769_comb;
  wire [7:0] p2_array_index_1076836_comb;
  wire [7:0] p2_array_index_1076837_comb;
  wire [7:0] p2_res7__8_comb;
  wire [7:0] p2_res7__520_comb;
  wire [7:0] p2_array_index_1076779_comb;
  wire [7:0] p2_array_index_1076780_comb;
  wire [7:0] p2_array_index_1076847_comb;
  wire [7:0] p2_array_index_1076848_comb;
  wire [7:0] p2_res7__9_comb;
  wire [7:0] p2_res7__521_comb;
  wire [7:0] p2_array_index_1076786_comb;
  wire [7:0] p2_array_index_1076787_comb;
  wire [7:0] p2_array_index_1076788_comb;
  wire [7:0] p2_array_index_1076789_comb;
  wire [7:0] p2_array_index_1076790_comb;
  wire [7:0] p2_array_index_1076791_comb;
  wire [7:0] p2_array_index_1076792_comb;
  wire [7:0] p2_array_index_1076793_comb;
  wire [7:0] p2_array_index_1076794_comb;
  wire [7:0] p2_array_index_1076854_comb;
  wire [7:0] p2_array_index_1076855_comb;
  wire [7:0] p2_array_index_1076856_comb;
  wire [7:0] p2_array_index_1076857_comb;
  wire [7:0] p2_array_index_1076858_comb;
  wire [7:0] p2_array_index_1076859_comb;
  wire [7:0] p2_array_index_1076860_comb;
  wire [7:0] p2_array_index_1076861_comb;
  wire [7:0] p2_array_index_1076862_comb;
  assign p2_array_index_1076729_comb = p1_literal_1076349[p1_res7__2];
  assign p2_array_index_1076730_comb = p1_literal_1076351[p1_res7__1];
  assign p2_array_index_1076731_comb = p1_literal_1076353[p1_res7];
  assign p2_array_index_1076732_comb = p1_literal_1076355[p1_array_index_1076346];
  assign p2_array_index_1076797_comb = p1_literal_1076349[p1_res7__514];
  assign p2_array_index_1076798_comb = p1_literal_1076351[p1_res7__513];
  assign p2_array_index_1076799_comb = p1_literal_1076353[p1_res7__512];
  assign p2_array_index_1076800_comb = p1_literal_1076355[p1_array_index_1076455];
  assign p2_res7__5_comb = p1_literal_1076345[p1_res7__4] ^ p1_literal_1076347[p1_res7__3] ^ p2_array_index_1076729_comb ^ p2_array_index_1076730_comb ^ p2_array_index_1076731_comb ^ p2_array_index_1076732_comb ^ p1_array_index_1076348 ^ p1_literal_1076358[p1_array_index_1076350] ^ p1_array_index_1076352 ^ p1_array_index_1076390 ^ p1_literal_1076353[p1_array_index_1076356] ^ p1_literal_1076351[p1_array_index_1076374] ^ p1_literal_1076349[p1_array_index_1076359] ^ p1_literal_1076347[p1_array_index_1076376] ^ p1_literal_1076345[p1_array_index_1076361] ^ p1_array_index_1076362;
  assign p2_res7__517_comb = p1_literal_1076345[p1_res7__516] ^ p1_literal_1076347[p1_res7__515] ^ p2_array_index_1076797_comb ^ p2_array_index_1076798_comb ^ p2_array_index_1076799_comb ^ p2_array_index_1076800_comb ^ p1_array_index_1076456 ^ p1_literal_1076358[p1_array_index_1076457] ^ p1_array_index_1076458 ^ p1_array_index_1076493 ^ p1_literal_1076353[p1_array_index_1076460] ^ p1_literal_1076351[p1_array_index_1076477] ^ p1_literal_1076349[p1_array_index_1076462] ^ p1_literal_1076347[p1_array_index_1076479] ^ p1_literal_1076345[p1_array_index_1076464] ^ p1_array_index_1076465;
  assign p2_array_index_1076743_comb = p1_literal_1076351[p1_res7__2];
  assign p2_array_index_1076744_comb = p1_literal_1076353[p1_res7__1];
  assign p2_array_index_1076745_comb = p1_literal_1076355[p1_res7];
  assign p2_array_index_1076811_comb = p1_literal_1076351[p1_res7__514];
  assign p2_array_index_1076812_comb = p1_literal_1076353[p1_res7__513];
  assign p2_array_index_1076813_comb = p1_literal_1076355[p1_res7__512];
  assign p2_res7__6_comb = p1_literal_1076345[p2_res7__5_comb] ^ p1_literal_1076347[p1_res7__4] ^ p1_literal_1076349[p1_res7__3] ^ p2_array_index_1076743_comb ^ p2_array_index_1076744_comb ^ p2_array_index_1076745_comb ^ p1_array_index_1076346 ^ p1_literal_1076358[p1_array_index_1076348] ^ p1_array_index_1076350 ^ p1_array_index_1076404 ^ p1_array_index_1076372 ^ p1_literal_1076351[p1_array_index_1076356] ^ p1_literal_1076349[p1_array_index_1076374] ^ p1_literal_1076347[p1_array_index_1076359] ^ p1_literal_1076345[p1_array_index_1076376] ^ p1_array_index_1076361;
  assign p2_res7__518_comb = p1_literal_1076345[p2_res7__517_comb] ^ p1_literal_1076347[p1_res7__516] ^ p1_literal_1076349[p1_res7__515] ^ p2_array_index_1076811_comb ^ p2_array_index_1076812_comb ^ p2_array_index_1076813_comb ^ p1_array_index_1076455 ^ p1_literal_1076358[p1_array_index_1076456] ^ p1_array_index_1076457 ^ p1_array_index_1076507 ^ p1_array_index_1076475 ^ p1_literal_1076351[p1_array_index_1076460] ^ p1_literal_1076349[p1_array_index_1076477] ^ p1_literal_1076347[p1_array_index_1076462] ^ p1_literal_1076345[p1_array_index_1076479] ^ p1_array_index_1076464;
  assign p2_array_index_1076755_comb = p1_literal_1076351[p1_res7__3];
  assign p2_array_index_1076756_comb = p1_literal_1076353[p1_res7__2];
  assign p2_array_index_1076757_comb = p1_literal_1076355[p1_res7__1];
  assign p2_array_index_1076823_comb = p1_literal_1076351[p1_res7__515];
  assign p2_array_index_1076824_comb = p1_literal_1076353[p1_res7__514];
  assign p2_array_index_1076825_comb = p1_literal_1076355[p1_res7__513];
  assign p2_res7__7_comb = p1_literal_1076345[p2_res7__6_comb] ^ p1_literal_1076347[p2_res7__5_comb] ^ p1_literal_1076349[p1_res7__4] ^ p2_array_index_1076755_comb ^ p2_array_index_1076756_comb ^ p2_array_index_1076757_comb ^ p1_res7 ^ p1_literal_1076358[p1_array_index_1076346] ^ p1_array_index_1076348 ^ p1_array_index_1076418 ^ p1_array_index_1076389 ^ p1_literal_1076351[p1_array_index_1076354] ^ p1_literal_1076349[p1_array_index_1076356] ^ p1_literal_1076347[p1_array_index_1076374] ^ p1_literal_1076345[p1_array_index_1076359] ^ p1_array_index_1076376;
  assign p2_res7__519_comb = p1_literal_1076345[p2_res7__518_comb] ^ p1_literal_1076347[p2_res7__517_comb] ^ p1_literal_1076349[p1_res7__516] ^ p2_array_index_1076823_comb ^ p2_array_index_1076824_comb ^ p2_array_index_1076825_comb ^ p1_res7__512 ^ p1_literal_1076358[p1_array_index_1076455] ^ p1_array_index_1076456 ^ p1_array_index_1076521 ^ p1_array_index_1076492 ^ p1_literal_1076351[p1_array_index_1076459] ^ p1_literal_1076349[p1_array_index_1076460] ^ p1_literal_1076347[p1_array_index_1076477] ^ p1_literal_1076345[p1_array_index_1076462] ^ p1_array_index_1076479;
  assign p2_array_index_1076768_comb = p1_literal_1076353[p1_res7__3];
  assign p2_array_index_1076769_comb = p1_literal_1076355[p1_res7__2];
  assign p2_array_index_1076836_comb = p1_literal_1076353[p1_res7__515];
  assign p2_array_index_1076837_comb = p1_literal_1076355[p1_res7__514];
  assign p2_res7__8_comb = p1_literal_1076345[p2_res7__7_comb] ^ p1_literal_1076347[p2_res7__6_comb] ^ p1_literal_1076349[p2_res7__5_comb] ^ p1_literal_1076351[p1_res7__4] ^ p2_array_index_1076768_comb ^ p2_array_index_1076769_comb ^ p1_res7__1 ^ p1_literal_1076358[p1_res7] ^ p1_array_index_1076346 ^ p1_array_index_1076432 ^ p1_array_index_1076403 ^ p1_array_index_1076371 ^ p1_literal_1076349[p1_array_index_1076354] ^ p1_literal_1076347[p1_array_index_1076356] ^ p1_literal_1076345[p1_array_index_1076374] ^ p1_array_index_1076359;
  assign p2_res7__520_comb = p1_literal_1076345[p2_res7__519_comb] ^ p1_literal_1076347[p2_res7__518_comb] ^ p1_literal_1076349[p2_res7__517_comb] ^ p1_literal_1076351[p1_res7__516] ^ p2_array_index_1076836_comb ^ p2_array_index_1076837_comb ^ p1_res7__513 ^ p1_literal_1076358[p1_res7__512] ^ p1_array_index_1076455 ^ p1_array_index_1076535 ^ p1_array_index_1076506 ^ p1_array_index_1076474 ^ p1_literal_1076349[p1_array_index_1076459] ^ p1_literal_1076347[p1_array_index_1076460] ^ p1_literal_1076345[p1_array_index_1076477] ^ p1_array_index_1076462;
  assign p2_array_index_1076779_comb = p1_literal_1076353[p1_res7__4];
  assign p2_array_index_1076780_comb = p1_literal_1076355[p1_res7__3];
  assign p2_array_index_1076847_comb = p1_literal_1076353[p1_res7__516];
  assign p2_array_index_1076848_comb = p1_literal_1076355[p1_res7__515];
  assign p2_res7__9_comb = p1_literal_1076345[p2_res7__8_comb] ^ p1_literal_1076347[p2_res7__7_comb] ^ p1_literal_1076349[p2_res7__6_comb] ^ p1_literal_1076351[p2_res7__5_comb] ^ p2_array_index_1076779_comb ^ p2_array_index_1076780_comb ^ p1_res7__2 ^ p1_literal_1076358[p1_res7__1] ^ p1_res7 ^ p2_array_index_1076732_comb ^ p1_array_index_1076417 ^ p1_array_index_1076388 ^ p1_literal_1076349[p1_array_index_1076352] ^ p1_literal_1076347[p1_array_index_1076354] ^ p1_literal_1076345[p1_array_index_1076356] ^ p1_array_index_1076374;
  assign p2_res7__521_comb = p1_literal_1076345[p2_res7__520_comb] ^ p1_literal_1076347[p2_res7__519_comb] ^ p1_literal_1076349[p2_res7__518_comb] ^ p1_literal_1076351[p2_res7__517_comb] ^ p2_array_index_1076847_comb ^ p2_array_index_1076848_comb ^ p1_res7__514 ^ p1_literal_1076358[p1_res7__513] ^ p1_res7__512 ^ p2_array_index_1076800_comb ^ p1_array_index_1076520 ^ p1_array_index_1076491 ^ p1_literal_1076349[p1_array_index_1076458] ^ p1_literal_1076347[p1_array_index_1076459] ^ p1_literal_1076345[p1_array_index_1076460] ^ p1_array_index_1076477;
  assign p2_array_index_1076786_comb = p1_literal_1076345[p2_res7__9_comb];
  assign p2_array_index_1076787_comb = p1_literal_1076347[p2_res7__8_comb];
  assign p2_array_index_1076788_comb = p1_literal_1076349[p2_res7__7_comb];
  assign p2_array_index_1076789_comb = p1_literal_1076351[p2_res7__6_comb];
  assign p2_array_index_1076790_comb = p1_literal_1076353[p2_res7__5_comb];
  assign p2_array_index_1076791_comb = p1_literal_1076355[p1_res7__4];
  assign p2_array_index_1076792_comb = p1_literal_1076358[p1_res7__2];
  assign p2_array_index_1076793_comb = p1_literal_1076347[p1_array_index_1076352];
  assign p2_array_index_1076794_comb = p1_literal_1076345[p1_array_index_1076354];
  assign p2_array_index_1076854_comb = p1_literal_1076345[p2_res7__521_comb];
  assign p2_array_index_1076855_comb = p1_literal_1076347[p2_res7__520_comb];
  assign p2_array_index_1076856_comb = p1_literal_1076349[p2_res7__519_comb];
  assign p2_array_index_1076857_comb = p1_literal_1076351[p2_res7__518_comb];
  assign p2_array_index_1076858_comb = p1_literal_1076353[p2_res7__517_comb];
  assign p2_array_index_1076859_comb = p1_literal_1076355[p1_res7__516];
  assign p2_array_index_1076860_comb = p1_literal_1076358[p1_res7__514];
  assign p2_array_index_1076861_comb = p1_literal_1076347[p1_array_index_1076458];
  assign p2_array_index_1076862_comb = p1_literal_1076345[p1_array_index_1076459];

  // Registers for pipe stage 2:
  reg [127:0] p2_bit_slice_1076328;
  reg [7:0] p2_array_index_1076346;
  reg [7:0] p2_array_index_1076348;
  reg [7:0] p2_array_index_1076350;
  reg [7:0] p2_array_index_1076352;
  reg [7:0] p2_array_index_1076354;
  reg [7:0] p2_array_index_1076356;
  reg [7:0] p2_array_index_1076368;
  reg [7:0] p2_array_index_1076369;
  reg [7:0] p2_array_index_1076370;
  reg [7:0] p2_res7;
  reg [7:0] p2_array_index_1076385;
  reg [7:0] p2_array_index_1076386;
  reg [7:0] p2_array_index_1076387;
  reg [7:0] p2_res7__1;
  reg [7:0] p2_array_index_1076400;
  reg [7:0] p2_array_index_1076401;
  reg [7:0] p2_array_index_1076402;
  reg [7:0] p2_res7__2;
  reg [7:0] p2_array_index_1076414;
  reg [7:0] p2_array_index_1076415;
  reg [7:0] p2_array_index_1076416;
  reg [7:0] p2_res7__3;
  reg [7:0] p2_array_index_1076429;
  reg [7:0] p2_array_index_1076430;
  reg [7:0] p2_array_index_1076431;
  reg [7:0] p2_res7__4;
  reg [7:0] p2_array_index_1076729;
  reg [7:0] p2_array_index_1076730;
  reg [7:0] p2_array_index_1076731;
  reg [7:0] p2_res7__5;
  reg [7:0] p2_array_index_1076743;
  reg [7:0] p2_array_index_1076744;
  reg [7:0] p2_array_index_1076745;
  reg [7:0] p2_res7__6;
  reg [7:0] p2_array_index_1076755;
  reg [7:0] p2_array_index_1076756;
  reg [7:0] p2_array_index_1076757;
  reg [7:0] p2_res7__7;
  reg [7:0] p2_array_index_1076768;
  reg [7:0] p2_array_index_1076769;
  reg [7:0] p2_res7__8;
  reg [7:0] p2_array_index_1076779;
  reg [7:0] p2_array_index_1076780;
  reg [7:0] p2_res7__9;
  reg [7:0] p2_array_index_1076786;
  reg [7:0] p2_array_index_1076787;
  reg [7:0] p2_array_index_1076788;
  reg [7:0] p2_array_index_1076789;
  reg [7:0] p2_array_index_1076790;
  reg [7:0] p2_array_index_1076791;
  reg [7:0] p2_array_index_1076792;
  reg [7:0] p2_array_index_1076793;
  reg [7:0] p2_array_index_1076794;
  reg [127:0] p2_bit_slice_1076440;
  reg [7:0] p2_array_index_1076455;
  reg [7:0] p2_array_index_1076456;
  reg [7:0] p2_array_index_1076457;
  reg [7:0] p2_array_index_1076458;
  reg [7:0] p2_array_index_1076459;
  reg [7:0] p2_array_index_1076460;
  reg [7:0] p2_array_index_1076471;
  reg [7:0] p2_array_index_1076472;
  reg [7:0] p2_array_index_1076473;
  reg [7:0] p2_res7__512;
  reg [7:0] p2_array_index_1076488;
  reg [7:0] p2_array_index_1076489;
  reg [7:0] p2_array_index_1076490;
  reg [7:0] p2_res7__513;
  reg [7:0] p2_array_index_1076503;
  reg [7:0] p2_array_index_1076504;
  reg [7:0] p2_array_index_1076505;
  reg [7:0] p2_res7__514;
  reg [7:0] p2_array_index_1076517;
  reg [7:0] p2_array_index_1076518;
  reg [7:0] p2_array_index_1076519;
  reg [7:0] p2_res7__515;
  reg [7:0] p2_array_index_1076532;
  reg [7:0] p2_array_index_1076533;
  reg [7:0] p2_array_index_1076534;
  reg [7:0] p2_res7__516;
  reg [7:0] p2_array_index_1076797;
  reg [7:0] p2_array_index_1076798;
  reg [7:0] p2_array_index_1076799;
  reg [7:0] p2_res7__517;
  reg [7:0] p2_array_index_1076811;
  reg [7:0] p2_array_index_1076812;
  reg [7:0] p2_array_index_1076813;
  reg [7:0] p2_res7__518;
  reg [7:0] p2_array_index_1076823;
  reg [7:0] p2_array_index_1076824;
  reg [7:0] p2_array_index_1076825;
  reg [7:0] p2_res7__519;
  reg [7:0] p2_array_index_1076836;
  reg [7:0] p2_array_index_1076837;
  reg [7:0] p2_res7__520;
  reg [7:0] p2_array_index_1076847;
  reg [7:0] p2_array_index_1076848;
  reg [7:0] p2_res7__521;
  reg [7:0] p2_array_index_1076854;
  reg [7:0] p2_array_index_1076855;
  reg [7:0] p2_array_index_1076856;
  reg [7:0] p2_array_index_1076857;
  reg [7:0] p2_array_index_1076858;
  reg [7:0] p2_array_index_1076859;
  reg [7:0] p2_array_index_1076860;
  reg [7:0] p2_array_index_1076861;
  reg [7:0] p2_array_index_1076862;
  reg [7:0] p3_arr[256];
  reg [7:0] p3_literal_1076345[256];
  reg [7:0] p3_literal_1076347[256];
  reg [7:0] p3_literal_1076349[256];
  reg [7:0] p3_literal_1076351[256];
  reg [7:0] p3_literal_1076353[256];
  reg [7:0] p3_literal_1076355[256];
  reg [7:0] p3_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p2_bit_slice_1076328 <= p1_bit_slice_1076328;
    p2_array_index_1076346 <= p1_array_index_1076346;
    p2_array_index_1076348 <= p1_array_index_1076348;
    p2_array_index_1076350 <= p1_array_index_1076350;
    p2_array_index_1076352 <= p1_array_index_1076352;
    p2_array_index_1076354 <= p1_array_index_1076354;
    p2_array_index_1076356 <= p1_array_index_1076356;
    p2_array_index_1076368 <= p1_array_index_1076368;
    p2_array_index_1076369 <= p1_array_index_1076369;
    p2_array_index_1076370 <= p1_array_index_1076370;
    p2_res7 <= p1_res7;
    p2_array_index_1076385 <= p1_array_index_1076385;
    p2_array_index_1076386 <= p1_array_index_1076386;
    p2_array_index_1076387 <= p1_array_index_1076387;
    p2_res7__1 <= p1_res7__1;
    p2_array_index_1076400 <= p1_array_index_1076400;
    p2_array_index_1076401 <= p1_array_index_1076401;
    p2_array_index_1076402 <= p1_array_index_1076402;
    p2_res7__2 <= p1_res7__2;
    p2_array_index_1076414 <= p1_array_index_1076414;
    p2_array_index_1076415 <= p1_array_index_1076415;
    p2_array_index_1076416 <= p1_array_index_1076416;
    p2_res7__3 <= p1_res7__3;
    p2_array_index_1076429 <= p1_array_index_1076429;
    p2_array_index_1076430 <= p1_array_index_1076430;
    p2_array_index_1076431 <= p1_array_index_1076431;
    p2_res7__4 <= p1_res7__4;
    p2_array_index_1076729 <= p2_array_index_1076729_comb;
    p2_array_index_1076730 <= p2_array_index_1076730_comb;
    p2_array_index_1076731 <= p2_array_index_1076731_comb;
    p2_res7__5 <= p2_res7__5_comb;
    p2_array_index_1076743 <= p2_array_index_1076743_comb;
    p2_array_index_1076744 <= p2_array_index_1076744_comb;
    p2_array_index_1076745 <= p2_array_index_1076745_comb;
    p2_res7__6 <= p2_res7__6_comb;
    p2_array_index_1076755 <= p2_array_index_1076755_comb;
    p2_array_index_1076756 <= p2_array_index_1076756_comb;
    p2_array_index_1076757 <= p2_array_index_1076757_comb;
    p2_res7__7 <= p2_res7__7_comb;
    p2_array_index_1076768 <= p2_array_index_1076768_comb;
    p2_array_index_1076769 <= p2_array_index_1076769_comb;
    p2_res7__8 <= p2_res7__8_comb;
    p2_array_index_1076779 <= p2_array_index_1076779_comb;
    p2_array_index_1076780 <= p2_array_index_1076780_comb;
    p2_res7__9 <= p2_res7__9_comb;
    p2_array_index_1076786 <= p2_array_index_1076786_comb;
    p2_array_index_1076787 <= p2_array_index_1076787_comb;
    p2_array_index_1076788 <= p2_array_index_1076788_comb;
    p2_array_index_1076789 <= p2_array_index_1076789_comb;
    p2_array_index_1076790 <= p2_array_index_1076790_comb;
    p2_array_index_1076791 <= p2_array_index_1076791_comb;
    p2_array_index_1076792 <= p2_array_index_1076792_comb;
    p2_array_index_1076793 <= p2_array_index_1076793_comb;
    p2_array_index_1076794 <= p2_array_index_1076794_comb;
    p2_bit_slice_1076440 <= p1_bit_slice_1076440;
    p2_array_index_1076455 <= p1_array_index_1076455;
    p2_array_index_1076456 <= p1_array_index_1076456;
    p2_array_index_1076457 <= p1_array_index_1076457;
    p2_array_index_1076458 <= p1_array_index_1076458;
    p2_array_index_1076459 <= p1_array_index_1076459;
    p2_array_index_1076460 <= p1_array_index_1076460;
    p2_array_index_1076471 <= p1_array_index_1076471;
    p2_array_index_1076472 <= p1_array_index_1076472;
    p2_array_index_1076473 <= p1_array_index_1076473;
    p2_res7__512 <= p1_res7__512;
    p2_array_index_1076488 <= p1_array_index_1076488;
    p2_array_index_1076489 <= p1_array_index_1076489;
    p2_array_index_1076490 <= p1_array_index_1076490;
    p2_res7__513 <= p1_res7__513;
    p2_array_index_1076503 <= p1_array_index_1076503;
    p2_array_index_1076504 <= p1_array_index_1076504;
    p2_array_index_1076505 <= p1_array_index_1076505;
    p2_res7__514 <= p1_res7__514;
    p2_array_index_1076517 <= p1_array_index_1076517;
    p2_array_index_1076518 <= p1_array_index_1076518;
    p2_array_index_1076519 <= p1_array_index_1076519;
    p2_res7__515 <= p1_res7__515;
    p2_array_index_1076532 <= p1_array_index_1076532;
    p2_array_index_1076533 <= p1_array_index_1076533;
    p2_array_index_1076534 <= p1_array_index_1076534;
    p2_res7__516 <= p1_res7__516;
    p2_array_index_1076797 <= p2_array_index_1076797_comb;
    p2_array_index_1076798 <= p2_array_index_1076798_comb;
    p2_array_index_1076799 <= p2_array_index_1076799_comb;
    p2_res7__517 <= p2_res7__517_comb;
    p2_array_index_1076811 <= p2_array_index_1076811_comb;
    p2_array_index_1076812 <= p2_array_index_1076812_comb;
    p2_array_index_1076813 <= p2_array_index_1076813_comb;
    p2_res7__518 <= p2_res7__518_comb;
    p2_array_index_1076823 <= p2_array_index_1076823_comb;
    p2_array_index_1076824 <= p2_array_index_1076824_comb;
    p2_array_index_1076825 <= p2_array_index_1076825_comb;
    p2_res7__519 <= p2_res7__519_comb;
    p2_array_index_1076836 <= p2_array_index_1076836_comb;
    p2_array_index_1076837 <= p2_array_index_1076837_comb;
    p2_res7__520 <= p2_res7__520_comb;
    p2_array_index_1076847 <= p2_array_index_1076847_comb;
    p2_array_index_1076848 <= p2_array_index_1076848_comb;
    p2_res7__521 <= p2_res7__521_comb;
    p2_array_index_1076854 <= p2_array_index_1076854_comb;
    p2_array_index_1076855 <= p2_array_index_1076855_comb;
    p2_array_index_1076856 <= p2_array_index_1076856_comb;
    p2_array_index_1076857 <= p2_array_index_1076857_comb;
    p2_array_index_1076858 <= p2_array_index_1076858_comb;
    p2_array_index_1076859 <= p2_array_index_1076859_comb;
    p2_array_index_1076860 <= p2_array_index_1076860_comb;
    p2_array_index_1076861 <= p2_array_index_1076861_comb;
    p2_array_index_1076862 <= p2_array_index_1076862_comb;
    p3_arr <= p2_arr;
    p3_literal_1076345 <= p2_literal_1076345;
    p3_literal_1076347 <= p2_literal_1076347;
    p3_literal_1076349 <= p2_literal_1076349;
    p3_literal_1076351 <= p2_literal_1076351;
    p3_literal_1076353 <= p2_literal_1076353;
    p3_literal_1076355 <= p2_literal_1076355;
    p3_literal_1076358 <= p2_literal_1076358;
  end

  // ===== Pipe stage 3:
  wire [7:0] p3_res7__522_comb;
  wire [7:0] p3_res7__10_comb;
  wire [7:0] p3_array_index_1077148_comb;
  wire [7:0] p3_array_index_1077101_comb;
  wire [7:0] p3_res7__523_comb;
  wire [7:0] p3_res7__11_comb;
  wire [7:0] p3_res7__524_comb;
  wire [7:0] p3_res7__12_comb;
  wire [7:0] p3_res7__525_comb;
  wire [7:0] p3_res7__13_comb;
  wire [7:0] p3_res7__526_comb;
  wire [7:0] p3_res7__14_comb;
  wire [7:0] p3_res7__527_comb;
  wire [7:0] p3_res7__15_comb;
  wire [127:0] p3_res__32_comb;
  wire [127:0] p3_res_comb;
  wire [127:0] p3_addedKey__33_comb;
  wire [127:0] p3_xor_1077141_comb;
  wire [7:0] p3_bit_slice_1077189_comb;
  wire [7:0] p3_bit_slice_1077190_comb;
  wire [7:0] p3_bit_slice_1077191_comb;
  wire [7:0] p3_bit_slice_1077192_comb;
  wire [7:0] p3_bit_slice_1077193_comb;
  wire [7:0] p3_bit_slice_1077194_comb;
  wire [7:0] p3_bit_slice_1077195_comb;
  wire [7:0] p3_bit_slice_1077196_comb;
  wire [7:0] p3_bit_slice_1077197_comb;
  wire [7:0] p3_bit_slice_1077198_comb;
  wire [7:0] p3_bit_slice_1077199_comb;
  wire [7:0] p3_bit_slice_1077200_comb;
  wire [7:0] p3_bit_slice_1077201_comb;
  wire [7:0] p3_bit_slice_1077202_comb;
  wire [7:0] p3_bit_slice_1077203_comb;
  wire [7:0] p3_bit_slice_1077204_comb;
  assign p3_res7__522_comb = p2_array_index_1076854 ^ p2_array_index_1076855 ^ p2_array_index_1076856 ^ p2_array_index_1076857 ^ p2_array_index_1076858 ^ p2_array_index_1076859 ^ p2_res7__515 ^ p2_array_index_1076860 ^ p2_res7__513 ^ p2_array_index_1076813 ^ p2_array_index_1076534 ^ p2_array_index_1076505 ^ p2_array_index_1076473 ^ p2_array_index_1076861 ^ p2_array_index_1076862 ^ p2_array_index_1076460;
  assign p3_res7__10_comb = p2_array_index_1076786 ^ p2_array_index_1076787 ^ p2_array_index_1076788 ^ p2_array_index_1076789 ^ p2_array_index_1076790 ^ p2_array_index_1076791 ^ p2_res7__3 ^ p2_array_index_1076792 ^ p2_res7__1 ^ p2_array_index_1076745 ^ p2_array_index_1076431 ^ p2_array_index_1076402 ^ p2_array_index_1076370 ^ p2_array_index_1076793 ^ p2_array_index_1076794 ^ p2_array_index_1076356;
  assign p3_array_index_1077148_comb = p2_literal_1076355[p2_res7__517];
  assign p3_array_index_1077101_comb = p2_literal_1076355[p2_res7__5];
  assign p3_res7__523_comb = p2_literal_1076345[p3_res7__522_comb] ^ p2_literal_1076347[p2_res7__521] ^ p2_literal_1076349[p2_res7__520] ^ p2_literal_1076351[p2_res7__519] ^ p2_literal_1076353[p2_res7__518] ^ p3_array_index_1077148_comb ^ p2_res7__516 ^ p2_literal_1076358[p2_res7__515] ^ p2_res7__514 ^ p2_array_index_1076825 ^ p2_array_index_1076799 ^ p2_array_index_1076519 ^ p2_array_index_1076490 ^ p2_literal_1076347[p2_array_index_1076457] ^ p2_literal_1076345[p2_array_index_1076458] ^ p2_array_index_1076459;
  assign p3_res7__11_comb = p2_literal_1076345[p3_res7__10_comb] ^ p2_literal_1076347[p2_res7__9] ^ p2_literal_1076349[p2_res7__8] ^ p2_literal_1076351[p2_res7__7] ^ p2_literal_1076353[p2_res7__6] ^ p3_array_index_1077101_comb ^ p2_res7__4 ^ p2_literal_1076358[p2_res7__3] ^ p2_res7__2 ^ p2_array_index_1076757 ^ p2_array_index_1076731 ^ p2_array_index_1076416 ^ p2_array_index_1076387 ^ p2_literal_1076347[p2_array_index_1076350] ^ p2_literal_1076345[p2_array_index_1076352] ^ p2_array_index_1076354;
  assign p3_res7__524_comb = p2_literal_1076345[p3_res7__523_comb] ^ p2_literal_1076347[p3_res7__522_comb] ^ p2_literal_1076349[p2_res7__521] ^ p2_literal_1076351[p2_res7__520] ^ p2_literal_1076353[p2_res7__519] ^ p2_literal_1076355[p2_res7__518] ^ p2_res7__517 ^ p2_literal_1076358[p2_res7__516] ^ p2_res7__515 ^ p2_array_index_1076837 ^ p2_array_index_1076812 ^ p2_array_index_1076533 ^ p2_array_index_1076504 ^ p2_array_index_1076472 ^ p2_literal_1076345[p2_array_index_1076457] ^ p2_array_index_1076458;
  assign p3_res7__12_comb = p2_literal_1076345[p3_res7__11_comb] ^ p2_literal_1076347[p3_res7__10_comb] ^ p2_literal_1076349[p2_res7__9] ^ p2_literal_1076351[p2_res7__8] ^ p2_literal_1076353[p2_res7__7] ^ p2_literal_1076355[p2_res7__6] ^ p2_res7__5 ^ p2_literal_1076358[p2_res7__4] ^ p2_res7__3 ^ p2_array_index_1076769 ^ p2_array_index_1076744 ^ p2_array_index_1076430 ^ p2_array_index_1076401 ^ p2_array_index_1076369 ^ p2_literal_1076345[p2_array_index_1076350] ^ p2_array_index_1076352;
  assign p3_res7__525_comb = p2_literal_1076345[p3_res7__524_comb] ^ p2_literal_1076347[p3_res7__523_comb] ^ p2_literal_1076349[p3_res7__522_comb] ^ p2_literal_1076351[p2_res7__521] ^ p2_literal_1076353[p2_res7__520] ^ p2_literal_1076355[p2_res7__519] ^ p2_res7__518 ^ p2_literal_1076358[p2_res7__517] ^ p2_res7__516 ^ p2_array_index_1076848 ^ p2_array_index_1076824 ^ p2_array_index_1076798 ^ p2_array_index_1076518 ^ p2_array_index_1076489 ^ p2_literal_1076345[p2_array_index_1076456] ^ p2_array_index_1076457;
  assign p3_res7__13_comb = p2_literal_1076345[p3_res7__12_comb] ^ p2_literal_1076347[p3_res7__11_comb] ^ p2_literal_1076349[p3_res7__10_comb] ^ p2_literal_1076351[p2_res7__9] ^ p2_literal_1076353[p2_res7__8] ^ p2_literal_1076355[p2_res7__7] ^ p2_res7__6 ^ p2_literal_1076358[p2_res7__5] ^ p2_res7__4 ^ p2_array_index_1076780 ^ p2_array_index_1076756 ^ p2_array_index_1076730 ^ p2_array_index_1076415 ^ p2_array_index_1076386 ^ p2_literal_1076345[p2_array_index_1076348] ^ p2_array_index_1076350;
  assign p3_res7__526_comb = p2_literal_1076345[p3_res7__525_comb] ^ p2_literal_1076347[p3_res7__524_comb] ^ p2_literal_1076349[p3_res7__523_comb] ^ p2_literal_1076351[p3_res7__522_comb] ^ p2_literal_1076353[p2_res7__521] ^ p2_literal_1076355[p2_res7__520] ^ p2_res7__519 ^ p2_literal_1076358[p2_res7__518] ^ p2_res7__517 ^ p2_array_index_1076859 ^ p2_array_index_1076836 ^ p2_array_index_1076811 ^ p2_array_index_1076532 ^ p2_array_index_1076503 ^ p2_array_index_1076471 ^ p2_array_index_1076456;
  assign p3_res7__14_comb = p2_literal_1076345[p3_res7__13_comb] ^ p2_literal_1076347[p3_res7__12_comb] ^ p2_literal_1076349[p3_res7__11_comb] ^ p2_literal_1076351[p3_res7__10_comb] ^ p2_literal_1076353[p2_res7__9] ^ p2_literal_1076355[p2_res7__8] ^ p2_res7__7 ^ p2_literal_1076358[p2_res7__6] ^ p2_res7__5 ^ p2_array_index_1076791 ^ p2_array_index_1076768 ^ p2_array_index_1076743 ^ p2_array_index_1076429 ^ p2_array_index_1076400 ^ p2_array_index_1076368 ^ p2_array_index_1076348;
  assign p3_res7__527_comb = p2_literal_1076345[p3_res7__526_comb] ^ p2_literal_1076347[p3_res7__525_comb] ^ p2_literal_1076349[p3_res7__524_comb] ^ p2_literal_1076351[p3_res7__523_comb] ^ p2_literal_1076353[p3_res7__522_comb] ^ p2_literal_1076355[p2_res7__521] ^ p2_res7__520 ^ p2_literal_1076358[p2_res7__519] ^ p2_res7__518 ^ p3_array_index_1077148_comb ^ p2_array_index_1076847 ^ p2_array_index_1076823 ^ p2_array_index_1076797 ^ p2_array_index_1076517 ^ p2_array_index_1076488 ^ p2_array_index_1076455;
  assign p3_res7__15_comb = p2_literal_1076345[p3_res7__14_comb] ^ p2_literal_1076347[p3_res7__13_comb] ^ p2_literal_1076349[p3_res7__12_comb] ^ p2_literal_1076351[p3_res7__11_comb] ^ p2_literal_1076353[p3_res7__10_comb] ^ p2_literal_1076355[p2_res7__9] ^ p2_res7__8 ^ p2_literal_1076358[p2_res7__7] ^ p2_res7__6 ^ p3_array_index_1077101_comb ^ p2_array_index_1076779 ^ p2_array_index_1076755 ^ p2_array_index_1076729 ^ p2_array_index_1076414 ^ p2_array_index_1076385 ^ p2_array_index_1076346;
  assign p3_res__32_comb = {p3_res7__527_comb, p3_res7__526_comb, p3_res7__525_comb, p3_res7__524_comb, p3_res7__523_comb, p3_res7__522_comb, p2_res7__521, p2_res7__520, p2_res7__519, p2_res7__518, p2_res7__517, p2_res7__516, p2_res7__515, p2_res7__514, p2_res7__513, p2_res7__512};
  assign p3_res_comb = {p3_res7__15_comb, p3_res7__14_comb, p3_res7__13_comb, p3_res7__12_comb, p3_res7__11_comb, p3_res7__10_comb, p2_res7__9, p2_res7__8, p2_res7__7, p2_res7__6, p2_res7__5, p2_res7__4, p2_res7__3, p2_res7__2, p2_res7__1, p2_res7};
  assign p3_addedKey__33_comb = p2_bit_slice_1076440 ^ p3_res__32_comb;
  assign p3_xor_1077141_comb = p3_res_comb ^ p2_bit_slice_1076440;
  assign p3_bit_slice_1077189_comb = p3_addedKey__33_comb[127:120];
  assign p3_bit_slice_1077190_comb = p3_addedKey__33_comb[119:112];
  assign p3_bit_slice_1077191_comb = p3_addedKey__33_comb[111:104];
  assign p3_bit_slice_1077192_comb = p3_addedKey__33_comb[103:96];
  assign p3_bit_slice_1077193_comb = p3_addedKey__33_comb[95:88];
  assign p3_bit_slice_1077194_comb = p3_addedKey__33_comb[87:80];
  assign p3_bit_slice_1077195_comb = p3_addedKey__33_comb[71:64];
  assign p3_bit_slice_1077196_comb = p3_addedKey__33_comb[55:48];
  assign p3_bit_slice_1077197_comb = p3_addedKey__33_comb[47:40];
  assign p3_bit_slice_1077198_comb = p3_addedKey__33_comb[39:32];
  assign p3_bit_slice_1077199_comb = p3_addedKey__33_comb[31:24];
  assign p3_bit_slice_1077200_comb = p3_addedKey__33_comb[23:16];
  assign p3_bit_slice_1077201_comb = p3_addedKey__33_comb[15:8];
  assign p3_bit_slice_1077202_comb = p3_addedKey__33_comb[79:72];
  assign p3_bit_slice_1077203_comb = p3_addedKey__33_comb[63:56];
  assign p3_bit_slice_1077204_comb = p3_addedKey__33_comb[7:0];

  // Registers for pipe stage 3:
  reg [127:0] p3_bit_slice_1076328;
  reg [127:0] p3_xor_1077141;
  reg [7:0] p3_bit_slice_1077189;
  reg [7:0] p3_bit_slice_1077190;
  reg [7:0] p3_bit_slice_1077191;
  reg [7:0] p3_bit_slice_1077192;
  reg [7:0] p3_bit_slice_1077193;
  reg [7:0] p3_bit_slice_1077194;
  reg [7:0] p3_bit_slice_1077195;
  reg [7:0] p3_bit_slice_1077196;
  reg [7:0] p3_bit_slice_1077197;
  reg [7:0] p3_bit_slice_1077198;
  reg [7:0] p3_bit_slice_1077199;
  reg [7:0] p3_bit_slice_1077200;
  reg [7:0] p3_bit_slice_1077201;
  reg [7:0] p3_bit_slice_1077202;
  reg [7:0] p3_bit_slice_1077203;
  reg [7:0] p3_bit_slice_1077204;
  reg [7:0] p4_arr[256];
  reg [7:0] p4_literal_1076345[256];
  reg [7:0] p4_literal_1076347[256];
  reg [7:0] p4_literal_1076349[256];
  reg [7:0] p4_literal_1076351[256];
  reg [7:0] p4_literal_1076353[256];
  reg [7:0] p4_literal_1076355[256];
  reg [7:0] p4_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p3_bit_slice_1076328 <= p2_bit_slice_1076328;
    p3_xor_1077141 <= p3_xor_1077141_comb;
    p3_bit_slice_1077189 <= p3_bit_slice_1077189_comb;
    p3_bit_slice_1077190 <= p3_bit_slice_1077190_comb;
    p3_bit_slice_1077191 <= p3_bit_slice_1077191_comb;
    p3_bit_slice_1077192 <= p3_bit_slice_1077192_comb;
    p3_bit_slice_1077193 <= p3_bit_slice_1077193_comb;
    p3_bit_slice_1077194 <= p3_bit_slice_1077194_comb;
    p3_bit_slice_1077195 <= p3_bit_slice_1077195_comb;
    p3_bit_slice_1077196 <= p3_bit_slice_1077196_comb;
    p3_bit_slice_1077197 <= p3_bit_slice_1077197_comb;
    p3_bit_slice_1077198 <= p3_bit_slice_1077198_comb;
    p3_bit_slice_1077199 <= p3_bit_slice_1077199_comb;
    p3_bit_slice_1077200 <= p3_bit_slice_1077200_comb;
    p3_bit_slice_1077201 <= p3_bit_slice_1077201_comb;
    p3_bit_slice_1077202 <= p3_bit_slice_1077202_comb;
    p3_bit_slice_1077203 <= p3_bit_slice_1077203_comb;
    p3_bit_slice_1077204 <= p3_bit_slice_1077204_comb;
    p4_arr <= p3_arr;
    p4_literal_1076345 <= p3_literal_1076345;
    p4_literal_1076347 <= p3_literal_1076347;
    p4_literal_1076349 <= p3_literal_1076349;
    p4_literal_1076351 <= p3_literal_1076351;
    p4_literal_1076353 <= p3_literal_1076353;
    p4_literal_1076355 <= p3_literal_1076355;
    p4_literal_1076358 <= p3_literal_1076358;
  end

  // ===== Pipe stage 4:
  wire [127:0] p4_addedKey__42_comb;
  wire [7:0] p4_array_index_1077272_comb;
  wire [7:0] p4_array_index_1077273_comb;
  wire [7:0] p4_array_index_1077274_comb;
  wire [7:0] p4_array_index_1077275_comb;
  wire [7:0] p4_array_index_1077276_comb;
  wire [7:0] p4_array_index_1077277_comb;
  wire [7:0] p4_array_index_1077279_comb;
  wire [7:0] p4_array_index_1077281_comb;
  wire [7:0] p4_array_index_1077282_comb;
  wire [7:0] p4_array_index_1077283_comb;
  wire [7:0] p4_array_index_1077284_comb;
  wire [7:0] p4_array_index_1077285_comb;
  wire [7:0] p4_array_index_1077286_comb;
  wire [7:0] p4_array_index_1077360_comb;
  wire [7:0] p4_array_index_1077361_comb;
  wire [7:0] p4_array_index_1077362_comb;
  wire [7:0] p4_array_index_1077363_comb;
  wire [7:0] p4_array_index_1077364_comb;
  wire [7:0] p4_array_index_1077365_comb;
  wire [7:0] p4_array_index_1077366_comb;
  wire [7:0] p4_array_index_1077367_comb;
  wire [7:0] p4_array_index_1077368_comb;
  wire [7:0] p4_array_index_1077369_comb;
  wire [7:0] p4_array_index_1077370_comb;
  wire [7:0] p4_array_index_1077371_comb;
  wire [7:0] p4_array_index_1077372_comb;
  wire [7:0] p4_array_index_1077288_comb;
  wire [7:0] p4_array_index_1077289_comb;
  wire [7:0] p4_array_index_1077290_comb;
  wire [7:0] p4_array_index_1077291_comb;
  wire [7:0] p4_array_index_1077292_comb;
  wire [7:0] p4_array_index_1077293_comb;
  wire [7:0] p4_array_index_1077294_comb;
  wire [7:0] p4_array_index_1077296_comb;
  wire [7:0] p4_array_index_1077373_comb;
  wire [7:0] p4_array_index_1077374_comb;
  wire [7:0] p4_array_index_1077375_comb;
  wire [7:0] p4_array_index_1077376_comb;
  wire [7:0] p4_array_index_1077377_comb;
  wire [7:0] p4_array_index_1077378_comb;
  wire [7:0] p4_array_index_1077379_comb;
  wire [7:0] p4_array_index_1077381_comb;
  wire [7:0] p4_res7__16_comb;
  wire [7:0] p4_res7__528_comb;
  wire [7:0] p4_array_index_1077305_comb;
  wire [7:0] p4_array_index_1077306_comb;
  wire [7:0] p4_array_index_1077307_comb;
  wire [7:0] p4_array_index_1077308_comb;
  wire [7:0] p4_array_index_1077309_comb;
  wire [7:0] p4_array_index_1077310_comb;
  wire [7:0] p4_array_index_1077390_comb;
  wire [7:0] p4_array_index_1077391_comb;
  wire [7:0] p4_array_index_1077392_comb;
  wire [7:0] p4_array_index_1077393_comb;
  wire [7:0] p4_array_index_1077394_comb;
  wire [7:0] p4_array_index_1077395_comb;
  wire [7:0] p4_res7__17_comb;
  wire [7:0] p4_res7__529_comb;
  wire [7:0] p4_array_index_1077320_comb;
  wire [7:0] p4_array_index_1077321_comb;
  wire [7:0] p4_array_index_1077322_comb;
  wire [7:0] p4_array_index_1077323_comb;
  wire [7:0] p4_array_index_1077324_comb;
  wire [7:0] p4_array_index_1077405_comb;
  wire [7:0] p4_array_index_1077406_comb;
  wire [7:0] p4_array_index_1077407_comb;
  wire [7:0] p4_array_index_1077408_comb;
  wire [7:0] p4_array_index_1077409_comb;
  wire [7:0] p4_res7__18_comb;
  wire [7:0] p4_res7__530_comb;
  wire [7:0] p4_array_index_1077334_comb;
  wire [7:0] p4_array_index_1077335_comb;
  wire [7:0] p4_array_index_1077336_comb;
  wire [7:0] p4_array_index_1077337_comb;
  wire [7:0] p4_array_index_1077338_comb;
  wire [7:0] p4_array_index_1077419_comb;
  wire [7:0] p4_array_index_1077420_comb;
  wire [7:0] p4_array_index_1077421_comb;
  wire [7:0] p4_array_index_1077422_comb;
  wire [7:0] p4_array_index_1077423_comb;
  wire [7:0] p4_res7__19_comb;
  wire [7:0] p4_res7__531_comb;
  wire [7:0] p4_array_index_1077349_comb;
  wire [7:0] p4_array_index_1077350_comb;
  wire [7:0] p4_array_index_1077351_comb;
  wire [7:0] p4_array_index_1077352_comb;
  wire [7:0] p4_array_index_1077434_comb;
  wire [7:0] p4_array_index_1077435_comb;
  wire [7:0] p4_array_index_1077436_comb;
  wire [7:0] p4_array_index_1077437_comb;
  wire [7:0] p4_res7__20_comb;
  wire [7:0] p4_res7__532_comb;
  assign p4_addedKey__42_comb = p3_xor_1077141 ^ 128'hdc87_ece4_d890_f4b3_ba4e_b920_79cb_eb02;
  assign p4_array_index_1077272_comb = p3_arr[p4_addedKey__42_comb[127:120]];
  assign p4_array_index_1077273_comb = p3_arr[p4_addedKey__42_comb[119:112]];
  assign p4_array_index_1077274_comb = p3_arr[p4_addedKey__42_comb[111:104]];
  assign p4_array_index_1077275_comb = p3_arr[p4_addedKey__42_comb[103:96]];
  assign p4_array_index_1077276_comb = p3_arr[p4_addedKey__42_comb[95:88]];
  assign p4_array_index_1077277_comb = p3_arr[p4_addedKey__42_comb[87:80]];
  assign p4_array_index_1077279_comb = p3_arr[p4_addedKey__42_comb[71:64]];
  assign p4_array_index_1077281_comb = p3_arr[p4_addedKey__42_comb[55:48]];
  assign p4_array_index_1077282_comb = p3_arr[p4_addedKey__42_comb[47:40]];
  assign p4_array_index_1077283_comb = p3_arr[p4_addedKey__42_comb[39:32]];
  assign p4_array_index_1077284_comb = p3_arr[p4_addedKey__42_comb[31:24]];
  assign p4_array_index_1077285_comb = p3_arr[p4_addedKey__42_comb[23:16]];
  assign p4_array_index_1077286_comb = p3_arr[p4_addedKey__42_comb[15:8]];
  assign p4_array_index_1077360_comb = p3_arr[p3_bit_slice_1077189];
  assign p4_array_index_1077361_comb = p3_arr[p3_bit_slice_1077190];
  assign p4_array_index_1077362_comb = p3_arr[p3_bit_slice_1077191];
  assign p4_array_index_1077363_comb = p3_arr[p3_bit_slice_1077192];
  assign p4_array_index_1077364_comb = p3_arr[p3_bit_slice_1077193];
  assign p4_array_index_1077365_comb = p3_arr[p3_bit_slice_1077194];
  assign p4_array_index_1077366_comb = p3_arr[p3_bit_slice_1077195];
  assign p4_array_index_1077367_comb = p3_arr[p3_bit_slice_1077196];
  assign p4_array_index_1077368_comb = p3_arr[p3_bit_slice_1077197];
  assign p4_array_index_1077369_comb = p3_arr[p3_bit_slice_1077198];
  assign p4_array_index_1077370_comb = p3_arr[p3_bit_slice_1077199];
  assign p4_array_index_1077371_comb = p3_arr[p3_bit_slice_1077200];
  assign p4_array_index_1077372_comb = p3_arr[p3_bit_slice_1077201];
  assign p4_array_index_1077288_comb = p3_literal_1076345[p4_array_index_1077272_comb];
  assign p4_array_index_1077289_comb = p3_literal_1076347[p4_array_index_1077273_comb];
  assign p4_array_index_1077290_comb = p3_literal_1076349[p4_array_index_1077274_comb];
  assign p4_array_index_1077291_comb = p3_literal_1076351[p4_array_index_1077275_comb];
  assign p4_array_index_1077292_comb = p3_literal_1076353[p4_array_index_1077276_comb];
  assign p4_array_index_1077293_comb = p3_literal_1076355[p4_array_index_1077277_comb];
  assign p4_array_index_1077294_comb = p3_arr[p4_addedKey__42_comb[79:72]];
  assign p4_array_index_1077296_comb = p3_arr[p4_addedKey__42_comb[63:56]];
  assign p4_array_index_1077373_comb = p3_literal_1076345[p4_array_index_1077360_comb];
  assign p4_array_index_1077374_comb = p3_literal_1076347[p4_array_index_1077361_comb];
  assign p4_array_index_1077375_comb = p3_literal_1076349[p4_array_index_1077362_comb];
  assign p4_array_index_1077376_comb = p3_literal_1076351[p4_array_index_1077363_comb];
  assign p4_array_index_1077377_comb = p3_literal_1076353[p4_array_index_1077364_comb];
  assign p4_array_index_1077378_comb = p3_literal_1076355[p4_array_index_1077365_comb];
  assign p4_array_index_1077379_comb = p3_arr[p3_bit_slice_1077202];
  assign p4_array_index_1077381_comb = p3_arr[p3_bit_slice_1077203];
  assign p4_res7__16_comb = p4_array_index_1077288_comb ^ p4_array_index_1077289_comb ^ p4_array_index_1077290_comb ^ p4_array_index_1077291_comb ^ p4_array_index_1077292_comb ^ p4_array_index_1077293_comb ^ p4_array_index_1077294_comb ^ p3_literal_1076358[p4_array_index_1077279_comb] ^ p4_array_index_1077296_comb ^ p3_literal_1076355[p4_array_index_1077281_comb] ^ p3_literal_1076353[p4_array_index_1077282_comb] ^ p3_literal_1076351[p4_array_index_1077283_comb] ^ p3_literal_1076349[p4_array_index_1077284_comb] ^ p3_literal_1076347[p4_array_index_1077285_comb] ^ p3_literal_1076345[p4_array_index_1077286_comb] ^ p3_arr[p4_addedKey__42_comb[7:0]];
  assign p4_res7__528_comb = p4_array_index_1077373_comb ^ p4_array_index_1077374_comb ^ p4_array_index_1077375_comb ^ p4_array_index_1077376_comb ^ p4_array_index_1077377_comb ^ p4_array_index_1077378_comb ^ p4_array_index_1077379_comb ^ p3_literal_1076358[p4_array_index_1077366_comb] ^ p4_array_index_1077381_comb ^ p3_literal_1076355[p4_array_index_1077367_comb] ^ p3_literal_1076353[p4_array_index_1077368_comb] ^ p3_literal_1076351[p4_array_index_1077369_comb] ^ p3_literal_1076349[p4_array_index_1077370_comb] ^ p3_literal_1076347[p4_array_index_1077371_comb] ^ p3_literal_1076345[p4_array_index_1077372_comb] ^ p3_arr[p3_bit_slice_1077204];
  assign p4_array_index_1077305_comb = p3_literal_1076345[p4_res7__16_comb];
  assign p4_array_index_1077306_comb = p3_literal_1076347[p4_array_index_1077272_comb];
  assign p4_array_index_1077307_comb = p3_literal_1076349[p4_array_index_1077273_comb];
  assign p4_array_index_1077308_comb = p3_literal_1076351[p4_array_index_1077274_comb];
  assign p4_array_index_1077309_comb = p3_literal_1076353[p4_array_index_1077275_comb];
  assign p4_array_index_1077310_comb = p3_literal_1076355[p4_array_index_1077276_comb];
  assign p4_array_index_1077390_comb = p3_literal_1076345[p4_res7__528_comb];
  assign p4_array_index_1077391_comb = p3_literal_1076347[p4_array_index_1077360_comb];
  assign p4_array_index_1077392_comb = p3_literal_1076349[p4_array_index_1077361_comb];
  assign p4_array_index_1077393_comb = p3_literal_1076351[p4_array_index_1077362_comb];
  assign p4_array_index_1077394_comb = p3_literal_1076353[p4_array_index_1077363_comb];
  assign p4_array_index_1077395_comb = p3_literal_1076355[p4_array_index_1077364_comb];
  assign p4_res7__17_comb = p4_array_index_1077305_comb ^ p4_array_index_1077306_comb ^ p4_array_index_1077307_comb ^ p4_array_index_1077308_comb ^ p4_array_index_1077309_comb ^ p4_array_index_1077310_comb ^ p4_array_index_1077277_comb ^ p3_literal_1076358[p4_array_index_1077294_comb] ^ p4_array_index_1077279_comb ^ p3_literal_1076355[p4_array_index_1077296_comb] ^ p3_literal_1076353[p4_array_index_1077281_comb] ^ p3_literal_1076351[p4_array_index_1077282_comb] ^ p3_literal_1076349[p4_array_index_1077283_comb] ^ p3_literal_1076347[p4_array_index_1077284_comb] ^ p3_literal_1076345[p4_array_index_1077285_comb] ^ p4_array_index_1077286_comb;
  assign p4_res7__529_comb = p4_array_index_1077390_comb ^ p4_array_index_1077391_comb ^ p4_array_index_1077392_comb ^ p4_array_index_1077393_comb ^ p4_array_index_1077394_comb ^ p4_array_index_1077395_comb ^ p4_array_index_1077365_comb ^ p3_literal_1076358[p4_array_index_1077379_comb] ^ p4_array_index_1077366_comb ^ p3_literal_1076355[p4_array_index_1077381_comb] ^ p3_literal_1076353[p4_array_index_1077367_comb] ^ p3_literal_1076351[p4_array_index_1077368_comb] ^ p3_literal_1076349[p4_array_index_1077369_comb] ^ p3_literal_1076347[p4_array_index_1077370_comb] ^ p3_literal_1076345[p4_array_index_1077371_comb] ^ p4_array_index_1077372_comb;
  assign p4_array_index_1077320_comb = p3_literal_1076347[p4_res7__16_comb];
  assign p4_array_index_1077321_comb = p3_literal_1076349[p4_array_index_1077272_comb];
  assign p4_array_index_1077322_comb = p3_literal_1076351[p4_array_index_1077273_comb];
  assign p4_array_index_1077323_comb = p3_literal_1076353[p4_array_index_1077274_comb];
  assign p4_array_index_1077324_comb = p3_literal_1076355[p4_array_index_1077275_comb];
  assign p4_array_index_1077405_comb = p3_literal_1076347[p4_res7__528_comb];
  assign p4_array_index_1077406_comb = p3_literal_1076349[p4_array_index_1077360_comb];
  assign p4_array_index_1077407_comb = p3_literal_1076351[p4_array_index_1077361_comb];
  assign p4_array_index_1077408_comb = p3_literal_1076353[p4_array_index_1077362_comb];
  assign p4_array_index_1077409_comb = p3_literal_1076355[p4_array_index_1077363_comb];
  assign p4_res7__18_comb = p3_literal_1076345[p4_res7__17_comb] ^ p4_array_index_1077320_comb ^ p4_array_index_1077321_comb ^ p4_array_index_1077322_comb ^ p4_array_index_1077323_comb ^ p4_array_index_1077324_comb ^ p4_array_index_1077276_comb ^ p3_literal_1076358[p4_array_index_1077277_comb] ^ p4_array_index_1077294_comb ^ p3_literal_1076355[p4_array_index_1077279_comb] ^ p3_literal_1076353[p4_array_index_1077296_comb] ^ p3_literal_1076351[p4_array_index_1077281_comb] ^ p3_literal_1076349[p4_array_index_1077282_comb] ^ p3_literal_1076347[p4_array_index_1077283_comb] ^ p3_literal_1076345[p4_array_index_1077284_comb] ^ p4_array_index_1077285_comb;
  assign p4_res7__530_comb = p3_literal_1076345[p4_res7__529_comb] ^ p4_array_index_1077405_comb ^ p4_array_index_1077406_comb ^ p4_array_index_1077407_comb ^ p4_array_index_1077408_comb ^ p4_array_index_1077409_comb ^ p4_array_index_1077364_comb ^ p3_literal_1076358[p4_array_index_1077365_comb] ^ p4_array_index_1077379_comb ^ p3_literal_1076355[p4_array_index_1077366_comb] ^ p3_literal_1076353[p4_array_index_1077381_comb] ^ p3_literal_1076351[p4_array_index_1077367_comb] ^ p3_literal_1076349[p4_array_index_1077368_comb] ^ p3_literal_1076347[p4_array_index_1077369_comb] ^ p3_literal_1076345[p4_array_index_1077370_comb] ^ p4_array_index_1077371_comb;
  assign p4_array_index_1077334_comb = p3_literal_1076347[p4_res7__17_comb];
  assign p4_array_index_1077335_comb = p3_literal_1076349[p4_res7__16_comb];
  assign p4_array_index_1077336_comb = p3_literal_1076351[p4_array_index_1077272_comb];
  assign p4_array_index_1077337_comb = p3_literal_1076353[p4_array_index_1077273_comb];
  assign p4_array_index_1077338_comb = p3_literal_1076355[p4_array_index_1077274_comb];
  assign p4_array_index_1077419_comb = p3_literal_1076347[p4_res7__529_comb];
  assign p4_array_index_1077420_comb = p3_literal_1076349[p4_res7__528_comb];
  assign p4_array_index_1077421_comb = p3_literal_1076351[p4_array_index_1077360_comb];
  assign p4_array_index_1077422_comb = p3_literal_1076353[p4_array_index_1077361_comb];
  assign p4_array_index_1077423_comb = p3_literal_1076355[p4_array_index_1077362_comb];
  assign p4_res7__19_comb = p3_literal_1076345[p4_res7__18_comb] ^ p4_array_index_1077334_comb ^ p4_array_index_1077335_comb ^ p4_array_index_1077336_comb ^ p4_array_index_1077337_comb ^ p4_array_index_1077338_comb ^ p4_array_index_1077275_comb ^ p3_literal_1076358[p4_array_index_1077276_comb] ^ p4_array_index_1077277_comb ^ p3_literal_1076355[p4_array_index_1077294_comb] ^ p3_literal_1076353[p4_array_index_1077279_comb] ^ p3_literal_1076351[p4_array_index_1077296_comb] ^ p3_literal_1076349[p4_array_index_1077281_comb] ^ p3_literal_1076347[p4_array_index_1077282_comb] ^ p3_literal_1076345[p4_array_index_1077283_comb] ^ p4_array_index_1077284_comb;
  assign p4_res7__531_comb = p3_literal_1076345[p4_res7__530_comb] ^ p4_array_index_1077419_comb ^ p4_array_index_1077420_comb ^ p4_array_index_1077421_comb ^ p4_array_index_1077422_comb ^ p4_array_index_1077423_comb ^ p4_array_index_1077363_comb ^ p3_literal_1076358[p4_array_index_1077364_comb] ^ p4_array_index_1077365_comb ^ p3_literal_1076355[p4_array_index_1077379_comb] ^ p3_literal_1076353[p4_array_index_1077366_comb] ^ p3_literal_1076351[p4_array_index_1077381_comb] ^ p3_literal_1076349[p4_array_index_1077367_comb] ^ p3_literal_1076347[p4_array_index_1077368_comb] ^ p3_literal_1076345[p4_array_index_1077369_comb] ^ p4_array_index_1077370_comb;
  assign p4_array_index_1077349_comb = p3_literal_1076349[p4_res7__17_comb];
  assign p4_array_index_1077350_comb = p3_literal_1076351[p4_res7__16_comb];
  assign p4_array_index_1077351_comb = p3_literal_1076353[p4_array_index_1077272_comb];
  assign p4_array_index_1077352_comb = p3_literal_1076355[p4_array_index_1077273_comb];
  assign p4_array_index_1077434_comb = p3_literal_1076349[p4_res7__529_comb];
  assign p4_array_index_1077435_comb = p3_literal_1076351[p4_res7__528_comb];
  assign p4_array_index_1077436_comb = p3_literal_1076353[p4_array_index_1077360_comb];
  assign p4_array_index_1077437_comb = p3_literal_1076355[p4_array_index_1077361_comb];
  assign p4_res7__20_comb = p3_literal_1076345[p4_res7__19_comb] ^ p3_literal_1076347[p4_res7__18_comb] ^ p4_array_index_1077349_comb ^ p4_array_index_1077350_comb ^ p4_array_index_1077351_comb ^ p4_array_index_1077352_comb ^ p4_array_index_1077274_comb ^ p3_literal_1076358[p4_array_index_1077275_comb] ^ p4_array_index_1077276_comb ^ p4_array_index_1077293_comb ^ p3_literal_1076353[p4_array_index_1077294_comb] ^ p3_literal_1076351[p4_array_index_1077279_comb] ^ p3_literal_1076349[p4_array_index_1077296_comb] ^ p3_literal_1076347[p4_array_index_1077281_comb] ^ p3_literal_1076345[p4_array_index_1077282_comb] ^ p4_array_index_1077283_comb;
  assign p4_res7__532_comb = p3_literal_1076345[p4_res7__531_comb] ^ p3_literal_1076347[p4_res7__530_comb] ^ p4_array_index_1077434_comb ^ p4_array_index_1077435_comb ^ p4_array_index_1077436_comb ^ p4_array_index_1077437_comb ^ p4_array_index_1077362_comb ^ p3_literal_1076358[p4_array_index_1077363_comb] ^ p4_array_index_1077364_comb ^ p4_array_index_1077378_comb ^ p3_literal_1076353[p4_array_index_1077379_comb] ^ p3_literal_1076351[p4_array_index_1077366_comb] ^ p3_literal_1076349[p4_array_index_1077381_comb] ^ p3_literal_1076347[p4_array_index_1077367_comb] ^ p3_literal_1076345[p4_array_index_1077368_comb] ^ p4_array_index_1077369_comb;

  // Registers for pipe stage 4:
  reg [127:0] p4_bit_slice_1076328;
  reg [127:0] p4_xor_1077141;
  reg [7:0] p4_array_index_1077272;
  reg [7:0] p4_array_index_1077273;
  reg [7:0] p4_array_index_1077274;
  reg [7:0] p4_array_index_1077275;
  reg [7:0] p4_array_index_1077276;
  reg [7:0] p4_array_index_1077277;
  reg [7:0] p4_array_index_1077279;
  reg [7:0] p4_array_index_1077281;
  reg [7:0] p4_array_index_1077282;
  reg [7:0] p4_array_index_1077288;
  reg [7:0] p4_array_index_1077289;
  reg [7:0] p4_array_index_1077290;
  reg [7:0] p4_array_index_1077291;
  reg [7:0] p4_array_index_1077292;
  reg [7:0] p4_array_index_1077294;
  reg [7:0] p4_array_index_1077296;
  reg [7:0] p4_res7__16;
  reg [7:0] p4_array_index_1077305;
  reg [7:0] p4_array_index_1077306;
  reg [7:0] p4_array_index_1077307;
  reg [7:0] p4_array_index_1077308;
  reg [7:0] p4_array_index_1077309;
  reg [7:0] p4_array_index_1077310;
  reg [7:0] p4_res7__17;
  reg [7:0] p4_array_index_1077320;
  reg [7:0] p4_array_index_1077321;
  reg [7:0] p4_array_index_1077322;
  reg [7:0] p4_array_index_1077323;
  reg [7:0] p4_array_index_1077324;
  reg [7:0] p4_res7__18;
  reg [7:0] p4_array_index_1077334;
  reg [7:0] p4_array_index_1077335;
  reg [7:0] p4_array_index_1077336;
  reg [7:0] p4_array_index_1077337;
  reg [7:0] p4_array_index_1077338;
  reg [7:0] p4_res7__19;
  reg [7:0] p4_array_index_1077349;
  reg [7:0] p4_array_index_1077350;
  reg [7:0] p4_array_index_1077351;
  reg [7:0] p4_array_index_1077352;
  reg [7:0] p4_res7__20;
  reg [7:0] p4_array_index_1077360;
  reg [7:0] p4_array_index_1077361;
  reg [7:0] p4_array_index_1077362;
  reg [7:0] p4_array_index_1077363;
  reg [7:0] p4_array_index_1077364;
  reg [7:0] p4_array_index_1077365;
  reg [7:0] p4_array_index_1077366;
  reg [7:0] p4_array_index_1077367;
  reg [7:0] p4_array_index_1077368;
  reg [7:0] p4_array_index_1077373;
  reg [7:0] p4_array_index_1077374;
  reg [7:0] p4_array_index_1077375;
  reg [7:0] p4_array_index_1077376;
  reg [7:0] p4_array_index_1077377;
  reg [7:0] p4_array_index_1077379;
  reg [7:0] p4_array_index_1077381;
  reg [7:0] p4_res7__528;
  reg [7:0] p4_array_index_1077390;
  reg [7:0] p4_array_index_1077391;
  reg [7:0] p4_array_index_1077392;
  reg [7:0] p4_array_index_1077393;
  reg [7:0] p4_array_index_1077394;
  reg [7:0] p4_array_index_1077395;
  reg [7:0] p4_res7__529;
  reg [7:0] p4_array_index_1077405;
  reg [7:0] p4_array_index_1077406;
  reg [7:0] p4_array_index_1077407;
  reg [7:0] p4_array_index_1077408;
  reg [7:0] p4_array_index_1077409;
  reg [7:0] p4_res7__530;
  reg [7:0] p4_array_index_1077419;
  reg [7:0] p4_array_index_1077420;
  reg [7:0] p4_array_index_1077421;
  reg [7:0] p4_array_index_1077422;
  reg [7:0] p4_array_index_1077423;
  reg [7:0] p4_res7__531;
  reg [7:0] p4_array_index_1077434;
  reg [7:0] p4_array_index_1077435;
  reg [7:0] p4_array_index_1077436;
  reg [7:0] p4_array_index_1077437;
  reg [7:0] p4_res7__532;
  reg [7:0] p5_arr[256];
  reg [7:0] p5_literal_1076345[256];
  reg [7:0] p5_literal_1076347[256];
  reg [7:0] p5_literal_1076349[256];
  reg [7:0] p5_literal_1076351[256];
  reg [7:0] p5_literal_1076353[256];
  reg [7:0] p5_literal_1076355[256];
  reg [7:0] p5_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p4_bit_slice_1076328 <= p3_bit_slice_1076328;
    p4_xor_1077141 <= p3_xor_1077141;
    p4_array_index_1077272 <= p4_array_index_1077272_comb;
    p4_array_index_1077273 <= p4_array_index_1077273_comb;
    p4_array_index_1077274 <= p4_array_index_1077274_comb;
    p4_array_index_1077275 <= p4_array_index_1077275_comb;
    p4_array_index_1077276 <= p4_array_index_1077276_comb;
    p4_array_index_1077277 <= p4_array_index_1077277_comb;
    p4_array_index_1077279 <= p4_array_index_1077279_comb;
    p4_array_index_1077281 <= p4_array_index_1077281_comb;
    p4_array_index_1077282 <= p4_array_index_1077282_comb;
    p4_array_index_1077288 <= p4_array_index_1077288_comb;
    p4_array_index_1077289 <= p4_array_index_1077289_comb;
    p4_array_index_1077290 <= p4_array_index_1077290_comb;
    p4_array_index_1077291 <= p4_array_index_1077291_comb;
    p4_array_index_1077292 <= p4_array_index_1077292_comb;
    p4_array_index_1077294 <= p4_array_index_1077294_comb;
    p4_array_index_1077296 <= p4_array_index_1077296_comb;
    p4_res7__16 <= p4_res7__16_comb;
    p4_array_index_1077305 <= p4_array_index_1077305_comb;
    p4_array_index_1077306 <= p4_array_index_1077306_comb;
    p4_array_index_1077307 <= p4_array_index_1077307_comb;
    p4_array_index_1077308 <= p4_array_index_1077308_comb;
    p4_array_index_1077309 <= p4_array_index_1077309_comb;
    p4_array_index_1077310 <= p4_array_index_1077310_comb;
    p4_res7__17 <= p4_res7__17_comb;
    p4_array_index_1077320 <= p4_array_index_1077320_comb;
    p4_array_index_1077321 <= p4_array_index_1077321_comb;
    p4_array_index_1077322 <= p4_array_index_1077322_comb;
    p4_array_index_1077323 <= p4_array_index_1077323_comb;
    p4_array_index_1077324 <= p4_array_index_1077324_comb;
    p4_res7__18 <= p4_res7__18_comb;
    p4_array_index_1077334 <= p4_array_index_1077334_comb;
    p4_array_index_1077335 <= p4_array_index_1077335_comb;
    p4_array_index_1077336 <= p4_array_index_1077336_comb;
    p4_array_index_1077337 <= p4_array_index_1077337_comb;
    p4_array_index_1077338 <= p4_array_index_1077338_comb;
    p4_res7__19 <= p4_res7__19_comb;
    p4_array_index_1077349 <= p4_array_index_1077349_comb;
    p4_array_index_1077350 <= p4_array_index_1077350_comb;
    p4_array_index_1077351 <= p4_array_index_1077351_comb;
    p4_array_index_1077352 <= p4_array_index_1077352_comb;
    p4_res7__20 <= p4_res7__20_comb;
    p4_array_index_1077360 <= p4_array_index_1077360_comb;
    p4_array_index_1077361 <= p4_array_index_1077361_comb;
    p4_array_index_1077362 <= p4_array_index_1077362_comb;
    p4_array_index_1077363 <= p4_array_index_1077363_comb;
    p4_array_index_1077364 <= p4_array_index_1077364_comb;
    p4_array_index_1077365 <= p4_array_index_1077365_comb;
    p4_array_index_1077366 <= p4_array_index_1077366_comb;
    p4_array_index_1077367 <= p4_array_index_1077367_comb;
    p4_array_index_1077368 <= p4_array_index_1077368_comb;
    p4_array_index_1077373 <= p4_array_index_1077373_comb;
    p4_array_index_1077374 <= p4_array_index_1077374_comb;
    p4_array_index_1077375 <= p4_array_index_1077375_comb;
    p4_array_index_1077376 <= p4_array_index_1077376_comb;
    p4_array_index_1077377 <= p4_array_index_1077377_comb;
    p4_array_index_1077379 <= p4_array_index_1077379_comb;
    p4_array_index_1077381 <= p4_array_index_1077381_comb;
    p4_res7__528 <= p4_res7__528_comb;
    p4_array_index_1077390 <= p4_array_index_1077390_comb;
    p4_array_index_1077391 <= p4_array_index_1077391_comb;
    p4_array_index_1077392 <= p4_array_index_1077392_comb;
    p4_array_index_1077393 <= p4_array_index_1077393_comb;
    p4_array_index_1077394 <= p4_array_index_1077394_comb;
    p4_array_index_1077395 <= p4_array_index_1077395_comb;
    p4_res7__529 <= p4_res7__529_comb;
    p4_array_index_1077405 <= p4_array_index_1077405_comb;
    p4_array_index_1077406 <= p4_array_index_1077406_comb;
    p4_array_index_1077407 <= p4_array_index_1077407_comb;
    p4_array_index_1077408 <= p4_array_index_1077408_comb;
    p4_array_index_1077409 <= p4_array_index_1077409_comb;
    p4_res7__530 <= p4_res7__530_comb;
    p4_array_index_1077419 <= p4_array_index_1077419_comb;
    p4_array_index_1077420 <= p4_array_index_1077420_comb;
    p4_array_index_1077421 <= p4_array_index_1077421_comb;
    p4_array_index_1077422 <= p4_array_index_1077422_comb;
    p4_array_index_1077423 <= p4_array_index_1077423_comb;
    p4_res7__531 <= p4_res7__531_comb;
    p4_array_index_1077434 <= p4_array_index_1077434_comb;
    p4_array_index_1077435 <= p4_array_index_1077435_comb;
    p4_array_index_1077436 <= p4_array_index_1077436_comb;
    p4_array_index_1077437 <= p4_array_index_1077437_comb;
    p4_res7__532 <= p4_res7__532_comb;
    p5_arr <= p4_arr;
    p5_literal_1076345 <= p4_literal_1076345;
    p5_literal_1076347 <= p4_literal_1076347;
    p5_literal_1076349 <= p4_literal_1076349;
    p5_literal_1076351 <= p4_literal_1076351;
    p5_literal_1076353 <= p4_literal_1076353;
    p5_literal_1076355 <= p4_literal_1076355;
    p5_literal_1076358 <= p4_literal_1076358;
  end

  // ===== Pipe stage 5:
  wire [7:0] p5_array_index_1077631_comb;
  wire [7:0] p5_array_index_1077632_comb;
  wire [7:0] p5_array_index_1077633_comb;
  wire [7:0] p5_array_index_1077634_comb;
  wire [7:0] p5_res7__21_comb;
  wire [7:0] p5_array_index_1077699_comb;
  wire [7:0] p5_array_index_1077700_comb;
  wire [7:0] p5_array_index_1077701_comb;
  wire [7:0] p5_array_index_1077702_comb;
  wire [7:0] p5_array_index_1077645_comb;
  wire [7:0] p5_array_index_1077646_comb;
  wire [7:0] p5_array_index_1077647_comb;
  wire [7:0] p5_res7__533_comb;
  wire [7:0] p5_res7__22_comb;
  wire [7:0] p5_array_index_1077713_comb;
  wire [7:0] p5_array_index_1077714_comb;
  wire [7:0] p5_array_index_1077715_comb;
  wire [7:0] p5_array_index_1077657_comb;
  wire [7:0] p5_array_index_1077658_comb;
  wire [7:0] p5_array_index_1077659_comb;
  wire [7:0] p5_res7__534_comb;
  wire [7:0] p5_res7__23_comb;
  wire [7:0] p5_array_index_1077725_comb;
  wire [7:0] p5_array_index_1077726_comb;
  wire [7:0] p5_array_index_1077727_comb;
  wire [7:0] p5_array_index_1077670_comb;
  wire [7:0] p5_array_index_1077671_comb;
  wire [7:0] p5_res7__535_comb;
  wire [7:0] p5_res7__24_comb;
  wire [7:0] p5_array_index_1077738_comb;
  wire [7:0] p5_array_index_1077739_comb;
  wire [7:0] p5_array_index_1077681_comb;
  wire [7:0] p5_array_index_1077682_comb;
  wire [7:0] p5_res7__536_comb;
  wire [7:0] p5_res7__25_comb;
  wire [7:0] p5_array_index_1077749_comb;
  wire [7:0] p5_array_index_1077750_comb;
  wire [7:0] p5_array_index_1077688_comb;
  wire [7:0] p5_array_index_1077689_comb;
  wire [7:0] p5_array_index_1077690_comb;
  wire [7:0] p5_array_index_1077691_comb;
  wire [7:0] p5_array_index_1077692_comb;
  wire [7:0] p5_array_index_1077693_comb;
  wire [7:0] p5_array_index_1077694_comb;
  wire [7:0] p5_array_index_1077695_comb;
  wire [7:0] p5_array_index_1077696_comb;
  wire [7:0] p5_res7__537_comb;
  assign p5_array_index_1077631_comb = p4_literal_1076349[p4_res7__18];
  assign p5_array_index_1077632_comb = p4_literal_1076351[p4_res7__17];
  assign p5_array_index_1077633_comb = p4_literal_1076353[p4_res7__16];
  assign p5_array_index_1077634_comb = p4_literal_1076355[p4_array_index_1077272];
  assign p5_res7__21_comb = p4_literal_1076345[p4_res7__20] ^ p4_literal_1076347[p4_res7__19] ^ p5_array_index_1077631_comb ^ p5_array_index_1077632_comb ^ p5_array_index_1077633_comb ^ p5_array_index_1077634_comb ^ p4_array_index_1077273 ^ p4_literal_1076358[p4_array_index_1077274] ^ p4_array_index_1077275 ^ p4_array_index_1077310 ^ p4_literal_1076353[p4_array_index_1077277] ^ p4_literal_1076351[p4_array_index_1077294] ^ p4_literal_1076349[p4_array_index_1077279] ^ p4_literal_1076347[p4_array_index_1077296] ^ p4_literal_1076345[p4_array_index_1077281] ^ p4_array_index_1077282;
  assign p5_array_index_1077699_comb = p4_literal_1076349[p4_res7__530];
  assign p5_array_index_1077700_comb = p4_literal_1076351[p4_res7__529];
  assign p5_array_index_1077701_comb = p4_literal_1076353[p4_res7__528];
  assign p5_array_index_1077702_comb = p4_literal_1076355[p4_array_index_1077360];
  assign p5_array_index_1077645_comb = p4_literal_1076351[p4_res7__18];
  assign p5_array_index_1077646_comb = p4_literal_1076353[p4_res7__17];
  assign p5_array_index_1077647_comb = p4_literal_1076355[p4_res7__16];
  assign p5_res7__533_comb = p4_literal_1076345[p4_res7__532] ^ p4_literal_1076347[p4_res7__531] ^ p5_array_index_1077699_comb ^ p5_array_index_1077700_comb ^ p5_array_index_1077701_comb ^ p5_array_index_1077702_comb ^ p4_array_index_1077361 ^ p4_literal_1076358[p4_array_index_1077362] ^ p4_array_index_1077363 ^ p4_array_index_1077395 ^ p4_literal_1076353[p4_array_index_1077365] ^ p4_literal_1076351[p4_array_index_1077379] ^ p4_literal_1076349[p4_array_index_1077366] ^ p4_literal_1076347[p4_array_index_1077381] ^ p4_literal_1076345[p4_array_index_1077367] ^ p4_array_index_1077368;
  assign p5_res7__22_comb = p4_literal_1076345[p5_res7__21_comb] ^ p4_literal_1076347[p4_res7__20] ^ p4_literal_1076349[p4_res7__19] ^ p5_array_index_1077645_comb ^ p5_array_index_1077646_comb ^ p5_array_index_1077647_comb ^ p4_array_index_1077272 ^ p4_literal_1076358[p4_array_index_1077273] ^ p4_array_index_1077274 ^ p4_array_index_1077324 ^ p4_array_index_1077292 ^ p4_literal_1076351[p4_array_index_1077277] ^ p4_literal_1076349[p4_array_index_1077294] ^ p4_literal_1076347[p4_array_index_1077279] ^ p4_literal_1076345[p4_array_index_1077296] ^ p4_array_index_1077281;
  assign p5_array_index_1077713_comb = p4_literal_1076351[p4_res7__530];
  assign p5_array_index_1077714_comb = p4_literal_1076353[p4_res7__529];
  assign p5_array_index_1077715_comb = p4_literal_1076355[p4_res7__528];
  assign p5_array_index_1077657_comb = p4_literal_1076351[p4_res7__19];
  assign p5_array_index_1077658_comb = p4_literal_1076353[p4_res7__18];
  assign p5_array_index_1077659_comb = p4_literal_1076355[p4_res7__17];
  assign p5_res7__534_comb = p4_literal_1076345[p5_res7__533_comb] ^ p4_literal_1076347[p4_res7__532] ^ p4_literal_1076349[p4_res7__531] ^ p5_array_index_1077713_comb ^ p5_array_index_1077714_comb ^ p5_array_index_1077715_comb ^ p4_array_index_1077360 ^ p4_literal_1076358[p4_array_index_1077361] ^ p4_array_index_1077362 ^ p4_array_index_1077409 ^ p4_array_index_1077377 ^ p4_literal_1076351[p4_array_index_1077365] ^ p4_literal_1076349[p4_array_index_1077379] ^ p4_literal_1076347[p4_array_index_1077366] ^ p4_literal_1076345[p4_array_index_1077381] ^ p4_array_index_1077367;
  assign p5_res7__23_comb = p4_literal_1076345[p5_res7__22_comb] ^ p4_literal_1076347[p5_res7__21_comb] ^ p4_literal_1076349[p4_res7__20] ^ p5_array_index_1077657_comb ^ p5_array_index_1077658_comb ^ p5_array_index_1077659_comb ^ p4_res7__16 ^ p4_literal_1076358[p4_array_index_1077272] ^ p4_array_index_1077273 ^ p4_array_index_1077338 ^ p4_array_index_1077309 ^ p4_literal_1076351[p4_array_index_1077276] ^ p4_literal_1076349[p4_array_index_1077277] ^ p4_literal_1076347[p4_array_index_1077294] ^ p4_literal_1076345[p4_array_index_1077279] ^ p4_array_index_1077296;
  assign p5_array_index_1077725_comb = p4_literal_1076351[p4_res7__531];
  assign p5_array_index_1077726_comb = p4_literal_1076353[p4_res7__530];
  assign p5_array_index_1077727_comb = p4_literal_1076355[p4_res7__529];
  assign p5_array_index_1077670_comb = p4_literal_1076353[p4_res7__19];
  assign p5_array_index_1077671_comb = p4_literal_1076355[p4_res7__18];
  assign p5_res7__535_comb = p4_literal_1076345[p5_res7__534_comb] ^ p4_literal_1076347[p5_res7__533_comb] ^ p4_literal_1076349[p4_res7__532] ^ p5_array_index_1077725_comb ^ p5_array_index_1077726_comb ^ p5_array_index_1077727_comb ^ p4_res7__528 ^ p4_literal_1076358[p4_array_index_1077360] ^ p4_array_index_1077361 ^ p4_array_index_1077423 ^ p4_array_index_1077394 ^ p4_literal_1076351[p4_array_index_1077364] ^ p4_literal_1076349[p4_array_index_1077365] ^ p4_literal_1076347[p4_array_index_1077379] ^ p4_literal_1076345[p4_array_index_1077366] ^ p4_array_index_1077381;
  assign p5_res7__24_comb = p4_literal_1076345[p5_res7__23_comb] ^ p4_literal_1076347[p5_res7__22_comb] ^ p4_literal_1076349[p5_res7__21_comb] ^ p4_literal_1076351[p4_res7__20] ^ p5_array_index_1077670_comb ^ p5_array_index_1077671_comb ^ p4_res7__17 ^ p4_literal_1076358[p4_res7__16] ^ p4_array_index_1077272 ^ p4_array_index_1077352 ^ p4_array_index_1077323 ^ p4_array_index_1077291 ^ p4_literal_1076349[p4_array_index_1077276] ^ p4_literal_1076347[p4_array_index_1077277] ^ p4_literal_1076345[p4_array_index_1077294] ^ p4_array_index_1077279;
  assign p5_array_index_1077738_comb = p4_literal_1076353[p4_res7__531];
  assign p5_array_index_1077739_comb = p4_literal_1076355[p4_res7__530];
  assign p5_array_index_1077681_comb = p4_literal_1076353[p4_res7__20];
  assign p5_array_index_1077682_comb = p4_literal_1076355[p4_res7__19];
  assign p5_res7__536_comb = p4_literal_1076345[p5_res7__535_comb] ^ p4_literal_1076347[p5_res7__534_comb] ^ p4_literal_1076349[p5_res7__533_comb] ^ p4_literal_1076351[p4_res7__532] ^ p5_array_index_1077738_comb ^ p5_array_index_1077739_comb ^ p4_res7__529 ^ p4_literal_1076358[p4_res7__528] ^ p4_array_index_1077360 ^ p4_array_index_1077437 ^ p4_array_index_1077408 ^ p4_array_index_1077376 ^ p4_literal_1076349[p4_array_index_1077364] ^ p4_literal_1076347[p4_array_index_1077365] ^ p4_literal_1076345[p4_array_index_1077379] ^ p4_array_index_1077366;
  assign p5_res7__25_comb = p4_literal_1076345[p5_res7__24_comb] ^ p4_literal_1076347[p5_res7__23_comb] ^ p4_literal_1076349[p5_res7__22_comb] ^ p4_literal_1076351[p5_res7__21_comb] ^ p5_array_index_1077681_comb ^ p5_array_index_1077682_comb ^ p4_res7__18 ^ p4_literal_1076358[p4_res7__17] ^ p4_res7__16 ^ p5_array_index_1077634_comb ^ p4_array_index_1077337 ^ p4_array_index_1077308 ^ p4_literal_1076349[p4_array_index_1077275] ^ p4_literal_1076347[p4_array_index_1077276] ^ p4_literal_1076345[p4_array_index_1077277] ^ p4_array_index_1077294;
  assign p5_array_index_1077749_comb = p4_literal_1076353[p4_res7__532];
  assign p5_array_index_1077750_comb = p4_literal_1076355[p4_res7__531];
  assign p5_array_index_1077688_comb = p4_literal_1076345[p5_res7__25_comb];
  assign p5_array_index_1077689_comb = p4_literal_1076347[p5_res7__24_comb];
  assign p5_array_index_1077690_comb = p4_literal_1076349[p5_res7__23_comb];
  assign p5_array_index_1077691_comb = p4_literal_1076351[p5_res7__22_comb];
  assign p5_array_index_1077692_comb = p4_literal_1076353[p5_res7__21_comb];
  assign p5_array_index_1077693_comb = p4_literal_1076355[p4_res7__20];
  assign p5_array_index_1077694_comb = p4_literal_1076358[p4_res7__18];
  assign p5_array_index_1077695_comb = p4_literal_1076347[p4_array_index_1077275];
  assign p5_array_index_1077696_comb = p4_literal_1076345[p4_array_index_1077276];
  assign p5_res7__537_comb = p4_literal_1076345[p5_res7__536_comb] ^ p4_literal_1076347[p5_res7__535_comb] ^ p4_literal_1076349[p5_res7__534_comb] ^ p4_literal_1076351[p5_res7__533_comb] ^ p5_array_index_1077749_comb ^ p5_array_index_1077750_comb ^ p4_res7__530 ^ p4_literal_1076358[p4_res7__529] ^ p4_res7__528 ^ p5_array_index_1077702_comb ^ p4_array_index_1077422 ^ p4_array_index_1077393 ^ p4_literal_1076349[p4_array_index_1077363] ^ p4_literal_1076347[p4_array_index_1077364] ^ p4_literal_1076345[p4_array_index_1077365] ^ p4_array_index_1077379;

  // Registers for pipe stage 5:
  reg [127:0] p5_bit_slice_1076328;
  reg [127:0] p5_xor_1077141;
  reg [7:0] p5_array_index_1077272;
  reg [7:0] p5_array_index_1077273;
  reg [7:0] p5_array_index_1077274;
  reg [7:0] p5_array_index_1077275;
  reg [7:0] p5_array_index_1077276;
  reg [7:0] p5_array_index_1077277;
  reg [7:0] p5_array_index_1077288;
  reg [7:0] p5_array_index_1077289;
  reg [7:0] p5_array_index_1077290;
  reg [7:0] p5_res7__16;
  reg [7:0] p5_array_index_1077305;
  reg [7:0] p5_array_index_1077306;
  reg [7:0] p5_array_index_1077307;
  reg [7:0] p5_res7__17;
  reg [7:0] p5_array_index_1077320;
  reg [7:0] p5_array_index_1077321;
  reg [7:0] p5_array_index_1077322;
  reg [7:0] p5_res7__18;
  reg [7:0] p5_array_index_1077334;
  reg [7:0] p5_array_index_1077335;
  reg [7:0] p5_array_index_1077336;
  reg [7:0] p5_res7__19;
  reg [7:0] p5_array_index_1077349;
  reg [7:0] p5_array_index_1077350;
  reg [7:0] p5_array_index_1077351;
  reg [7:0] p5_res7__20;
  reg [7:0] p5_array_index_1077631;
  reg [7:0] p5_array_index_1077632;
  reg [7:0] p5_array_index_1077633;
  reg [7:0] p5_res7__21;
  reg [7:0] p5_array_index_1077645;
  reg [7:0] p5_array_index_1077646;
  reg [7:0] p5_array_index_1077647;
  reg [7:0] p5_res7__22;
  reg [7:0] p5_array_index_1077657;
  reg [7:0] p5_array_index_1077658;
  reg [7:0] p5_array_index_1077659;
  reg [7:0] p5_res7__23;
  reg [7:0] p5_array_index_1077670;
  reg [7:0] p5_array_index_1077671;
  reg [7:0] p5_res7__24;
  reg [7:0] p5_array_index_1077681;
  reg [7:0] p5_array_index_1077682;
  reg [7:0] p5_res7__25;
  reg [7:0] p5_array_index_1077688;
  reg [7:0] p5_array_index_1077689;
  reg [7:0] p5_array_index_1077690;
  reg [7:0] p5_array_index_1077691;
  reg [7:0] p5_array_index_1077692;
  reg [7:0] p5_array_index_1077693;
  reg [7:0] p5_array_index_1077694;
  reg [7:0] p5_array_index_1077695;
  reg [7:0] p5_array_index_1077696;
  reg [7:0] p5_array_index_1077360;
  reg [7:0] p5_array_index_1077361;
  reg [7:0] p5_array_index_1077362;
  reg [7:0] p5_array_index_1077363;
  reg [7:0] p5_array_index_1077364;
  reg [7:0] p5_array_index_1077365;
  reg [7:0] p5_array_index_1077373;
  reg [7:0] p5_array_index_1077374;
  reg [7:0] p5_array_index_1077375;
  reg [7:0] p5_res7__528;
  reg [7:0] p5_array_index_1077390;
  reg [7:0] p5_array_index_1077391;
  reg [7:0] p5_array_index_1077392;
  reg [7:0] p5_res7__529;
  reg [7:0] p5_array_index_1077405;
  reg [7:0] p5_array_index_1077406;
  reg [7:0] p5_array_index_1077407;
  reg [7:0] p5_res7__530;
  reg [7:0] p5_array_index_1077419;
  reg [7:0] p5_array_index_1077420;
  reg [7:0] p5_array_index_1077421;
  reg [7:0] p5_res7__531;
  reg [7:0] p5_array_index_1077434;
  reg [7:0] p5_array_index_1077435;
  reg [7:0] p5_array_index_1077436;
  reg [7:0] p5_res7__532;
  reg [7:0] p5_array_index_1077699;
  reg [7:0] p5_array_index_1077700;
  reg [7:0] p5_array_index_1077701;
  reg [7:0] p5_res7__533;
  reg [7:0] p5_array_index_1077713;
  reg [7:0] p5_array_index_1077714;
  reg [7:0] p5_array_index_1077715;
  reg [7:0] p5_res7__534;
  reg [7:0] p5_array_index_1077725;
  reg [7:0] p5_array_index_1077726;
  reg [7:0] p5_array_index_1077727;
  reg [7:0] p5_res7__535;
  reg [7:0] p5_array_index_1077738;
  reg [7:0] p5_array_index_1077739;
  reg [7:0] p5_res7__536;
  reg [7:0] p5_array_index_1077749;
  reg [7:0] p5_array_index_1077750;
  reg [7:0] p5_res7__537;
  reg [7:0] p6_arr[256];
  reg [7:0] p6_literal_1076345[256];
  reg [7:0] p6_literal_1076347[256];
  reg [7:0] p6_literal_1076349[256];
  reg [7:0] p6_literal_1076351[256];
  reg [7:0] p6_literal_1076353[256];
  reg [7:0] p6_literal_1076355[256];
  reg [7:0] p6_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p5_bit_slice_1076328 <= p4_bit_slice_1076328;
    p5_xor_1077141 <= p4_xor_1077141;
    p5_array_index_1077272 <= p4_array_index_1077272;
    p5_array_index_1077273 <= p4_array_index_1077273;
    p5_array_index_1077274 <= p4_array_index_1077274;
    p5_array_index_1077275 <= p4_array_index_1077275;
    p5_array_index_1077276 <= p4_array_index_1077276;
    p5_array_index_1077277 <= p4_array_index_1077277;
    p5_array_index_1077288 <= p4_array_index_1077288;
    p5_array_index_1077289 <= p4_array_index_1077289;
    p5_array_index_1077290 <= p4_array_index_1077290;
    p5_res7__16 <= p4_res7__16;
    p5_array_index_1077305 <= p4_array_index_1077305;
    p5_array_index_1077306 <= p4_array_index_1077306;
    p5_array_index_1077307 <= p4_array_index_1077307;
    p5_res7__17 <= p4_res7__17;
    p5_array_index_1077320 <= p4_array_index_1077320;
    p5_array_index_1077321 <= p4_array_index_1077321;
    p5_array_index_1077322 <= p4_array_index_1077322;
    p5_res7__18 <= p4_res7__18;
    p5_array_index_1077334 <= p4_array_index_1077334;
    p5_array_index_1077335 <= p4_array_index_1077335;
    p5_array_index_1077336 <= p4_array_index_1077336;
    p5_res7__19 <= p4_res7__19;
    p5_array_index_1077349 <= p4_array_index_1077349;
    p5_array_index_1077350 <= p4_array_index_1077350;
    p5_array_index_1077351 <= p4_array_index_1077351;
    p5_res7__20 <= p4_res7__20;
    p5_array_index_1077631 <= p5_array_index_1077631_comb;
    p5_array_index_1077632 <= p5_array_index_1077632_comb;
    p5_array_index_1077633 <= p5_array_index_1077633_comb;
    p5_res7__21 <= p5_res7__21_comb;
    p5_array_index_1077645 <= p5_array_index_1077645_comb;
    p5_array_index_1077646 <= p5_array_index_1077646_comb;
    p5_array_index_1077647 <= p5_array_index_1077647_comb;
    p5_res7__22 <= p5_res7__22_comb;
    p5_array_index_1077657 <= p5_array_index_1077657_comb;
    p5_array_index_1077658 <= p5_array_index_1077658_comb;
    p5_array_index_1077659 <= p5_array_index_1077659_comb;
    p5_res7__23 <= p5_res7__23_comb;
    p5_array_index_1077670 <= p5_array_index_1077670_comb;
    p5_array_index_1077671 <= p5_array_index_1077671_comb;
    p5_res7__24 <= p5_res7__24_comb;
    p5_array_index_1077681 <= p5_array_index_1077681_comb;
    p5_array_index_1077682 <= p5_array_index_1077682_comb;
    p5_res7__25 <= p5_res7__25_comb;
    p5_array_index_1077688 <= p5_array_index_1077688_comb;
    p5_array_index_1077689 <= p5_array_index_1077689_comb;
    p5_array_index_1077690 <= p5_array_index_1077690_comb;
    p5_array_index_1077691 <= p5_array_index_1077691_comb;
    p5_array_index_1077692 <= p5_array_index_1077692_comb;
    p5_array_index_1077693 <= p5_array_index_1077693_comb;
    p5_array_index_1077694 <= p5_array_index_1077694_comb;
    p5_array_index_1077695 <= p5_array_index_1077695_comb;
    p5_array_index_1077696 <= p5_array_index_1077696_comb;
    p5_array_index_1077360 <= p4_array_index_1077360;
    p5_array_index_1077361 <= p4_array_index_1077361;
    p5_array_index_1077362 <= p4_array_index_1077362;
    p5_array_index_1077363 <= p4_array_index_1077363;
    p5_array_index_1077364 <= p4_array_index_1077364;
    p5_array_index_1077365 <= p4_array_index_1077365;
    p5_array_index_1077373 <= p4_array_index_1077373;
    p5_array_index_1077374 <= p4_array_index_1077374;
    p5_array_index_1077375 <= p4_array_index_1077375;
    p5_res7__528 <= p4_res7__528;
    p5_array_index_1077390 <= p4_array_index_1077390;
    p5_array_index_1077391 <= p4_array_index_1077391;
    p5_array_index_1077392 <= p4_array_index_1077392;
    p5_res7__529 <= p4_res7__529;
    p5_array_index_1077405 <= p4_array_index_1077405;
    p5_array_index_1077406 <= p4_array_index_1077406;
    p5_array_index_1077407 <= p4_array_index_1077407;
    p5_res7__530 <= p4_res7__530;
    p5_array_index_1077419 <= p4_array_index_1077419;
    p5_array_index_1077420 <= p4_array_index_1077420;
    p5_array_index_1077421 <= p4_array_index_1077421;
    p5_res7__531 <= p4_res7__531;
    p5_array_index_1077434 <= p4_array_index_1077434;
    p5_array_index_1077435 <= p4_array_index_1077435;
    p5_array_index_1077436 <= p4_array_index_1077436;
    p5_res7__532 <= p4_res7__532;
    p5_array_index_1077699 <= p5_array_index_1077699_comb;
    p5_array_index_1077700 <= p5_array_index_1077700_comb;
    p5_array_index_1077701 <= p5_array_index_1077701_comb;
    p5_res7__533 <= p5_res7__533_comb;
    p5_array_index_1077713 <= p5_array_index_1077713_comb;
    p5_array_index_1077714 <= p5_array_index_1077714_comb;
    p5_array_index_1077715 <= p5_array_index_1077715_comb;
    p5_res7__534 <= p5_res7__534_comb;
    p5_array_index_1077725 <= p5_array_index_1077725_comb;
    p5_array_index_1077726 <= p5_array_index_1077726_comb;
    p5_array_index_1077727 <= p5_array_index_1077727_comb;
    p5_res7__535 <= p5_res7__535_comb;
    p5_array_index_1077738 <= p5_array_index_1077738_comb;
    p5_array_index_1077739 <= p5_array_index_1077739_comb;
    p5_res7__536 <= p5_res7__536_comb;
    p5_array_index_1077749 <= p5_array_index_1077749_comb;
    p5_array_index_1077750 <= p5_array_index_1077750_comb;
    p5_res7__537 <= p5_res7__537_comb;
    p6_arr <= p5_arr;
    p6_literal_1076345 <= p5_literal_1076345;
    p6_literal_1076347 <= p5_literal_1076347;
    p6_literal_1076349 <= p5_literal_1076349;
    p6_literal_1076351 <= p5_literal_1076351;
    p6_literal_1076353 <= p5_literal_1076353;
    p6_literal_1076355 <= p5_literal_1076355;
    p6_literal_1076358 <= p5_literal_1076358;
  end

  // ===== Pipe stage 6:
  wire [7:0] p6_res7__26_comb;
  wire [7:0] p6_array_index_1077976_comb;
  wire [7:0] p6_res7__27_comb;
  wire [7:0] p6_array_index_1078022_comb;
  wire [7:0] p6_res7__28_comb;
  wire [7:0] p6_res7__538_comb;
  wire [7:0] p6_array_index_1078032_comb;
  wire [7:0] p6_res7__29_comb;
  wire [7:0] p6_res7__539_comb;
  wire [7:0] p6_res7__30_comb;
  wire [7:0] p6_res7__540_comb;
  wire [7:0] p6_res7__31_comb;
  wire [7:0] p6_res7__541_comb;
  wire [127:0] p6_res__1_comb;
  wire [127:0] p6_xor_1078016_comb;
  wire [7:0] p6_res7__542_comb;
  assign p6_res7__26_comb = p5_array_index_1077688 ^ p5_array_index_1077689 ^ p5_array_index_1077690 ^ p5_array_index_1077691 ^ p5_array_index_1077692 ^ p5_array_index_1077693 ^ p5_res7__19 ^ p5_array_index_1077694 ^ p5_res7__17 ^ p5_array_index_1077647 ^ p5_array_index_1077351 ^ p5_array_index_1077322 ^ p5_array_index_1077290 ^ p5_array_index_1077695 ^ p5_array_index_1077696 ^ p5_array_index_1077277;
  assign p6_array_index_1077976_comb = p5_literal_1076355[p5_res7__21];
  assign p6_res7__27_comb = p5_literal_1076345[p6_res7__26_comb] ^ p5_literal_1076347[p5_res7__25] ^ p5_literal_1076349[p5_res7__24] ^ p5_literal_1076351[p5_res7__23] ^ p5_literal_1076353[p5_res7__22] ^ p6_array_index_1077976_comb ^ p5_res7__20 ^ p5_literal_1076358[p5_res7__19] ^ p5_res7__18 ^ p5_array_index_1077659 ^ p5_array_index_1077633 ^ p5_array_index_1077336 ^ p5_array_index_1077307 ^ p5_literal_1076347[p5_array_index_1077274] ^ p5_literal_1076345[p5_array_index_1077275] ^ p5_array_index_1077276;
  assign p6_array_index_1078022_comb = p5_literal_1076355[p5_res7__532];
  assign p6_res7__28_comb = p5_literal_1076345[p6_res7__27_comb] ^ p5_literal_1076347[p6_res7__26_comb] ^ p5_literal_1076349[p5_res7__25] ^ p5_literal_1076351[p5_res7__24] ^ p5_literal_1076353[p5_res7__23] ^ p5_literal_1076355[p5_res7__22] ^ p5_res7__21 ^ p5_literal_1076358[p5_res7__20] ^ p5_res7__19 ^ p5_array_index_1077671 ^ p5_array_index_1077646 ^ p5_array_index_1077350 ^ p5_array_index_1077321 ^ p5_array_index_1077289 ^ p5_literal_1076345[p5_array_index_1077274] ^ p5_array_index_1077275;
  assign p6_res7__538_comb = p5_literal_1076345[p5_res7__537] ^ p5_literal_1076347[p5_res7__536] ^ p5_literal_1076349[p5_res7__535] ^ p5_literal_1076351[p5_res7__534] ^ p5_literal_1076353[p5_res7__533] ^ p6_array_index_1078022_comb ^ p5_res7__531 ^ p5_literal_1076358[p5_res7__530] ^ p5_res7__529 ^ p5_array_index_1077715 ^ p5_array_index_1077436 ^ p5_array_index_1077407 ^ p5_array_index_1077375 ^ p5_literal_1076347[p5_array_index_1077363] ^ p5_literal_1076345[p5_array_index_1077364] ^ p5_array_index_1077365;
  assign p6_array_index_1078032_comb = p5_literal_1076355[p5_res7__533];
  assign p6_res7__29_comb = p5_literal_1076345[p6_res7__28_comb] ^ p5_literal_1076347[p6_res7__27_comb] ^ p5_literal_1076349[p6_res7__26_comb] ^ p5_literal_1076351[p5_res7__25] ^ p5_literal_1076353[p5_res7__24] ^ p5_literal_1076355[p5_res7__23] ^ p5_res7__22 ^ p5_literal_1076358[p5_res7__21] ^ p5_res7__20 ^ p5_array_index_1077682 ^ p5_array_index_1077658 ^ p5_array_index_1077632 ^ p5_array_index_1077335 ^ p5_array_index_1077306 ^ p5_literal_1076345[p5_array_index_1077273] ^ p5_array_index_1077274;
  assign p6_res7__539_comb = p5_literal_1076345[p6_res7__538_comb] ^ p5_literal_1076347[p5_res7__537] ^ p5_literal_1076349[p5_res7__536] ^ p5_literal_1076351[p5_res7__535] ^ p5_literal_1076353[p5_res7__534] ^ p6_array_index_1078032_comb ^ p5_res7__532 ^ p5_literal_1076358[p5_res7__531] ^ p5_res7__530 ^ p5_array_index_1077727 ^ p5_array_index_1077701 ^ p5_array_index_1077421 ^ p5_array_index_1077392 ^ p5_literal_1076347[p5_array_index_1077362] ^ p5_literal_1076345[p5_array_index_1077363] ^ p5_array_index_1077364;
  assign p6_res7__30_comb = p5_literal_1076345[p6_res7__29_comb] ^ p5_literal_1076347[p6_res7__28_comb] ^ p5_literal_1076349[p6_res7__27_comb] ^ p5_literal_1076351[p6_res7__26_comb] ^ p5_literal_1076353[p5_res7__25] ^ p5_literal_1076355[p5_res7__24] ^ p5_res7__23 ^ p5_literal_1076358[p5_res7__22] ^ p5_res7__21 ^ p5_array_index_1077693 ^ p5_array_index_1077670 ^ p5_array_index_1077645 ^ p5_array_index_1077349 ^ p5_array_index_1077320 ^ p5_array_index_1077288 ^ p5_array_index_1077273;
  assign p6_res7__540_comb = p5_literal_1076345[p6_res7__539_comb] ^ p5_literal_1076347[p6_res7__538_comb] ^ p5_literal_1076349[p5_res7__537] ^ p5_literal_1076351[p5_res7__536] ^ p5_literal_1076353[p5_res7__535] ^ p5_literal_1076355[p5_res7__534] ^ p5_res7__533 ^ p5_literal_1076358[p5_res7__532] ^ p5_res7__531 ^ p5_array_index_1077739 ^ p5_array_index_1077714 ^ p5_array_index_1077435 ^ p5_array_index_1077406 ^ p5_array_index_1077374 ^ p5_literal_1076345[p5_array_index_1077362] ^ p5_array_index_1077363;
  assign p6_res7__31_comb = p5_literal_1076345[p6_res7__30_comb] ^ p5_literal_1076347[p6_res7__29_comb] ^ p5_literal_1076349[p6_res7__28_comb] ^ p5_literal_1076351[p6_res7__27_comb] ^ p5_literal_1076353[p6_res7__26_comb] ^ p5_literal_1076355[p5_res7__25] ^ p5_res7__24 ^ p5_literal_1076358[p5_res7__23] ^ p5_res7__22 ^ p6_array_index_1077976_comb ^ p5_array_index_1077681 ^ p5_array_index_1077657 ^ p5_array_index_1077631 ^ p5_array_index_1077334 ^ p5_array_index_1077305 ^ p5_array_index_1077272;
  assign p6_res7__541_comb = p5_literal_1076345[p6_res7__540_comb] ^ p5_literal_1076347[p6_res7__539_comb] ^ p5_literal_1076349[p6_res7__538_comb] ^ p5_literal_1076351[p5_res7__537] ^ p5_literal_1076353[p5_res7__536] ^ p5_literal_1076355[p5_res7__535] ^ p5_res7__534 ^ p5_literal_1076358[p5_res7__533] ^ p5_res7__532 ^ p5_array_index_1077750 ^ p5_array_index_1077726 ^ p5_array_index_1077700 ^ p5_array_index_1077420 ^ p5_array_index_1077391 ^ p5_literal_1076345[p5_array_index_1077361] ^ p5_array_index_1077362;
  assign p6_res__1_comb = {p6_res7__31_comb, p6_res7__30_comb, p6_res7__29_comb, p6_res7__28_comb, p6_res7__27_comb, p6_res7__26_comb, p5_res7__25, p5_res7__24, p5_res7__23, p5_res7__22, p5_res7__21, p5_res7__20, p5_res7__19, p5_res7__18, p5_res7__17, p5_res7__16};
  assign p6_xor_1078016_comb = p6_res__1_comb ^ p5_bit_slice_1076328;
  assign p6_res7__542_comb = p5_literal_1076345[p6_res7__541_comb] ^ p5_literal_1076347[p6_res7__540_comb] ^ p5_literal_1076349[p6_res7__539_comb] ^ p5_literal_1076351[p6_res7__538_comb] ^ p5_literal_1076353[p5_res7__537] ^ p5_literal_1076355[p5_res7__536] ^ p5_res7__535 ^ p5_literal_1076358[p5_res7__534] ^ p5_res7__533 ^ p6_array_index_1078022_comb ^ p5_array_index_1077738 ^ p5_array_index_1077713 ^ p5_array_index_1077434 ^ p5_array_index_1077405 ^ p5_array_index_1077373 ^ p5_array_index_1077361;

  // Registers for pipe stage 6:
  reg [127:0] p6_xor_1077141;
  reg [127:0] p6_xor_1078016;
  reg [7:0] p6_array_index_1077360;
  reg [7:0] p6_res7__528;
  reg [7:0] p6_array_index_1077390;
  reg [7:0] p6_res7__529;
  reg [7:0] p6_res7__530;
  reg [7:0] p6_array_index_1077419;
  reg [7:0] p6_res7__531;
  reg [7:0] p6_res7__532;
  reg [7:0] p6_array_index_1077699;
  reg [7:0] p6_res7__533;
  reg [7:0] p6_res7__534;
  reg [7:0] p6_array_index_1077725;
  reg [7:0] p6_res7__535;
  reg [7:0] p6_res7__536;
  reg [7:0] p6_array_index_1077749;
  reg [7:0] p6_res7__537;
  reg [7:0] p6_res7__538;
  reg [7:0] p6_array_index_1078032;
  reg [7:0] p6_res7__539;
  reg [7:0] p6_res7__540;
  reg [7:0] p6_res7__541;
  reg [7:0] p6_res7__542;
  reg [7:0] p7_arr[256];
  reg [7:0] p7_literal_1076345[256];
  reg [7:0] p7_literal_1076347[256];
  reg [7:0] p7_literal_1076349[256];
  reg [7:0] p7_literal_1076351[256];
  reg [7:0] p7_literal_1076353[256];
  reg [7:0] p7_literal_1076355[256];
  reg [7:0] p7_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p6_xor_1077141 <= p5_xor_1077141;
    p6_xor_1078016 <= p6_xor_1078016_comb;
    p6_array_index_1077360 <= p5_array_index_1077360;
    p6_res7__528 <= p5_res7__528;
    p6_array_index_1077390 <= p5_array_index_1077390;
    p6_res7__529 <= p5_res7__529;
    p6_res7__530 <= p5_res7__530;
    p6_array_index_1077419 <= p5_array_index_1077419;
    p6_res7__531 <= p5_res7__531;
    p6_res7__532 <= p5_res7__532;
    p6_array_index_1077699 <= p5_array_index_1077699;
    p6_res7__533 <= p5_res7__533;
    p6_res7__534 <= p5_res7__534;
    p6_array_index_1077725 <= p5_array_index_1077725;
    p6_res7__535 <= p5_res7__535;
    p6_res7__536 <= p5_res7__536;
    p6_array_index_1077749 <= p5_array_index_1077749;
    p6_res7__537 <= p5_res7__537;
    p6_res7__538 <= p6_res7__538_comb;
    p6_array_index_1078032 <= p6_array_index_1078032_comb;
    p6_res7__539 <= p6_res7__539_comb;
    p6_res7__540 <= p6_res7__540_comb;
    p6_res7__541 <= p6_res7__541_comb;
    p6_res7__542 <= p6_res7__542_comb;
    p7_arr <= p6_arr;
    p7_literal_1076345 <= p6_literal_1076345;
    p7_literal_1076347 <= p6_literal_1076347;
    p7_literal_1076349 <= p6_literal_1076349;
    p7_literal_1076351 <= p6_literal_1076351;
    p7_literal_1076353 <= p6_literal_1076353;
    p7_literal_1076355 <= p6_literal_1076355;
    p7_literal_1076358 <= p6_literal_1076358;
  end

  // ===== Pipe stage 7:
  wire [127:0] p7_addedKey__43_comb;
  wire [7:0] p7_array_index_1078142_comb;
  wire [7:0] p7_array_index_1078143_comb;
  wire [7:0] p7_array_index_1078144_comb;
  wire [7:0] p7_array_index_1078145_comb;
  wire [7:0] p7_array_index_1078146_comb;
  wire [7:0] p7_array_index_1078147_comb;
  wire [7:0] p7_array_index_1078149_comb;
  wire [7:0] p7_array_index_1078151_comb;
  wire [7:0] p7_array_index_1078152_comb;
  wire [7:0] p7_array_index_1078153_comb;
  wire [7:0] p7_array_index_1078154_comb;
  wire [7:0] p7_array_index_1078155_comb;
  wire [7:0] p7_array_index_1078156_comb;
  wire [7:0] p7_array_index_1078158_comb;
  wire [7:0] p7_array_index_1078159_comb;
  wire [7:0] p7_array_index_1078160_comb;
  wire [7:0] p7_array_index_1078161_comb;
  wire [7:0] p7_array_index_1078162_comb;
  wire [7:0] p7_array_index_1078163_comb;
  wire [7:0] p7_array_index_1078164_comb;
  wire [7:0] p7_array_index_1078166_comb;
  wire [7:0] p7_res7__32_comb;
  wire [7:0] p7_array_index_1078175_comb;
  wire [7:0] p7_array_index_1078176_comb;
  wire [7:0] p7_array_index_1078177_comb;
  wire [7:0] p7_array_index_1078178_comb;
  wire [7:0] p7_array_index_1078179_comb;
  wire [7:0] p7_array_index_1078180_comb;
  wire [7:0] p7_res7__33_comb;
  wire [7:0] p7_array_index_1078190_comb;
  wire [7:0] p7_array_index_1078191_comb;
  wire [7:0] p7_array_index_1078192_comb;
  wire [7:0] p7_array_index_1078193_comb;
  wire [7:0] p7_array_index_1078194_comb;
  wire [7:0] p7_res7__34_comb;
  wire [7:0] p7_array_index_1078204_comb;
  wire [7:0] p7_array_index_1078205_comb;
  wire [7:0] p7_array_index_1078206_comb;
  wire [7:0] p7_array_index_1078207_comb;
  wire [7:0] p7_array_index_1078208_comb;
  wire [7:0] p7_res7__35_comb;
  wire [7:0] p7_array_index_1078219_comb;
  wire [7:0] p7_array_index_1078220_comb;
  wire [7:0] p7_array_index_1078221_comb;
  wire [7:0] p7_array_index_1078222_comb;
  wire [7:0] p7_res7__543_comb;
  wire [7:0] p7_res7__36_comb;
  wire [127:0] p7_res__33_comb;
  assign p7_addedKey__43_comb = p6_xor_1078016 ^ 128'hb225_9a96_b4d8_8e0b_e769_0430_a44f_7f03;
  assign p7_array_index_1078142_comb = p6_arr[p7_addedKey__43_comb[127:120]];
  assign p7_array_index_1078143_comb = p6_arr[p7_addedKey__43_comb[119:112]];
  assign p7_array_index_1078144_comb = p6_arr[p7_addedKey__43_comb[111:104]];
  assign p7_array_index_1078145_comb = p6_arr[p7_addedKey__43_comb[103:96]];
  assign p7_array_index_1078146_comb = p6_arr[p7_addedKey__43_comb[95:88]];
  assign p7_array_index_1078147_comb = p6_arr[p7_addedKey__43_comb[87:80]];
  assign p7_array_index_1078149_comb = p6_arr[p7_addedKey__43_comb[71:64]];
  assign p7_array_index_1078151_comb = p6_arr[p7_addedKey__43_comb[55:48]];
  assign p7_array_index_1078152_comb = p6_arr[p7_addedKey__43_comb[47:40]];
  assign p7_array_index_1078153_comb = p6_arr[p7_addedKey__43_comb[39:32]];
  assign p7_array_index_1078154_comb = p6_arr[p7_addedKey__43_comb[31:24]];
  assign p7_array_index_1078155_comb = p6_arr[p7_addedKey__43_comb[23:16]];
  assign p7_array_index_1078156_comb = p6_arr[p7_addedKey__43_comb[15:8]];
  assign p7_array_index_1078158_comb = p6_literal_1076345[p7_array_index_1078142_comb];
  assign p7_array_index_1078159_comb = p6_literal_1076347[p7_array_index_1078143_comb];
  assign p7_array_index_1078160_comb = p6_literal_1076349[p7_array_index_1078144_comb];
  assign p7_array_index_1078161_comb = p6_literal_1076351[p7_array_index_1078145_comb];
  assign p7_array_index_1078162_comb = p6_literal_1076353[p7_array_index_1078146_comb];
  assign p7_array_index_1078163_comb = p6_literal_1076355[p7_array_index_1078147_comb];
  assign p7_array_index_1078164_comb = p6_arr[p7_addedKey__43_comb[79:72]];
  assign p7_array_index_1078166_comb = p6_arr[p7_addedKey__43_comb[63:56]];
  assign p7_res7__32_comb = p7_array_index_1078158_comb ^ p7_array_index_1078159_comb ^ p7_array_index_1078160_comb ^ p7_array_index_1078161_comb ^ p7_array_index_1078162_comb ^ p7_array_index_1078163_comb ^ p7_array_index_1078164_comb ^ p6_literal_1076358[p7_array_index_1078149_comb] ^ p7_array_index_1078166_comb ^ p6_literal_1076355[p7_array_index_1078151_comb] ^ p6_literal_1076353[p7_array_index_1078152_comb] ^ p6_literal_1076351[p7_array_index_1078153_comb] ^ p6_literal_1076349[p7_array_index_1078154_comb] ^ p6_literal_1076347[p7_array_index_1078155_comb] ^ p6_literal_1076345[p7_array_index_1078156_comb] ^ p6_arr[p7_addedKey__43_comb[7:0]];
  assign p7_array_index_1078175_comb = p6_literal_1076345[p7_res7__32_comb];
  assign p7_array_index_1078176_comb = p6_literal_1076347[p7_array_index_1078142_comb];
  assign p7_array_index_1078177_comb = p6_literal_1076349[p7_array_index_1078143_comb];
  assign p7_array_index_1078178_comb = p6_literal_1076351[p7_array_index_1078144_comb];
  assign p7_array_index_1078179_comb = p6_literal_1076353[p7_array_index_1078145_comb];
  assign p7_array_index_1078180_comb = p6_literal_1076355[p7_array_index_1078146_comb];
  assign p7_res7__33_comb = p7_array_index_1078175_comb ^ p7_array_index_1078176_comb ^ p7_array_index_1078177_comb ^ p7_array_index_1078178_comb ^ p7_array_index_1078179_comb ^ p7_array_index_1078180_comb ^ p7_array_index_1078147_comb ^ p6_literal_1076358[p7_array_index_1078164_comb] ^ p7_array_index_1078149_comb ^ p6_literal_1076355[p7_array_index_1078166_comb] ^ p6_literal_1076353[p7_array_index_1078151_comb] ^ p6_literal_1076351[p7_array_index_1078152_comb] ^ p6_literal_1076349[p7_array_index_1078153_comb] ^ p6_literal_1076347[p7_array_index_1078154_comb] ^ p6_literal_1076345[p7_array_index_1078155_comb] ^ p7_array_index_1078156_comb;
  assign p7_array_index_1078190_comb = p6_literal_1076347[p7_res7__32_comb];
  assign p7_array_index_1078191_comb = p6_literal_1076349[p7_array_index_1078142_comb];
  assign p7_array_index_1078192_comb = p6_literal_1076351[p7_array_index_1078143_comb];
  assign p7_array_index_1078193_comb = p6_literal_1076353[p7_array_index_1078144_comb];
  assign p7_array_index_1078194_comb = p6_literal_1076355[p7_array_index_1078145_comb];
  assign p7_res7__34_comb = p6_literal_1076345[p7_res7__33_comb] ^ p7_array_index_1078190_comb ^ p7_array_index_1078191_comb ^ p7_array_index_1078192_comb ^ p7_array_index_1078193_comb ^ p7_array_index_1078194_comb ^ p7_array_index_1078146_comb ^ p6_literal_1076358[p7_array_index_1078147_comb] ^ p7_array_index_1078164_comb ^ p6_literal_1076355[p7_array_index_1078149_comb] ^ p6_literal_1076353[p7_array_index_1078166_comb] ^ p6_literal_1076351[p7_array_index_1078151_comb] ^ p6_literal_1076349[p7_array_index_1078152_comb] ^ p6_literal_1076347[p7_array_index_1078153_comb] ^ p6_literal_1076345[p7_array_index_1078154_comb] ^ p7_array_index_1078155_comb;
  assign p7_array_index_1078204_comb = p6_literal_1076347[p7_res7__33_comb];
  assign p7_array_index_1078205_comb = p6_literal_1076349[p7_res7__32_comb];
  assign p7_array_index_1078206_comb = p6_literal_1076351[p7_array_index_1078142_comb];
  assign p7_array_index_1078207_comb = p6_literal_1076353[p7_array_index_1078143_comb];
  assign p7_array_index_1078208_comb = p6_literal_1076355[p7_array_index_1078144_comb];
  assign p7_res7__35_comb = p6_literal_1076345[p7_res7__34_comb] ^ p7_array_index_1078204_comb ^ p7_array_index_1078205_comb ^ p7_array_index_1078206_comb ^ p7_array_index_1078207_comb ^ p7_array_index_1078208_comb ^ p7_array_index_1078145_comb ^ p6_literal_1076358[p7_array_index_1078146_comb] ^ p7_array_index_1078147_comb ^ p6_literal_1076355[p7_array_index_1078164_comb] ^ p6_literal_1076353[p7_array_index_1078149_comb] ^ p6_literal_1076351[p7_array_index_1078166_comb] ^ p6_literal_1076349[p7_array_index_1078151_comb] ^ p6_literal_1076347[p7_array_index_1078152_comb] ^ p6_literal_1076345[p7_array_index_1078153_comb] ^ p7_array_index_1078154_comb;
  assign p7_array_index_1078219_comb = p6_literal_1076349[p7_res7__33_comb];
  assign p7_array_index_1078220_comb = p6_literal_1076351[p7_res7__32_comb];
  assign p7_array_index_1078221_comb = p6_literal_1076353[p7_array_index_1078142_comb];
  assign p7_array_index_1078222_comb = p6_literal_1076355[p7_array_index_1078143_comb];
  assign p7_res7__543_comb = p6_literal_1076345[p6_res7__542] ^ p6_literal_1076347[p6_res7__541] ^ p6_literal_1076349[p6_res7__540] ^ p6_literal_1076351[p6_res7__539] ^ p6_literal_1076353[p6_res7__538] ^ p6_literal_1076355[p6_res7__537] ^ p6_res7__536 ^ p6_literal_1076358[p6_res7__535] ^ p6_res7__534 ^ p6_array_index_1078032 ^ p6_array_index_1077749 ^ p6_array_index_1077725 ^ p6_array_index_1077699 ^ p6_array_index_1077419 ^ p6_array_index_1077390 ^ p6_array_index_1077360;
  assign p7_res7__36_comb = p6_literal_1076345[p7_res7__35_comb] ^ p6_literal_1076347[p7_res7__34_comb] ^ p7_array_index_1078219_comb ^ p7_array_index_1078220_comb ^ p7_array_index_1078221_comb ^ p7_array_index_1078222_comb ^ p7_array_index_1078144_comb ^ p6_literal_1076358[p7_array_index_1078145_comb] ^ p7_array_index_1078146_comb ^ p7_array_index_1078163_comb ^ p6_literal_1076353[p7_array_index_1078164_comb] ^ p6_literal_1076351[p7_array_index_1078149_comb] ^ p6_literal_1076349[p7_array_index_1078166_comb] ^ p6_literal_1076347[p7_array_index_1078151_comb] ^ p6_literal_1076345[p7_array_index_1078152_comb] ^ p7_array_index_1078153_comb;
  assign p7_res__33_comb = {p7_res7__543_comb, p6_res7__542, p6_res7__541, p6_res7__540, p6_res7__539, p6_res7__538, p6_res7__537, p6_res7__536, p6_res7__535, p6_res7__534, p6_res7__533, p6_res7__532, p6_res7__531, p6_res7__530, p6_res7__529, p6_res7__528};

  // Registers for pipe stage 7:
  reg [127:0] p7_xor_1077141;
  reg [127:0] p7_xor_1078016;
  reg [7:0] p7_array_index_1078142;
  reg [7:0] p7_array_index_1078143;
  reg [7:0] p7_array_index_1078144;
  reg [7:0] p7_array_index_1078145;
  reg [7:0] p7_array_index_1078146;
  reg [7:0] p7_array_index_1078147;
  reg [7:0] p7_array_index_1078149;
  reg [7:0] p7_array_index_1078151;
  reg [7:0] p7_array_index_1078152;
  reg [7:0] p7_array_index_1078158;
  reg [7:0] p7_array_index_1078159;
  reg [7:0] p7_array_index_1078160;
  reg [7:0] p7_array_index_1078161;
  reg [7:0] p7_array_index_1078162;
  reg [7:0] p7_array_index_1078164;
  reg [7:0] p7_array_index_1078166;
  reg [7:0] p7_res7__32;
  reg [7:0] p7_array_index_1078175;
  reg [7:0] p7_array_index_1078176;
  reg [7:0] p7_array_index_1078177;
  reg [7:0] p7_array_index_1078178;
  reg [7:0] p7_array_index_1078179;
  reg [7:0] p7_array_index_1078180;
  reg [7:0] p7_res7__33;
  reg [7:0] p7_array_index_1078190;
  reg [7:0] p7_array_index_1078191;
  reg [7:0] p7_array_index_1078192;
  reg [7:0] p7_array_index_1078193;
  reg [7:0] p7_array_index_1078194;
  reg [7:0] p7_res7__34;
  reg [7:0] p7_array_index_1078204;
  reg [7:0] p7_array_index_1078205;
  reg [7:0] p7_array_index_1078206;
  reg [7:0] p7_array_index_1078207;
  reg [7:0] p7_array_index_1078208;
  reg [7:0] p7_res7__35;
  reg [7:0] p7_array_index_1078219;
  reg [7:0] p7_array_index_1078220;
  reg [7:0] p7_array_index_1078221;
  reg [7:0] p7_array_index_1078222;
  reg [7:0] p7_res7__36;
  reg [127:0] p7_res__33;
  reg [7:0] p8_arr[256];
  reg [7:0] p8_literal_1076345[256];
  reg [7:0] p8_literal_1076347[256];
  reg [7:0] p8_literal_1076349[256];
  reg [7:0] p8_literal_1076351[256];
  reg [7:0] p8_literal_1076353[256];
  reg [7:0] p8_literal_1076355[256];
  reg [7:0] p8_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p7_xor_1077141 <= p6_xor_1077141;
    p7_xor_1078016 <= p6_xor_1078016;
    p7_array_index_1078142 <= p7_array_index_1078142_comb;
    p7_array_index_1078143 <= p7_array_index_1078143_comb;
    p7_array_index_1078144 <= p7_array_index_1078144_comb;
    p7_array_index_1078145 <= p7_array_index_1078145_comb;
    p7_array_index_1078146 <= p7_array_index_1078146_comb;
    p7_array_index_1078147 <= p7_array_index_1078147_comb;
    p7_array_index_1078149 <= p7_array_index_1078149_comb;
    p7_array_index_1078151 <= p7_array_index_1078151_comb;
    p7_array_index_1078152 <= p7_array_index_1078152_comb;
    p7_array_index_1078158 <= p7_array_index_1078158_comb;
    p7_array_index_1078159 <= p7_array_index_1078159_comb;
    p7_array_index_1078160 <= p7_array_index_1078160_comb;
    p7_array_index_1078161 <= p7_array_index_1078161_comb;
    p7_array_index_1078162 <= p7_array_index_1078162_comb;
    p7_array_index_1078164 <= p7_array_index_1078164_comb;
    p7_array_index_1078166 <= p7_array_index_1078166_comb;
    p7_res7__32 <= p7_res7__32_comb;
    p7_array_index_1078175 <= p7_array_index_1078175_comb;
    p7_array_index_1078176 <= p7_array_index_1078176_comb;
    p7_array_index_1078177 <= p7_array_index_1078177_comb;
    p7_array_index_1078178 <= p7_array_index_1078178_comb;
    p7_array_index_1078179 <= p7_array_index_1078179_comb;
    p7_array_index_1078180 <= p7_array_index_1078180_comb;
    p7_res7__33 <= p7_res7__33_comb;
    p7_array_index_1078190 <= p7_array_index_1078190_comb;
    p7_array_index_1078191 <= p7_array_index_1078191_comb;
    p7_array_index_1078192 <= p7_array_index_1078192_comb;
    p7_array_index_1078193 <= p7_array_index_1078193_comb;
    p7_array_index_1078194 <= p7_array_index_1078194_comb;
    p7_res7__34 <= p7_res7__34_comb;
    p7_array_index_1078204 <= p7_array_index_1078204_comb;
    p7_array_index_1078205 <= p7_array_index_1078205_comb;
    p7_array_index_1078206 <= p7_array_index_1078206_comb;
    p7_array_index_1078207 <= p7_array_index_1078207_comb;
    p7_array_index_1078208 <= p7_array_index_1078208_comb;
    p7_res7__35 <= p7_res7__35_comb;
    p7_array_index_1078219 <= p7_array_index_1078219_comb;
    p7_array_index_1078220 <= p7_array_index_1078220_comb;
    p7_array_index_1078221 <= p7_array_index_1078221_comb;
    p7_array_index_1078222 <= p7_array_index_1078222_comb;
    p7_res7__36 <= p7_res7__36_comb;
    p7_res__33 <= p7_res__33_comb;
    p8_arr <= p7_arr;
    p8_literal_1076345 <= p7_literal_1076345;
    p8_literal_1076347 <= p7_literal_1076347;
    p8_literal_1076349 <= p7_literal_1076349;
    p8_literal_1076351 <= p7_literal_1076351;
    p8_literal_1076353 <= p7_literal_1076353;
    p8_literal_1076355 <= p7_literal_1076355;
    p8_literal_1076358 <= p7_literal_1076358;
  end

  // ===== Pipe stage 8:
  wire [7:0] p8_array_index_1078345_comb;
  wire [7:0] p8_array_index_1078346_comb;
  wire [7:0] p8_array_index_1078347_comb;
  wire [7:0] p8_array_index_1078348_comb;
  wire [7:0] p8_res7__37_comb;
  wire [7:0] p8_array_index_1078359_comb;
  wire [7:0] p8_array_index_1078360_comb;
  wire [7:0] p8_array_index_1078361_comb;
  wire [7:0] p8_res7__38_comb;
  wire [7:0] p8_array_index_1078371_comb;
  wire [7:0] p8_array_index_1078372_comb;
  wire [7:0] p8_array_index_1078373_comb;
  wire [7:0] p8_res7__39_comb;
  wire [7:0] p8_array_index_1078384_comb;
  wire [7:0] p8_array_index_1078385_comb;
  wire [7:0] p8_res7__40_comb;
  wire [7:0] p8_array_index_1078395_comb;
  wire [7:0] p8_array_index_1078396_comb;
  wire [7:0] p8_res7__41_comb;
  wire [7:0] p8_array_index_1078402_comb;
  wire [7:0] p8_array_index_1078403_comb;
  wire [7:0] p8_array_index_1078404_comb;
  wire [7:0] p8_array_index_1078405_comb;
  wire [7:0] p8_array_index_1078406_comb;
  wire [7:0] p8_array_index_1078407_comb;
  wire [7:0] p8_array_index_1078408_comb;
  wire [7:0] p8_array_index_1078409_comb;
  wire [7:0] p8_array_index_1078410_comb;
  assign p8_array_index_1078345_comb = p7_literal_1076349[p7_res7__34];
  assign p8_array_index_1078346_comb = p7_literal_1076351[p7_res7__33];
  assign p8_array_index_1078347_comb = p7_literal_1076353[p7_res7__32];
  assign p8_array_index_1078348_comb = p7_literal_1076355[p7_array_index_1078142];
  assign p8_res7__37_comb = p7_literal_1076345[p7_res7__36] ^ p7_literal_1076347[p7_res7__35] ^ p8_array_index_1078345_comb ^ p8_array_index_1078346_comb ^ p8_array_index_1078347_comb ^ p8_array_index_1078348_comb ^ p7_array_index_1078143 ^ p7_literal_1076358[p7_array_index_1078144] ^ p7_array_index_1078145 ^ p7_array_index_1078180 ^ p7_literal_1076353[p7_array_index_1078147] ^ p7_literal_1076351[p7_array_index_1078164] ^ p7_literal_1076349[p7_array_index_1078149] ^ p7_literal_1076347[p7_array_index_1078166] ^ p7_literal_1076345[p7_array_index_1078151] ^ p7_array_index_1078152;
  assign p8_array_index_1078359_comb = p7_literal_1076351[p7_res7__34];
  assign p8_array_index_1078360_comb = p7_literal_1076353[p7_res7__33];
  assign p8_array_index_1078361_comb = p7_literal_1076355[p7_res7__32];
  assign p8_res7__38_comb = p7_literal_1076345[p8_res7__37_comb] ^ p7_literal_1076347[p7_res7__36] ^ p7_literal_1076349[p7_res7__35] ^ p8_array_index_1078359_comb ^ p8_array_index_1078360_comb ^ p8_array_index_1078361_comb ^ p7_array_index_1078142 ^ p7_literal_1076358[p7_array_index_1078143] ^ p7_array_index_1078144 ^ p7_array_index_1078194 ^ p7_array_index_1078162 ^ p7_literal_1076351[p7_array_index_1078147] ^ p7_literal_1076349[p7_array_index_1078164] ^ p7_literal_1076347[p7_array_index_1078149] ^ p7_literal_1076345[p7_array_index_1078166] ^ p7_array_index_1078151;
  assign p8_array_index_1078371_comb = p7_literal_1076351[p7_res7__35];
  assign p8_array_index_1078372_comb = p7_literal_1076353[p7_res7__34];
  assign p8_array_index_1078373_comb = p7_literal_1076355[p7_res7__33];
  assign p8_res7__39_comb = p7_literal_1076345[p8_res7__38_comb] ^ p7_literal_1076347[p8_res7__37_comb] ^ p7_literal_1076349[p7_res7__36] ^ p8_array_index_1078371_comb ^ p8_array_index_1078372_comb ^ p8_array_index_1078373_comb ^ p7_res7__32 ^ p7_literal_1076358[p7_array_index_1078142] ^ p7_array_index_1078143 ^ p7_array_index_1078208 ^ p7_array_index_1078179 ^ p7_literal_1076351[p7_array_index_1078146] ^ p7_literal_1076349[p7_array_index_1078147] ^ p7_literal_1076347[p7_array_index_1078164] ^ p7_literal_1076345[p7_array_index_1078149] ^ p7_array_index_1078166;
  assign p8_array_index_1078384_comb = p7_literal_1076353[p7_res7__35];
  assign p8_array_index_1078385_comb = p7_literal_1076355[p7_res7__34];
  assign p8_res7__40_comb = p7_literal_1076345[p8_res7__39_comb] ^ p7_literal_1076347[p8_res7__38_comb] ^ p7_literal_1076349[p8_res7__37_comb] ^ p7_literal_1076351[p7_res7__36] ^ p8_array_index_1078384_comb ^ p8_array_index_1078385_comb ^ p7_res7__33 ^ p7_literal_1076358[p7_res7__32] ^ p7_array_index_1078142 ^ p7_array_index_1078222 ^ p7_array_index_1078193 ^ p7_array_index_1078161 ^ p7_literal_1076349[p7_array_index_1078146] ^ p7_literal_1076347[p7_array_index_1078147] ^ p7_literal_1076345[p7_array_index_1078164] ^ p7_array_index_1078149;
  assign p8_array_index_1078395_comb = p7_literal_1076353[p7_res7__36];
  assign p8_array_index_1078396_comb = p7_literal_1076355[p7_res7__35];
  assign p8_res7__41_comb = p7_literal_1076345[p8_res7__40_comb] ^ p7_literal_1076347[p8_res7__39_comb] ^ p7_literal_1076349[p8_res7__38_comb] ^ p7_literal_1076351[p8_res7__37_comb] ^ p8_array_index_1078395_comb ^ p8_array_index_1078396_comb ^ p7_res7__34 ^ p7_literal_1076358[p7_res7__33] ^ p7_res7__32 ^ p8_array_index_1078348_comb ^ p7_array_index_1078207 ^ p7_array_index_1078178 ^ p7_literal_1076349[p7_array_index_1078145] ^ p7_literal_1076347[p7_array_index_1078146] ^ p7_literal_1076345[p7_array_index_1078147] ^ p7_array_index_1078164;
  assign p8_array_index_1078402_comb = p7_literal_1076345[p8_res7__41_comb];
  assign p8_array_index_1078403_comb = p7_literal_1076347[p8_res7__40_comb];
  assign p8_array_index_1078404_comb = p7_literal_1076349[p8_res7__39_comb];
  assign p8_array_index_1078405_comb = p7_literal_1076351[p8_res7__38_comb];
  assign p8_array_index_1078406_comb = p7_literal_1076353[p8_res7__37_comb];
  assign p8_array_index_1078407_comb = p7_literal_1076355[p7_res7__36];
  assign p8_array_index_1078408_comb = p7_literal_1076358[p7_res7__34];
  assign p8_array_index_1078409_comb = p7_literal_1076347[p7_array_index_1078145];
  assign p8_array_index_1078410_comb = p7_literal_1076345[p7_array_index_1078146];

  // Registers for pipe stage 8:
  reg [127:0] p8_xor_1077141;
  reg [127:0] p8_xor_1078016;
  reg [7:0] p8_array_index_1078142;
  reg [7:0] p8_array_index_1078143;
  reg [7:0] p8_array_index_1078144;
  reg [7:0] p8_array_index_1078145;
  reg [7:0] p8_array_index_1078146;
  reg [7:0] p8_array_index_1078147;
  reg [7:0] p8_array_index_1078158;
  reg [7:0] p8_array_index_1078159;
  reg [7:0] p8_array_index_1078160;
  reg [7:0] p8_res7__32;
  reg [7:0] p8_array_index_1078175;
  reg [7:0] p8_array_index_1078176;
  reg [7:0] p8_array_index_1078177;
  reg [7:0] p8_res7__33;
  reg [7:0] p8_array_index_1078190;
  reg [7:0] p8_array_index_1078191;
  reg [7:0] p8_array_index_1078192;
  reg [7:0] p8_res7__34;
  reg [7:0] p8_array_index_1078204;
  reg [7:0] p8_array_index_1078205;
  reg [7:0] p8_array_index_1078206;
  reg [7:0] p8_res7__35;
  reg [7:0] p8_array_index_1078219;
  reg [7:0] p8_array_index_1078220;
  reg [7:0] p8_array_index_1078221;
  reg [7:0] p8_res7__36;
  reg [7:0] p8_array_index_1078345;
  reg [7:0] p8_array_index_1078346;
  reg [7:0] p8_array_index_1078347;
  reg [7:0] p8_res7__37;
  reg [7:0] p8_array_index_1078359;
  reg [7:0] p8_array_index_1078360;
  reg [7:0] p8_array_index_1078361;
  reg [7:0] p8_res7__38;
  reg [7:0] p8_array_index_1078371;
  reg [7:0] p8_array_index_1078372;
  reg [7:0] p8_array_index_1078373;
  reg [7:0] p8_res7__39;
  reg [7:0] p8_array_index_1078384;
  reg [7:0] p8_array_index_1078385;
  reg [7:0] p8_res7__40;
  reg [7:0] p8_array_index_1078395;
  reg [7:0] p8_array_index_1078396;
  reg [7:0] p8_res7__41;
  reg [7:0] p8_array_index_1078402;
  reg [7:0] p8_array_index_1078403;
  reg [7:0] p8_array_index_1078404;
  reg [7:0] p8_array_index_1078405;
  reg [7:0] p8_array_index_1078406;
  reg [7:0] p8_array_index_1078407;
  reg [7:0] p8_array_index_1078408;
  reg [7:0] p8_array_index_1078409;
  reg [7:0] p8_array_index_1078410;
  reg [127:0] p8_res__33;
  reg [7:0] p9_arr[256];
  reg [7:0] p9_literal_1076345[256];
  reg [7:0] p9_literal_1076347[256];
  reg [7:0] p9_literal_1076349[256];
  reg [7:0] p9_literal_1076351[256];
  reg [7:0] p9_literal_1076353[256];
  reg [7:0] p9_literal_1076355[256];
  reg [7:0] p9_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p8_xor_1077141 <= p7_xor_1077141;
    p8_xor_1078016 <= p7_xor_1078016;
    p8_array_index_1078142 <= p7_array_index_1078142;
    p8_array_index_1078143 <= p7_array_index_1078143;
    p8_array_index_1078144 <= p7_array_index_1078144;
    p8_array_index_1078145 <= p7_array_index_1078145;
    p8_array_index_1078146 <= p7_array_index_1078146;
    p8_array_index_1078147 <= p7_array_index_1078147;
    p8_array_index_1078158 <= p7_array_index_1078158;
    p8_array_index_1078159 <= p7_array_index_1078159;
    p8_array_index_1078160 <= p7_array_index_1078160;
    p8_res7__32 <= p7_res7__32;
    p8_array_index_1078175 <= p7_array_index_1078175;
    p8_array_index_1078176 <= p7_array_index_1078176;
    p8_array_index_1078177 <= p7_array_index_1078177;
    p8_res7__33 <= p7_res7__33;
    p8_array_index_1078190 <= p7_array_index_1078190;
    p8_array_index_1078191 <= p7_array_index_1078191;
    p8_array_index_1078192 <= p7_array_index_1078192;
    p8_res7__34 <= p7_res7__34;
    p8_array_index_1078204 <= p7_array_index_1078204;
    p8_array_index_1078205 <= p7_array_index_1078205;
    p8_array_index_1078206 <= p7_array_index_1078206;
    p8_res7__35 <= p7_res7__35;
    p8_array_index_1078219 <= p7_array_index_1078219;
    p8_array_index_1078220 <= p7_array_index_1078220;
    p8_array_index_1078221 <= p7_array_index_1078221;
    p8_res7__36 <= p7_res7__36;
    p8_array_index_1078345 <= p8_array_index_1078345_comb;
    p8_array_index_1078346 <= p8_array_index_1078346_comb;
    p8_array_index_1078347 <= p8_array_index_1078347_comb;
    p8_res7__37 <= p8_res7__37_comb;
    p8_array_index_1078359 <= p8_array_index_1078359_comb;
    p8_array_index_1078360 <= p8_array_index_1078360_comb;
    p8_array_index_1078361 <= p8_array_index_1078361_comb;
    p8_res7__38 <= p8_res7__38_comb;
    p8_array_index_1078371 <= p8_array_index_1078371_comb;
    p8_array_index_1078372 <= p8_array_index_1078372_comb;
    p8_array_index_1078373 <= p8_array_index_1078373_comb;
    p8_res7__39 <= p8_res7__39_comb;
    p8_array_index_1078384 <= p8_array_index_1078384_comb;
    p8_array_index_1078385 <= p8_array_index_1078385_comb;
    p8_res7__40 <= p8_res7__40_comb;
    p8_array_index_1078395 <= p8_array_index_1078395_comb;
    p8_array_index_1078396 <= p8_array_index_1078396_comb;
    p8_res7__41 <= p8_res7__41_comb;
    p8_array_index_1078402 <= p8_array_index_1078402_comb;
    p8_array_index_1078403 <= p8_array_index_1078403_comb;
    p8_array_index_1078404 <= p8_array_index_1078404_comb;
    p8_array_index_1078405 <= p8_array_index_1078405_comb;
    p8_array_index_1078406 <= p8_array_index_1078406_comb;
    p8_array_index_1078407 <= p8_array_index_1078407_comb;
    p8_array_index_1078408 <= p8_array_index_1078408_comb;
    p8_array_index_1078409 <= p8_array_index_1078409_comb;
    p8_array_index_1078410 <= p8_array_index_1078410_comb;
    p8_res__33 <= p7_res__33;
    p9_arr <= p8_arr;
    p9_literal_1076345 <= p8_literal_1076345;
    p9_literal_1076347 <= p8_literal_1076347;
    p9_literal_1076349 <= p8_literal_1076349;
    p9_literal_1076351 <= p8_literal_1076351;
    p9_literal_1076353 <= p8_literal_1076353;
    p9_literal_1076355 <= p8_literal_1076355;
    p9_literal_1076358 <= p8_literal_1076358;
  end

  // ===== Pipe stage 9:
  wire [7:0] p9_res7__42_comb;
  wire [7:0] p9_array_index_1078545_comb;
  wire [7:0] p9_res7__43_comb;
  wire [7:0] p9_res7__44_comb;
  wire [7:0] p9_res7__45_comb;
  wire [7:0] p9_res7__46_comb;
  wire [7:0] p9_res7__47_comb;
  wire [127:0] p9_res__2_comb;
  wire [127:0] p9_xor_1078585_comb;
  assign p9_res7__42_comb = p8_array_index_1078402 ^ p8_array_index_1078403 ^ p8_array_index_1078404 ^ p8_array_index_1078405 ^ p8_array_index_1078406 ^ p8_array_index_1078407 ^ p8_res7__35 ^ p8_array_index_1078408 ^ p8_res7__33 ^ p8_array_index_1078361 ^ p8_array_index_1078221 ^ p8_array_index_1078192 ^ p8_array_index_1078160 ^ p8_array_index_1078409 ^ p8_array_index_1078410 ^ p8_array_index_1078147;
  assign p9_array_index_1078545_comb = p8_literal_1076355[p8_res7__37];
  assign p9_res7__43_comb = p8_literal_1076345[p9_res7__42_comb] ^ p8_literal_1076347[p8_res7__41] ^ p8_literal_1076349[p8_res7__40] ^ p8_literal_1076351[p8_res7__39] ^ p8_literal_1076353[p8_res7__38] ^ p9_array_index_1078545_comb ^ p8_res7__36 ^ p8_literal_1076358[p8_res7__35] ^ p8_res7__34 ^ p8_array_index_1078373 ^ p8_array_index_1078347 ^ p8_array_index_1078206 ^ p8_array_index_1078177 ^ p8_literal_1076347[p8_array_index_1078144] ^ p8_literal_1076345[p8_array_index_1078145] ^ p8_array_index_1078146;
  assign p9_res7__44_comb = p8_literal_1076345[p9_res7__43_comb] ^ p8_literal_1076347[p9_res7__42_comb] ^ p8_literal_1076349[p8_res7__41] ^ p8_literal_1076351[p8_res7__40] ^ p8_literal_1076353[p8_res7__39] ^ p8_literal_1076355[p8_res7__38] ^ p8_res7__37 ^ p8_literal_1076358[p8_res7__36] ^ p8_res7__35 ^ p8_array_index_1078385 ^ p8_array_index_1078360 ^ p8_array_index_1078220 ^ p8_array_index_1078191 ^ p8_array_index_1078159 ^ p8_literal_1076345[p8_array_index_1078144] ^ p8_array_index_1078145;
  assign p9_res7__45_comb = p8_literal_1076345[p9_res7__44_comb] ^ p8_literal_1076347[p9_res7__43_comb] ^ p8_literal_1076349[p9_res7__42_comb] ^ p8_literal_1076351[p8_res7__41] ^ p8_literal_1076353[p8_res7__40] ^ p8_literal_1076355[p8_res7__39] ^ p8_res7__38 ^ p8_literal_1076358[p8_res7__37] ^ p8_res7__36 ^ p8_array_index_1078396 ^ p8_array_index_1078372 ^ p8_array_index_1078346 ^ p8_array_index_1078205 ^ p8_array_index_1078176 ^ p8_literal_1076345[p8_array_index_1078143] ^ p8_array_index_1078144;
  assign p9_res7__46_comb = p8_literal_1076345[p9_res7__45_comb] ^ p8_literal_1076347[p9_res7__44_comb] ^ p8_literal_1076349[p9_res7__43_comb] ^ p8_literal_1076351[p9_res7__42_comb] ^ p8_literal_1076353[p8_res7__41] ^ p8_literal_1076355[p8_res7__40] ^ p8_res7__39 ^ p8_literal_1076358[p8_res7__38] ^ p8_res7__37 ^ p8_array_index_1078407 ^ p8_array_index_1078384 ^ p8_array_index_1078359 ^ p8_array_index_1078219 ^ p8_array_index_1078190 ^ p8_array_index_1078158 ^ p8_array_index_1078143;
  assign p9_res7__47_comb = p8_literal_1076345[p9_res7__46_comb] ^ p8_literal_1076347[p9_res7__45_comb] ^ p8_literal_1076349[p9_res7__44_comb] ^ p8_literal_1076351[p9_res7__43_comb] ^ p8_literal_1076353[p9_res7__42_comb] ^ p8_literal_1076355[p8_res7__41] ^ p8_res7__40 ^ p8_literal_1076358[p8_res7__39] ^ p8_res7__38 ^ p9_array_index_1078545_comb ^ p8_array_index_1078395 ^ p8_array_index_1078371 ^ p8_array_index_1078345 ^ p8_array_index_1078204 ^ p8_array_index_1078175 ^ p8_array_index_1078142;
  assign p9_res__2_comb = {p9_res7__47_comb, p9_res7__46_comb, p9_res7__45_comb, p9_res7__44_comb, p9_res7__43_comb, p9_res7__42_comb, p8_res7__41, p8_res7__40, p8_res7__39, p8_res7__38, p8_res7__37, p8_res7__36, p8_res7__35, p8_res7__34, p8_res7__33, p8_res7__32};
  assign p9_xor_1078585_comb = p9_res__2_comb ^ p8_xor_1077141;

  // Registers for pipe stage 9:
  reg [127:0] p9_xor_1078016;
  reg [127:0] p9_xor_1078585;
  reg [127:0] p9_res__33;
  reg [7:0] p10_arr[256];
  reg [7:0] p10_literal_1076345[256];
  reg [7:0] p10_literal_1076347[256];
  reg [7:0] p10_literal_1076349[256];
  reg [7:0] p10_literal_1076351[256];
  reg [7:0] p10_literal_1076353[256];
  reg [7:0] p10_literal_1076355[256];
  reg [7:0] p10_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p9_xor_1078016 <= p8_xor_1078016;
    p9_xor_1078585 <= p9_xor_1078585_comb;
    p9_res__33 <= p8_res__33;
    p10_arr <= p9_arr;
    p10_literal_1076345 <= p9_literal_1076345;
    p10_literal_1076347 <= p9_literal_1076347;
    p10_literal_1076349 <= p9_literal_1076349;
    p10_literal_1076351 <= p9_literal_1076351;
    p10_literal_1076353 <= p9_literal_1076353;
    p10_literal_1076355 <= p9_literal_1076355;
    p10_literal_1076358 <= p9_literal_1076358;
  end

  // ===== Pipe stage 10:
  wire [127:0] p10_addedKey__44_comb;
  wire [7:0] p10_array_index_1078623_comb;
  wire [7:0] p10_array_index_1078624_comb;
  wire [7:0] p10_array_index_1078625_comb;
  wire [7:0] p10_array_index_1078626_comb;
  wire [7:0] p10_array_index_1078627_comb;
  wire [7:0] p10_array_index_1078628_comb;
  wire [7:0] p10_array_index_1078630_comb;
  wire [7:0] p10_array_index_1078632_comb;
  wire [7:0] p10_array_index_1078633_comb;
  wire [7:0] p10_array_index_1078634_comb;
  wire [7:0] p10_array_index_1078635_comb;
  wire [7:0] p10_array_index_1078636_comb;
  wire [7:0] p10_array_index_1078637_comb;
  wire [7:0] p10_array_index_1078639_comb;
  wire [7:0] p10_array_index_1078640_comb;
  wire [7:0] p10_array_index_1078641_comb;
  wire [7:0] p10_array_index_1078642_comb;
  wire [7:0] p10_array_index_1078643_comb;
  wire [7:0] p10_array_index_1078644_comb;
  wire [7:0] p10_array_index_1078645_comb;
  wire [7:0] p10_array_index_1078647_comb;
  wire [7:0] p10_res7__48_comb;
  wire [7:0] p10_array_index_1078656_comb;
  wire [7:0] p10_array_index_1078657_comb;
  wire [7:0] p10_array_index_1078658_comb;
  wire [7:0] p10_array_index_1078659_comb;
  wire [7:0] p10_array_index_1078660_comb;
  wire [7:0] p10_array_index_1078661_comb;
  wire [7:0] p10_res7__49_comb;
  wire [7:0] p10_array_index_1078671_comb;
  wire [7:0] p10_array_index_1078672_comb;
  wire [7:0] p10_array_index_1078673_comb;
  wire [7:0] p10_array_index_1078674_comb;
  wire [7:0] p10_array_index_1078675_comb;
  wire [7:0] p10_res7__50_comb;
  wire [7:0] p10_array_index_1078685_comb;
  wire [7:0] p10_array_index_1078686_comb;
  wire [7:0] p10_array_index_1078687_comb;
  wire [7:0] p10_array_index_1078688_comb;
  wire [7:0] p10_array_index_1078689_comb;
  wire [7:0] p10_res7__51_comb;
  wire [7:0] p10_array_index_1078700_comb;
  wire [7:0] p10_array_index_1078701_comb;
  wire [7:0] p10_array_index_1078702_comb;
  wire [7:0] p10_array_index_1078703_comb;
  wire [7:0] p10_res7__52_comb;
  assign p10_addedKey__44_comb = p9_xor_1078585 ^ 128'h7bcd_1b0b_73e3_2ba5_b79c_b140_f255_1504;
  assign p10_array_index_1078623_comb = p9_arr[p10_addedKey__44_comb[127:120]];
  assign p10_array_index_1078624_comb = p9_arr[p10_addedKey__44_comb[119:112]];
  assign p10_array_index_1078625_comb = p9_arr[p10_addedKey__44_comb[111:104]];
  assign p10_array_index_1078626_comb = p9_arr[p10_addedKey__44_comb[103:96]];
  assign p10_array_index_1078627_comb = p9_arr[p10_addedKey__44_comb[95:88]];
  assign p10_array_index_1078628_comb = p9_arr[p10_addedKey__44_comb[87:80]];
  assign p10_array_index_1078630_comb = p9_arr[p10_addedKey__44_comb[71:64]];
  assign p10_array_index_1078632_comb = p9_arr[p10_addedKey__44_comb[55:48]];
  assign p10_array_index_1078633_comb = p9_arr[p10_addedKey__44_comb[47:40]];
  assign p10_array_index_1078634_comb = p9_arr[p10_addedKey__44_comb[39:32]];
  assign p10_array_index_1078635_comb = p9_arr[p10_addedKey__44_comb[31:24]];
  assign p10_array_index_1078636_comb = p9_arr[p10_addedKey__44_comb[23:16]];
  assign p10_array_index_1078637_comb = p9_arr[p10_addedKey__44_comb[15:8]];
  assign p10_array_index_1078639_comb = p9_literal_1076345[p10_array_index_1078623_comb];
  assign p10_array_index_1078640_comb = p9_literal_1076347[p10_array_index_1078624_comb];
  assign p10_array_index_1078641_comb = p9_literal_1076349[p10_array_index_1078625_comb];
  assign p10_array_index_1078642_comb = p9_literal_1076351[p10_array_index_1078626_comb];
  assign p10_array_index_1078643_comb = p9_literal_1076353[p10_array_index_1078627_comb];
  assign p10_array_index_1078644_comb = p9_literal_1076355[p10_array_index_1078628_comb];
  assign p10_array_index_1078645_comb = p9_arr[p10_addedKey__44_comb[79:72]];
  assign p10_array_index_1078647_comb = p9_arr[p10_addedKey__44_comb[63:56]];
  assign p10_res7__48_comb = p10_array_index_1078639_comb ^ p10_array_index_1078640_comb ^ p10_array_index_1078641_comb ^ p10_array_index_1078642_comb ^ p10_array_index_1078643_comb ^ p10_array_index_1078644_comb ^ p10_array_index_1078645_comb ^ p9_literal_1076358[p10_array_index_1078630_comb] ^ p10_array_index_1078647_comb ^ p9_literal_1076355[p10_array_index_1078632_comb] ^ p9_literal_1076353[p10_array_index_1078633_comb] ^ p9_literal_1076351[p10_array_index_1078634_comb] ^ p9_literal_1076349[p10_array_index_1078635_comb] ^ p9_literal_1076347[p10_array_index_1078636_comb] ^ p9_literal_1076345[p10_array_index_1078637_comb] ^ p9_arr[p10_addedKey__44_comb[7:0]];
  assign p10_array_index_1078656_comb = p9_literal_1076345[p10_res7__48_comb];
  assign p10_array_index_1078657_comb = p9_literal_1076347[p10_array_index_1078623_comb];
  assign p10_array_index_1078658_comb = p9_literal_1076349[p10_array_index_1078624_comb];
  assign p10_array_index_1078659_comb = p9_literal_1076351[p10_array_index_1078625_comb];
  assign p10_array_index_1078660_comb = p9_literal_1076353[p10_array_index_1078626_comb];
  assign p10_array_index_1078661_comb = p9_literal_1076355[p10_array_index_1078627_comb];
  assign p10_res7__49_comb = p10_array_index_1078656_comb ^ p10_array_index_1078657_comb ^ p10_array_index_1078658_comb ^ p10_array_index_1078659_comb ^ p10_array_index_1078660_comb ^ p10_array_index_1078661_comb ^ p10_array_index_1078628_comb ^ p9_literal_1076358[p10_array_index_1078645_comb] ^ p10_array_index_1078630_comb ^ p9_literal_1076355[p10_array_index_1078647_comb] ^ p9_literal_1076353[p10_array_index_1078632_comb] ^ p9_literal_1076351[p10_array_index_1078633_comb] ^ p9_literal_1076349[p10_array_index_1078634_comb] ^ p9_literal_1076347[p10_array_index_1078635_comb] ^ p9_literal_1076345[p10_array_index_1078636_comb] ^ p10_array_index_1078637_comb;
  assign p10_array_index_1078671_comb = p9_literal_1076347[p10_res7__48_comb];
  assign p10_array_index_1078672_comb = p9_literal_1076349[p10_array_index_1078623_comb];
  assign p10_array_index_1078673_comb = p9_literal_1076351[p10_array_index_1078624_comb];
  assign p10_array_index_1078674_comb = p9_literal_1076353[p10_array_index_1078625_comb];
  assign p10_array_index_1078675_comb = p9_literal_1076355[p10_array_index_1078626_comb];
  assign p10_res7__50_comb = p9_literal_1076345[p10_res7__49_comb] ^ p10_array_index_1078671_comb ^ p10_array_index_1078672_comb ^ p10_array_index_1078673_comb ^ p10_array_index_1078674_comb ^ p10_array_index_1078675_comb ^ p10_array_index_1078627_comb ^ p9_literal_1076358[p10_array_index_1078628_comb] ^ p10_array_index_1078645_comb ^ p9_literal_1076355[p10_array_index_1078630_comb] ^ p9_literal_1076353[p10_array_index_1078647_comb] ^ p9_literal_1076351[p10_array_index_1078632_comb] ^ p9_literal_1076349[p10_array_index_1078633_comb] ^ p9_literal_1076347[p10_array_index_1078634_comb] ^ p9_literal_1076345[p10_array_index_1078635_comb] ^ p10_array_index_1078636_comb;
  assign p10_array_index_1078685_comb = p9_literal_1076347[p10_res7__49_comb];
  assign p10_array_index_1078686_comb = p9_literal_1076349[p10_res7__48_comb];
  assign p10_array_index_1078687_comb = p9_literal_1076351[p10_array_index_1078623_comb];
  assign p10_array_index_1078688_comb = p9_literal_1076353[p10_array_index_1078624_comb];
  assign p10_array_index_1078689_comb = p9_literal_1076355[p10_array_index_1078625_comb];
  assign p10_res7__51_comb = p9_literal_1076345[p10_res7__50_comb] ^ p10_array_index_1078685_comb ^ p10_array_index_1078686_comb ^ p10_array_index_1078687_comb ^ p10_array_index_1078688_comb ^ p10_array_index_1078689_comb ^ p10_array_index_1078626_comb ^ p9_literal_1076358[p10_array_index_1078627_comb] ^ p10_array_index_1078628_comb ^ p9_literal_1076355[p10_array_index_1078645_comb] ^ p9_literal_1076353[p10_array_index_1078630_comb] ^ p9_literal_1076351[p10_array_index_1078647_comb] ^ p9_literal_1076349[p10_array_index_1078632_comb] ^ p9_literal_1076347[p10_array_index_1078633_comb] ^ p9_literal_1076345[p10_array_index_1078634_comb] ^ p10_array_index_1078635_comb;
  assign p10_array_index_1078700_comb = p9_literal_1076349[p10_res7__49_comb];
  assign p10_array_index_1078701_comb = p9_literal_1076351[p10_res7__48_comb];
  assign p10_array_index_1078702_comb = p9_literal_1076353[p10_array_index_1078623_comb];
  assign p10_array_index_1078703_comb = p9_literal_1076355[p10_array_index_1078624_comb];
  assign p10_res7__52_comb = p9_literal_1076345[p10_res7__51_comb] ^ p9_literal_1076347[p10_res7__50_comb] ^ p10_array_index_1078700_comb ^ p10_array_index_1078701_comb ^ p10_array_index_1078702_comb ^ p10_array_index_1078703_comb ^ p10_array_index_1078625_comb ^ p9_literal_1076358[p10_array_index_1078626_comb] ^ p10_array_index_1078627_comb ^ p10_array_index_1078644_comb ^ p9_literal_1076353[p10_array_index_1078645_comb] ^ p9_literal_1076351[p10_array_index_1078630_comb] ^ p9_literal_1076349[p10_array_index_1078647_comb] ^ p9_literal_1076347[p10_array_index_1078632_comb] ^ p9_literal_1076345[p10_array_index_1078633_comb] ^ p10_array_index_1078634_comb;

  // Registers for pipe stage 10:
  reg [127:0] p10_xor_1078016;
  reg [127:0] p10_xor_1078585;
  reg [7:0] p10_array_index_1078623;
  reg [7:0] p10_array_index_1078624;
  reg [7:0] p10_array_index_1078625;
  reg [7:0] p10_array_index_1078626;
  reg [7:0] p10_array_index_1078627;
  reg [7:0] p10_array_index_1078628;
  reg [7:0] p10_array_index_1078630;
  reg [7:0] p10_array_index_1078632;
  reg [7:0] p10_array_index_1078633;
  reg [7:0] p10_array_index_1078639;
  reg [7:0] p10_array_index_1078640;
  reg [7:0] p10_array_index_1078641;
  reg [7:0] p10_array_index_1078642;
  reg [7:0] p10_array_index_1078643;
  reg [7:0] p10_array_index_1078645;
  reg [7:0] p10_array_index_1078647;
  reg [7:0] p10_res7__48;
  reg [7:0] p10_array_index_1078656;
  reg [7:0] p10_array_index_1078657;
  reg [7:0] p10_array_index_1078658;
  reg [7:0] p10_array_index_1078659;
  reg [7:0] p10_array_index_1078660;
  reg [7:0] p10_array_index_1078661;
  reg [7:0] p10_res7__49;
  reg [7:0] p10_array_index_1078671;
  reg [7:0] p10_array_index_1078672;
  reg [7:0] p10_array_index_1078673;
  reg [7:0] p10_array_index_1078674;
  reg [7:0] p10_array_index_1078675;
  reg [7:0] p10_res7__50;
  reg [7:0] p10_array_index_1078685;
  reg [7:0] p10_array_index_1078686;
  reg [7:0] p10_array_index_1078687;
  reg [7:0] p10_array_index_1078688;
  reg [7:0] p10_array_index_1078689;
  reg [7:0] p10_res7__51;
  reg [7:0] p10_array_index_1078700;
  reg [7:0] p10_array_index_1078701;
  reg [7:0] p10_array_index_1078702;
  reg [7:0] p10_array_index_1078703;
  reg [7:0] p10_res7__52;
  reg [127:0] p10_res__33;
  reg [7:0] p11_arr[256];
  reg [7:0] p11_literal_1076345[256];
  reg [7:0] p11_literal_1076347[256];
  reg [7:0] p11_literal_1076349[256];
  reg [7:0] p11_literal_1076351[256];
  reg [7:0] p11_literal_1076353[256];
  reg [7:0] p11_literal_1076355[256];
  reg [7:0] p11_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p10_xor_1078016 <= p9_xor_1078016;
    p10_xor_1078585 <= p9_xor_1078585;
    p10_array_index_1078623 <= p10_array_index_1078623_comb;
    p10_array_index_1078624 <= p10_array_index_1078624_comb;
    p10_array_index_1078625 <= p10_array_index_1078625_comb;
    p10_array_index_1078626 <= p10_array_index_1078626_comb;
    p10_array_index_1078627 <= p10_array_index_1078627_comb;
    p10_array_index_1078628 <= p10_array_index_1078628_comb;
    p10_array_index_1078630 <= p10_array_index_1078630_comb;
    p10_array_index_1078632 <= p10_array_index_1078632_comb;
    p10_array_index_1078633 <= p10_array_index_1078633_comb;
    p10_array_index_1078639 <= p10_array_index_1078639_comb;
    p10_array_index_1078640 <= p10_array_index_1078640_comb;
    p10_array_index_1078641 <= p10_array_index_1078641_comb;
    p10_array_index_1078642 <= p10_array_index_1078642_comb;
    p10_array_index_1078643 <= p10_array_index_1078643_comb;
    p10_array_index_1078645 <= p10_array_index_1078645_comb;
    p10_array_index_1078647 <= p10_array_index_1078647_comb;
    p10_res7__48 <= p10_res7__48_comb;
    p10_array_index_1078656 <= p10_array_index_1078656_comb;
    p10_array_index_1078657 <= p10_array_index_1078657_comb;
    p10_array_index_1078658 <= p10_array_index_1078658_comb;
    p10_array_index_1078659 <= p10_array_index_1078659_comb;
    p10_array_index_1078660 <= p10_array_index_1078660_comb;
    p10_array_index_1078661 <= p10_array_index_1078661_comb;
    p10_res7__49 <= p10_res7__49_comb;
    p10_array_index_1078671 <= p10_array_index_1078671_comb;
    p10_array_index_1078672 <= p10_array_index_1078672_comb;
    p10_array_index_1078673 <= p10_array_index_1078673_comb;
    p10_array_index_1078674 <= p10_array_index_1078674_comb;
    p10_array_index_1078675 <= p10_array_index_1078675_comb;
    p10_res7__50 <= p10_res7__50_comb;
    p10_array_index_1078685 <= p10_array_index_1078685_comb;
    p10_array_index_1078686 <= p10_array_index_1078686_comb;
    p10_array_index_1078687 <= p10_array_index_1078687_comb;
    p10_array_index_1078688 <= p10_array_index_1078688_comb;
    p10_array_index_1078689 <= p10_array_index_1078689_comb;
    p10_res7__51 <= p10_res7__51_comb;
    p10_array_index_1078700 <= p10_array_index_1078700_comb;
    p10_array_index_1078701 <= p10_array_index_1078701_comb;
    p10_array_index_1078702 <= p10_array_index_1078702_comb;
    p10_array_index_1078703 <= p10_array_index_1078703_comb;
    p10_res7__52 <= p10_res7__52_comb;
    p10_res__33 <= p9_res__33;
    p11_arr <= p10_arr;
    p11_literal_1076345 <= p10_literal_1076345;
    p11_literal_1076347 <= p10_literal_1076347;
    p11_literal_1076349 <= p10_literal_1076349;
    p11_literal_1076351 <= p10_literal_1076351;
    p11_literal_1076353 <= p10_literal_1076353;
    p11_literal_1076355 <= p10_literal_1076355;
    p11_literal_1076358 <= p10_literal_1076358;
  end

  // ===== Pipe stage 11:
  wire [7:0] p11_array_index_1078817_comb;
  wire [7:0] p11_array_index_1078818_comb;
  wire [7:0] p11_array_index_1078819_comb;
  wire [7:0] p11_array_index_1078820_comb;
  wire [7:0] p11_res7__53_comb;
  wire [7:0] p11_array_index_1078831_comb;
  wire [7:0] p11_array_index_1078832_comb;
  wire [7:0] p11_array_index_1078833_comb;
  wire [7:0] p11_res7__54_comb;
  wire [7:0] p11_array_index_1078843_comb;
  wire [7:0] p11_array_index_1078844_comb;
  wire [7:0] p11_array_index_1078845_comb;
  wire [7:0] p11_res7__55_comb;
  wire [7:0] p11_array_index_1078856_comb;
  wire [7:0] p11_array_index_1078857_comb;
  wire [7:0] p11_res7__56_comb;
  wire [7:0] p11_array_index_1078867_comb;
  wire [7:0] p11_array_index_1078868_comb;
  wire [7:0] p11_res7__57_comb;
  wire [7:0] p11_array_index_1078874_comb;
  wire [7:0] p11_array_index_1078875_comb;
  wire [7:0] p11_array_index_1078876_comb;
  wire [7:0] p11_array_index_1078877_comb;
  wire [7:0] p11_array_index_1078878_comb;
  wire [7:0] p11_array_index_1078879_comb;
  wire [7:0] p11_array_index_1078880_comb;
  wire [7:0] p11_array_index_1078881_comb;
  wire [7:0] p11_array_index_1078882_comb;
  assign p11_array_index_1078817_comb = p10_literal_1076349[p10_res7__50];
  assign p11_array_index_1078818_comb = p10_literal_1076351[p10_res7__49];
  assign p11_array_index_1078819_comb = p10_literal_1076353[p10_res7__48];
  assign p11_array_index_1078820_comb = p10_literal_1076355[p10_array_index_1078623];
  assign p11_res7__53_comb = p10_literal_1076345[p10_res7__52] ^ p10_literal_1076347[p10_res7__51] ^ p11_array_index_1078817_comb ^ p11_array_index_1078818_comb ^ p11_array_index_1078819_comb ^ p11_array_index_1078820_comb ^ p10_array_index_1078624 ^ p10_literal_1076358[p10_array_index_1078625] ^ p10_array_index_1078626 ^ p10_array_index_1078661 ^ p10_literal_1076353[p10_array_index_1078628] ^ p10_literal_1076351[p10_array_index_1078645] ^ p10_literal_1076349[p10_array_index_1078630] ^ p10_literal_1076347[p10_array_index_1078647] ^ p10_literal_1076345[p10_array_index_1078632] ^ p10_array_index_1078633;
  assign p11_array_index_1078831_comb = p10_literal_1076351[p10_res7__50];
  assign p11_array_index_1078832_comb = p10_literal_1076353[p10_res7__49];
  assign p11_array_index_1078833_comb = p10_literal_1076355[p10_res7__48];
  assign p11_res7__54_comb = p10_literal_1076345[p11_res7__53_comb] ^ p10_literal_1076347[p10_res7__52] ^ p10_literal_1076349[p10_res7__51] ^ p11_array_index_1078831_comb ^ p11_array_index_1078832_comb ^ p11_array_index_1078833_comb ^ p10_array_index_1078623 ^ p10_literal_1076358[p10_array_index_1078624] ^ p10_array_index_1078625 ^ p10_array_index_1078675 ^ p10_array_index_1078643 ^ p10_literal_1076351[p10_array_index_1078628] ^ p10_literal_1076349[p10_array_index_1078645] ^ p10_literal_1076347[p10_array_index_1078630] ^ p10_literal_1076345[p10_array_index_1078647] ^ p10_array_index_1078632;
  assign p11_array_index_1078843_comb = p10_literal_1076351[p10_res7__51];
  assign p11_array_index_1078844_comb = p10_literal_1076353[p10_res7__50];
  assign p11_array_index_1078845_comb = p10_literal_1076355[p10_res7__49];
  assign p11_res7__55_comb = p10_literal_1076345[p11_res7__54_comb] ^ p10_literal_1076347[p11_res7__53_comb] ^ p10_literal_1076349[p10_res7__52] ^ p11_array_index_1078843_comb ^ p11_array_index_1078844_comb ^ p11_array_index_1078845_comb ^ p10_res7__48 ^ p10_literal_1076358[p10_array_index_1078623] ^ p10_array_index_1078624 ^ p10_array_index_1078689 ^ p10_array_index_1078660 ^ p10_literal_1076351[p10_array_index_1078627] ^ p10_literal_1076349[p10_array_index_1078628] ^ p10_literal_1076347[p10_array_index_1078645] ^ p10_literal_1076345[p10_array_index_1078630] ^ p10_array_index_1078647;
  assign p11_array_index_1078856_comb = p10_literal_1076353[p10_res7__51];
  assign p11_array_index_1078857_comb = p10_literal_1076355[p10_res7__50];
  assign p11_res7__56_comb = p10_literal_1076345[p11_res7__55_comb] ^ p10_literal_1076347[p11_res7__54_comb] ^ p10_literal_1076349[p11_res7__53_comb] ^ p10_literal_1076351[p10_res7__52] ^ p11_array_index_1078856_comb ^ p11_array_index_1078857_comb ^ p10_res7__49 ^ p10_literal_1076358[p10_res7__48] ^ p10_array_index_1078623 ^ p10_array_index_1078703 ^ p10_array_index_1078674 ^ p10_array_index_1078642 ^ p10_literal_1076349[p10_array_index_1078627] ^ p10_literal_1076347[p10_array_index_1078628] ^ p10_literal_1076345[p10_array_index_1078645] ^ p10_array_index_1078630;
  assign p11_array_index_1078867_comb = p10_literal_1076353[p10_res7__52];
  assign p11_array_index_1078868_comb = p10_literal_1076355[p10_res7__51];
  assign p11_res7__57_comb = p10_literal_1076345[p11_res7__56_comb] ^ p10_literal_1076347[p11_res7__55_comb] ^ p10_literal_1076349[p11_res7__54_comb] ^ p10_literal_1076351[p11_res7__53_comb] ^ p11_array_index_1078867_comb ^ p11_array_index_1078868_comb ^ p10_res7__50 ^ p10_literal_1076358[p10_res7__49] ^ p10_res7__48 ^ p11_array_index_1078820_comb ^ p10_array_index_1078688 ^ p10_array_index_1078659 ^ p10_literal_1076349[p10_array_index_1078626] ^ p10_literal_1076347[p10_array_index_1078627] ^ p10_literal_1076345[p10_array_index_1078628] ^ p10_array_index_1078645;
  assign p11_array_index_1078874_comb = p10_literal_1076345[p11_res7__57_comb];
  assign p11_array_index_1078875_comb = p10_literal_1076347[p11_res7__56_comb];
  assign p11_array_index_1078876_comb = p10_literal_1076349[p11_res7__55_comb];
  assign p11_array_index_1078877_comb = p10_literal_1076351[p11_res7__54_comb];
  assign p11_array_index_1078878_comb = p10_literal_1076353[p11_res7__53_comb];
  assign p11_array_index_1078879_comb = p10_literal_1076355[p10_res7__52];
  assign p11_array_index_1078880_comb = p10_literal_1076358[p10_res7__50];
  assign p11_array_index_1078881_comb = p10_literal_1076347[p10_array_index_1078626];
  assign p11_array_index_1078882_comb = p10_literal_1076345[p10_array_index_1078627];

  // Registers for pipe stage 11:
  reg [127:0] p11_xor_1078016;
  reg [127:0] p11_xor_1078585;
  reg [7:0] p11_array_index_1078623;
  reg [7:0] p11_array_index_1078624;
  reg [7:0] p11_array_index_1078625;
  reg [7:0] p11_array_index_1078626;
  reg [7:0] p11_array_index_1078627;
  reg [7:0] p11_array_index_1078628;
  reg [7:0] p11_array_index_1078639;
  reg [7:0] p11_array_index_1078640;
  reg [7:0] p11_array_index_1078641;
  reg [7:0] p11_res7__48;
  reg [7:0] p11_array_index_1078656;
  reg [7:0] p11_array_index_1078657;
  reg [7:0] p11_array_index_1078658;
  reg [7:0] p11_res7__49;
  reg [7:0] p11_array_index_1078671;
  reg [7:0] p11_array_index_1078672;
  reg [7:0] p11_array_index_1078673;
  reg [7:0] p11_res7__50;
  reg [7:0] p11_array_index_1078685;
  reg [7:0] p11_array_index_1078686;
  reg [7:0] p11_array_index_1078687;
  reg [7:0] p11_res7__51;
  reg [7:0] p11_array_index_1078700;
  reg [7:0] p11_array_index_1078701;
  reg [7:0] p11_array_index_1078702;
  reg [7:0] p11_res7__52;
  reg [7:0] p11_array_index_1078817;
  reg [7:0] p11_array_index_1078818;
  reg [7:0] p11_array_index_1078819;
  reg [7:0] p11_res7__53;
  reg [7:0] p11_array_index_1078831;
  reg [7:0] p11_array_index_1078832;
  reg [7:0] p11_array_index_1078833;
  reg [7:0] p11_res7__54;
  reg [7:0] p11_array_index_1078843;
  reg [7:0] p11_array_index_1078844;
  reg [7:0] p11_array_index_1078845;
  reg [7:0] p11_res7__55;
  reg [7:0] p11_array_index_1078856;
  reg [7:0] p11_array_index_1078857;
  reg [7:0] p11_res7__56;
  reg [7:0] p11_array_index_1078867;
  reg [7:0] p11_array_index_1078868;
  reg [7:0] p11_res7__57;
  reg [7:0] p11_array_index_1078874;
  reg [7:0] p11_array_index_1078875;
  reg [7:0] p11_array_index_1078876;
  reg [7:0] p11_array_index_1078877;
  reg [7:0] p11_array_index_1078878;
  reg [7:0] p11_array_index_1078879;
  reg [7:0] p11_array_index_1078880;
  reg [7:0] p11_array_index_1078881;
  reg [7:0] p11_array_index_1078882;
  reg [127:0] p11_res__33;
  reg [7:0] p12_arr[256];
  reg [7:0] p12_literal_1076345[256];
  reg [7:0] p12_literal_1076347[256];
  reg [7:0] p12_literal_1076349[256];
  reg [7:0] p12_literal_1076351[256];
  reg [7:0] p12_literal_1076353[256];
  reg [7:0] p12_literal_1076355[256];
  reg [7:0] p12_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p11_xor_1078016 <= p10_xor_1078016;
    p11_xor_1078585 <= p10_xor_1078585;
    p11_array_index_1078623 <= p10_array_index_1078623;
    p11_array_index_1078624 <= p10_array_index_1078624;
    p11_array_index_1078625 <= p10_array_index_1078625;
    p11_array_index_1078626 <= p10_array_index_1078626;
    p11_array_index_1078627 <= p10_array_index_1078627;
    p11_array_index_1078628 <= p10_array_index_1078628;
    p11_array_index_1078639 <= p10_array_index_1078639;
    p11_array_index_1078640 <= p10_array_index_1078640;
    p11_array_index_1078641 <= p10_array_index_1078641;
    p11_res7__48 <= p10_res7__48;
    p11_array_index_1078656 <= p10_array_index_1078656;
    p11_array_index_1078657 <= p10_array_index_1078657;
    p11_array_index_1078658 <= p10_array_index_1078658;
    p11_res7__49 <= p10_res7__49;
    p11_array_index_1078671 <= p10_array_index_1078671;
    p11_array_index_1078672 <= p10_array_index_1078672;
    p11_array_index_1078673 <= p10_array_index_1078673;
    p11_res7__50 <= p10_res7__50;
    p11_array_index_1078685 <= p10_array_index_1078685;
    p11_array_index_1078686 <= p10_array_index_1078686;
    p11_array_index_1078687 <= p10_array_index_1078687;
    p11_res7__51 <= p10_res7__51;
    p11_array_index_1078700 <= p10_array_index_1078700;
    p11_array_index_1078701 <= p10_array_index_1078701;
    p11_array_index_1078702 <= p10_array_index_1078702;
    p11_res7__52 <= p10_res7__52;
    p11_array_index_1078817 <= p11_array_index_1078817_comb;
    p11_array_index_1078818 <= p11_array_index_1078818_comb;
    p11_array_index_1078819 <= p11_array_index_1078819_comb;
    p11_res7__53 <= p11_res7__53_comb;
    p11_array_index_1078831 <= p11_array_index_1078831_comb;
    p11_array_index_1078832 <= p11_array_index_1078832_comb;
    p11_array_index_1078833 <= p11_array_index_1078833_comb;
    p11_res7__54 <= p11_res7__54_comb;
    p11_array_index_1078843 <= p11_array_index_1078843_comb;
    p11_array_index_1078844 <= p11_array_index_1078844_comb;
    p11_array_index_1078845 <= p11_array_index_1078845_comb;
    p11_res7__55 <= p11_res7__55_comb;
    p11_array_index_1078856 <= p11_array_index_1078856_comb;
    p11_array_index_1078857 <= p11_array_index_1078857_comb;
    p11_res7__56 <= p11_res7__56_comb;
    p11_array_index_1078867 <= p11_array_index_1078867_comb;
    p11_array_index_1078868 <= p11_array_index_1078868_comb;
    p11_res7__57 <= p11_res7__57_comb;
    p11_array_index_1078874 <= p11_array_index_1078874_comb;
    p11_array_index_1078875 <= p11_array_index_1078875_comb;
    p11_array_index_1078876 <= p11_array_index_1078876_comb;
    p11_array_index_1078877 <= p11_array_index_1078877_comb;
    p11_array_index_1078878 <= p11_array_index_1078878_comb;
    p11_array_index_1078879 <= p11_array_index_1078879_comb;
    p11_array_index_1078880 <= p11_array_index_1078880_comb;
    p11_array_index_1078881 <= p11_array_index_1078881_comb;
    p11_array_index_1078882 <= p11_array_index_1078882_comb;
    p11_res__33 <= p10_res__33;
    p12_arr <= p11_arr;
    p12_literal_1076345 <= p11_literal_1076345;
    p12_literal_1076347 <= p11_literal_1076347;
    p12_literal_1076349 <= p11_literal_1076349;
    p12_literal_1076351 <= p11_literal_1076351;
    p12_literal_1076353 <= p11_literal_1076353;
    p12_literal_1076355 <= p11_literal_1076355;
    p12_literal_1076358 <= p11_literal_1076358;
  end

  // ===== Pipe stage 12:
  wire [7:0] p12_res7__58_comb;
  wire [7:0] p12_array_index_1079017_comb;
  wire [7:0] p12_res7__59_comb;
  wire [7:0] p12_res7__60_comb;
  wire [7:0] p12_res7__61_comb;
  wire [7:0] p12_res7__62_comb;
  wire [7:0] p12_res7__63_comb;
  wire [127:0] p12_res__3_comb;
  wire [127:0] p12_xor_1079057_comb;
  assign p12_res7__58_comb = p11_array_index_1078874 ^ p11_array_index_1078875 ^ p11_array_index_1078876 ^ p11_array_index_1078877 ^ p11_array_index_1078878 ^ p11_array_index_1078879 ^ p11_res7__51 ^ p11_array_index_1078880 ^ p11_res7__49 ^ p11_array_index_1078833 ^ p11_array_index_1078702 ^ p11_array_index_1078673 ^ p11_array_index_1078641 ^ p11_array_index_1078881 ^ p11_array_index_1078882 ^ p11_array_index_1078628;
  assign p12_array_index_1079017_comb = p11_literal_1076355[p11_res7__53];
  assign p12_res7__59_comb = p11_literal_1076345[p12_res7__58_comb] ^ p11_literal_1076347[p11_res7__57] ^ p11_literal_1076349[p11_res7__56] ^ p11_literal_1076351[p11_res7__55] ^ p11_literal_1076353[p11_res7__54] ^ p12_array_index_1079017_comb ^ p11_res7__52 ^ p11_literal_1076358[p11_res7__51] ^ p11_res7__50 ^ p11_array_index_1078845 ^ p11_array_index_1078819 ^ p11_array_index_1078687 ^ p11_array_index_1078658 ^ p11_literal_1076347[p11_array_index_1078625] ^ p11_literal_1076345[p11_array_index_1078626] ^ p11_array_index_1078627;
  assign p12_res7__60_comb = p11_literal_1076345[p12_res7__59_comb] ^ p11_literal_1076347[p12_res7__58_comb] ^ p11_literal_1076349[p11_res7__57] ^ p11_literal_1076351[p11_res7__56] ^ p11_literal_1076353[p11_res7__55] ^ p11_literal_1076355[p11_res7__54] ^ p11_res7__53 ^ p11_literal_1076358[p11_res7__52] ^ p11_res7__51 ^ p11_array_index_1078857 ^ p11_array_index_1078832 ^ p11_array_index_1078701 ^ p11_array_index_1078672 ^ p11_array_index_1078640 ^ p11_literal_1076345[p11_array_index_1078625] ^ p11_array_index_1078626;
  assign p12_res7__61_comb = p11_literal_1076345[p12_res7__60_comb] ^ p11_literal_1076347[p12_res7__59_comb] ^ p11_literal_1076349[p12_res7__58_comb] ^ p11_literal_1076351[p11_res7__57] ^ p11_literal_1076353[p11_res7__56] ^ p11_literal_1076355[p11_res7__55] ^ p11_res7__54 ^ p11_literal_1076358[p11_res7__53] ^ p11_res7__52 ^ p11_array_index_1078868 ^ p11_array_index_1078844 ^ p11_array_index_1078818 ^ p11_array_index_1078686 ^ p11_array_index_1078657 ^ p11_literal_1076345[p11_array_index_1078624] ^ p11_array_index_1078625;
  assign p12_res7__62_comb = p11_literal_1076345[p12_res7__61_comb] ^ p11_literal_1076347[p12_res7__60_comb] ^ p11_literal_1076349[p12_res7__59_comb] ^ p11_literal_1076351[p12_res7__58_comb] ^ p11_literal_1076353[p11_res7__57] ^ p11_literal_1076355[p11_res7__56] ^ p11_res7__55 ^ p11_literal_1076358[p11_res7__54] ^ p11_res7__53 ^ p11_array_index_1078879 ^ p11_array_index_1078856 ^ p11_array_index_1078831 ^ p11_array_index_1078700 ^ p11_array_index_1078671 ^ p11_array_index_1078639 ^ p11_array_index_1078624;
  assign p12_res7__63_comb = p11_literal_1076345[p12_res7__62_comb] ^ p11_literal_1076347[p12_res7__61_comb] ^ p11_literal_1076349[p12_res7__60_comb] ^ p11_literal_1076351[p12_res7__59_comb] ^ p11_literal_1076353[p12_res7__58_comb] ^ p11_literal_1076355[p11_res7__57] ^ p11_res7__56 ^ p11_literal_1076358[p11_res7__55] ^ p11_res7__54 ^ p12_array_index_1079017_comb ^ p11_array_index_1078867 ^ p11_array_index_1078843 ^ p11_array_index_1078817 ^ p11_array_index_1078685 ^ p11_array_index_1078656 ^ p11_array_index_1078623;
  assign p12_res__3_comb = {p12_res7__63_comb, p12_res7__62_comb, p12_res7__61_comb, p12_res7__60_comb, p12_res7__59_comb, p12_res7__58_comb, p11_res7__57, p11_res7__56, p11_res7__55, p11_res7__54, p11_res7__53, p11_res7__52, p11_res7__51, p11_res7__50, p11_res7__49, p11_res7__48};
  assign p12_xor_1079057_comb = p12_res__3_comb ^ p11_xor_1078016;

  // Registers for pipe stage 12:
  reg [127:0] p12_xor_1078585;
  reg [127:0] p12_xor_1079057;
  reg [127:0] p12_res__33;
  reg [7:0] p13_arr[256];
  reg [7:0] p13_literal_1076345[256];
  reg [7:0] p13_literal_1076347[256];
  reg [7:0] p13_literal_1076349[256];
  reg [7:0] p13_literal_1076351[256];
  reg [7:0] p13_literal_1076353[256];
  reg [7:0] p13_literal_1076355[256];
  reg [7:0] p13_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p12_xor_1078585 <= p11_xor_1078585;
    p12_xor_1079057 <= p12_xor_1079057_comb;
    p12_res__33 <= p11_res__33;
    p13_arr <= p12_arr;
    p13_literal_1076345 <= p12_literal_1076345;
    p13_literal_1076347 <= p12_literal_1076347;
    p13_literal_1076349 <= p12_literal_1076349;
    p13_literal_1076351 <= p12_literal_1076351;
    p13_literal_1076353 <= p12_literal_1076353;
    p13_literal_1076355 <= p12_literal_1076355;
    p13_literal_1076358 <= p12_literal_1076358;
  end

  // ===== Pipe stage 13:
  wire [127:0] p13_addedKey__45_comb;
  wire [7:0] p13_array_index_1079095_comb;
  wire [7:0] p13_array_index_1079096_comb;
  wire [7:0] p13_array_index_1079097_comb;
  wire [7:0] p13_array_index_1079098_comb;
  wire [7:0] p13_array_index_1079099_comb;
  wire [7:0] p13_array_index_1079100_comb;
  wire [7:0] p13_array_index_1079102_comb;
  wire [7:0] p13_array_index_1079104_comb;
  wire [7:0] p13_array_index_1079105_comb;
  wire [7:0] p13_array_index_1079106_comb;
  wire [7:0] p13_array_index_1079107_comb;
  wire [7:0] p13_array_index_1079108_comb;
  wire [7:0] p13_array_index_1079109_comb;
  wire [7:0] p13_array_index_1079111_comb;
  wire [7:0] p13_array_index_1079112_comb;
  wire [7:0] p13_array_index_1079113_comb;
  wire [7:0] p13_array_index_1079114_comb;
  wire [7:0] p13_array_index_1079115_comb;
  wire [7:0] p13_array_index_1079116_comb;
  wire [7:0] p13_array_index_1079117_comb;
  wire [7:0] p13_array_index_1079119_comb;
  wire [7:0] p13_res7__64_comb;
  wire [7:0] p13_array_index_1079128_comb;
  wire [7:0] p13_array_index_1079129_comb;
  wire [7:0] p13_array_index_1079130_comb;
  wire [7:0] p13_array_index_1079131_comb;
  wire [7:0] p13_array_index_1079132_comb;
  wire [7:0] p13_array_index_1079133_comb;
  wire [7:0] p13_res7__65_comb;
  wire [7:0] p13_array_index_1079143_comb;
  wire [7:0] p13_array_index_1079144_comb;
  wire [7:0] p13_array_index_1079145_comb;
  wire [7:0] p13_array_index_1079146_comb;
  wire [7:0] p13_array_index_1079147_comb;
  wire [7:0] p13_res7__66_comb;
  wire [7:0] p13_array_index_1079157_comb;
  wire [7:0] p13_array_index_1079158_comb;
  wire [7:0] p13_array_index_1079159_comb;
  wire [7:0] p13_array_index_1079160_comb;
  wire [7:0] p13_array_index_1079161_comb;
  wire [7:0] p13_res7__67_comb;
  wire [7:0] p13_array_index_1079172_comb;
  wire [7:0] p13_array_index_1079173_comb;
  wire [7:0] p13_array_index_1079174_comb;
  wire [7:0] p13_array_index_1079175_comb;
  wire [7:0] p13_res7__68_comb;
  assign p13_addedKey__45_comb = p12_xor_1079057 ^ 128'h156f_6d79_1fab_511d_eabb_0c50_2fd1_8105;
  assign p13_array_index_1079095_comb = p12_arr[p13_addedKey__45_comb[127:120]];
  assign p13_array_index_1079096_comb = p12_arr[p13_addedKey__45_comb[119:112]];
  assign p13_array_index_1079097_comb = p12_arr[p13_addedKey__45_comb[111:104]];
  assign p13_array_index_1079098_comb = p12_arr[p13_addedKey__45_comb[103:96]];
  assign p13_array_index_1079099_comb = p12_arr[p13_addedKey__45_comb[95:88]];
  assign p13_array_index_1079100_comb = p12_arr[p13_addedKey__45_comb[87:80]];
  assign p13_array_index_1079102_comb = p12_arr[p13_addedKey__45_comb[71:64]];
  assign p13_array_index_1079104_comb = p12_arr[p13_addedKey__45_comb[55:48]];
  assign p13_array_index_1079105_comb = p12_arr[p13_addedKey__45_comb[47:40]];
  assign p13_array_index_1079106_comb = p12_arr[p13_addedKey__45_comb[39:32]];
  assign p13_array_index_1079107_comb = p12_arr[p13_addedKey__45_comb[31:24]];
  assign p13_array_index_1079108_comb = p12_arr[p13_addedKey__45_comb[23:16]];
  assign p13_array_index_1079109_comb = p12_arr[p13_addedKey__45_comb[15:8]];
  assign p13_array_index_1079111_comb = p12_literal_1076345[p13_array_index_1079095_comb];
  assign p13_array_index_1079112_comb = p12_literal_1076347[p13_array_index_1079096_comb];
  assign p13_array_index_1079113_comb = p12_literal_1076349[p13_array_index_1079097_comb];
  assign p13_array_index_1079114_comb = p12_literal_1076351[p13_array_index_1079098_comb];
  assign p13_array_index_1079115_comb = p12_literal_1076353[p13_array_index_1079099_comb];
  assign p13_array_index_1079116_comb = p12_literal_1076355[p13_array_index_1079100_comb];
  assign p13_array_index_1079117_comb = p12_arr[p13_addedKey__45_comb[79:72]];
  assign p13_array_index_1079119_comb = p12_arr[p13_addedKey__45_comb[63:56]];
  assign p13_res7__64_comb = p13_array_index_1079111_comb ^ p13_array_index_1079112_comb ^ p13_array_index_1079113_comb ^ p13_array_index_1079114_comb ^ p13_array_index_1079115_comb ^ p13_array_index_1079116_comb ^ p13_array_index_1079117_comb ^ p12_literal_1076358[p13_array_index_1079102_comb] ^ p13_array_index_1079119_comb ^ p12_literal_1076355[p13_array_index_1079104_comb] ^ p12_literal_1076353[p13_array_index_1079105_comb] ^ p12_literal_1076351[p13_array_index_1079106_comb] ^ p12_literal_1076349[p13_array_index_1079107_comb] ^ p12_literal_1076347[p13_array_index_1079108_comb] ^ p12_literal_1076345[p13_array_index_1079109_comb] ^ p12_arr[p13_addedKey__45_comb[7:0]];
  assign p13_array_index_1079128_comb = p12_literal_1076345[p13_res7__64_comb];
  assign p13_array_index_1079129_comb = p12_literal_1076347[p13_array_index_1079095_comb];
  assign p13_array_index_1079130_comb = p12_literal_1076349[p13_array_index_1079096_comb];
  assign p13_array_index_1079131_comb = p12_literal_1076351[p13_array_index_1079097_comb];
  assign p13_array_index_1079132_comb = p12_literal_1076353[p13_array_index_1079098_comb];
  assign p13_array_index_1079133_comb = p12_literal_1076355[p13_array_index_1079099_comb];
  assign p13_res7__65_comb = p13_array_index_1079128_comb ^ p13_array_index_1079129_comb ^ p13_array_index_1079130_comb ^ p13_array_index_1079131_comb ^ p13_array_index_1079132_comb ^ p13_array_index_1079133_comb ^ p13_array_index_1079100_comb ^ p12_literal_1076358[p13_array_index_1079117_comb] ^ p13_array_index_1079102_comb ^ p12_literal_1076355[p13_array_index_1079119_comb] ^ p12_literal_1076353[p13_array_index_1079104_comb] ^ p12_literal_1076351[p13_array_index_1079105_comb] ^ p12_literal_1076349[p13_array_index_1079106_comb] ^ p12_literal_1076347[p13_array_index_1079107_comb] ^ p12_literal_1076345[p13_array_index_1079108_comb] ^ p13_array_index_1079109_comb;
  assign p13_array_index_1079143_comb = p12_literal_1076347[p13_res7__64_comb];
  assign p13_array_index_1079144_comb = p12_literal_1076349[p13_array_index_1079095_comb];
  assign p13_array_index_1079145_comb = p12_literal_1076351[p13_array_index_1079096_comb];
  assign p13_array_index_1079146_comb = p12_literal_1076353[p13_array_index_1079097_comb];
  assign p13_array_index_1079147_comb = p12_literal_1076355[p13_array_index_1079098_comb];
  assign p13_res7__66_comb = p12_literal_1076345[p13_res7__65_comb] ^ p13_array_index_1079143_comb ^ p13_array_index_1079144_comb ^ p13_array_index_1079145_comb ^ p13_array_index_1079146_comb ^ p13_array_index_1079147_comb ^ p13_array_index_1079099_comb ^ p12_literal_1076358[p13_array_index_1079100_comb] ^ p13_array_index_1079117_comb ^ p12_literal_1076355[p13_array_index_1079102_comb] ^ p12_literal_1076353[p13_array_index_1079119_comb] ^ p12_literal_1076351[p13_array_index_1079104_comb] ^ p12_literal_1076349[p13_array_index_1079105_comb] ^ p12_literal_1076347[p13_array_index_1079106_comb] ^ p12_literal_1076345[p13_array_index_1079107_comb] ^ p13_array_index_1079108_comb;
  assign p13_array_index_1079157_comb = p12_literal_1076347[p13_res7__65_comb];
  assign p13_array_index_1079158_comb = p12_literal_1076349[p13_res7__64_comb];
  assign p13_array_index_1079159_comb = p12_literal_1076351[p13_array_index_1079095_comb];
  assign p13_array_index_1079160_comb = p12_literal_1076353[p13_array_index_1079096_comb];
  assign p13_array_index_1079161_comb = p12_literal_1076355[p13_array_index_1079097_comb];
  assign p13_res7__67_comb = p12_literal_1076345[p13_res7__66_comb] ^ p13_array_index_1079157_comb ^ p13_array_index_1079158_comb ^ p13_array_index_1079159_comb ^ p13_array_index_1079160_comb ^ p13_array_index_1079161_comb ^ p13_array_index_1079098_comb ^ p12_literal_1076358[p13_array_index_1079099_comb] ^ p13_array_index_1079100_comb ^ p12_literal_1076355[p13_array_index_1079117_comb] ^ p12_literal_1076353[p13_array_index_1079102_comb] ^ p12_literal_1076351[p13_array_index_1079119_comb] ^ p12_literal_1076349[p13_array_index_1079104_comb] ^ p12_literal_1076347[p13_array_index_1079105_comb] ^ p12_literal_1076345[p13_array_index_1079106_comb] ^ p13_array_index_1079107_comb;
  assign p13_array_index_1079172_comb = p12_literal_1076349[p13_res7__65_comb];
  assign p13_array_index_1079173_comb = p12_literal_1076351[p13_res7__64_comb];
  assign p13_array_index_1079174_comb = p12_literal_1076353[p13_array_index_1079095_comb];
  assign p13_array_index_1079175_comb = p12_literal_1076355[p13_array_index_1079096_comb];
  assign p13_res7__68_comb = p12_literal_1076345[p13_res7__67_comb] ^ p12_literal_1076347[p13_res7__66_comb] ^ p13_array_index_1079172_comb ^ p13_array_index_1079173_comb ^ p13_array_index_1079174_comb ^ p13_array_index_1079175_comb ^ p13_array_index_1079097_comb ^ p12_literal_1076358[p13_array_index_1079098_comb] ^ p13_array_index_1079099_comb ^ p13_array_index_1079116_comb ^ p12_literal_1076353[p13_array_index_1079117_comb] ^ p12_literal_1076351[p13_array_index_1079102_comb] ^ p12_literal_1076349[p13_array_index_1079119_comb] ^ p12_literal_1076347[p13_array_index_1079104_comb] ^ p12_literal_1076345[p13_array_index_1079105_comb] ^ p13_array_index_1079106_comb;

  // Registers for pipe stage 13:
  reg [127:0] p13_xor_1078585;
  reg [127:0] p13_xor_1079057;
  reg [7:0] p13_array_index_1079095;
  reg [7:0] p13_array_index_1079096;
  reg [7:0] p13_array_index_1079097;
  reg [7:0] p13_array_index_1079098;
  reg [7:0] p13_array_index_1079099;
  reg [7:0] p13_array_index_1079100;
  reg [7:0] p13_array_index_1079102;
  reg [7:0] p13_array_index_1079104;
  reg [7:0] p13_array_index_1079105;
  reg [7:0] p13_array_index_1079111;
  reg [7:0] p13_array_index_1079112;
  reg [7:0] p13_array_index_1079113;
  reg [7:0] p13_array_index_1079114;
  reg [7:0] p13_array_index_1079115;
  reg [7:0] p13_array_index_1079117;
  reg [7:0] p13_array_index_1079119;
  reg [7:0] p13_res7__64;
  reg [7:0] p13_array_index_1079128;
  reg [7:0] p13_array_index_1079129;
  reg [7:0] p13_array_index_1079130;
  reg [7:0] p13_array_index_1079131;
  reg [7:0] p13_array_index_1079132;
  reg [7:0] p13_array_index_1079133;
  reg [7:0] p13_res7__65;
  reg [7:0] p13_array_index_1079143;
  reg [7:0] p13_array_index_1079144;
  reg [7:0] p13_array_index_1079145;
  reg [7:0] p13_array_index_1079146;
  reg [7:0] p13_array_index_1079147;
  reg [7:0] p13_res7__66;
  reg [7:0] p13_array_index_1079157;
  reg [7:0] p13_array_index_1079158;
  reg [7:0] p13_array_index_1079159;
  reg [7:0] p13_array_index_1079160;
  reg [7:0] p13_array_index_1079161;
  reg [7:0] p13_res7__67;
  reg [7:0] p13_array_index_1079172;
  reg [7:0] p13_array_index_1079173;
  reg [7:0] p13_array_index_1079174;
  reg [7:0] p13_array_index_1079175;
  reg [7:0] p13_res7__68;
  reg [127:0] p13_res__33;
  reg [7:0] p14_arr[256];
  reg [7:0] p14_literal_1076345[256];
  reg [7:0] p14_literal_1076347[256];
  reg [7:0] p14_literal_1076349[256];
  reg [7:0] p14_literal_1076351[256];
  reg [7:0] p14_literal_1076353[256];
  reg [7:0] p14_literal_1076355[256];
  reg [7:0] p14_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p13_xor_1078585 <= p12_xor_1078585;
    p13_xor_1079057 <= p12_xor_1079057;
    p13_array_index_1079095 <= p13_array_index_1079095_comb;
    p13_array_index_1079096 <= p13_array_index_1079096_comb;
    p13_array_index_1079097 <= p13_array_index_1079097_comb;
    p13_array_index_1079098 <= p13_array_index_1079098_comb;
    p13_array_index_1079099 <= p13_array_index_1079099_comb;
    p13_array_index_1079100 <= p13_array_index_1079100_comb;
    p13_array_index_1079102 <= p13_array_index_1079102_comb;
    p13_array_index_1079104 <= p13_array_index_1079104_comb;
    p13_array_index_1079105 <= p13_array_index_1079105_comb;
    p13_array_index_1079111 <= p13_array_index_1079111_comb;
    p13_array_index_1079112 <= p13_array_index_1079112_comb;
    p13_array_index_1079113 <= p13_array_index_1079113_comb;
    p13_array_index_1079114 <= p13_array_index_1079114_comb;
    p13_array_index_1079115 <= p13_array_index_1079115_comb;
    p13_array_index_1079117 <= p13_array_index_1079117_comb;
    p13_array_index_1079119 <= p13_array_index_1079119_comb;
    p13_res7__64 <= p13_res7__64_comb;
    p13_array_index_1079128 <= p13_array_index_1079128_comb;
    p13_array_index_1079129 <= p13_array_index_1079129_comb;
    p13_array_index_1079130 <= p13_array_index_1079130_comb;
    p13_array_index_1079131 <= p13_array_index_1079131_comb;
    p13_array_index_1079132 <= p13_array_index_1079132_comb;
    p13_array_index_1079133 <= p13_array_index_1079133_comb;
    p13_res7__65 <= p13_res7__65_comb;
    p13_array_index_1079143 <= p13_array_index_1079143_comb;
    p13_array_index_1079144 <= p13_array_index_1079144_comb;
    p13_array_index_1079145 <= p13_array_index_1079145_comb;
    p13_array_index_1079146 <= p13_array_index_1079146_comb;
    p13_array_index_1079147 <= p13_array_index_1079147_comb;
    p13_res7__66 <= p13_res7__66_comb;
    p13_array_index_1079157 <= p13_array_index_1079157_comb;
    p13_array_index_1079158 <= p13_array_index_1079158_comb;
    p13_array_index_1079159 <= p13_array_index_1079159_comb;
    p13_array_index_1079160 <= p13_array_index_1079160_comb;
    p13_array_index_1079161 <= p13_array_index_1079161_comb;
    p13_res7__67 <= p13_res7__67_comb;
    p13_array_index_1079172 <= p13_array_index_1079172_comb;
    p13_array_index_1079173 <= p13_array_index_1079173_comb;
    p13_array_index_1079174 <= p13_array_index_1079174_comb;
    p13_array_index_1079175 <= p13_array_index_1079175_comb;
    p13_res7__68 <= p13_res7__68_comb;
    p13_res__33 <= p12_res__33;
    p14_arr <= p13_arr;
    p14_literal_1076345 <= p13_literal_1076345;
    p14_literal_1076347 <= p13_literal_1076347;
    p14_literal_1076349 <= p13_literal_1076349;
    p14_literal_1076351 <= p13_literal_1076351;
    p14_literal_1076353 <= p13_literal_1076353;
    p14_literal_1076355 <= p13_literal_1076355;
    p14_literal_1076358 <= p13_literal_1076358;
  end

  // ===== Pipe stage 14:
  wire [7:0] p14_array_index_1079289_comb;
  wire [7:0] p14_array_index_1079290_comb;
  wire [7:0] p14_array_index_1079291_comb;
  wire [7:0] p14_array_index_1079292_comb;
  wire [7:0] p14_res7__69_comb;
  wire [7:0] p14_array_index_1079303_comb;
  wire [7:0] p14_array_index_1079304_comb;
  wire [7:0] p14_array_index_1079305_comb;
  wire [7:0] p14_res7__70_comb;
  wire [7:0] p14_array_index_1079315_comb;
  wire [7:0] p14_array_index_1079316_comb;
  wire [7:0] p14_array_index_1079317_comb;
  wire [7:0] p14_res7__71_comb;
  wire [7:0] p14_array_index_1079328_comb;
  wire [7:0] p14_array_index_1079329_comb;
  wire [7:0] p14_res7__72_comb;
  wire [7:0] p14_array_index_1079339_comb;
  wire [7:0] p14_array_index_1079340_comb;
  wire [7:0] p14_res7__73_comb;
  wire [7:0] p14_array_index_1079346_comb;
  wire [7:0] p14_array_index_1079347_comb;
  wire [7:0] p14_array_index_1079348_comb;
  wire [7:0] p14_array_index_1079349_comb;
  wire [7:0] p14_array_index_1079350_comb;
  wire [7:0] p14_array_index_1079351_comb;
  wire [7:0] p14_array_index_1079352_comb;
  wire [7:0] p14_array_index_1079353_comb;
  wire [7:0] p14_array_index_1079354_comb;
  assign p14_array_index_1079289_comb = p13_literal_1076349[p13_res7__66];
  assign p14_array_index_1079290_comb = p13_literal_1076351[p13_res7__65];
  assign p14_array_index_1079291_comb = p13_literal_1076353[p13_res7__64];
  assign p14_array_index_1079292_comb = p13_literal_1076355[p13_array_index_1079095];
  assign p14_res7__69_comb = p13_literal_1076345[p13_res7__68] ^ p13_literal_1076347[p13_res7__67] ^ p14_array_index_1079289_comb ^ p14_array_index_1079290_comb ^ p14_array_index_1079291_comb ^ p14_array_index_1079292_comb ^ p13_array_index_1079096 ^ p13_literal_1076358[p13_array_index_1079097] ^ p13_array_index_1079098 ^ p13_array_index_1079133 ^ p13_literal_1076353[p13_array_index_1079100] ^ p13_literal_1076351[p13_array_index_1079117] ^ p13_literal_1076349[p13_array_index_1079102] ^ p13_literal_1076347[p13_array_index_1079119] ^ p13_literal_1076345[p13_array_index_1079104] ^ p13_array_index_1079105;
  assign p14_array_index_1079303_comb = p13_literal_1076351[p13_res7__66];
  assign p14_array_index_1079304_comb = p13_literal_1076353[p13_res7__65];
  assign p14_array_index_1079305_comb = p13_literal_1076355[p13_res7__64];
  assign p14_res7__70_comb = p13_literal_1076345[p14_res7__69_comb] ^ p13_literal_1076347[p13_res7__68] ^ p13_literal_1076349[p13_res7__67] ^ p14_array_index_1079303_comb ^ p14_array_index_1079304_comb ^ p14_array_index_1079305_comb ^ p13_array_index_1079095 ^ p13_literal_1076358[p13_array_index_1079096] ^ p13_array_index_1079097 ^ p13_array_index_1079147 ^ p13_array_index_1079115 ^ p13_literal_1076351[p13_array_index_1079100] ^ p13_literal_1076349[p13_array_index_1079117] ^ p13_literal_1076347[p13_array_index_1079102] ^ p13_literal_1076345[p13_array_index_1079119] ^ p13_array_index_1079104;
  assign p14_array_index_1079315_comb = p13_literal_1076351[p13_res7__67];
  assign p14_array_index_1079316_comb = p13_literal_1076353[p13_res7__66];
  assign p14_array_index_1079317_comb = p13_literal_1076355[p13_res7__65];
  assign p14_res7__71_comb = p13_literal_1076345[p14_res7__70_comb] ^ p13_literal_1076347[p14_res7__69_comb] ^ p13_literal_1076349[p13_res7__68] ^ p14_array_index_1079315_comb ^ p14_array_index_1079316_comb ^ p14_array_index_1079317_comb ^ p13_res7__64 ^ p13_literal_1076358[p13_array_index_1079095] ^ p13_array_index_1079096 ^ p13_array_index_1079161 ^ p13_array_index_1079132 ^ p13_literal_1076351[p13_array_index_1079099] ^ p13_literal_1076349[p13_array_index_1079100] ^ p13_literal_1076347[p13_array_index_1079117] ^ p13_literal_1076345[p13_array_index_1079102] ^ p13_array_index_1079119;
  assign p14_array_index_1079328_comb = p13_literal_1076353[p13_res7__67];
  assign p14_array_index_1079329_comb = p13_literal_1076355[p13_res7__66];
  assign p14_res7__72_comb = p13_literal_1076345[p14_res7__71_comb] ^ p13_literal_1076347[p14_res7__70_comb] ^ p13_literal_1076349[p14_res7__69_comb] ^ p13_literal_1076351[p13_res7__68] ^ p14_array_index_1079328_comb ^ p14_array_index_1079329_comb ^ p13_res7__65 ^ p13_literal_1076358[p13_res7__64] ^ p13_array_index_1079095 ^ p13_array_index_1079175 ^ p13_array_index_1079146 ^ p13_array_index_1079114 ^ p13_literal_1076349[p13_array_index_1079099] ^ p13_literal_1076347[p13_array_index_1079100] ^ p13_literal_1076345[p13_array_index_1079117] ^ p13_array_index_1079102;
  assign p14_array_index_1079339_comb = p13_literal_1076353[p13_res7__68];
  assign p14_array_index_1079340_comb = p13_literal_1076355[p13_res7__67];
  assign p14_res7__73_comb = p13_literal_1076345[p14_res7__72_comb] ^ p13_literal_1076347[p14_res7__71_comb] ^ p13_literal_1076349[p14_res7__70_comb] ^ p13_literal_1076351[p14_res7__69_comb] ^ p14_array_index_1079339_comb ^ p14_array_index_1079340_comb ^ p13_res7__66 ^ p13_literal_1076358[p13_res7__65] ^ p13_res7__64 ^ p14_array_index_1079292_comb ^ p13_array_index_1079160 ^ p13_array_index_1079131 ^ p13_literal_1076349[p13_array_index_1079098] ^ p13_literal_1076347[p13_array_index_1079099] ^ p13_literal_1076345[p13_array_index_1079100] ^ p13_array_index_1079117;
  assign p14_array_index_1079346_comb = p13_literal_1076345[p14_res7__73_comb];
  assign p14_array_index_1079347_comb = p13_literal_1076347[p14_res7__72_comb];
  assign p14_array_index_1079348_comb = p13_literal_1076349[p14_res7__71_comb];
  assign p14_array_index_1079349_comb = p13_literal_1076351[p14_res7__70_comb];
  assign p14_array_index_1079350_comb = p13_literal_1076353[p14_res7__69_comb];
  assign p14_array_index_1079351_comb = p13_literal_1076355[p13_res7__68];
  assign p14_array_index_1079352_comb = p13_literal_1076358[p13_res7__66];
  assign p14_array_index_1079353_comb = p13_literal_1076347[p13_array_index_1079098];
  assign p14_array_index_1079354_comb = p13_literal_1076345[p13_array_index_1079099];

  // Registers for pipe stage 14:
  reg [127:0] p14_xor_1078585;
  reg [127:0] p14_xor_1079057;
  reg [7:0] p14_array_index_1079095;
  reg [7:0] p14_array_index_1079096;
  reg [7:0] p14_array_index_1079097;
  reg [7:0] p14_array_index_1079098;
  reg [7:0] p14_array_index_1079099;
  reg [7:0] p14_array_index_1079100;
  reg [7:0] p14_array_index_1079111;
  reg [7:0] p14_array_index_1079112;
  reg [7:0] p14_array_index_1079113;
  reg [7:0] p14_res7__64;
  reg [7:0] p14_array_index_1079128;
  reg [7:0] p14_array_index_1079129;
  reg [7:0] p14_array_index_1079130;
  reg [7:0] p14_res7__65;
  reg [7:0] p14_array_index_1079143;
  reg [7:0] p14_array_index_1079144;
  reg [7:0] p14_array_index_1079145;
  reg [7:0] p14_res7__66;
  reg [7:0] p14_array_index_1079157;
  reg [7:0] p14_array_index_1079158;
  reg [7:0] p14_array_index_1079159;
  reg [7:0] p14_res7__67;
  reg [7:0] p14_array_index_1079172;
  reg [7:0] p14_array_index_1079173;
  reg [7:0] p14_array_index_1079174;
  reg [7:0] p14_res7__68;
  reg [7:0] p14_array_index_1079289;
  reg [7:0] p14_array_index_1079290;
  reg [7:0] p14_array_index_1079291;
  reg [7:0] p14_res7__69;
  reg [7:0] p14_array_index_1079303;
  reg [7:0] p14_array_index_1079304;
  reg [7:0] p14_array_index_1079305;
  reg [7:0] p14_res7__70;
  reg [7:0] p14_array_index_1079315;
  reg [7:0] p14_array_index_1079316;
  reg [7:0] p14_array_index_1079317;
  reg [7:0] p14_res7__71;
  reg [7:0] p14_array_index_1079328;
  reg [7:0] p14_array_index_1079329;
  reg [7:0] p14_res7__72;
  reg [7:0] p14_array_index_1079339;
  reg [7:0] p14_array_index_1079340;
  reg [7:0] p14_res7__73;
  reg [7:0] p14_array_index_1079346;
  reg [7:0] p14_array_index_1079347;
  reg [7:0] p14_array_index_1079348;
  reg [7:0] p14_array_index_1079349;
  reg [7:0] p14_array_index_1079350;
  reg [7:0] p14_array_index_1079351;
  reg [7:0] p14_array_index_1079352;
  reg [7:0] p14_array_index_1079353;
  reg [7:0] p14_array_index_1079354;
  reg [127:0] p14_res__33;
  reg [7:0] p15_arr[256];
  reg [7:0] p15_literal_1076345[256];
  reg [7:0] p15_literal_1076347[256];
  reg [7:0] p15_literal_1076349[256];
  reg [7:0] p15_literal_1076351[256];
  reg [7:0] p15_literal_1076353[256];
  reg [7:0] p15_literal_1076355[256];
  reg [7:0] p15_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p14_xor_1078585 <= p13_xor_1078585;
    p14_xor_1079057 <= p13_xor_1079057;
    p14_array_index_1079095 <= p13_array_index_1079095;
    p14_array_index_1079096 <= p13_array_index_1079096;
    p14_array_index_1079097 <= p13_array_index_1079097;
    p14_array_index_1079098 <= p13_array_index_1079098;
    p14_array_index_1079099 <= p13_array_index_1079099;
    p14_array_index_1079100 <= p13_array_index_1079100;
    p14_array_index_1079111 <= p13_array_index_1079111;
    p14_array_index_1079112 <= p13_array_index_1079112;
    p14_array_index_1079113 <= p13_array_index_1079113;
    p14_res7__64 <= p13_res7__64;
    p14_array_index_1079128 <= p13_array_index_1079128;
    p14_array_index_1079129 <= p13_array_index_1079129;
    p14_array_index_1079130 <= p13_array_index_1079130;
    p14_res7__65 <= p13_res7__65;
    p14_array_index_1079143 <= p13_array_index_1079143;
    p14_array_index_1079144 <= p13_array_index_1079144;
    p14_array_index_1079145 <= p13_array_index_1079145;
    p14_res7__66 <= p13_res7__66;
    p14_array_index_1079157 <= p13_array_index_1079157;
    p14_array_index_1079158 <= p13_array_index_1079158;
    p14_array_index_1079159 <= p13_array_index_1079159;
    p14_res7__67 <= p13_res7__67;
    p14_array_index_1079172 <= p13_array_index_1079172;
    p14_array_index_1079173 <= p13_array_index_1079173;
    p14_array_index_1079174 <= p13_array_index_1079174;
    p14_res7__68 <= p13_res7__68;
    p14_array_index_1079289 <= p14_array_index_1079289_comb;
    p14_array_index_1079290 <= p14_array_index_1079290_comb;
    p14_array_index_1079291 <= p14_array_index_1079291_comb;
    p14_res7__69 <= p14_res7__69_comb;
    p14_array_index_1079303 <= p14_array_index_1079303_comb;
    p14_array_index_1079304 <= p14_array_index_1079304_comb;
    p14_array_index_1079305 <= p14_array_index_1079305_comb;
    p14_res7__70 <= p14_res7__70_comb;
    p14_array_index_1079315 <= p14_array_index_1079315_comb;
    p14_array_index_1079316 <= p14_array_index_1079316_comb;
    p14_array_index_1079317 <= p14_array_index_1079317_comb;
    p14_res7__71 <= p14_res7__71_comb;
    p14_array_index_1079328 <= p14_array_index_1079328_comb;
    p14_array_index_1079329 <= p14_array_index_1079329_comb;
    p14_res7__72 <= p14_res7__72_comb;
    p14_array_index_1079339 <= p14_array_index_1079339_comb;
    p14_array_index_1079340 <= p14_array_index_1079340_comb;
    p14_res7__73 <= p14_res7__73_comb;
    p14_array_index_1079346 <= p14_array_index_1079346_comb;
    p14_array_index_1079347 <= p14_array_index_1079347_comb;
    p14_array_index_1079348 <= p14_array_index_1079348_comb;
    p14_array_index_1079349 <= p14_array_index_1079349_comb;
    p14_array_index_1079350 <= p14_array_index_1079350_comb;
    p14_array_index_1079351 <= p14_array_index_1079351_comb;
    p14_array_index_1079352 <= p14_array_index_1079352_comb;
    p14_array_index_1079353 <= p14_array_index_1079353_comb;
    p14_array_index_1079354 <= p14_array_index_1079354_comb;
    p14_res__33 <= p13_res__33;
    p15_arr <= p14_arr;
    p15_literal_1076345 <= p14_literal_1076345;
    p15_literal_1076347 <= p14_literal_1076347;
    p15_literal_1076349 <= p14_literal_1076349;
    p15_literal_1076351 <= p14_literal_1076351;
    p15_literal_1076353 <= p14_literal_1076353;
    p15_literal_1076355 <= p14_literal_1076355;
    p15_literal_1076358 <= p14_literal_1076358;
  end

  // ===== Pipe stage 15:
  wire [7:0] p15_res7__74_comb;
  wire [7:0] p15_array_index_1079489_comb;
  wire [7:0] p15_res7__75_comb;
  wire [7:0] p15_res7__76_comb;
  wire [7:0] p15_res7__77_comb;
  wire [7:0] p15_res7__78_comb;
  wire [7:0] p15_res7__79_comb;
  wire [127:0] p15_res__4_comb;
  wire [127:0] p15_xor_1079529_comb;
  assign p15_res7__74_comb = p14_array_index_1079346 ^ p14_array_index_1079347 ^ p14_array_index_1079348 ^ p14_array_index_1079349 ^ p14_array_index_1079350 ^ p14_array_index_1079351 ^ p14_res7__67 ^ p14_array_index_1079352 ^ p14_res7__65 ^ p14_array_index_1079305 ^ p14_array_index_1079174 ^ p14_array_index_1079145 ^ p14_array_index_1079113 ^ p14_array_index_1079353 ^ p14_array_index_1079354 ^ p14_array_index_1079100;
  assign p15_array_index_1079489_comb = p14_literal_1076355[p14_res7__69];
  assign p15_res7__75_comb = p14_literal_1076345[p15_res7__74_comb] ^ p14_literal_1076347[p14_res7__73] ^ p14_literal_1076349[p14_res7__72] ^ p14_literal_1076351[p14_res7__71] ^ p14_literal_1076353[p14_res7__70] ^ p15_array_index_1079489_comb ^ p14_res7__68 ^ p14_literal_1076358[p14_res7__67] ^ p14_res7__66 ^ p14_array_index_1079317 ^ p14_array_index_1079291 ^ p14_array_index_1079159 ^ p14_array_index_1079130 ^ p14_literal_1076347[p14_array_index_1079097] ^ p14_literal_1076345[p14_array_index_1079098] ^ p14_array_index_1079099;
  assign p15_res7__76_comb = p14_literal_1076345[p15_res7__75_comb] ^ p14_literal_1076347[p15_res7__74_comb] ^ p14_literal_1076349[p14_res7__73] ^ p14_literal_1076351[p14_res7__72] ^ p14_literal_1076353[p14_res7__71] ^ p14_literal_1076355[p14_res7__70] ^ p14_res7__69 ^ p14_literal_1076358[p14_res7__68] ^ p14_res7__67 ^ p14_array_index_1079329 ^ p14_array_index_1079304 ^ p14_array_index_1079173 ^ p14_array_index_1079144 ^ p14_array_index_1079112 ^ p14_literal_1076345[p14_array_index_1079097] ^ p14_array_index_1079098;
  assign p15_res7__77_comb = p14_literal_1076345[p15_res7__76_comb] ^ p14_literal_1076347[p15_res7__75_comb] ^ p14_literal_1076349[p15_res7__74_comb] ^ p14_literal_1076351[p14_res7__73] ^ p14_literal_1076353[p14_res7__72] ^ p14_literal_1076355[p14_res7__71] ^ p14_res7__70 ^ p14_literal_1076358[p14_res7__69] ^ p14_res7__68 ^ p14_array_index_1079340 ^ p14_array_index_1079316 ^ p14_array_index_1079290 ^ p14_array_index_1079158 ^ p14_array_index_1079129 ^ p14_literal_1076345[p14_array_index_1079096] ^ p14_array_index_1079097;
  assign p15_res7__78_comb = p14_literal_1076345[p15_res7__77_comb] ^ p14_literal_1076347[p15_res7__76_comb] ^ p14_literal_1076349[p15_res7__75_comb] ^ p14_literal_1076351[p15_res7__74_comb] ^ p14_literal_1076353[p14_res7__73] ^ p14_literal_1076355[p14_res7__72] ^ p14_res7__71 ^ p14_literal_1076358[p14_res7__70] ^ p14_res7__69 ^ p14_array_index_1079351 ^ p14_array_index_1079328 ^ p14_array_index_1079303 ^ p14_array_index_1079172 ^ p14_array_index_1079143 ^ p14_array_index_1079111 ^ p14_array_index_1079096;
  assign p15_res7__79_comb = p14_literal_1076345[p15_res7__78_comb] ^ p14_literal_1076347[p15_res7__77_comb] ^ p14_literal_1076349[p15_res7__76_comb] ^ p14_literal_1076351[p15_res7__75_comb] ^ p14_literal_1076353[p15_res7__74_comb] ^ p14_literal_1076355[p14_res7__73] ^ p14_res7__72 ^ p14_literal_1076358[p14_res7__71] ^ p14_res7__70 ^ p15_array_index_1079489_comb ^ p14_array_index_1079339 ^ p14_array_index_1079315 ^ p14_array_index_1079289 ^ p14_array_index_1079157 ^ p14_array_index_1079128 ^ p14_array_index_1079095;
  assign p15_res__4_comb = {p15_res7__79_comb, p15_res7__78_comb, p15_res7__77_comb, p15_res7__76_comb, p15_res7__75_comb, p15_res7__74_comb, p14_res7__73, p14_res7__72, p14_res7__71, p14_res7__70, p14_res7__69, p14_res7__68, p14_res7__67, p14_res7__66, p14_res7__65, p14_res7__64};
  assign p15_xor_1079529_comb = p15_res__4_comb ^ p14_xor_1078585;

  // Registers for pipe stage 15:
  reg [127:0] p15_xor_1079057;
  reg [127:0] p15_xor_1079529;
  reg [127:0] p15_res__33;
  reg [7:0] p16_arr[256];
  reg [7:0] p16_literal_1076345[256];
  reg [7:0] p16_literal_1076347[256];
  reg [7:0] p16_literal_1076349[256];
  reg [7:0] p16_literal_1076351[256];
  reg [7:0] p16_literal_1076353[256];
  reg [7:0] p16_literal_1076355[256];
  reg [7:0] p16_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p15_xor_1079057 <= p14_xor_1079057;
    p15_xor_1079529 <= p15_xor_1079529_comb;
    p15_res__33 <= p14_res__33;
    p16_arr <= p15_arr;
    p16_literal_1076345 <= p15_literal_1076345;
    p16_literal_1076347 <= p15_literal_1076347;
    p16_literal_1076349 <= p15_literal_1076349;
    p16_literal_1076351 <= p15_literal_1076351;
    p16_literal_1076353 <= p15_literal_1076353;
    p16_literal_1076355 <= p15_literal_1076355;
    p16_literal_1076358 <= p15_literal_1076358;
  end

  // ===== Pipe stage 16:
  wire [127:0] p16_addedKey__46_comb;
  wire [7:0] p16_array_index_1079567_comb;
  wire [7:0] p16_array_index_1079568_comb;
  wire [7:0] p16_array_index_1079569_comb;
  wire [7:0] p16_array_index_1079570_comb;
  wire [7:0] p16_array_index_1079571_comb;
  wire [7:0] p16_array_index_1079572_comb;
  wire [7:0] p16_array_index_1079574_comb;
  wire [7:0] p16_array_index_1079576_comb;
  wire [7:0] p16_array_index_1079577_comb;
  wire [7:0] p16_array_index_1079578_comb;
  wire [7:0] p16_array_index_1079579_comb;
  wire [7:0] p16_array_index_1079580_comb;
  wire [7:0] p16_array_index_1079581_comb;
  wire [7:0] p16_array_index_1079583_comb;
  wire [7:0] p16_array_index_1079584_comb;
  wire [7:0] p16_array_index_1079585_comb;
  wire [7:0] p16_array_index_1079586_comb;
  wire [7:0] p16_array_index_1079587_comb;
  wire [7:0] p16_array_index_1079588_comb;
  wire [7:0] p16_array_index_1079589_comb;
  wire [7:0] p16_array_index_1079591_comb;
  wire [7:0] p16_res7__80_comb;
  wire [7:0] p16_array_index_1079600_comb;
  wire [7:0] p16_array_index_1079601_comb;
  wire [7:0] p16_array_index_1079602_comb;
  wire [7:0] p16_array_index_1079603_comb;
  wire [7:0] p16_array_index_1079604_comb;
  wire [7:0] p16_array_index_1079605_comb;
  wire [7:0] p16_res7__81_comb;
  wire [7:0] p16_array_index_1079615_comb;
  wire [7:0] p16_array_index_1079616_comb;
  wire [7:0] p16_array_index_1079617_comb;
  wire [7:0] p16_array_index_1079618_comb;
  wire [7:0] p16_array_index_1079619_comb;
  wire [7:0] p16_res7__82_comb;
  wire [7:0] p16_array_index_1079629_comb;
  wire [7:0] p16_array_index_1079630_comb;
  wire [7:0] p16_array_index_1079631_comb;
  wire [7:0] p16_array_index_1079632_comb;
  wire [7:0] p16_array_index_1079633_comb;
  wire [7:0] p16_res7__83_comb;
  wire [7:0] p16_array_index_1079644_comb;
  wire [7:0] p16_array_index_1079645_comb;
  wire [7:0] p16_array_index_1079646_comb;
  wire [7:0] p16_array_index_1079647_comb;
  wire [7:0] p16_res7__84_comb;
  assign p16_addedKey__46_comb = p15_xor_1079529 ^ 128'ha74a_f7ef_ab73_df16_0dd2_0860_8b9e_fe06;
  assign p16_array_index_1079567_comb = p15_arr[p16_addedKey__46_comb[127:120]];
  assign p16_array_index_1079568_comb = p15_arr[p16_addedKey__46_comb[119:112]];
  assign p16_array_index_1079569_comb = p15_arr[p16_addedKey__46_comb[111:104]];
  assign p16_array_index_1079570_comb = p15_arr[p16_addedKey__46_comb[103:96]];
  assign p16_array_index_1079571_comb = p15_arr[p16_addedKey__46_comb[95:88]];
  assign p16_array_index_1079572_comb = p15_arr[p16_addedKey__46_comb[87:80]];
  assign p16_array_index_1079574_comb = p15_arr[p16_addedKey__46_comb[71:64]];
  assign p16_array_index_1079576_comb = p15_arr[p16_addedKey__46_comb[55:48]];
  assign p16_array_index_1079577_comb = p15_arr[p16_addedKey__46_comb[47:40]];
  assign p16_array_index_1079578_comb = p15_arr[p16_addedKey__46_comb[39:32]];
  assign p16_array_index_1079579_comb = p15_arr[p16_addedKey__46_comb[31:24]];
  assign p16_array_index_1079580_comb = p15_arr[p16_addedKey__46_comb[23:16]];
  assign p16_array_index_1079581_comb = p15_arr[p16_addedKey__46_comb[15:8]];
  assign p16_array_index_1079583_comb = p15_literal_1076345[p16_array_index_1079567_comb];
  assign p16_array_index_1079584_comb = p15_literal_1076347[p16_array_index_1079568_comb];
  assign p16_array_index_1079585_comb = p15_literal_1076349[p16_array_index_1079569_comb];
  assign p16_array_index_1079586_comb = p15_literal_1076351[p16_array_index_1079570_comb];
  assign p16_array_index_1079587_comb = p15_literal_1076353[p16_array_index_1079571_comb];
  assign p16_array_index_1079588_comb = p15_literal_1076355[p16_array_index_1079572_comb];
  assign p16_array_index_1079589_comb = p15_arr[p16_addedKey__46_comb[79:72]];
  assign p16_array_index_1079591_comb = p15_arr[p16_addedKey__46_comb[63:56]];
  assign p16_res7__80_comb = p16_array_index_1079583_comb ^ p16_array_index_1079584_comb ^ p16_array_index_1079585_comb ^ p16_array_index_1079586_comb ^ p16_array_index_1079587_comb ^ p16_array_index_1079588_comb ^ p16_array_index_1079589_comb ^ p15_literal_1076358[p16_array_index_1079574_comb] ^ p16_array_index_1079591_comb ^ p15_literal_1076355[p16_array_index_1079576_comb] ^ p15_literal_1076353[p16_array_index_1079577_comb] ^ p15_literal_1076351[p16_array_index_1079578_comb] ^ p15_literal_1076349[p16_array_index_1079579_comb] ^ p15_literal_1076347[p16_array_index_1079580_comb] ^ p15_literal_1076345[p16_array_index_1079581_comb] ^ p15_arr[p16_addedKey__46_comb[7:0]];
  assign p16_array_index_1079600_comb = p15_literal_1076345[p16_res7__80_comb];
  assign p16_array_index_1079601_comb = p15_literal_1076347[p16_array_index_1079567_comb];
  assign p16_array_index_1079602_comb = p15_literal_1076349[p16_array_index_1079568_comb];
  assign p16_array_index_1079603_comb = p15_literal_1076351[p16_array_index_1079569_comb];
  assign p16_array_index_1079604_comb = p15_literal_1076353[p16_array_index_1079570_comb];
  assign p16_array_index_1079605_comb = p15_literal_1076355[p16_array_index_1079571_comb];
  assign p16_res7__81_comb = p16_array_index_1079600_comb ^ p16_array_index_1079601_comb ^ p16_array_index_1079602_comb ^ p16_array_index_1079603_comb ^ p16_array_index_1079604_comb ^ p16_array_index_1079605_comb ^ p16_array_index_1079572_comb ^ p15_literal_1076358[p16_array_index_1079589_comb] ^ p16_array_index_1079574_comb ^ p15_literal_1076355[p16_array_index_1079591_comb] ^ p15_literal_1076353[p16_array_index_1079576_comb] ^ p15_literal_1076351[p16_array_index_1079577_comb] ^ p15_literal_1076349[p16_array_index_1079578_comb] ^ p15_literal_1076347[p16_array_index_1079579_comb] ^ p15_literal_1076345[p16_array_index_1079580_comb] ^ p16_array_index_1079581_comb;
  assign p16_array_index_1079615_comb = p15_literal_1076347[p16_res7__80_comb];
  assign p16_array_index_1079616_comb = p15_literal_1076349[p16_array_index_1079567_comb];
  assign p16_array_index_1079617_comb = p15_literal_1076351[p16_array_index_1079568_comb];
  assign p16_array_index_1079618_comb = p15_literal_1076353[p16_array_index_1079569_comb];
  assign p16_array_index_1079619_comb = p15_literal_1076355[p16_array_index_1079570_comb];
  assign p16_res7__82_comb = p15_literal_1076345[p16_res7__81_comb] ^ p16_array_index_1079615_comb ^ p16_array_index_1079616_comb ^ p16_array_index_1079617_comb ^ p16_array_index_1079618_comb ^ p16_array_index_1079619_comb ^ p16_array_index_1079571_comb ^ p15_literal_1076358[p16_array_index_1079572_comb] ^ p16_array_index_1079589_comb ^ p15_literal_1076355[p16_array_index_1079574_comb] ^ p15_literal_1076353[p16_array_index_1079591_comb] ^ p15_literal_1076351[p16_array_index_1079576_comb] ^ p15_literal_1076349[p16_array_index_1079577_comb] ^ p15_literal_1076347[p16_array_index_1079578_comb] ^ p15_literal_1076345[p16_array_index_1079579_comb] ^ p16_array_index_1079580_comb;
  assign p16_array_index_1079629_comb = p15_literal_1076347[p16_res7__81_comb];
  assign p16_array_index_1079630_comb = p15_literal_1076349[p16_res7__80_comb];
  assign p16_array_index_1079631_comb = p15_literal_1076351[p16_array_index_1079567_comb];
  assign p16_array_index_1079632_comb = p15_literal_1076353[p16_array_index_1079568_comb];
  assign p16_array_index_1079633_comb = p15_literal_1076355[p16_array_index_1079569_comb];
  assign p16_res7__83_comb = p15_literal_1076345[p16_res7__82_comb] ^ p16_array_index_1079629_comb ^ p16_array_index_1079630_comb ^ p16_array_index_1079631_comb ^ p16_array_index_1079632_comb ^ p16_array_index_1079633_comb ^ p16_array_index_1079570_comb ^ p15_literal_1076358[p16_array_index_1079571_comb] ^ p16_array_index_1079572_comb ^ p15_literal_1076355[p16_array_index_1079589_comb] ^ p15_literal_1076353[p16_array_index_1079574_comb] ^ p15_literal_1076351[p16_array_index_1079591_comb] ^ p15_literal_1076349[p16_array_index_1079576_comb] ^ p15_literal_1076347[p16_array_index_1079577_comb] ^ p15_literal_1076345[p16_array_index_1079578_comb] ^ p16_array_index_1079579_comb;
  assign p16_array_index_1079644_comb = p15_literal_1076349[p16_res7__81_comb];
  assign p16_array_index_1079645_comb = p15_literal_1076351[p16_res7__80_comb];
  assign p16_array_index_1079646_comb = p15_literal_1076353[p16_array_index_1079567_comb];
  assign p16_array_index_1079647_comb = p15_literal_1076355[p16_array_index_1079568_comb];
  assign p16_res7__84_comb = p15_literal_1076345[p16_res7__83_comb] ^ p15_literal_1076347[p16_res7__82_comb] ^ p16_array_index_1079644_comb ^ p16_array_index_1079645_comb ^ p16_array_index_1079646_comb ^ p16_array_index_1079647_comb ^ p16_array_index_1079569_comb ^ p15_literal_1076358[p16_array_index_1079570_comb] ^ p16_array_index_1079571_comb ^ p16_array_index_1079588_comb ^ p15_literal_1076353[p16_array_index_1079589_comb] ^ p15_literal_1076351[p16_array_index_1079574_comb] ^ p15_literal_1076349[p16_array_index_1079591_comb] ^ p15_literal_1076347[p16_array_index_1079576_comb] ^ p15_literal_1076345[p16_array_index_1079577_comb] ^ p16_array_index_1079578_comb;

  // Registers for pipe stage 16:
  reg [127:0] p16_xor_1079057;
  reg [127:0] p16_xor_1079529;
  reg [7:0] p16_array_index_1079567;
  reg [7:0] p16_array_index_1079568;
  reg [7:0] p16_array_index_1079569;
  reg [7:0] p16_array_index_1079570;
  reg [7:0] p16_array_index_1079571;
  reg [7:0] p16_array_index_1079572;
  reg [7:0] p16_array_index_1079574;
  reg [7:0] p16_array_index_1079576;
  reg [7:0] p16_array_index_1079577;
  reg [7:0] p16_array_index_1079583;
  reg [7:0] p16_array_index_1079584;
  reg [7:0] p16_array_index_1079585;
  reg [7:0] p16_array_index_1079586;
  reg [7:0] p16_array_index_1079587;
  reg [7:0] p16_array_index_1079589;
  reg [7:0] p16_array_index_1079591;
  reg [7:0] p16_res7__80;
  reg [7:0] p16_array_index_1079600;
  reg [7:0] p16_array_index_1079601;
  reg [7:0] p16_array_index_1079602;
  reg [7:0] p16_array_index_1079603;
  reg [7:0] p16_array_index_1079604;
  reg [7:0] p16_array_index_1079605;
  reg [7:0] p16_res7__81;
  reg [7:0] p16_array_index_1079615;
  reg [7:0] p16_array_index_1079616;
  reg [7:0] p16_array_index_1079617;
  reg [7:0] p16_array_index_1079618;
  reg [7:0] p16_array_index_1079619;
  reg [7:0] p16_res7__82;
  reg [7:0] p16_array_index_1079629;
  reg [7:0] p16_array_index_1079630;
  reg [7:0] p16_array_index_1079631;
  reg [7:0] p16_array_index_1079632;
  reg [7:0] p16_array_index_1079633;
  reg [7:0] p16_res7__83;
  reg [7:0] p16_array_index_1079644;
  reg [7:0] p16_array_index_1079645;
  reg [7:0] p16_array_index_1079646;
  reg [7:0] p16_array_index_1079647;
  reg [7:0] p16_res7__84;
  reg [127:0] p16_res__33;
  reg [7:0] p17_arr[256];
  reg [7:0] p17_literal_1076345[256];
  reg [7:0] p17_literal_1076347[256];
  reg [7:0] p17_literal_1076349[256];
  reg [7:0] p17_literal_1076351[256];
  reg [7:0] p17_literal_1076353[256];
  reg [7:0] p17_literal_1076355[256];
  reg [7:0] p17_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p16_xor_1079057 <= p15_xor_1079057;
    p16_xor_1079529 <= p15_xor_1079529;
    p16_array_index_1079567 <= p16_array_index_1079567_comb;
    p16_array_index_1079568 <= p16_array_index_1079568_comb;
    p16_array_index_1079569 <= p16_array_index_1079569_comb;
    p16_array_index_1079570 <= p16_array_index_1079570_comb;
    p16_array_index_1079571 <= p16_array_index_1079571_comb;
    p16_array_index_1079572 <= p16_array_index_1079572_comb;
    p16_array_index_1079574 <= p16_array_index_1079574_comb;
    p16_array_index_1079576 <= p16_array_index_1079576_comb;
    p16_array_index_1079577 <= p16_array_index_1079577_comb;
    p16_array_index_1079583 <= p16_array_index_1079583_comb;
    p16_array_index_1079584 <= p16_array_index_1079584_comb;
    p16_array_index_1079585 <= p16_array_index_1079585_comb;
    p16_array_index_1079586 <= p16_array_index_1079586_comb;
    p16_array_index_1079587 <= p16_array_index_1079587_comb;
    p16_array_index_1079589 <= p16_array_index_1079589_comb;
    p16_array_index_1079591 <= p16_array_index_1079591_comb;
    p16_res7__80 <= p16_res7__80_comb;
    p16_array_index_1079600 <= p16_array_index_1079600_comb;
    p16_array_index_1079601 <= p16_array_index_1079601_comb;
    p16_array_index_1079602 <= p16_array_index_1079602_comb;
    p16_array_index_1079603 <= p16_array_index_1079603_comb;
    p16_array_index_1079604 <= p16_array_index_1079604_comb;
    p16_array_index_1079605 <= p16_array_index_1079605_comb;
    p16_res7__81 <= p16_res7__81_comb;
    p16_array_index_1079615 <= p16_array_index_1079615_comb;
    p16_array_index_1079616 <= p16_array_index_1079616_comb;
    p16_array_index_1079617 <= p16_array_index_1079617_comb;
    p16_array_index_1079618 <= p16_array_index_1079618_comb;
    p16_array_index_1079619 <= p16_array_index_1079619_comb;
    p16_res7__82 <= p16_res7__82_comb;
    p16_array_index_1079629 <= p16_array_index_1079629_comb;
    p16_array_index_1079630 <= p16_array_index_1079630_comb;
    p16_array_index_1079631 <= p16_array_index_1079631_comb;
    p16_array_index_1079632 <= p16_array_index_1079632_comb;
    p16_array_index_1079633 <= p16_array_index_1079633_comb;
    p16_res7__83 <= p16_res7__83_comb;
    p16_array_index_1079644 <= p16_array_index_1079644_comb;
    p16_array_index_1079645 <= p16_array_index_1079645_comb;
    p16_array_index_1079646 <= p16_array_index_1079646_comb;
    p16_array_index_1079647 <= p16_array_index_1079647_comb;
    p16_res7__84 <= p16_res7__84_comb;
    p16_res__33 <= p15_res__33;
    p17_arr <= p16_arr;
    p17_literal_1076345 <= p16_literal_1076345;
    p17_literal_1076347 <= p16_literal_1076347;
    p17_literal_1076349 <= p16_literal_1076349;
    p17_literal_1076351 <= p16_literal_1076351;
    p17_literal_1076353 <= p16_literal_1076353;
    p17_literal_1076355 <= p16_literal_1076355;
    p17_literal_1076358 <= p16_literal_1076358;
  end

  // ===== Pipe stage 17:
  wire [7:0] p17_array_index_1079761_comb;
  wire [7:0] p17_array_index_1079762_comb;
  wire [7:0] p17_array_index_1079763_comb;
  wire [7:0] p17_array_index_1079764_comb;
  wire [7:0] p17_res7__85_comb;
  wire [7:0] p17_array_index_1079775_comb;
  wire [7:0] p17_array_index_1079776_comb;
  wire [7:0] p17_array_index_1079777_comb;
  wire [7:0] p17_res7__86_comb;
  wire [7:0] p17_array_index_1079787_comb;
  wire [7:0] p17_array_index_1079788_comb;
  wire [7:0] p17_array_index_1079789_comb;
  wire [7:0] p17_res7__87_comb;
  wire [7:0] p17_array_index_1079800_comb;
  wire [7:0] p17_array_index_1079801_comb;
  wire [7:0] p17_res7__88_comb;
  wire [7:0] p17_array_index_1079811_comb;
  wire [7:0] p17_array_index_1079812_comb;
  wire [7:0] p17_res7__89_comb;
  wire [7:0] p17_array_index_1079818_comb;
  wire [7:0] p17_array_index_1079819_comb;
  wire [7:0] p17_array_index_1079820_comb;
  wire [7:0] p17_array_index_1079821_comb;
  wire [7:0] p17_array_index_1079822_comb;
  wire [7:0] p17_array_index_1079823_comb;
  wire [7:0] p17_array_index_1079824_comb;
  wire [7:0] p17_array_index_1079825_comb;
  wire [7:0] p17_array_index_1079826_comb;
  assign p17_array_index_1079761_comb = p16_literal_1076349[p16_res7__82];
  assign p17_array_index_1079762_comb = p16_literal_1076351[p16_res7__81];
  assign p17_array_index_1079763_comb = p16_literal_1076353[p16_res7__80];
  assign p17_array_index_1079764_comb = p16_literal_1076355[p16_array_index_1079567];
  assign p17_res7__85_comb = p16_literal_1076345[p16_res7__84] ^ p16_literal_1076347[p16_res7__83] ^ p17_array_index_1079761_comb ^ p17_array_index_1079762_comb ^ p17_array_index_1079763_comb ^ p17_array_index_1079764_comb ^ p16_array_index_1079568 ^ p16_literal_1076358[p16_array_index_1079569] ^ p16_array_index_1079570 ^ p16_array_index_1079605 ^ p16_literal_1076353[p16_array_index_1079572] ^ p16_literal_1076351[p16_array_index_1079589] ^ p16_literal_1076349[p16_array_index_1079574] ^ p16_literal_1076347[p16_array_index_1079591] ^ p16_literal_1076345[p16_array_index_1079576] ^ p16_array_index_1079577;
  assign p17_array_index_1079775_comb = p16_literal_1076351[p16_res7__82];
  assign p17_array_index_1079776_comb = p16_literal_1076353[p16_res7__81];
  assign p17_array_index_1079777_comb = p16_literal_1076355[p16_res7__80];
  assign p17_res7__86_comb = p16_literal_1076345[p17_res7__85_comb] ^ p16_literal_1076347[p16_res7__84] ^ p16_literal_1076349[p16_res7__83] ^ p17_array_index_1079775_comb ^ p17_array_index_1079776_comb ^ p17_array_index_1079777_comb ^ p16_array_index_1079567 ^ p16_literal_1076358[p16_array_index_1079568] ^ p16_array_index_1079569 ^ p16_array_index_1079619 ^ p16_array_index_1079587 ^ p16_literal_1076351[p16_array_index_1079572] ^ p16_literal_1076349[p16_array_index_1079589] ^ p16_literal_1076347[p16_array_index_1079574] ^ p16_literal_1076345[p16_array_index_1079591] ^ p16_array_index_1079576;
  assign p17_array_index_1079787_comb = p16_literal_1076351[p16_res7__83];
  assign p17_array_index_1079788_comb = p16_literal_1076353[p16_res7__82];
  assign p17_array_index_1079789_comb = p16_literal_1076355[p16_res7__81];
  assign p17_res7__87_comb = p16_literal_1076345[p17_res7__86_comb] ^ p16_literal_1076347[p17_res7__85_comb] ^ p16_literal_1076349[p16_res7__84] ^ p17_array_index_1079787_comb ^ p17_array_index_1079788_comb ^ p17_array_index_1079789_comb ^ p16_res7__80 ^ p16_literal_1076358[p16_array_index_1079567] ^ p16_array_index_1079568 ^ p16_array_index_1079633 ^ p16_array_index_1079604 ^ p16_literal_1076351[p16_array_index_1079571] ^ p16_literal_1076349[p16_array_index_1079572] ^ p16_literal_1076347[p16_array_index_1079589] ^ p16_literal_1076345[p16_array_index_1079574] ^ p16_array_index_1079591;
  assign p17_array_index_1079800_comb = p16_literal_1076353[p16_res7__83];
  assign p17_array_index_1079801_comb = p16_literal_1076355[p16_res7__82];
  assign p17_res7__88_comb = p16_literal_1076345[p17_res7__87_comb] ^ p16_literal_1076347[p17_res7__86_comb] ^ p16_literal_1076349[p17_res7__85_comb] ^ p16_literal_1076351[p16_res7__84] ^ p17_array_index_1079800_comb ^ p17_array_index_1079801_comb ^ p16_res7__81 ^ p16_literal_1076358[p16_res7__80] ^ p16_array_index_1079567 ^ p16_array_index_1079647 ^ p16_array_index_1079618 ^ p16_array_index_1079586 ^ p16_literal_1076349[p16_array_index_1079571] ^ p16_literal_1076347[p16_array_index_1079572] ^ p16_literal_1076345[p16_array_index_1079589] ^ p16_array_index_1079574;
  assign p17_array_index_1079811_comb = p16_literal_1076353[p16_res7__84];
  assign p17_array_index_1079812_comb = p16_literal_1076355[p16_res7__83];
  assign p17_res7__89_comb = p16_literal_1076345[p17_res7__88_comb] ^ p16_literal_1076347[p17_res7__87_comb] ^ p16_literal_1076349[p17_res7__86_comb] ^ p16_literal_1076351[p17_res7__85_comb] ^ p17_array_index_1079811_comb ^ p17_array_index_1079812_comb ^ p16_res7__82 ^ p16_literal_1076358[p16_res7__81] ^ p16_res7__80 ^ p17_array_index_1079764_comb ^ p16_array_index_1079632 ^ p16_array_index_1079603 ^ p16_literal_1076349[p16_array_index_1079570] ^ p16_literal_1076347[p16_array_index_1079571] ^ p16_literal_1076345[p16_array_index_1079572] ^ p16_array_index_1079589;
  assign p17_array_index_1079818_comb = p16_literal_1076345[p17_res7__89_comb];
  assign p17_array_index_1079819_comb = p16_literal_1076347[p17_res7__88_comb];
  assign p17_array_index_1079820_comb = p16_literal_1076349[p17_res7__87_comb];
  assign p17_array_index_1079821_comb = p16_literal_1076351[p17_res7__86_comb];
  assign p17_array_index_1079822_comb = p16_literal_1076353[p17_res7__85_comb];
  assign p17_array_index_1079823_comb = p16_literal_1076355[p16_res7__84];
  assign p17_array_index_1079824_comb = p16_literal_1076358[p16_res7__82];
  assign p17_array_index_1079825_comb = p16_literal_1076347[p16_array_index_1079570];
  assign p17_array_index_1079826_comb = p16_literal_1076345[p16_array_index_1079571];

  // Registers for pipe stage 17:
  reg [127:0] p17_xor_1079057;
  reg [127:0] p17_xor_1079529;
  reg [7:0] p17_array_index_1079567;
  reg [7:0] p17_array_index_1079568;
  reg [7:0] p17_array_index_1079569;
  reg [7:0] p17_array_index_1079570;
  reg [7:0] p17_array_index_1079571;
  reg [7:0] p17_array_index_1079572;
  reg [7:0] p17_array_index_1079583;
  reg [7:0] p17_array_index_1079584;
  reg [7:0] p17_array_index_1079585;
  reg [7:0] p17_res7__80;
  reg [7:0] p17_array_index_1079600;
  reg [7:0] p17_array_index_1079601;
  reg [7:0] p17_array_index_1079602;
  reg [7:0] p17_res7__81;
  reg [7:0] p17_array_index_1079615;
  reg [7:0] p17_array_index_1079616;
  reg [7:0] p17_array_index_1079617;
  reg [7:0] p17_res7__82;
  reg [7:0] p17_array_index_1079629;
  reg [7:0] p17_array_index_1079630;
  reg [7:0] p17_array_index_1079631;
  reg [7:0] p17_res7__83;
  reg [7:0] p17_array_index_1079644;
  reg [7:0] p17_array_index_1079645;
  reg [7:0] p17_array_index_1079646;
  reg [7:0] p17_res7__84;
  reg [7:0] p17_array_index_1079761;
  reg [7:0] p17_array_index_1079762;
  reg [7:0] p17_array_index_1079763;
  reg [7:0] p17_res7__85;
  reg [7:0] p17_array_index_1079775;
  reg [7:0] p17_array_index_1079776;
  reg [7:0] p17_array_index_1079777;
  reg [7:0] p17_res7__86;
  reg [7:0] p17_array_index_1079787;
  reg [7:0] p17_array_index_1079788;
  reg [7:0] p17_array_index_1079789;
  reg [7:0] p17_res7__87;
  reg [7:0] p17_array_index_1079800;
  reg [7:0] p17_array_index_1079801;
  reg [7:0] p17_res7__88;
  reg [7:0] p17_array_index_1079811;
  reg [7:0] p17_array_index_1079812;
  reg [7:0] p17_res7__89;
  reg [7:0] p17_array_index_1079818;
  reg [7:0] p17_array_index_1079819;
  reg [7:0] p17_array_index_1079820;
  reg [7:0] p17_array_index_1079821;
  reg [7:0] p17_array_index_1079822;
  reg [7:0] p17_array_index_1079823;
  reg [7:0] p17_array_index_1079824;
  reg [7:0] p17_array_index_1079825;
  reg [7:0] p17_array_index_1079826;
  reg [127:0] p17_res__33;
  reg [7:0] p18_arr[256];
  reg [7:0] p18_literal_1076345[256];
  reg [7:0] p18_literal_1076347[256];
  reg [7:0] p18_literal_1076349[256];
  reg [7:0] p18_literal_1076351[256];
  reg [7:0] p18_literal_1076353[256];
  reg [7:0] p18_literal_1076355[256];
  reg [7:0] p18_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p17_xor_1079057 <= p16_xor_1079057;
    p17_xor_1079529 <= p16_xor_1079529;
    p17_array_index_1079567 <= p16_array_index_1079567;
    p17_array_index_1079568 <= p16_array_index_1079568;
    p17_array_index_1079569 <= p16_array_index_1079569;
    p17_array_index_1079570 <= p16_array_index_1079570;
    p17_array_index_1079571 <= p16_array_index_1079571;
    p17_array_index_1079572 <= p16_array_index_1079572;
    p17_array_index_1079583 <= p16_array_index_1079583;
    p17_array_index_1079584 <= p16_array_index_1079584;
    p17_array_index_1079585 <= p16_array_index_1079585;
    p17_res7__80 <= p16_res7__80;
    p17_array_index_1079600 <= p16_array_index_1079600;
    p17_array_index_1079601 <= p16_array_index_1079601;
    p17_array_index_1079602 <= p16_array_index_1079602;
    p17_res7__81 <= p16_res7__81;
    p17_array_index_1079615 <= p16_array_index_1079615;
    p17_array_index_1079616 <= p16_array_index_1079616;
    p17_array_index_1079617 <= p16_array_index_1079617;
    p17_res7__82 <= p16_res7__82;
    p17_array_index_1079629 <= p16_array_index_1079629;
    p17_array_index_1079630 <= p16_array_index_1079630;
    p17_array_index_1079631 <= p16_array_index_1079631;
    p17_res7__83 <= p16_res7__83;
    p17_array_index_1079644 <= p16_array_index_1079644;
    p17_array_index_1079645 <= p16_array_index_1079645;
    p17_array_index_1079646 <= p16_array_index_1079646;
    p17_res7__84 <= p16_res7__84;
    p17_array_index_1079761 <= p17_array_index_1079761_comb;
    p17_array_index_1079762 <= p17_array_index_1079762_comb;
    p17_array_index_1079763 <= p17_array_index_1079763_comb;
    p17_res7__85 <= p17_res7__85_comb;
    p17_array_index_1079775 <= p17_array_index_1079775_comb;
    p17_array_index_1079776 <= p17_array_index_1079776_comb;
    p17_array_index_1079777 <= p17_array_index_1079777_comb;
    p17_res7__86 <= p17_res7__86_comb;
    p17_array_index_1079787 <= p17_array_index_1079787_comb;
    p17_array_index_1079788 <= p17_array_index_1079788_comb;
    p17_array_index_1079789 <= p17_array_index_1079789_comb;
    p17_res7__87 <= p17_res7__87_comb;
    p17_array_index_1079800 <= p17_array_index_1079800_comb;
    p17_array_index_1079801 <= p17_array_index_1079801_comb;
    p17_res7__88 <= p17_res7__88_comb;
    p17_array_index_1079811 <= p17_array_index_1079811_comb;
    p17_array_index_1079812 <= p17_array_index_1079812_comb;
    p17_res7__89 <= p17_res7__89_comb;
    p17_array_index_1079818 <= p17_array_index_1079818_comb;
    p17_array_index_1079819 <= p17_array_index_1079819_comb;
    p17_array_index_1079820 <= p17_array_index_1079820_comb;
    p17_array_index_1079821 <= p17_array_index_1079821_comb;
    p17_array_index_1079822 <= p17_array_index_1079822_comb;
    p17_array_index_1079823 <= p17_array_index_1079823_comb;
    p17_array_index_1079824 <= p17_array_index_1079824_comb;
    p17_array_index_1079825 <= p17_array_index_1079825_comb;
    p17_array_index_1079826 <= p17_array_index_1079826_comb;
    p17_res__33 <= p16_res__33;
    p18_arr <= p17_arr;
    p18_literal_1076345 <= p17_literal_1076345;
    p18_literal_1076347 <= p17_literal_1076347;
    p18_literal_1076349 <= p17_literal_1076349;
    p18_literal_1076351 <= p17_literal_1076351;
    p18_literal_1076353 <= p17_literal_1076353;
    p18_literal_1076355 <= p17_literal_1076355;
    p18_literal_1076358 <= p17_literal_1076358;
  end

  // ===== Pipe stage 18:
  wire [7:0] p18_res7__90_comb;
  wire [7:0] p18_array_index_1079961_comb;
  wire [7:0] p18_res7__91_comb;
  wire [7:0] p18_res7__92_comb;
  wire [7:0] p18_res7__93_comb;
  wire [7:0] p18_res7__94_comb;
  wire [7:0] p18_res7__95_comb;
  wire [127:0] p18_res__5_comb;
  wire [127:0] p18_xor_1080001_comb;
  assign p18_res7__90_comb = p17_array_index_1079818 ^ p17_array_index_1079819 ^ p17_array_index_1079820 ^ p17_array_index_1079821 ^ p17_array_index_1079822 ^ p17_array_index_1079823 ^ p17_res7__83 ^ p17_array_index_1079824 ^ p17_res7__81 ^ p17_array_index_1079777 ^ p17_array_index_1079646 ^ p17_array_index_1079617 ^ p17_array_index_1079585 ^ p17_array_index_1079825 ^ p17_array_index_1079826 ^ p17_array_index_1079572;
  assign p18_array_index_1079961_comb = p17_literal_1076355[p17_res7__85];
  assign p18_res7__91_comb = p17_literal_1076345[p18_res7__90_comb] ^ p17_literal_1076347[p17_res7__89] ^ p17_literal_1076349[p17_res7__88] ^ p17_literal_1076351[p17_res7__87] ^ p17_literal_1076353[p17_res7__86] ^ p18_array_index_1079961_comb ^ p17_res7__84 ^ p17_literal_1076358[p17_res7__83] ^ p17_res7__82 ^ p17_array_index_1079789 ^ p17_array_index_1079763 ^ p17_array_index_1079631 ^ p17_array_index_1079602 ^ p17_literal_1076347[p17_array_index_1079569] ^ p17_literal_1076345[p17_array_index_1079570] ^ p17_array_index_1079571;
  assign p18_res7__92_comb = p17_literal_1076345[p18_res7__91_comb] ^ p17_literal_1076347[p18_res7__90_comb] ^ p17_literal_1076349[p17_res7__89] ^ p17_literal_1076351[p17_res7__88] ^ p17_literal_1076353[p17_res7__87] ^ p17_literal_1076355[p17_res7__86] ^ p17_res7__85 ^ p17_literal_1076358[p17_res7__84] ^ p17_res7__83 ^ p17_array_index_1079801 ^ p17_array_index_1079776 ^ p17_array_index_1079645 ^ p17_array_index_1079616 ^ p17_array_index_1079584 ^ p17_literal_1076345[p17_array_index_1079569] ^ p17_array_index_1079570;
  assign p18_res7__93_comb = p17_literal_1076345[p18_res7__92_comb] ^ p17_literal_1076347[p18_res7__91_comb] ^ p17_literal_1076349[p18_res7__90_comb] ^ p17_literal_1076351[p17_res7__89] ^ p17_literal_1076353[p17_res7__88] ^ p17_literal_1076355[p17_res7__87] ^ p17_res7__86 ^ p17_literal_1076358[p17_res7__85] ^ p17_res7__84 ^ p17_array_index_1079812 ^ p17_array_index_1079788 ^ p17_array_index_1079762 ^ p17_array_index_1079630 ^ p17_array_index_1079601 ^ p17_literal_1076345[p17_array_index_1079568] ^ p17_array_index_1079569;
  assign p18_res7__94_comb = p17_literal_1076345[p18_res7__93_comb] ^ p17_literal_1076347[p18_res7__92_comb] ^ p17_literal_1076349[p18_res7__91_comb] ^ p17_literal_1076351[p18_res7__90_comb] ^ p17_literal_1076353[p17_res7__89] ^ p17_literal_1076355[p17_res7__88] ^ p17_res7__87 ^ p17_literal_1076358[p17_res7__86] ^ p17_res7__85 ^ p17_array_index_1079823 ^ p17_array_index_1079800 ^ p17_array_index_1079775 ^ p17_array_index_1079644 ^ p17_array_index_1079615 ^ p17_array_index_1079583 ^ p17_array_index_1079568;
  assign p18_res7__95_comb = p17_literal_1076345[p18_res7__94_comb] ^ p17_literal_1076347[p18_res7__93_comb] ^ p17_literal_1076349[p18_res7__92_comb] ^ p17_literal_1076351[p18_res7__91_comb] ^ p17_literal_1076353[p18_res7__90_comb] ^ p17_literal_1076355[p17_res7__89] ^ p17_res7__88 ^ p17_literal_1076358[p17_res7__87] ^ p17_res7__86 ^ p18_array_index_1079961_comb ^ p17_array_index_1079811 ^ p17_array_index_1079787 ^ p17_array_index_1079761 ^ p17_array_index_1079629 ^ p17_array_index_1079600 ^ p17_array_index_1079567;
  assign p18_res__5_comb = {p18_res7__95_comb, p18_res7__94_comb, p18_res7__93_comb, p18_res7__92_comb, p18_res7__91_comb, p18_res7__90_comb, p17_res7__89, p17_res7__88, p17_res7__87, p17_res7__86, p17_res7__85, p17_res7__84, p17_res7__83, p17_res7__82, p17_res7__81, p17_res7__80};
  assign p18_xor_1080001_comb = p18_res__5_comb ^ p17_xor_1079057;

  // Registers for pipe stage 18:
  reg [127:0] p18_xor_1079529;
  reg [127:0] p18_xor_1080001;
  reg [127:0] p18_res__33;
  reg [7:0] p19_arr[256];
  reg [7:0] p19_literal_1076345[256];
  reg [7:0] p19_literal_1076347[256];
  reg [7:0] p19_literal_1076349[256];
  reg [7:0] p19_literal_1076351[256];
  reg [7:0] p19_literal_1076353[256];
  reg [7:0] p19_literal_1076355[256];
  reg [7:0] p19_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p18_xor_1079529 <= p17_xor_1079529;
    p18_xor_1080001 <= p18_xor_1080001_comb;
    p18_res__33 <= p17_res__33;
    p19_arr <= p18_arr;
    p19_literal_1076345 <= p18_literal_1076345;
    p19_literal_1076347 <= p18_literal_1076347;
    p19_literal_1076349 <= p18_literal_1076349;
    p19_literal_1076351 <= p18_literal_1076351;
    p19_literal_1076353 <= p18_literal_1076353;
    p19_literal_1076355 <= p18_literal_1076355;
    p19_literal_1076358 <= p18_literal_1076358;
  end

  // ===== Pipe stage 19:
  wire [127:0] p19_addedKey__47_comb;
  wire [7:0] p19_array_index_1080039_comb;
  wire [7:0] p19_array_index_1080040_comb;
  wire [7:0] p19_array_index_1080041_comb;
  wire [7:0] p19_array_index_1080042_comb;
  wire [7:0] p19_array_index_1080043_comb;
  wire [7:0] p19_array_index_1080044_comb;
  wire [7:0] p19_array_index_1080046_comb;
  wire [7:0] p19_array_index_1080048_comb;
  wire [7:0] p19_array_index_1080049_comb;
  wire [7:0] p19_array_index_1080050_comb;
  wire [7:0] p19_array_index_1080051_comb;
  wire [7:0] p19_array_index_1080052_comb;
  wire [7:0] p19_array_index_1080053_comb;
  wire [7:0] p19_array_index_1080055_comb;
  wire [7:0] p19_array_index_1080056_comb;
  wire [7:0] p19_array_index_1080057_comb;
  wire [7:0] p19_array_index_1080058_comb;
  wire [7:0] p19_array_index_1080059_comb;
  wire [7:0] p19_array_index_1080060_comb;
  wire [7:0] p19_array_index_1080061_comb;
  wire [7:0] p19_array_index_1080063_comb;
  wire [7:0] p19_res7__96_comb;
  wire [7:0] p19_array_index_1080072_comb;
  wire [7:0] p19_array_index_1080073_comb;
  wire [7:0] p19_array_index_1080074_comb;
  wire [7:0] p19_array_index_1080075_comb;
  wire [7:0] p19_array_index_1080076_comb;
  wire [7:0] p19_array_index_1080077_comb;
  wire [7:0] p19_res7__97_comb;
  wire [7:0] p19_array_index_1080087_comb;
  wire [7:0] p19_array_index_1080088_comb;
  wire [7:0] p19_array_index_1080089_comb;
  wire [7:0] p19_array_index_1080090_comb;
  wire [7:0] p19_array_index_1080091_comb;
  wire [7:0] p19_res7__98_comb;
  wire [7:0] p19_array_index_1080101_comb;
  wire [7:0] p19_array_index_1080102_comb;
  wire [7:0] p19_array_index_1080103_comb;
  wire [7:0] p19_array_index_1080104_comb;
  wire [7:0] p19_array_index_1080105_comb;
  wire [7:0] p19_res7__99_comb;
  wire [7:0] p19_array_index_1080116_comb;
  wire [7:0] p19_array_index_1080117_comb;
  wire [7:0] p19_array_index_1080118_comb;
  wire [7:0] p19_array_index_1080119_comb;
  wire [7:0] p19_res7__100_comb;
  assign p19_addedKey__47_comb = p18_xor_1080001 ^ 128'hc9e8_819d_c73b_a5ae_50f5_b570_561a_6a07;
  assign p19_array_index_1080039_comb = p18_arr[p19_addedKey__47_comb[127:120]];
  assign p19_array_index_1080040_comb = p18_arr[p19_addedKey__47_comb[119:112]];
  assign p19_array_index_1080041_comb = p18_arr[p19_addedKey__47_comb[111:104]];
  assign p19_array_index_1080042_comb = p18_arr[p19_addedKey__47_comb[103:96]];
  assign p19_array_index_1080043_comb = p18_arr[p19_addedKey__47_comb[95:88]];
  assign p19_array_index_1080044_comb = p18_arr[p19_addedKey__47_comb[87:80]];
  assign p19_array_index_1080046_comb = p18_arr[p19_addedKey__47_comb[71:64]];
  assign p19_array_index_1080048_comb = p18_arr[p19_addedKey__47_comb[55:48]];
  assign p19_array_index_1080049_comb = p18_arr[p19_addedKey__47_comb[47:40]];
  assign p19_array_index_1080050_comb = p18_arr[p19_addedKey__47_comb[39:32]];
  assign p19_array_index_1080051_comb = p18_arr[p19_addedKey__47_comb[31:24]];
  assign p19_array_index_1080052_comb = p18_arr[p19_addedKey__47_comb[23:16]];
  assign p19_array_index_1080053_comb = p18_arr[p19_addedKey__47_comb[15:8]];
  assign p19_array_index_1080055_comb = p18_literal_1076345[p19_array_index_1080039_comb];
  assign p19_array_index_1080056_comb = p18_literal_1076347[p19_array_index_1080040_comb];
  assign p19_array_index_1080057_comb = p18_literal_1076349[p19_array_index_1080041_comb];
  assign p19_array_index_1080058_comb = p18_literal_1076351[p19_array_index_1080042_comb];
  assign p19_array_index_1080059_comb = p18_literal_1076353[p19_array_index_1080043_comb];
  assign p19_array_index_1080060_comb = p18_literal_1076355[p19_array_index_1080044_comb];
  assign p19_array_index_1080061_comb = p18_arr[p19_addedKey__47_comb[79:72]];
  assign p19_array_index_1080063_comb = p18_arr[p19_addedKey__47_comb[63:56]];
  assign p19_res7__96_comb = p19_array_index_1080055_comb ^ p19_array_index_1080056_comb ^ p19_array_index_1080057_comb ^ p19_array_index_1080058_comb ^ p19_array_index_1080059_comb ^ p19_array_index_1080060_comb ^ p19_array_index_1080061_comb ^ p18_literal_1076358[p19_array_index_1080046_comb] ^ p19_array_index_1080063_comb ^ p18_literal_1076355[p19_array_index_1080048_comb] ^ p18_literal_1076353[p19_array_index_1080049_comb] ^ p18_literal_1076351[p19_array_index_1080050_comb] ^ p18_literal_1076349[p19_array_index_1080051_comb] ^ p18_literal_1076347[p19_array_index_1080052_comb] ^ p18_literal_1076345[p19_array_index_1080053_comb] ^ p18_arr[p19_addedKey__47_comb[7:0]];
  assign p19_array_index_1080072_comb = p18_literal_1076345[p19_res7__96_comb];
  assign p19_array_index_1080073_comb = p18_literal_1076347[p19_array_index_1080039_comb];
  assign p19_array_index_1080074_comb = p18_literal_1076349[p19_array_index_1080040_comb];
  assign p19_array_index_1080075_comb = p18_literal_1076351[p19_array_index_1080041_comb];
  assign p19_array_index_1080076_comb = p18_literal_1076353[p19_array_index_1080042_comb];
  assign p19_array_index_1080077_comb = p18_literal_1076355[p19_array_index_1080043_comb];
  assign p19_res7__97_comb = p19_array_index_1080072_comb ^ p19_array_index_1080073_comb ^ p19_array_index_1080074_comb ^ p19_array_index_1080075_comb ^ p19_array_index_1080076_comb ^ p19_array_index_1080077_comb ^ p19_array_index_1080044_comb ^ p18_literal_1076358[p19_array_index_1080061_comb] ^ p19_array_index_1080046_comb ^ p18_literal_1076355[p19_array_index_1080063_comb] ^ p18_literal_1076353[p19_array_index_1080048_comb] ^ p18_literal_1076351[p19_array_index_1080049_comb] ^ p18_literal_1076349[p19_array_index_1080050_comb] ^ p18_literal_1076347[p19_array_index_1080051_comb] ^ p18_literal_1076345[p19_array_index_1080052_comb] ^ p19_array_index_1080053_comb;
  assign p19_array_index_1080087_comb = p18_literal_1076347[p19_res7__96_comb];
  assign p19_array_index_1080088_comb = p18_literal_1076349[p19_array_index_1080039_comb];
  assign p19_array_index_1080089_comb = p18_literal_1076351[p19_array_index_1080040_comb];
  assign p19_array_index_1080090_comb = p18_literal_1076353[p19_array_index_1080041_comb];
  assign p19_array_index_1080091_comb = p18_literal_1076355[p19_array_index_1080042_comb];
  assign p19_res7__98_comb = p18_literal_1076345[p19_res7__97_comb] ^ p19_array_index_1080087_comb ^ p19_array_index_1080088_comb ^ p19_array_index_1080089_comb ^ p19_array_index_1080090_comb ^ p19_array_index_1080091_comb ^ p19_array_index_1080043_comb ^ p18_literal_1076358[p19_array_index_1080044_comb] ^ p19_array_index_1080061_comb ^ p18_literal_1076355[p19_array_index_1080046_comb] ^ p18_literal_1076353[p19_array_index_1080063_comb] ^ p18_literal_1076351[p19_array_index_1080048_comb] ^ p18_literal_1076349[p19_array_index_1080049_comb] ^ p18_literal_1076347[p19_array_index_1080050_comb] ^ p18_literal_1076345[p19_array_index_1080051_comb] ^ p19_array_index_1080052_comb;
  assign p19_array_index_1080101_comb = p18_literal_1076347[p19_res7__97_comb];
  assign p19_array_index_1080102_comb = p18_literal_1076349[p19_res7__96_comb];
  assign p19_array_index_1080103_comb = p18_literal_1076351[p19_array_index_1080039_comb];
  assign p19_array_index_1080104_comb = p18_literal_1076353[p19_array_index_1080040_comb];
  assign p19_array_index_1080105_comb = p18_literal_1076355[p19_array_index_1080041_comb];
  assign p19_res7__99_comb = p18_literal_1076345[p19_res7__98_comb] ^ p19_array_index_1080101_comb ^ p19_array_index_1080102_comb ^ p19_array_index_1080103_comb ^ p19_array_index_1080104_comb ^ p19_array_index_1080105_comb ^ p19_array_index_1080042_comb ^ p18_literal_1076358[p19_array_index_1080043_comb] ^ p19_array_index_1080044_comb ^ p18_literal_1076355[p19_array_index_1080061_comb] ^ p18_literal_1076353[p19_array_index_1080046_comb] ^ p18_literal_1076351[p19_array_index_1080063_comb] ^ p18_literal_1076349[p19_array_index_1080048_comb] ^ p18_literal_1076347[p19_array_index_1080049_comb] ^ p18_literal_1076345[p19_array_index_1080050_comb] ^ p19_array_index_1080051_comb;
  assign p19_array_index_1080116_comb = p18_literal_1076349[p19_res7__97_comb];
  assign p19_array_index_1080117_comb = p18_literal_1076351[p19_res7__96_comb];
  assign p19_array_index_1080118_comb = p18_literal_1076353[p19_array_index_1080039_comb];
  assign p19_array_index_1080119_comb = p18_literal_1076355[p19_array_index_1080040_comb];
  assign p19_res7__100_comb = p18_literal_1076345[p19_res7__99_comb] ^ p18_literal_1076347[p19_res7__98_comb] ^ p19_array_index_1080116_comb ^ p19_array_index_1080117_comb ^ p19_array_index_1080118_comb ^ p19_array_index_1080119_comb ^ p19_array_index_1080041_comb ^ p18_literal_1076358[p19_array_index_1080042_comb] ^ p19_array_index_1080043_comb ^ p19_array_index_1080060_comb ^ p18_literal_1076353[p19_array_index_1080061_comb] ^ p18_literal_1076351[p19_array_index_1080046_comb] ^ p18_literal_1076349[p19_array_index_1080063_comb] ^ p18_literal_1076347[p19_array_index_1080048_comb] ^ p18_literal_1076345[p19_array_index_1080049_comb] ^ p19_array_index_1080050_comb;

  // Registers for pipe stage 19:
  reg [127:0] p19_xor_1079529;
  reg [127:0] p19_xor_1080001;
  reg [7:0] p19_array_index_1080039;
  reg [7:0] p19_array_index_1080040;
  reg [7:0] p19_array_index_1080041;
  reg [7:0] p19_array_index_1080042;
  reg [7:0] p19_array_index_1080043;
  reg [7:0] p19_array_index_1080044;
  reg [7:0] p19_array_index_1080046;
  reg [7:0] p19_array_index_1080048;
  reg [7:0] p19_array_index_1080049;
  reg [7:0] p19_array_index_1080055;
  reg [7:0] p19_array_index_1080056;
  reg [7:0] p19_array_index_1080057;
  reg [7:0] p19_array_index_1080058;
  reg [7:0] p19_array_index_1080059;
  reg [7:0] p19_array_index_1080061;
  reg [7:0] p19_array_index_1080063;
  reg [7:0] p19_res7__96;
  reg [7:0] p19_array_index_1080072;
  reg [7:0] p19_array_index_1080073;
  reg [7:0] p19_array_index_1080074;
  reg [7:0] p19_array_index_1080075;
  reg [7:0] p19_array_index_1080076;
  reg [7:0] p19_array_index_1080077;
  reg [7:0] p19_res7__97;
  reg [7:0] p19_array_index_1080087;
  reg [7:0] p19_array_index_1080088;
  reg [7:0] p19_array_index_1080089;
  reg [7:0] p19_array_index_1080090;
  reg [7:0] p19_array_index_1080091;
  reg [7:0] p19_res7__98;
  reg [7:0] p19_array_index_1080101;
  reg [7:0] p19_array_index_1080102;
  reg [7:0] p19_array_index_1080103;
  reg [7:0] p19_array_index_1080104;
  reg [7:0] p19_array_index_1080105;
  reg [7:0] p19_res7__99;
  reg [7:0] p19_array_index_1080116;
  reg [7:0] p19_array_index_1080117;
  reg [7:0] p19_array_index_1080118;
  reg [7:0] p19_array_index_1080119;
  reg [7:0] p19_res7__100;
  reg [127:0] p19_res__33;
  reg [7:0] p20_arr[256];
  reg [7:0] p20_literal_1076345[256];
  reg [7:0] p20_literal_1076347[256];
  reg [7:0] p20_literal_1076349[256];
  reg [7:0] p20_literal_1076351[256];
  reg [7:0] p20_literal_1076353[256];
  reg [7:0] p20_literal_1076355[256];
  reg [7:0] p20_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p19_xor_1079529 <= p18_xor_1079529;
    p19_xor_1080001 <= p18_xor_1080001;
    p19_array_index_1080039 <= p19_array_index_1080039_comb;
    p19_array_index_1080040 <= p19_array_index_1080040_comb;
    p19_array_index_1080041 <= p19_array_index_1080041_comb;
    p19_array_index_1080042 <= p19_array_index_1080042_comb;
    p19_array_index_1080043 <= p19_array_index_1080043_comb;
    p19_array_index_1080044 <= p19_array_index_1080044_comb;
    p19_array_index_1080046 <= p19_array_index_1080046_comb;
    p19_array_index_1080048 <= p19_array_index_1080048_comb;
    p19_array_index_1080049 <= p19_array_index_1080049_comb;
    p19_array_index_1080055 <= p19_array_index_1080055_comb;
    p19_array_index_1080056 <= p19_array_index_1080056_comb;
    p19_array_index_1080057 <= p19_array_index_1080057_comb;
    p19_array_index_1080058 <= p19_array_index_1080058_comb;
    p19_array_index_1080059 <= p19_array_index_1080059_comb;
    p19_array_index_1080061 <= p19_array_index_1080061_comb;
    p19_array_index_1080063 <= p19_array_index_1080063_comb;
    p19_res7__96 <= p19_res7__96_comb;
    p19_array_index_1080072 <= p19_array_index_1080072_comb;
    p19_array_index_1080073 <= p19_array_index_1080073_comb;
    p19_array_index_1080074 <= p19_array_index_1080074_comb;
    p19_array_index_1080075 <= p19_array_index_1080075_comb;
    p19_array_index_1080076 <= p19_array_index_1080076_comb;
    p19_array_index_1080077 <= p19_array_index_1080077_comb;
    p19_res7__97 <= p19_res7__97_comb;
    p19_array_index_1080087 <= p19_array_index_1080087_comb;
    p19_array_index_1080088 <= p19_array_index_1080088_comb;
    p19_array_index_1080089 <= p19_array_index_1080089_comb;
    p19_array_index_1080090 <= p19_array_index_1080090_comb;
    p19_array_index_1080091 <= p19_array_index_1080091_comb;
    p19_res7__98 <= p19_res7__98_comb;
    p19_array_index_1080101 <= p19_array_index_1080101_comb;
    p19_array_index_1080102 <= p19_array_index_1080102_comb;
    p19_array_index_1080103 <= p19_array_index_1080103_comb;
    p19_array_index_1080104 <= p19_array_index_1080104_comb;
    p19_array_index_1080105 <= p19_array_index_1080105_comb;
    p19_res7__99 <= p19_res7__99_comb;
    p19_array_index_1080116 <= p19_array_index_1080116_comb;
    p19_array_index_1080117 <= p19_array_index_1080117_comb;
    p19_array_index_1080118 <= p19_array_index_1080118_comb;
    p19_array_index_1080119 <= p19_array_index_1080119_comb;
    p19_res7__100 <= p19_res7__100_comb;
    p19_res__33 <= p18_res__33;
    p20_arr <= p19_arr;
    p20_literal_1076345 <= p19_literal_1076345;
    p20_literal_1076347 <= p19_literal_1076347;
    p20_literal_1076349 <= p19_literal_1076349;
    p20_literal_1076351 <= p19_literal_1076351;
    p20_literal_1076353 <= p19_literal_1076353;
    p20_literal_1076355 <= p19_literal_1076355;
    p20_literal_1076358 <= p19_literal_1076358;
  end

  // ===== Pipe stage 20:
  wire [7:0] p20_array_index_1080233_comb;
  wire [7:0] p20_array_index_1080234_comb;
  wire [7:0] p20_array_index_1080235_comb;
  wire [7:0] p20_array_index_1080236_comb;
  wire [7:0] p20_res7__101_comb;
  wire [7:0] p20_array_index_1080247_comb;
  wire [7:0] p20_array_index_1080248_comb;
  wire [7:0] p20_array_index_1080249_comb;
  wire [7:0] p20_res7__102_comb;
  wire [7:0] p20_array_index_1080259_comb;
  wire [7:0] p20_array_index_1080260_comb;
  wire [7:0] p20_array_index_1080261_comb;
  wire [7:0] p20_res7__103_comb;
  wire [7:0] p20_array_index_1080272_comb;
  wire [7:0] p20_array_index_1080273_comb;
  wire [7:0] p20_res7__104_comb;
  wire [7:0] p20_array_index_1080283_comb;
  wire [7:0] p20_array_index_1080284_comb;
  wire [7:0] p20_res7__105_comb;
  wire [7:0] p20_array_index_1080290_comb;
  wire [7:0] p20_array_index_1080291_comb;
  wire [7:0] p20_array_index_1080292_comb;
  wire [7:0] p20_array_index_1080293_comb;
  wire [7:0] p20_array_index_1080294_comb;
  wire [7:0] p20_array_index_1080295_comb;
  wire [7:0] p20_array_index_1080296_comb;
  wire [7:0] p20_array_index_1080297_comb;
  wire [7:0] p20_array_index_1080298_comb;
  assign p20_array_index_1080233_comb = p19_literal_1076349[p19_res7__98];
  assign p20_array_index_1080234_comb = p19_literal_1076351[p19_res7__97];
  assign p20_array_index_1080235_comb = p19_literal_1076353[p19_res7__96];
  assign p20_array_index_1080236_comb = p19_literal_1076355[p19_array_index_1080039];
  assign p20_res7__101_comb = p19_literal_1076345[p19_res7__100] ^ p19_literal_1076347[p19_res7__99] ^ p20_array_index_1080233_comb ^ p20_array_index_1080234_comb ^ p20_array_index_1080235_comb ^ p20_array_index_1080236_comb ^ p19_array_index_1080040 ^ p19_literal_1076358[p19_array_index_1080041] ^ p19_array_index_1080042 ^ p19_array_index_1080077 ^ p19_literal_1076353[p19_array_index_1080044] ^ p19_literal_1076351[p19_array_index_1080061] ^ p19_literal_1076349[p19_array_index_1080046] ^ p19_literal_1076347[p19_array_index_1080063] ^ p19_literal_1076345[p19_array_index_1080048] ^ p19_array_index_1080049;
  assign p20_array_index_1080247_comb = p19_literal_1076351[p19_res7__98];
  assign p20_array_index_1080248_comb = p19_literal_1076353[p19_res7__97];
  assign p20_array_index_1080249_comb = p19_literal_1076355[p19_res7__96];
  assign p20_res7__102_comb = p19_literal_1076345[p20_res7__101_comb] ^ p19_literal_1076347[p19_res7__100] ^ p19_literal_1076349[p19_res7__99] ^ p20_array_index_1080247_comb ^ p20_array_index_1080248_comb ^ p20_array_index_1080249_comb ^ p19_array_index_1080039 ^ p19_literal_1076358[p19_array_index_1080040] ^ p19_array_index_1080041 ^ p19_array_index_1080091 ^ p19_array_index_1080059 ^ p19_literal_1076351[p19_array_index_1080044] ^ p19_literal_1076349[p19_array_index_1080061] ^ p19_literal_1076347[p19_array_index_1080046] ^ p19_literal_1076345[p19_array_index_1080063] ^ p19_array_index_1080048;
  assign p20_array_index_1080259_comb = p19_literal_1076351[p19_res7__99];
  assign p20_array_index_1080260_comb = p19_literal_1076353[p19_res7__98];
  assign p20_array_index_1080261_comb = p19_literal_1076355[p19_res7__97];
  assign p20_res7__103_comb = p19_literal_1076345[p20_res7__102_comb] ^ p19_literal_1076347[p20_res7__101_comb] ^ p19_literal_1076349[p19_res7__100] ^ p20_array_index_1080259_comb ^ p20_array_index_1080260_comb ^ p20_array_index_1080261_comb ^ p19_res7__96 ^ p19_literal_1076358[p19_array_index_1080039] ^ p19_array_index_1080040 ^ p19_array_index_1080105 ^ p19_array_index_1080076 ^ p19_literal_1076351[p19_array_index_1080043] ^ p19_literal_1076349[p19_array_index_1080044] ^ p19_literal_1076347[p19_array_index_1080061] ^ p19_literal_1076345[p19_array_index_1080046] ^ p19_array_index_1080063;
  assign p20_array_index_1080272_comb = p19_literal_1076353[p19_res7__99];
  assign p20_array_index_1080273_comb = p19_literal_1076355[p19_res7__98];
  assign p20_res7__104_comb = p19_literal_1076345[p20_res7__103_comb] ^ p19_literal_1076347[p20_res7__102_comb] ^ p19_literal_1076349[p20_res7__101_comb] ^ p19_literal_1076351[p19_res7__100] ^ p20_array_index_1080272_comb ^ p20_array_index_1080273_comb ^ p19_res7__97 ^ p19_literal_1076358[p19_res7__96] ^ p19_array_index_1080039 ^ p19_array_index_1080119 ^ p19_array_index_1080090 ^ p19_array_index_1080058 ^ p19_literal_1076349[p19_array_index_1080043] ^ p19_literal_1076347[p19_array_index_1080044] ^ p19_literal_1076345[p19_array_index_1080061] ^ p19_array_index_1080046;
  assign p20_array_index_1080283_comb = p19_literal_1076353[p19_res7__100];
  assign p20_array_index_1080284_comb = p19_literal_1076355[p19_res7__99];
  assign p20_res7__105_comb = p19_literal_1076345[p20_res7__104_comb] ^ p19_literal_1076347[p20_res7__103_comb] ^ p19_literal_1076349[p20_res7__102_comb] ^ p19_literal_1076351[p20_res7__101_comb] ^ p20_array_index_1080283_comb ^ p20_array_index_1080284_comb ^ p19_res7__98 ^ p19_literal_1076358[p19_res7__97] ^ p19_res7__96 ^ p20_array_index_1080236_comb ^ p19_array_index_1080104 ^ p19_array_index_1080075 ^ p19_literal_1076349[p19_array_index_1080042] ^ p19_literal_1076347[p19_array_index_1080043] ^ p19_literal_1076345[p19_array_index_1080044] ^ p19_array_index_1080061;
  assign p20_array_index_1080290_comb = p19_literal_1076345[p20_res7__105_comb];
  assign p20_array_index_1080291_comb = p19_literal_1076347[p20_res7__104_comb];
  assign p20_array_index_1080292_comb = p19_literal_1076349[p20_res7__103_comb];
  assign p20_array_index_1080293_comb = p19_literal_1076351[p20_res7__102_comb];
  assign p20_array_index_1080294_comb = p19_literal_1076353[p20_res7__101_comb];
  assign p20_array_index_1080295_comb = p19_literal_1076355[p19_res7__100];
  assign p20_array_index_1080296_comb = p19_literal_1076358[p19_res7__98];
  assign p20_array_index_1080297_comb = p19_literal_1076347[p19_array_index_1080042];
  assign p20_array_index_1080298_comb = p19_literal_1076345[p19_array_index_1080043];

  // Registers for pipe stage 20:
  reg [127:0] p20_xor_1079529;
  reg [127:0] p20_xor_1080001;
  reg [7:0] p20_array_index_1080039;
  reg [7:0] p20_array_index_1080040;
  reg [7:0] p20_array_index_1080041;
  reg [7:0] p20_array_index_1080042;
  reg [7:0] p20_array_index_1080043;
  reg [7:0] p20_array_index_1080044;
  reg [7:0] p20_array_index_1080055;
  reg [7:0] p20_array_index_1080056;
  reg [7:0] p20_array_index_1080057;
  reg [7:0] p20_res7__96;
  reg [7:0] p20_array_index_1080072;
  reg [7:0] p20_array_index_1080073;
  reg [7:0] p20_array_index_1080074;
  reg [7:0] p20_res7__97;
  reg [7:0] p20_array_index_1080087;
  reg [7:0] p20_array_index_1080088;
  reg [7:0] p20_array_index_1080089;
  reg [7:0] p20_res7__98;
  reg [7:0] p20_array_index_1080101;
  reg [7:0] p20_array_index_1080102;
  reg [7:0] p20_array_index_1080103;
  reg [7:0] p20_res7__99;
  reg [7:0] p20_array_index_1080116;
  reg [7:0] p20_array_index_1080117;
  reg [7:0] p20_array_index_1080118;
  reg [7:0] p20_res7__100;
  reg [7:0] p20_array_index_1080233;
  reg [7:0] p20_array_index_1080234;
  reg [7:0] p20_array_index_1080235;
  reg [7:0] p20_res7__101;
  reg [7:0] p20_array_index_1080247;
  reg [7:0] p20_array_index_1080248;
  reg [7:0] p20_array_index_1080249;
  reg [7:0] p20_res7__102;
  reg [7:0] p20_array_index_1080259;
  reg [7:0] p20_array_index_1080260;
  reg [7:0] p20_array_index_1080261;
  reg [7:0] p20_res7__103;
  reg [7:0] p20_array_index_1080272;
  reg [7:0] p20_array_index_1080273;
  reg [7:0] p20_res7__104;
  reg [7:0] p20_array_index_1080283;
  reg [7:0] p20_array_index_1080284;
  reg [7:0] p20_res7__105;
  reg [7:0] p20_array_index_1080290;
  reg [7:0] p20_array_index_1080291;
  reg [7:0] p20_array_index_1080292;
  reg [7:0] p20_array_index_1080293;
  reg [7:0] p20_array_index_1080294;
  reg [7:0] p20_array_index_1080295;
  reg [7:0] p20_array_index_1080296;
  reg [7:0] p20_array_index_1080297;
  reg [7:0] p20_array_index_1080298;
  reg [127:0] p20_res__33;
  reg [7:0] p21_arr[256];
  reg [7:0] p21_literal_1076345[256];
  reg [7:0] p21_literal_1076347[256];
  reg [7:0] p21_literal_1076349[256];
  reg [7:0] p21_literal_1076351[256];
  reg [7:0] p21_literal_1076353[256];
  reg [7:0] p21_literal_1076355[256];
  reg [7:0] p21_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p20_xor_1079529 <= p19_xor_1079529;
    p20_xor_1080001 <= p19_xor_1080001;
    p20_array_index_1080039 <= p19_array_index_1080039;
    p20_array_index_1080040 <= p19_array_index_1080040;
    p20_array_index_1080041 <= p19_array_index_1080041;
    p20_array_index_1080042 <= p19_array_index_1080042;
    p20_array_index_1080043 <= p19_array_index_1080043;
    p20_array_index_1080044 <= p19_array_index_1080044;
    p20_array_index_1080055 <= p19_array_index_1080055;
    p20_array_index_1080056 <= p19_array_index_1080056;
    p20_array_index_1080057 <= p19_array_index_1080057;
    p20_res7__96 <= p19_res7__96;
    p20_array_index_1080072 <= p19_array_index_1080072;
    p20_array_index_1080073 <= p19_array_index_1080073;
    p20_array_index_1080074 <= p19_array_index_1080074;
    p20_res7__97 <= p19_res7__97;
    p20_array_index_1080087 <= p19_array_index_1080087;
    p20_array_index_1080088 <= p19_array_index_1080088;
    p20_array_index_1080089 <= p19_array_index_1080089;
    p20_res7__98 <= p19_res7__98;
    p20_array_index_1080101 <= p19_array_index_1080101;
    p20_array_index_1080102 <= p19_array_index_1080102;
    p20_array_index_1080103 <= p19_array_index_1080103;
    p20_res7__99 <= p19_res7__99;
    p20_array_index_1080116 <= p19_array_index_1080116;
    p20_array_index_1080117 <= p19_array_index_1080117;
    p20_array_index_1080118 <= p19_array_index_1080118;
    p20_res7__100 <= p19_res7__100;
    p20_array_index_1080233 <= p20_array_index_1080233_comb;
    p20_array_index_1080234 <= p20_array_index_1080234_comb;
    p20_array_index_1080235 <= p20_array_index_1080235_comb;
    p20_res7__101 <= p20_res7__101_comb;
    p20_array_index_1080247 <= p20_array_index_1080247_comb;
    p20_array_index_1080248 <= p20_array_index_1080248_comb;
    p20_array_index_1080249 <= p20_array_index_1080249_comb;
    p20_res7__102 <= p20_res7__102_comb;
    p20_array_index_1080259 <= p20_array_index_1080259_comb;
    p20_array_index_1080260 <= p20_array_index_1080260_comb;
    p20_array_index_1080261 <= p20_array_index_1080261_comb;
    p20_res7__103 <= p20_res7__103_comb;
    p20_array_index_1080272 <= p20_array_index_1080272_comb;
    p20_array_index_1080273 <= p20_array_index_1080273_comb;
    p20_res7__104 <= p20_res7__104_comb;
    p20_array_index_1080283 <= p20_array_index_1080283_comb;
    p20_array_index_1080284 <= p20_array_index_1080284_comb;
    p20_res7__105 <= p20_res7__105_comb;
    p20_array_index_1080290 <= p20_array_index_1080290_comb;
    p20_array_index_1080291 <= p20_array_index_1080291_comb;
    p20_array_index_1080292 <= p20_array_index_1080292_comb;
    p20_array_index_1080293 <= p20_array_index_1080293_comb;
    p20_array_index_1080294 <= p20_array_index_1080294_comb;
    p20_array_index_1080295 <= p20_array_index_1080295_comb;
    p20_array_index_1080296 <= p20_array_index_1080296_comb;
    p20_array_index_1080297 <= p20_array_index_1080297_comb;
    p20_array_index_1080298 <= p20_array_index_1080298_comb;
    p20_res__33 <= p19_res__33;
    p21_arr <= p20_arr;
    p21_literal_1076345 <= p20_literal_1076345;
    p21_literal_1076347 <= p20_literal_1076347;
    p21_literal_1076349 <= p20_literal_1076349;
    p21_literal_1076351 <= p20_literal_1076351;
    p21_literal_1076353 <= p20_literal_1076353;
    p21_literal_1076355 <= p20_literal_1076355;
    p21_literal_1076358 <= p20_literal_1076358;
  end

  // ===== Pipe stage 21:
  wire [7:0] p21_res7__106_comb;
  wire [7:0] p21_array_index_1080433_comb;
  wire [7:0] p21_res7__107_comb;
  wire [7:0] p21_res7__108_comb;
  wire [7:0] p21_res7__109_comb;
  wire [7:0] p21_res7__110_comb;
  wire [7:0] p21_res7__111_comb;
  wire [127:0] p21_res__6_comb;
  wire [127:0] p21_k3_comb;
  assign p21_res7__106_comb = p20_array_index_1080290 ^ p20_array_index_1080291 ^ p20_array_index_1080292 ^ p20_array_index_1080293 ^ p20_array_index_1080294 ^ p20_array_index_1080295 ^ p20_res7__99 ^ p20_array_index_1080296 ^ p20_res7__97 ^ p20_array_index_1080249 ^ p20_array_index_1080118 ^ p20_array_index_1080089 ^ p20_array_index_1080057 ^ p20_array_index_1080297 ^ p20_array_index_1080298 ^ p20_array_index_1080044;
  assign p21_array_index_1080433_comb = p20_literal_1076355[p20_res7__101];
  assign p21_res7__107_comb = p20_literal_1076345[p21_res7__106_comb] ^ p20_literal_1076347[p20_res7__105] ^ p20_literal_1076349[p20_res7__104] ^ p20_literal_1076351[p20_res7__103] ^ p20_literal_1076353[p20_res7__102] ^ p21_array_index_1080433_comb ^ p20_res7__100 ^ p20_literal_1076358[p20_res7__99] ^ p20_res7__98 ^ p20_array_index_1080261 ^ p20_array_index_1080235 ^ p20_array_index_1080103 ^ p20_array_index_1080074 ^ p20_literal_1076347[p20_array_index_1080041] ^ p20_literal_1076345[p20_array_index_1080042] ^ p20_array_index_1080043;
  assign p21_res7__108_comb = p20_literal_1076345[p21_res7__107_comb] ^ p20_literal_1076347[p21_res7__106_comb] ^ p20_literal_1076349[p20_res7__105] ^ p20_literal_1076351[p20_res7__104] ^ p20_literal_1076353[p20_res7__103] ^ p20_literal_1076355[p20_res7__102] ^ p20_res7__101 ^ p20_literal_1076358[p20_res7__100] ^ p20_res7__99 ^ p20_array_index_1080273 ^ p20_array_index_1080248 ^ p20_array_index_1080117 ^ p20_array_index_1080088 ^ p20_array_index_1080056 ^ p20_literal_1076345[p20_array_index_1080041] ^ p20_array_index_1080042;
  assign p21_res7__109_comb = p20_literal_1076345[p21_res7__108_comb] ^ p20_literal_1076347[p21_res7__107_comb] ^ p20_literal_1076349[p21_res7__106_comb] ^ p20_literal_1076351[p20_res7__105] ^ p20_literal_1076353[p20_res7__104] ^ p20_literal_1076355[p20_res7__103] ^ p20_res7__102 ^ p20_literal_1076358[p20_res7__101] ^ p20_res7__100 ^ p20_array_index_1080284 ^ p20_array_index_1080260 ^ p20_array_index_1080234 ^ p20_array_index_1080102 ^ p20_array_index_1080073 ^ p20_literal_1076345[p20_array_index_1080040] ^ p20_array_index_1080041;
  assign p21_res7__110_comb = p20_literal_1076345[p21_res7__109_comb] ^ p20_literal_1076347[p21_res7__108_comb] ^ p20_literal_1076349[p21_res7__107_comb] ^ p20_literal_1076351[p21_res7__106_comb] ^ p20_literal_1076353[p20_res7__105] ^ p20_literal_1076355[p20_res7__104] ^ p20_res7__103 ^ p20_literal_1076358[p20_res7__102] ^ p20_res7__101 ^ p20_array_index_1080295 ^ p20_array_index_1080272 ^ p20_array_index_1080247 ^ p20_array_index_1080116 ^ p20_array_index_1080087 ^ p20_array_index_1080055 ^ p20_array_index_1080040;
  assign p21_res7__111_comb = p20_literal_1076345[p21_res7__110_comb] ^ p20_literal_1076347[p21_res7__109_comb] ^ p20_literal_1076349[p21_res7__108_comb] ^ p20_literal_1076351[p21_res7__107_comb] ^ p20_literal_1076353[p21_res7__106_comb] ^ p20_literal_1076355[p20_res7__105] ^ p20_res7__104 ^ p20_literal_1076358[p20_res7__103] ^ p20_res7__102 ^ p21_array_index_1080433_comb ^ p20_array_index_1080283 ^ p20_array_index_1080259 ^ p20_array_index_1080233 ^ p20_array_index_1080101 ^ p20_array_index_1080072 ^ p20_array_index_1080039;
  assign p21_res__6_comb = {p21_res7__111_comb, p21_res7__110_comb, p21_res7__109_comb, p21_res7__108_comb, p21_res7__107_comb, p21_res7__106_comb, p20_res7__105, p20_res7__104, p20_res7__103, p20_res7__102, p20_res7__101, p20_res7__100, p20_res7__99, p20_res7__98, p20_res7__97, p20_res7__96};
  assign p21_k3_comb = p21_res__6_comb ^ p20_xor_1079529;

  // Registers for pipe stage 21:
  reg [127:0] p21_xor_1080001;
  reg [127:0] p21_k3;
  reg [127:0] p21_res__33;
  reg [7:0] p22_arr[256];
  reg [7:0] p22_literal_1076345[256];
  reg [7:0] p22_literal_1076347[256];
  reg [7:0] p22_literal_1076349[256];
  reg [7:0] p22_literal_1076351[256];
  reg [7:0] p22_literal_1076353[256];
  reg [7:0] p22_literal_1076355[256];
  reg [7:0] p22_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p21_xor_1080001 <= p20_xor_1080001;
    p21_k3 <= p21_k3_comb;
    p21_res__33 <= p20_res__33;
    p22_arr <= p21_arr;
    p22_literal_1076345 <= p21_literal_1076345;
    p22_literal_1076347 <= p21_literal_1076347;
    p22_literal_1076349 <= p21_literal_1076349;
    p22_literal_1076351 <= p21_literal_1076351;
    p22_literal_1076353 <= p21_literal_1076353;
    p22_literal_1076355 <= p21_literal_1076355;
    p22_literal_1076358 <= p21_literal_1076358;
  end

  // ===== Pipe stage 22:
  wire [127:0] p22_addedKey__48_comb;
  wire [7:0] p22_array_index_1080511_comb;
  wire [7:0] p22_array_index_1080512_comb;
  wire [7:0] p22_array_index_1080513_comb;
  wire [7:0] p22_array_index_1080514_comb;
  wire [7:0] p22_array_index_1080515_comb;
  wire [7:0] p22_array_index_1080516_comb;
  wire [7:0] p22_array_index_1080518_comb;
  wire [7:0] p22_array_index_1080520_comb;
  wire [7:0] p22_array_index_1080521_comb;
  wire [7:0] p22_array_index_1080522_comb;
  wire [7:0] p22_array_index_1080523_comb;
  wire [7:0] p22_array_index_1080524_comb;
  wire [7:0] p22_array_index_1080525_comb;
  wire [7:0] p22_array_index_1080527_comb;
  wire [7:0] p22_array_index_1080528_comb;
  wire [7:0] p22_array_index_1080529_comb;
  wire [7:0] p22_array_index_1080530_comb;
  wire [7:0] p22_array_index_1080531_comb;
  wire [7:0] p22_array_index_1080532_comb;
  wire [7:0] p22_array_index_1080533_comb;
  wire [7:0] p22_array_index_1080535_comb;
  wire [7:0] p22_res7__112_comb;
  wire [7:0] p22_array_index_1080544_comb;
  wire [7:0] p22_array_index_1080545_comb;
  wire [7:0] p22_array_index_1080546_comb;
  wire [7:0] p22_array_index_1080547_comb;
  wire [7:0] p22_array_index_1080548_comb;
  wire [7:0] p22_array_index_1080549_comb;
  wire [7:0] p22_res7__113_comb;
  wire [7:0] p22_array_index_1080559_comb;
  wire [7:0] p22_array_index_1080560_comb;
  wire [7:0] p22_array_index_1080561_comb;
  wire [7:0] p22_array_index_1080562_comb;
  wire [7:0] p22_array_index_1080563_comb;
  wire [7:0] p22_res7__114_comb;
  wire [7:0] p22_array_index_1080573_comb;
  wire [7:0] p22_array_index_1080574_comb;
  wire [7:0] p22_array_index_1080575_comb;
  wire [7:0] p22_array_index_1080576_comb;
  wire [7:0] p22_array_index_1080577_comb;
  wire [7:0] p22_res7__115_comb;
  wire [7:0] p22_array_index_1080588_comb;
  wire [7:0] p22_array_index_1080589_comb;
  wire [7:0] p22_array_index_1080590_comb;
  wire [7:0] p22_array_index_1080591_comb;
  wire [7:0] p22_res7__116_comb;
  assign p22_addedKey__48_comb = p21_k3 ^ 128'hf659_3616_e605_5689_adfb_a180_27aa_2a08;
  assign p22_array_index_1080511_comb = p21_arr[p22_addedKey__48_comb[127:120]];
  assign p22_array_index_1080512_comb = p21_arr[p22_addedKey__48_comb[119:112]];
  assign p22_array_index_1080513_comb = p21_arr[p22_addedKey__48_comb[111:104]];
  assign p22_array_index_1080514_comb = p21_arr[p22_addedKey__48_comb[103:96]];
  assign p22_array_index_1080515_comb = p21_arr[p22_addedKey__48_comb[95:88]];
  assign p22_array_index_1080516_comb = p21_arr[p22_addedKey__48_comb[87:80]];
  assign p22_array_index_1080518_comb = p21_arr[p22_addedKey__48_comb[71:64]];
  assign p22_array_index_1080520_comb = p21_arr[p22_addedKey__48_comb[55:48]];
  assign p22_array_index_1080521_comb = p21_arr[p22_addedKey__48_comb[47:40]];
  assign p22_array_index_1080522_comb = p21_arr[p22_addedKey__48_comb[39:32]];
  assign p22_array_index_1080523_comb = p21_arr[p22_addedKey__48_comb[31:24]];
  assign p22_array_index_1080524_comb = p21_arr[p22_addedKey__48_comb[23:16]];
  assign p22_array_index_1080525_comb = p21_arr[p22_addedKey__48_comb[15:8]];
  assign p22_array_index_1080527_comb = p21_literal_1076345[p22_array_index_1080511_comb];
  assign p22_array_index_1080528_comb = p21_literal_1076347[p22_array_index_1080512_comb];
  assign p22_array_index_1080529_comb = p21_literal_1076349[p22_array_index_1080513_comb];
  assign p22_array_index_1080530_comb = p21_literal_1076351[p22_array_index_1080514_comb];
  assign p22_array_index_1080531_comb = p21_literal_1076353[p22_array_index_1080515_comb];
  assign p22_array_index_1080532_comb = p21_literal_1076355[p22_array_index_1080516_comb];
  assign p22_array_index_1080533_comb = p21_arr[p22_addedKey__48_comb[79:72]];
  assign p22_array_index_1080535_comb = p21_arr[p22_addedKey__48_comb[63:56]];
  assign p22_res7__112_comb = p22_array_index_1080527_comb ^ p22_array_index_1080528_comb ^ p22_array_index_1080529_comb ^ p22_array_index_1080530_comb ^ p22_array_index_1080531_comb ^ p22_array_index_1080532_comb ^ p22_array_index_1080533_comb ^ p21_literal_1076358[p22_array_index_1080518_comb] ^ p22_array_index_1080535_comb ^ p21_literal_1076355[p22_array_index_1080520_comb] ^ p21_literal_1076353[p22_array_index_1080521_comb] ^ p21_literal_1076351[p22_array_index_1080522_comb] ^ p21_literal_1076349[p22_array_index_1080523_comb] ^ p21_literal_1076347[p22_array_index_1080524_comb] ^ p21_literal_1076345[p22_array_index_1080525_comb] ^ p21_arr[p22_addedKey__48_comb[7:0]];
  assign p22_array_index_1080544_comb = p21_literal_1076345[p22_res7__112_comb];
  assign p22_array_index_1080545_comb = p21_literal_1076347[p22_array_index_1080511_comb];
  assign p22_array_index_1080546_comb = p21_literal_1076349[p22_array_index_1080512_comb];
  assign p22_array_index_1080547_comb = p21_literal_1076351[p22_array_index_1080513_comb];
  assign p22_array_index_1080548_comb = p21_literal_1076353[p22_array_index_1080514_comb];
  assign p22_array_index_1080549_comb = p21_literal_1076355[p22_array_index_1080515_comb];
  assign p22_res7__113_comb = p22_array_index_1080544_comb ^ p22_array_index_1080545_comb ^ p22_array_index_1080546_comb ^ p22_array_index_1080547_comb ^ p22_array_index_1080548_comb ^ p22_array_index_1080549_comb ^ p22_array_index_1080516_comb ^ p21_literal_1076358[p22_array_index_1080533_comb] ^ p22_array_index_1080518_comb ^ p21_literal_1076355[p22_array_index_1080535_comb] ^ p21_literal_1076353[p22_array_index_1080520_comb] ^ p21_literal_1076351[p22_array_index_1080521_comb] ^ p21_literal_1076349[p22_array_index_1080522_comb] ^ p21_literal_1076347[p22_array_index_1080523_comb] ^ p21_literal_1076345[p22_array_index_1080524_comb] ^ p22_array_index_1080525_comb;
  assign p22_array_index_1080559_comb = p21_literal_1076347[p22_res7__112_comb];
  assign p22_array_index_1080560_comb = p21_literal_1076349[p22_array_index_1080511_comb];
  assign p22_array_index_1080561_comb = p21_literal_1076351[p22_array_index_1080512_comb];
  assign p22_array_index_1080562_comb = p21_literal_1076353[p22_array_index_1080513_comb];
  assign p22_array_index_1080563_comb = p21_literal_1076355[p22_array_index_1080514_comb];
  assign p22_res7__114_comb = p21_literal_1076345[p22_res7__113_comb] ^ p22_array_index_1080559_comb ^ p22_array_index_1080560_comb ^ p22_array_index_1080561_comb ^ p22_array_index_1080562_comb ^ p22_array_index_1080563_comb ^ p22_array_index_1080515_comb ^ p21_literal_1076358[p22_array_index_1080516_comb] ^ p22_array_index_1080533_comb ^ p21_literal_1076355[p22_array_index_1080518_comb] ^ p21_literal_1076353[p22_array_index_1080535_comb] ^ p21_literal_1076351[p22_array_index_1080520_comb] ^ p21_literal_1076349[p22_array_index_1080521_comb] ^ p21_literal_1076347[p22_array_index_1080522_comb] ^ p21_literal_1076345[p22_array_index_1080523_comb] ^ p22_array_index_1080524_comb;
  assign p22_array_index_1080573_comb = p21_literal_1076347[p22_res7__113_comb];
  assign p22_array_index_1080574_comb = p21_literal_1076349[p22_res7__112_comb];
  assign p22_array_index_1080575_comb = p21_literal_1076351[p22_array_index_1080511_comb];
  assign p22_array_index_1080576_comb = p21_literal_1076353[p22_array_index_1080512_comb];
  assign p22_array_index_1080577_comb = p21_literal_1076355[p22_array_index_1080513_comb];
  assign p22_res7__115_comb = p21_literal_1076345[p22_res7__114_comb] ^ p22_array_index_1080573_comb ^ p22_array_index_1080574_comb ^ p22_array_index_1080575_comb ^ p22_array_index_1080576_comb ^ p22_array_index_1080577_comb ^ p22_array_index_1080514_comb ^ p21_literal_1076358[p22_array_index_1080515_comb] ^ p22_array_index_1080516_comb ^ p21_literal_1076355[p22_array_index_1080533_comb] ^ p21_literal_1076353[p22_array_index_1080518_comb] ^ p21_literal_1076351[p22_array_index_1080535_comb] ^ p21_literal_1076349[p22_array_index_1080520_comb] ^ p21_literal_1076347[p22_array_index_1080521_comb] ^ p21_literal_1076345[p22_array_index_1080522_comb] ^ p22_array_index_1080523_comb;
  assign p22_array_index_1080588_comb = p21_literal_1076349[p22_res7__113_comb];
  assign p22_array_index_1080589_comb = p21_literal_1076351[p22_res7__112_comb];
  assign p22_array_index_1080590_comb = p21_literal_1076353[p22_array_index_1080511_comb];
  assign p22_array_index_1080591_comb = p21_literal_1076355[p22_array_index_1080512_comb];
  assign p22_res7__116_comb = p21_literal_1076345[p22_res7__115_comb] ^ p21_literal_1076347[p22_res7__114_comb] ^ p22_array_index_1080588_comb ^ p22_array_index_1080589_comb ^ p22_array_index_1080590_comb ^ p22_array_index_1080591_comb ^ p22_array_index_1080513_comb ^ p21_literal_1076358[p22_array_index_1080514_comb] ^ p22_array_index_1080515_comb ^ p22_array_index_1080532_comb ^ p21_literal_1076353[p22_array_index_1080533_comb] ^ p21_literal_1076351[p22_array_index_1080518_comb] ^ p21_literal_1076349[p22_array_index_1080535_comb] ^ p21_literal_1076347[p22_array_index_1080520_comb] ^ p21_literal_1076345[p22_array_index_1080521_comb] ^ p22_array_index_1080522_comb;

  // Registers for pipe stage 22:
  reg [127:0] p22_xor_1080001;
  reg [127:0] p22_k3;
  reg [7:0] p22_array_index_1080511;
  reg [7:0] p22_array_index_1080512;
  reg [7:0] p22_array_index_1080513;
  reg [7:0] p22_array_index_1080514;
  reg [7:0] p22_array_index_1080515;
  reg [7:0] p22_array_index_1080516;
  reg [7:0] p22_array_index_1080518;
  reg [7:0] p22_array_index_1080520;
  reg [7:0] p22_array_index_1080521;
  reg [7:0] p22_array_index_1080527;
  reg [7:0] p22_array_index_1080528;
  reg [7:0] p22_array_index_1080529;
  reg [7:0] p22_array_index_1080530;
  reg [7:0] p22_array_index_1080531;
  reg [7:0] p22_array_index_1080533;
  reg [7:0] p22_array_index_1080535;
  reg [7:0] p22_res7__112;
  reg [7:0] p22_array_index_1080544;
  reg [7:0] p22_array_index_1080545;
  reg [7:0] p22_array_index_1080546;
  reg [7:0] p22_array_index_1080547;
  reg [7:0] p22_array_index_1080548;
  reg [7:0] p22_array_index_1080549;
  reg [7:0] p22_res7__113;
  reg [7:0] p22_array_index_1080559;
  reg [7:0] p22_array_index_1080560;
  reg [7:0] p22_array_index_1080561;
  reg [7:0] p22_array_index_1080562;
  reg [7:0] p22_array_index_1080563;
  reg [7:0] p22_res7__114;
  reg [7:0] p22_array_index_1080573;
  reg [7:0] p22_array_index_1080574;
  reg [7:0] p22_array_index_1080575;
  reg [7:0] p22_array_index_1080576;
  reg [7:0] p22_array_index_1080577;
  reg [7:0] p22_res7__115;
  reg [7:0] p22_array_index_1080588;
  reg [7:0] p22_array_index_1080589;
  reg [7:0] p22_array_index_1080590;
  reg [7:0] p22_array_index_1080591;
  reg [7:0] p22_res7__116;
  reg [127:0] p22_res__33;
  reg [7:0] p23_arr[256];
  reg [7:0] p23_literal_1076345[256];
  reg [7:0] p23_literal_1076347[256];
  reg [7:0] p23_literal_1076349[256];
  reg [7:0] p23_literal_1076351[256];
  reg [7:0] p23_literal_1076353[256];
  reg [7:0] p23_literal_1076355[256];
  reg [7:0] p23_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p22_xor_1080001 <= p21_xor_1080001;
    p22_k3 <= p21_k3;
    p22_array_index_1080511 <= p22_array_index_1080511_comb;
    p22_array_index_1080512 <= p22_array_index_1080512_comb;
    p22_array_index_1080513 <= p22_array_index_1080513_comb;
    p22_array_index_1080514 <= p22_array_index_1080514_comb;
    p22_array_index_1080515 <= p22_array_index_1080515_comb;
    p22_array_index_1080516 <= p22_array_index_1080516_comb;
    p22_array_index_1080518 <= p22_array_index_1080518_comb;
    p22_array_index_1080520 <= p22_array_index_1080520_comb;
    p22_array_index_1080521 <= p22_array_index_1080521_comb;
    p22_array_index_1080527 <= p22_array_index_1080527_comb;
    p22_array_index_1080528 <= p22_array_index_1080528_comb;
    p22_array_index_1080529 <= p22_array_index_1080529_comb;
    p22_array_index_1080530 <= p22_array_index_1080530_comb;
    p22_array_index_1080531 <= p22_array_index_1080531_comb;
    p22_array_index_1080533 <= p22_array_index_1080533_comb;
    p22_array_index_1080535 <= p22_array_index_1080535_comb;
    p22_res7__112 <= p22_res7__112_comb;
    p22_array_index_1080544 <= p22_array_index_1080544_comb;
    p22_array_index_1080545 <= p22_array_index_1080545_comb;
    p22_array_index_1080546 <= p22_array_index_1080546_comb;
    p22_array_index_1080547 <= p22_array_index_1080547_comb;
    p22_array_index_1080548 <= p22_array_index_1080548_comb;
    p22_array_index_1080549 <= p22_array_index_1080549_comb;
    p22_res7__113 <= p22_res7__113_comb;
    p22_array_index_1080559 <= p22_array_index_1080559_comb;
    p22_array_index_1080560 <= p22_array_index_1080560_comb;
    p22_array_index_1080561 <= p22_array_index_1080561_comb;
    p22_array_index_1080562 <= p22_array_index_1080562_comb;
    p22_array_index_1080563 <= p22_array_index_1080563_comb;
    p22_res7__114 <= p22_res7__114_comb;
    p22_array_index_1080573 <= p22_array_index_1080573_comb;
    p22_array_index_1080574 <= p22_array_index_1080574_comb;
    p22_array_index_1080575 <= p22_array_index_1080575_comb;
    p22_array_index_1080576 <= p22_array_index_1080576_comb;
    p22_array_index_1080577 <= p22_array_index_1080577_comb;
    p22_res7__115 <= p22_res7__115_comb;
    p22_array_index_1080588 <= p22_array_index_1080588_comb;
    p22_array_index_1080589 <= p22_array_index_1080589_comb;
    p22_array_index_1080590 <= p22_array_index_1080590_comb;
    p22_array_index_1080591 <= p22_array_index_1080591_comb;
    p22_res7__116 <= p22_res7__116_comb;
    p22_res__33 <= p21_res__33;
    p23_arr <= p22_arr;
    p23_literal_1076345 <= p22_literal_1076345;
    p23_literal_1076347 <= p22_literal_1076347;
    p23_literal_1076349 <= p22_literal_1076349;
    p23_literal_1076351 <= p22_literal_1076351;
    p23_literal_1076353 <= p22_literal_1076353;
    p23_literal_1076355 <= p22_literal_1076355;
    p23_literal_1076358 <= p22_literal_1076358;
  end

  // ===== Pipe stage 23:
  wire [7:0] p23_array_index_1080705_comb;
  wire [7:0] p23_array_index_1080706_comb;
  wire [7:0] p23_array_index_1080707_comb;
  wire [7:0] p23_array_index_1080708_comb;
  wire [7:0] p23_res7__117_comb;
  wire [7:0] p23_array_index_1080719_comb;
  wire [7:0] p23_array_index_1080720_comb;
  wire [7:0] p23_array_index_1080721_comb;
  wire [7:0] p23_res7__118_comb;
  wire [7:0] p23_array_index_1080731_comb;
  wire [7:0] p23_array_index_1080732_comb;
  wire [7:0] p23_array_index_1080733_comb;
  wire [7:0] p23_res7__119_comb;
  wire [7:0] p23_array_index_1080744_comb;
  wire [7:0] p23_array_index_1080745_comb;
  wire [7:0] p23_res7__120_comb;
  wire [7:0] p23_array_index_1080755_comb;
  wire [7:0] p23_array_index_1080756_comb;
  wire [7:0] p23_res7__121_comb;
  wire [7:0] p23_array_index_1080762_comb;
  wire [7:0] p23_array_index_1080763_comb;
  wire [7:0] p23_array_index_1080764_comb;
  wire [7:0] p23_array_index_1080765_comb;
  wire [7:0] p23_array_index_1080766_comb;
  wire [7:0] p23_array_index_1080767_comb;
  wire [7:0] p23_array_index_1080768_comb;
  wire [7:0] p23_array_index_1080769_comb;
  wire [7:0] p23_array_index_1080770_comb;
  assign p23_array_index_1080705_comb = p22_literal_1076349[p22_res7__114];
  assign p23_array_index_1080706_comb = p22_literal_1076351[p22_res7__113];
  assign p23_array_index_1080707_comb = p22_literal_1076353[p22_res7__112];
  assign p23_array_index_1080708_comb = p22_literal_1076355[p22_array_index_1080511];
  assign p23_res7__117_comb = p22_literal_1076345[p22_res7__116] ^ p22_literal_1076347[p22_res7__115] ^ p23_array_index_1080705_comb ^ p23_array_index_1080706_comb ^ p23_array_index_1080707_comb ^ p23_array_index_1080708_comb ^ p22_array_index_1080512 ^ p22_literal_1076358[p22_array_index_1080513] ^ p22_array_index_1080514 ^ p22_array_index_1080549 ^ p22_literal_1076353[p22_array_index_1080516] ^ p22_literal_1076351[p22_array_index_1080533] ^ p22_literal_1076349[p22_array_index_1080518] ^ p22_literal_1076347[p22_array_index_1080535] ^ p22_literal_1076345[p22_array_index_1080520] ^ p22_array_index_1080521;
  assign p23_array_index_1080719_comb = p22_literal_1076351[p22_res7__114];
  assign p23_array_index_1080720_comb = p22_literal_1076353[p22_res7__113];
  assign p23_array_index_1080721_comb = p22_literal_1076355[p22_res7__112];
  assign p23_res7__118_comb = p22_literal_1076345[p23_res7__117_comb] ^ p22_literal_1076347[p22_res7__116] ^ p22_literal_1076349[p22_res7__115] ^ p23_array_index_1080719_comb ^ p23_array_index_1080720_comb ^ p23_array_index_1080721_comb ^ p22_array_index_1080511 ^ p22_literal_1076358[p22_array_index_1080512] ^ p22_array_index_1080513 ^ p22_array_index_1080563 ^ p22_array_index_1080531 ^ p22_literal_1076351[p22_array_index_1080516] ^ p22_literal_1076349[p22_array_index_1080533] ^ p22_literal_1076347[p22_array_index_1080518] ^ p22_literal_1076345[p22_array_index_1080535] ^ p22_array_index_1080520;
  assign p23_array_index_1080731_comb = p22_literal_1076351[p22_res7__115];
  assign p23_array_index_1080732_comb = p22_literal_1076353[p22_res7__114];
  assign p23_array_index_1080733_comb = p22_literal_1076355[p22_res7__113];
  assign p23_res7__119_comb = p22_literal_1076345[p23_res7__118_comb] ^ p22_literal_1076347[p23_res7__117_comb] ^ p22_literal_1076349[p22_res7__116] ^ p23_array_index_1080731_comb ^ p23_array_index_1080732_comb ^ p23_array_index_1080733_comb ^ p22_res7__112 ^ p22_literal_1076358[p22_array_index_1080511] ^ p22_array_index_1080512 ^ p22_array_index_1080577 ^ p22_array_index_1080548 ^ p22_literal_1076351[p22_array_index_1080515] ^ p22_literal_1076349[p22_array_index_1080516] ^ p22_literal_1076347[p22_array_index_1080533] ^ p22_literal_1076345[p22_array_index_1080518] ^ p22_array_index_1080535;
  assign p23_array_index_1080744_comb = p22_literal_1076353[p22_res7__115];
  assign p23_array_index_1080745_comb = p22_literal_1076355[p22_res7__114];
  assign p23_res7__120_comb = p22_literal_1076345[p23_res7__119_comb] ^ p22_literal_1076347[p23_res7__118_comb] ^ p22_literal_1076349[p23_res7__117_comb] ^ p22_literal_1076351[p22_res7__116] ^ p23_array_index_1080744_comb ^ p23_array_index_1080745_comb ^ p22_res7__113 ^ p22_literal_1076358[p22_res7__112] ^ p22_array_index_1080511 ^ p22_array_index_1080591 ^ p22_array_index_1080562 ^ p22_array_index_1080530 ^ p22_literal_1076349[p22_array_index_1080515] ^ p22_literal_1076347[p22_array_index_1080516] ^ p22_literal_1076345[p22_array_index_1080533] ^ p22_array_index_1080518;
  assign p23_array_index_1080755_comb = p22_literal_1076353[p22_res7__116];
  assign p23_array_index_1080756_comb = p22_literal_1076355[p22_res7__115];
  assign p23_res7__121_comb = p22_literal_1076345[p23_res7__120_comb] ^ p22_literal_1076347[p23_res7__119_comb] ^ p22_literal_1076349[p23_res7__118_comb] ^ p22_literal_1076351[p23_res7__117_comb] ^ p23_array_index_1080755_comb ^ p23_array_index_1080756_comb ^ p22_res7__114 ^ p22_literal_1076358[p22_res7__113] ^ p22_res7__112 ^ p23_array_index_1080708_comb ^ p22_array_index_1080576 ^ p22_array_index_1080547 ^ p22_literal_1076349[p22_array_index_1080514] ^ p22_literal_1076347[p22_array_index_1080515] ^ p22_literal_1076345[p22_array_index_1080516] ^ p22_array_index_1080533;
  assign p23_array_index_1080762_comb = p22_literal_1076345[p23_res7__121_comb];
  assign p23_array_index_1080763_comb = p22_literal_1076347[p23_res7__120_comb];
  assign p23_array_index_1080764_comb = p22_literal_1076349[p23_res7__119_comb];
  assign p23_array_index_1080765_comb = p22_literal_1076351[p23_res7__118_comb];
  assign p23_array_index_1080766_comb = p22_literal_1076353[p23_res7__117_comb];
  assign p23_array_index_1080767_comb = p22_literal_1076355[p22_res7__116];
  assign p23_array_index_1080768_comb = p22_literal_1076358[p22_res7__114];
  assign p23_array_index_1080769_comb = p22_literal_1076347[p22_array_index_1080514];
  assign p23_array_index_1080770_comb = p22_literal_1076345[p22_array_index_1080515];

  // Registers for pipe stage 23:
  reg [127:0] p23_xor_1080001;
  reg [127:0] p23_k3;
  reg [7:0] p23_array_index_1080511;
  reg [7:0] p23_array_index_1080512;
  reg [7:0] p23_array_index_1080513;
  reg [7:0] p23_array_index_1080514;
  reg [7:0] p23_array_index_1080515;
  reg [7:0] p23_array_index_1080516;
  reg [7:0] p23_array_index_1080527;
  reg [7:0] p23_array_index_1080528;
  reg [7:0] p23_array_index_1080529;
  reg [7:0] p23_res7__112;
  reg [7:0] p23_array_index_1080544;
  reg [7:0] p23_array_index_1080545;
  reg [7:0] p23_array_index_1080546;
  reg [7:0] p23_res7__113;
  reg [7:0] p23_array_index_1080559;
  reg [7:0] p23_array_index_1080560;
  reg [7:0] p23_array_index_1080561;
  reg [7:0] p23_res7__114;
  reg [7:0] p23_array_index_1080573;
  reg [7:0] p23_array_index_1080574;
  reg [7:0] p23_array_index_1080575;
  reg [7:0] p23_res7__115;
  reg [7:0] p23_array_index_1080588;
  reg [7:0] p23_array_index_1080589;
  reg [7:0] p23_array_index_1080590;
  reg [7:0] p23_res7__116;
  reg [7:0] p23_array_index_1080705;
  reg [7:0] p23_array_index_1080706;
  reg [7:0] p23_array_index_1080707;
  reg [7:0] p23_res7__117;
  reg [7:0] p23_array_index_1080719;
  reg [7:0] p23_array_index_1080720;
  reg [7:0] p23_array_index_1080721;
  reg [7:0] p23_res7__118;
  reg [7:0] p23_array_index_1080731;
  reg [7:0] p23_array_index_1080732;
  reg [7:0] p23_array_index_1080733;
  reg [7:0] p23_res7__119;
  reg [7:0] p23_array_index_1080744;
  reg [7:0] p23_array_index_1080745;
  reg [7:0] p23_res7__120;
  reg [7:0] p23_array_index_1080755;
  reg [7:0] p23_array_index_1080756;
  reg [7:0] p23_res7__121;
  reg [7:0] p23_array_index_1080762;
  reg [7:0] p23_array_index_1080763;
  reg [7:0] p23_array_index_1080764;
  reg [7:0] p23_array_index_1080765;
  reg [7:0] p23_array_index_1080766;
  reg [7:0] p23_array_index_1080767;
  reg [7:0] p23_array_index_1080768;
  reg [7:0] p23_array_index_1080769;
  reg [7:0] p23_array_index_1080770;
  reg [127:0] p23_res__33;
  reg [7:0] p24_arr[256];
  reg [7:0] p24_literal_1076345[256];
  reg [7:0] p24_literal_1076347[256];
  reg [7:0] p24_literal_1076349[256];
  reg [7:0] p24_literal_1076351[256];
  reg [7:0] p24_literal_1076353[256];
  reg [7:0] p24_literal_1076355[256];
  reg [7:0] p24_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p23_xor_1080001 <= p22_xor_1080001;
    p23_k3 <= p22_k3;
    p23_array_index_1080511 <= p22_array_index_1080511;
    p23_array_index_1080512 <= p22_array_index_1080512;
    p23_array_index_1080513 <= p22_array_index_1080513;
    p23_array_index_1080514 <= p22_array_index_1080514;
    p23_array_index_1080515 <= p22_array_index_1080515;
    p23_array_index_1080516 <= p22_array_index_1080516;
    p23_array_index_1080527 <= p22_array_index_1080527;
    p23_array_index_1080528 <= p22_array_index_1080528;
    p23_array_index_1080529 <= p22_array_index_1080529;
    p23_res7__112 <= p22_res7__112;
    p23_array_index_1080544 <= p22_array_index_1080544;
    p23_array_index_1080545 <= p22_array_index_1080545;
    p23_array_index_1080546 <= p22_array_index_1080546;
    p23_res7__113 <= p22_res7__113;
    p23_array_index_1080559 <= p22_array_index_1080559;
    p23_array_index_1080560 <= p22_array_index_1080560;
    p23_array_index_1080561 <= p22_array_index_1080561;
    p23_res7__114 <= p22_res7__114;
    p23_array_index_1080573 <= p22_array_index_1080573;
    p23_array_index_1080574 <= p22_array_index_1080574;
    p23_array_index_1080575 <= p22_array_index_1080575;
    p23_res7__115 <= p22_res7__115;
    p23_array_index_1080588 <= p22_array_index_1080588;
    p23_array_index_1080589 <= p22_array_index_1080589;
    p23_array_index_1080590 <= p22_array_index_1080590;
    p23_res7__116 <= p22_res7__116;
    p23_array_index_1080705 <= p23_array_index_1080705_comb;
    p23_array_index_1080706 <= p23_array_index_1080706_comb;
    p23_array_index_1080707 <= p23_array_index_1080707_comb;
    p23_res7__117 <= p23_res7__117_comb;
    p23_array_index_1080719 <= p23_array_index_1080719_comb;
    p23_array_index_1080720 <= p23_array_index_1080720_comb;
    p23_array_index_1080721 <= p23_array_index_1080721_comb;
    p23_res7__118 <= p23_res7__118_comb;
    p23_array_index_1080731 <= p23_array_index_1080731_comb;
    p23_array_index_1080732 <= p23_array_index_1080732_comb;
    p23_array_index_1080733 <= p23_array_index_1080733_comb;
    p23_res7__119 <= p23_res7__119_comb;
    p23_array_index_1080744 <= p23_array_index_1080744_comb;
    p23_array_index_1080745 <= p23_array_index_1080745_comb;
    p23_res7__120 <= p23_res7__120_comb;
    p23_array_index_1080755 <= p23_array_index_1080755_comb;
    p23_array_index_1080756 <= p23_array_index_1080756_comb;
    p23_res7__121 <= p23_res7__121_comb;
    p23_array_index_1080762 <= p23_array_index_1080762_comb;
    p23_array_index_1080763 <= p23_array_index_1080763_comb;
    p23_array_index_1080764 <= p23_array_index_1080764_comb;
    p23_array_index_1080765 <= p23_array_index_1080765_comb;
    p23_array_index_1080766 <= p23_array_index_1080766_comb;
    p23_array_index_1080767 <= p23_array_index_1080767_comb;
    p23_array_index_1080768 <= p23_array_index_1080768_comb;
    p23_array_index_1080769 <= p23_array_index_1080769_comb;
    p23_array_index_1080770 <= p23_array_index_1080770_comb;
    p23_res__33 <= p22_res__33;
    p24_arr <= p23_arr;
    p24_literal_1076345 <= p23_literal_1076345;
    p24_literal_1076347 <= p23_literal_1076347;
    p24_literal_1076349 <= p23_literal_1076349;
    p24_literal_1076351 <= p23_literal_1076351;
    p24_literal_1076353 <= p23_literal_1076353;
    p24_literal_1076355 <= p23_literal_1076355;
    p24_literal_1076358 <= p23_literal_1076358;
  end

  // ===== Pipe stage 24:
  wire [7:0] p24_res7__122_comb;
  wire [7:0] p24_array_index_1080905_comb;
  wire [7:0] p24_res7__123_comb;
  wire [7:0] p24_res7__124_comb;
  wire [7:0] p24_res7__125_comb;
  wire [7:0] p24_res7__126_comb;
  wire [7:0] p24_res7__127_comb;
  wire [127:0] p24_res__7_comb;
  wire [127:0] p24_k2_comb;
  wire [127:0] p24_addedKey__34_comb;
  wire [7:0] p24_bit_slice_1080947_comb;
  wire [7:0] p24_bit_slice_1080948_comb;
  wire [7:0] p24_bit_slice_1080949_comb;
  wire [7:0] p24_bit_slice_1080950_comb;
  wire [7:0] p24_bit_slice_1080951_comb;
  wire [7:0] p24_bit_slice_1080952_comb;
  wire [7:0] p24_bit_slice_1080953_comb;
  wire [7:0] p24_bit_slice_1080954_comb;
  wire [7:0] p24_bit_slice_1080955_comb;
  wire [7:0] p24_bit_slice_1080956_comb;
  wire [7:0] p24_bit_slice_1080957_comb;
  wire [7:0] p24_bit_slice_1080958_comb;
  wire [7:0] p24_bit_slice_1080959_comb;
  wire [7:0] p24_bit_slice_1080960_comb;
  wire [7:0] p24_bit_slice_1080961_comb;
  wire [7:0] p24_bit_slice_1080962_comb;
  assign p24_res7__122_comb = p23_array_index_1080762 ^ p23_array_index_1080763 ^ p23_array_index_1080764 ^ p23_array_index_1080765 ^ p23_array_index_1080766 ^ p23_array_index_1080767 ^ p23_res7__115 ^ p23_array_index_1080768 ^ p23_res7__113 ^ p23_array_index_1080721 ^ p23_array_index_1080590 ^ p23_array_index_1080561 ^ p23_array_index_1080529 ^ p23_array_index_1080769 ^ p23_array_index_1080770 ^ p23_array_index_1080516;
  assign p24_array_index_1080905_comb = p23_literal_1076355[p23_res7__117];
  assign p24_res7__123_comb = p23_literal_1076345[p24_res7__122_comb] ^ p23_literal_1076347[p23_res7__121] ^ p23_literal_1076349[p23_res7__120] ^ p23_literal_1076351[p23_res7__119] ^ p23_literal_1076353[p23_res7__118] ^ p24_array_index_1080905_comb ^ p23_res7__116 ^ p23_literal_1076358[p23_res7__115] ^ p23_res7__114 ^ p23_array_index_1080733 ^ p23_array_index_1080707 ^ p23_array_index_1080575 ^ p23_array_index_1080546 ^ p23_literal_1076347[p23_array_index_1080513] ^ p23_literal_1076345[p23_array_index_1080514] ^ p23_array_index_1080515;
  assign p24_res7__124_comb = p23_literal_1076345[p24_res7__123_comb] ^ p23_literal_1076347[p24_res7__122_comb] ^ p23_literal_1076349[p23_res7__121] ^ p23_literal_1076351[p23_res7__120] ^ p23_literal_1076353[p23_res7__119] ^ p23_literal_1076355[p23_res7__118] ^ p23_res7__117 ^ p23_literal_1076358[p23_res7__116] ^ p23_res7__115 ^ p23_array_index_1080745 ^ p23_array_index_1080720 ^ p23_array_index_1080589 ^ p23_array_index_1080560 ^ p23_array_index_1080528 ^ p23_literal_1076345[p23_array_index_1080513] ^ p23_array_index_1080514;
  assign p24_res7__125_comb = p23_literal_1076345[p24_res7__124_comb] ^ p23_literal_1076347[p24_res7__123_comb] ^ p23_literal_1076349[p24_res7__122_comb] ^ p23_literal_1076351[p23_res7__121] ^ p23_literal_1076353[p23_res7__120] ^ p23_literal_1076355[p23_res7__119] ^ p23_res7__118 ^ p23_literal_1076358[p23_res7__117] ^ p23_res7__116 ^ p23_array_index_1080756 ^ p23_array_index_1080732 ^ p23_array_index_1080706 ^ p23_array_index_1080574 ^ p23_array_index_1080545 ^ p23_literal_1076345[p23_array_index_1080512] ^ p23_array_index_1080513;
  assign p24_res7__126_comb = p23_literal_1076345[p24_res7__125_comb] ^ p23_literal_1076347[p24_res7__124_comb] ^ p23_literal_1076349[p24_res7__123_comb] ^ p23_literal_1076351[p24_res7__122_comb] ^ p23_literal_1076353[p23_res7__121] ^ p23_literal_1076355[p23_res7__120] ^ p23_res7__119 ^ p23_literal_1076358[p23_res7__118] ^ p23_res7__117 ^ p23_array_index_1080767 ^ p23_array_index_1080744 ^ p23_array_index_1080719 ^ p23_array_index_1080588 ^ p23_array_index_1080559 ^ p23_array_index_1080527 ^ p23_array_index_1080512;
  assign p24_res7__127_comb = p23_literal_1076345[p24_res7__126_comb] ^ p23_literal_1076347[p24_res7__125_comb] ^ p23_literal_1076349[p24_res7__124_comb] ^ p23_literal_1076351[p24_res7__123_comb] ^ p23_literal_1076353[p24_res7__122_comb] ^ p23_literal_1076355[p23_res7__121] ^ p23_res7__120 ^ p23_literal_1076358[p23_res7__119] ^ p23_res7__118 ^ p24_array_index_1080905_comb ^ p23_array_index_1080755 ^ p23_array_index_1080731 ^ p23_array_index_1080705 ^ p23_array_index_1080573 ^ p23_array_index_1080544 ^ p23_array_index_1080511;
  assign p24_res__7_comb = {p24_res7__127_comb, p24_res7__126_comb, p24_res7__125_comb, p24_res7__124_comb, p24_res7__123_comb, p24_res7__122_comb, p23_res7__121, p23_res7__120, p23_res7__119, p23_res7__118, p23_res7__117, p23_res7__116, p23_res7__115, p23_res7__114, p23_res7__113, p23_res7__112};
  assign p24_k2_comb = p24_res__7_comb ^ p23_xor_1080001;
  assign p24_addedKey__34_comb = p24_k2_comb ^ p23_res__33;
  assign p24_bit_slice_1080947_comb = p24_addedKey__34_comb[127:120];
  assign p24_bit_slice_1080948_comb = p24_addedKey__34_comb[119:112];
  assign p24_bit_slice_1080949_comb = p24_addedKey__34_comb[111:104];
  assign p24_bit_slice_1080950_comb = p24_addedKey__34_comb[103:96];
  assign p24_bit_slice_1080951_comb = p24_addedKey__34_comb[95:88];
  assign p24_bit_slice_1080952_comb = p24_addedKey__34_comb[87:80];
  assign p24_bit_slice_1080953_comb = p24_addedKey__34_comb[71:64];
  assign p24_bit_slice_1080954_comb = p24_addedKey__34_comb[55:48];
  assign p24_bit_slice_1080955_comb = p24_addedKey__34_comb[47:40];
  assign p24_bit_slice_1080956_comb = p24_addedKey__34_comb[39:32];
  assign p24_bit_slice_1080957_comb = p24_addedKey__34_comb[31:24];
  assign p24_bit_slice_1080958_comb = p24_addedKey__34_comb[23:16];
  assign p24_bit_slice_1080959_comb = p24_addedKey__34_comb[15:8];
  assign p24_bit_slice_1080960_comb = p24_addedKey__34_comb[79:72];
  assign p24_bit_slice_1080961_comb = p24_addedKey__34_comb[63:56];
  assign p24_bit_slice_1080962_comb = p24_addedKey__34_comb[7:0];

  // Registers for pipe stage 24:
  reg [127:0] p24_k3;
  reg [127:0] p24_k2;
  reg [7:0] p24_bit_slice_1080947;
  reg [7:0] p24_bit_slice_1080948;
  reg [7:0] p24_bit_slice_1080949;
  reg [7:0] p24_bit_slice_1080950;
  reg [7:0] p24_bit_slice_1080951;
  reg [7:0] p24_bit_slice_1080952;
  reg [7:0] p24_bit_slice_1080953;
  reg [7:0] p24_bit_slice_1080954;
  reg [7:0] p24_bit_slice_1080955;
  reg [7:0] p24_bit_slice_1080956;
  reg [7:0] p24_bit_slice_1080957;
  reg [7:0] p24_bit_slice_1080958;
  reg [7:0] p24_bit_slice_1080959;
  reg [7:0] p24_bit_slice_1080960;
  reg [7:0] p24_bit_slice_1080961;
  reg [7:0] p24_bit_slice_1080962;
  reg [7:0] p25_arr[256];
  reg [7:0] p25_literal_1076345[256];
  reg [7:0] p25_literal_1076347[256];
  reg [7:0] p25_literal_1076349[256];
  reg [7:0] p25_literal_1076351[256];
  reg [7:0] p25_literal_1076353[256];
  reg [7:0] p25_literal_1076355[256];
  reg [7:0] p25_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p24_k3 <= p23_k3;
    p24_k2 <= p24_k2_comb;
    p24_bit_slice_1080947 <= p24_bit_slice_1080947_comb;
    p24_bit_slice_1080948 <= p24_bit_slice_1080948_comb;
    p24_bit_slice_1080949 <= p24_bit_slice_1080949_comb;
    p24_bit_slice_1080950 <= p24_bit_slice_1080950_comb;
    p24_bit_slice_1080951 <= p24_bit_slice_1080951_comb;
    p24_bit_slice_1080952 <= p24_bit_slice_1080952_comb;
    p24_bit_slice_1080953 <= p24_bit_slice_1080953_comb;
    p24_bit_slice_1080954 <= p24_bit_slice_1080954_comb;
    p24_bit_slice_1080955 <= p24_bit_slice_1080955_comb;
    p24_bit_slice_1080956 <= p24_bit_slice_1080956_comb;
    p24_bit_slice_1080957 <= p24_bit_slice_1080957_comb;
    p24_bit_slice_1080958 <= p24_bit_slice_1080958_comb;
    p24_bit_slice_1080959 <= p24_bit_slice_1080959_comb;
    p24_bit_slice_1080960 <= p24_bit_slice_1080960_comb;
    p24_bit_slice_1080961 <= p24_bit_slice_1080961_comb;
    p24_bit_slice_1080962 <= p24_bit_slice_1080962_comb;
    p25_arr <= p24_arr;
    p25_literal_1076345 <= p24_literal_1076345;
    p25_literal_1076347 <= p24_literal_1076347;
    p25_literal_1076349 <= p24_literal_1076349;
    p25_literal_1076351 <= p24_literal_1076351;
    p25_literal_1076353 <= p24_literal_1076353;
    p25_literal_1076355 <= p24_literal_1076355;
    p25_literal_1076358 <= p24_literal_1076358;
  end

  // ===== Pipe stage 25:
  wire [127:0] p25_addedKey__49_comb;
  wire [7:0] p25_array_index_1081030_comb;
  wire [7:0] p25_array_index_1081031_comb;
  wire [7:0] p25_array_index_1081032_comb;
  wire [7:0] p25_array_index_1081033_comb;
  wire [7:0] p25_array_index_1081034_comb;
  wire [7:0] p25_array_index_1081035_comb;
  wire [7:0] p25_array_index_1081037_comb;
  wire [7:0] p25_array_index_1081039_comb;
  wire [7:0] p25_array_index_1081040_comb;
  wire [7:0] p25_array_index_1081041_comb;
  wire [7:0] p25_array_index_1081042_comb;
  wire [7:0] p25_array_index_1081043_comb;
  wire [7:0] p25_array_index_1081044_comb;
  wire [7:0] p25_array_index_1081118_comb;
  wire [7:0] p25_array_index_1081119_comb;
  wire [7:0] p25_array_index_1081120_comb;
  wire [7:0] p25_array_index_1081121_comb;
  wire [7:0] p25_array_index_1081122_comb;
  wire [7:0] p25_array_index_1081123_comb;
  wire [7:0] p25_array_index_1081124_comb;
  wire [7:0] p25_array_index_1081125_comb;
  wire [7:0] p25_array_index_1081126_comb;
  wire [7:0] p25_array_index_1081127_comb;
  wire [7:0] p25_array_index_1081128_comb;
  wire [7:0] p25_array_index_1081129_comb;
  wire [7:0] p25_array_index_1081130_comb;
  wire [7:0] p25_array_index_1081046_comb;
  wire [7:0] p25_array_index_1081047_comb;
  wire [7:0] p25_array_index_1081048_comb;
  wire [7:0] p25_array_index_1081049_comb;
  wire [7:0] p25_array_index_1081050_comb;
  wire [7:0] p25_array_index_1081051_comb;
  wire [7:0] p25_array_index_1081052_comb;
  wire [7:0] p25_array_index_1081054_comb;
  wire [7:0] p25_array_index_1081131_comb;
  wire [7:0] p25_array_index_1081132_comb;
  wire [7:0] p25_array_index_1081133_comb;
  wire [7:0] p25_array_index_1081134_comb;
  wire [7:0] p25_array_index_1081135_comb;
  wire [7:0] p25_array_index_1081136_comb;
  wire [7:0] p25_array_index_1081137_comb;
  wire [7:0] p25_array_index_1081139_comb;
  wire [7:0] p25_res7__128_comb;
  wire [7:0] p25_res7__544_comb;
  wire [7:0] p25_array_index_1081063_comb;
  wire [7:0] p25_array_index_1081064_comb;
  wire [7:0] p25_array_index_1081065_comb;
  wire [7:0] p25_array_index_1081066_comb;
  wire [7:0] p25_array_index_1081067_comb;
  wire [7:0] p25_array_index_1081068_comb;
  wire [7:0] p25_array_index_1081148_comb;
  wire [7:0] p25_array_index_1081149_comb;
  wire [7:0] p25_array_index_1081150_comb;
  wire [7:0] p25_array_index_1081151_comb;
  wire [7:0] p25_array_index_1081152_comb;
  wire [7:0] p25_array_index_1081153_comb;
  wire [7:0] p25_res7__129_comb;
  wire [7:0] p25_res7__545_comb;
  wire [7:0] p25_array_index_1081078_comb;
  wire [7:0] p25_array_index_1081079_comb;
  wire [7:0] p25_array_index_1081080_comb;
  wire [7:0] p25_array_index_1081081_comb;
  wire [7:0] p25_array_index_1081082_comb;
  wire [7:0] p25_array_index_1081163_comb;
  wire [7:0] p25_array_index_1081164_comb;
  wire [7:0] p25_array_index_1081165_comb;
  wire [7:0] p25_array_index_1081166_comb;
  wire [7:0] p25_array_index_1081167_comb;
  wire [7:0] p25_res7__130_comb;
  wire [7:0] p25_res7__546_comb;
  wire [7:0] p25_array_index_1081092_comb;
  wire [7:0] p25_array_index_1081093_comb;
  wire [7:0] p25_array_index_1081094_comb;
  wire [7:0] p25_array_index_1081095_comb;
  wire [7:0] p25_array_index_1081096_comb;
  wire [7:0] p25_array_index_1081177_comb;
  wire [7:0] p25_array_index_1081178_comb;
  wire [7:0] p25_array_index_1081179_comb;
  wire [7:0] p25_array_index_1081180_comb;
  wire [7:0] p25_array_index_1081181_comb;
  wire [7:0] p25_res7__131_comb;
  wire [7:0] p25_res7__547_comb;
  wire [7:0] p25_array_index_1081107_comb;
  wire [7:0] p25_array_index_1081108_comb;
  wire [7:0] p25_array_index_1081109_comb;
  wire [7:0] p25_array_index_1081110_comb;
  wire [7:0] p25_array_index_1081192_comb;
  wire [7:0] p25_array_index_1081193_comb;
  wire [7:0] p25_array_index_1081194_comb;
  wire [7:0] p25_array_index_1081195_comb;
  wire [7:0] p25_res7__132_comb;
  wire [7:0] p25_res7__548_comb;
  assign p25_addedKey__49_comb = p24_k2 ^ 128'h98fb_4064_8a4d_2c31_f0dc_1c90_fa2e_be09;
  assign p25_array_index_1081030_comb = p24_arr[p25_addedKey__49_comb[127:120]];
  assign p25_array_index_1081031_comb = p24_arr[p25_addedKey__49_comb[119:112]];
  assign p25_array_index_1081032_comb = p24_arr[p25_addedKey__49_comb[111:104]];
  assign p25_array_index_1081033_comb = p24_arr[p25_addedKey__49_comb[103:96]];
  assign p25_array_index_1081034_comb = p24_arr[p25_addedKey__49_comb[95:88]];
  assign p25_array_index_1081035_comb = p24_arr[p25_addedKey__49_comb[87:80]];
  assign p25_array_index_1081037_comb = p24_arr[p25_addedKey__49_comb[71:64]];
  assign p25_array_index_1081039_comb = p24_arr[p25_addedKey__49_comb[55:48]];
  assign p25_array_index_1081040_comb = p24_arr[p25_addedKey__49_comb[47:40]];
  assign p25_array_index_1081041_comb = p24_arr[p25_addedKey__49_comb[39:32]];
  assign p25_array_index_1081042_comb = p24_arr[p25_addedKey__49_comb[31:24]];
  assign p25_array_index_1081043_comb = p24_arr[p25_addedKey__49_comb[23:16]];
  assign p25_array_index_1081044_comb = p24_arr[p25_addedKey__49_comb[15:8]];
  assign p25_array_index_1081118_comb = p24_arr[p24_bit_slice_1080947];
  assign p25_array_index_1081119_comb = p24_arr[p24_bit_slice_1080948];
  assign p25_array_index_1081120_comb = p24_arr[p24_bit_slice_1080949];
  assign p25_array_index_1081121_comb = p24_arr[p24_bit_slice_1080950];
  assign p25_array_index_1081122_comb = p24_arr[p24_bit_slice_1080951];
  assign p25_array_index_1081123_comb = p24_arr[p24_bit_slice_1080952];
  assign p25_array_index_1081124_comb = p24_arr[p24_bit_slice_1080953];
  assign p25_array_index_1081125_comb = p24_arr[p24_bit_slice_1080954];
  assign p25_array_index_1081126_comb = p24_arr[p24_bit_slice_1080955];
  assign p25_array_index_1081127_comb = p24_arr[p24_bit_slice_1080956];
  assign p25_array_index_1081128_comb = p24_arr[p24_bit_slice_1080957];
  assign p25_array_index_1081129_comb = p24_arr[p24_bit_slice_1080958];
  assign p25_array_index_1081130_comb = p24_arr[p24_bit_slice_1080959];
  assign p25_array_index_1081046_comb = p24_literal_1076345[p25_array_index_1081030_comb];
  assign p25_array_index_1081047_comb = p24_literal_1076347[p25_array_index_1081031_comb];
  assign p25_array_index_1081048_comb = p24_literal_1076349[p25_array_index_1081032_comb];
  assign p25_array_index_1081049_comb = p24_literal_1076351[p25_array_index_1081033_comb];
  assign p25_array_index_1081050_comb = p24_literal_1076353[p25_array_index_1081034_comb];
  assign p25_array_index_1081051_comb = p24_literal_1076355[p25_array_index_1081035_comb];
  assign p25_array_index_1081052_comb = p24_arr[p25_addedKey__49_comb[79:72]];
  assign p25_array_index_1081054_comb = p24_arr[p25_addedKey__49_comb[63:56]];
  assign p25_array_index_1081131_comb = p24_literal_1076345[p25_array_index_1081118_comb];
  assign p25_array_index_1081132_comb = p24_literal_1076347[p25_array_index_1081119_comb];
  assign p25_array_index_1081133_comb = p24_literal_1076349[p25_array_index_1081120_comb];
  assign p25_array_index_1081134_comb = p24_literal_1076351[p25_array_index_1081121_comb];
  assign p25_array_index_1081135_comb = p24_literal_1076353[p25_array_index_1081122_comb];
  assign p25_array_index_1081136_comb = p24_literal_1076355[p25_array_index_1081123_comb];
  assign p25_array_index_1081137_comb = p24_arr[p24_bit_slice_1080960];
  assign p25_array_index_1081139_comb = p24_arr[p24_bit_slice_1080961];
  assign p25_res7__128_comb = p25_array_index_1081046_comb ^ p25_array_index_1081047_comb ^ p25_array_index_1081048_comb ^ p25_array_index_1081049_comb ^ p25_array_index_1081050_comb ^ p25_array_index_1081051_comb ^ p25_array_index_1081052_comb ^ p24_literal_1076358[p25_array_index_1081037_comb] ^ p25_array_index_1081054_comb ^ p24_literal_1076355[p25_array_index_1081039_comb] ^ p24_literal_1076353[p25_array_index_1081040_comb] ^ p24_literal_1076351[p25_array_index_1081041_comb] ^ p24_literal_1076349[p25_array_index_1081042_comb] ^ p24_literal_1076347[p25_array_index_1081043_comb] ^ p24_literal_1076345[p25_array_index_1081044_comb] ^ p24_arr[p25_addedKey__49_comb[7:0]];
  assign p25_res7__544_comb = p25_array_index_1081131_comb ^ p25_array_index_1081132_comb ^ p25_array_index_1081133_comb ^ p25_array_index_1081134_comb ^ p25_array_index_1081135_comb ^ p25_array_index_1081136_comb ^ p25_array_index_1081137_comb ^ p24_literal_1076358[p25_array_index_1081124_comb] ^ p25_array_index_1081139_comb ^ p24_literal_1076355[p25_array_index_1081125_comb] ^ p24_literal_1076353[p25_array_index_1081126_comb] ^ p24_literal_1076351[p25_array_index_1081127_comb] ^ p24_literal_1076349[p25_array_index_1081128_comb] ^ p24_literal_1076347[p25_array_index_1081129_comb] ^ p24_literal_1076345[p25_array_index_1081130_comb] ^ p24_arr[p24_bit_slice_1080962];
  assign p25_array_index_1081063_comb = p24_literal_1076345[p25_res7__128_comb];
  assign p25_array_index_1081064_comb = p24_literal_1076347[p25_array_index_1081030_comb];
  assign p25_array_index_1081065_comb = p24_literal_1076349[p25_array_index_1081031_comb];
  assign p25_array_index_1081066_comb = p24_literal_1076351[p25_array_index_1081032_comb];
  assign p25_array_index_1081067_comb = p24_literal_1076353[p25_array_index_1081033_comb];
  assign p25_array_index_1081068_comb = p24_literal_1076355[p25_array_index_1081034_comb];
  assign p25_array_index_1081148_comb = p24_literal_1076345[p25_res7__544_comb];
  assign p25_array_index_1081149_comb = p24_literal_1076347[p25_array_index_1081118_comb];
  assign p25_array_index_1081150_comb = p24_literal_1076349[p25_array_index_1081119_comb];
  assign p25_array_index_1081151_comb = p24_literal_1076351[p25_array_index_1081120_comb];
  assign p25_array_index_1081152_comb = p24_literal_1076353[p25_array_index_1081121_comb];
  assign p25_array_index_1081153_comb = p24_literal_1076355[p25_array_index_1081122_comb];
  assign p25_res7__129_comb = p25_array_index_1081063_comb ^ p25_array_index_1081064_comb ^ p25_array_index_1081065_comb ^ p25_array_index_1081066_comb ^ p25_array_index_1081067_comb ^ p25_array_index_1081068_comb ^ p25_array_index_1081035_comb ^ p24_literal_1076358[p25_array_index_1081052_comb] ^ p25_array_index_1081037_comb ^ p24_literal_1076355[p25_array_index_1081054_comb] ^ p24_literal_1076353[p25_array_index_1081039_comb] ^ p24_literal_1076351[p25_array_index_1081040_comb] ^ p24_literal_1076349[p25_array_index_1081041_comb] ^ p24_literal_1076347[p25_array_index_1081042_comb] ^ p24_literal_1076345[p25_array_index_1081043_comb] ^ p25_array_index_1081044_comb;
  assign p25_res7__545_comb = p25_array_index_1081148_comb ^ p25_array_index_1081149_comb ^ p25_array_index_1081150_comb ^ p25_array_index_1081151_comb ^ p25_array_index_1081152_comb ^ p25_array_index_1081153_comb ^ p25_array_index_1081123_comb ^ p24_literal_1076358[p25_array_index_1081137_comb] ^ p25_array_index_1081124_comb ^ p24_literal_1076355[p25_array_index_1081139_comb] ^ p24_literal_1076353[p25_array_index_1081125_comb] ^ p24_literal_1076351[p25_array_index_1081126_comb] ^ p24_literal_1076349[p25_array_index_1081127_comb] ^ p24_literal_1076347[p25_array_index_1081128_comb] ^ p24_literal_1076345[p25_array_index_1081129_comb] ^ p25_array_index_1081130_comb;
  assign p25_array_index_1081078_comb = p24_literal_1076347[p25_res7__128_comb];
  assign p25_array_index_1081079_comb = p24_literal_1076349[p25_array_index_1081030_comb];
  assign p25_array_index_1081080_comb = p24_literal_1076351[p25_array_index_1081031_comb];
  assign p25_array_index_1081081_comb = p24_literal_1076353[p25_array_index_1081032_comb];
  assign p25_array_index_1081082_comb = p24_literal_1076355[p25_array_index_1081033_comb];
  assign p25_array_index_1081163_comb = p24_literal_1076347[p25_res7__544_comb];
  assign p25_array_index_1081164_comb = p24_literal_1076349[p25_array_index_1081118_comb];
  assign p25_array_index_1081165_comb = p24_literal_1076351[p25_array_index_1081119_comb];
  assign p25_array_index_1081166_comb = p24_literal_1076353[p25_array_index_1081120_comb];
  assign p25_array_index_1081167_comb = p24_literal_1076355[p25_array_index_1081121_comb];
  assign p25_res7__130_comb = p24_literal_1076345[p25_res7__129_comb] ^ p25_array_index_1081078_comb ^ p25_array_index_1081079_comb ^ p25_array_index_1081080_comb ^ p25_array_index_1081081_comb ^ p25_array_index_1081082_comb ^ p25_array_index_1081034_comb ^ p24_literal_1076358[p25_array_index_1081035_comb] ^ p25_array_index_1081052_comb ^ p24_literal_1076355[p25_array_index_1081037_comb] ^ p24_literal_1076353[p25_array_index_1081054_comb] ^ p24_literal_1076351[p25_array_index_1081039_comb] ^ p24_literal_1076349[p25_array_index_1081040_comb] ^ p24_literal_1076347[p25_array_index_1081041_comb] ^ p24_literal_1076345[p25_array_index_1081042_comb] ^ p25_array_index_1081043_comb;
  assign p25_res7__546_comb = p24_literal_1076345[p25_res7__545_comb] ^ p25_array_index_1081163_comb ^ p25_array_index_1081164_comb ^ p25_array_index_1081165_comb ^ p25_array_index_1081166_comb ^ p25_array_index_1081167_comb ^ p25_array_index_1081122_comb ^ p24_literal_1076358[p25_array_index_1081123_comb] ^ p25_array_index_1081137_comb ^ p24_literal_1076355[p25_array_index_1081124_comb] ^ p24_literal_1076353[p25_array_index_1081139_comb] ^ p24_literal_1076351[p25_array_index_1081125_comb] ^ p24_literal_1076349[p25_array_index_1081126_comb] ^ p24_literal_1076347[p25_array_index_1081127_comb] ^ p24_literal_1076345[p25_array_index_1081128_comb] ^ p25_array_index_1081129_comb;
  assign p25_array_index_1081092_comb = p24_literal_1076347[p25_res7__129_comb];
  assign p25_array_index_1081093_comb = p24_literal_1076349[p25_res7__128_comb];
  assign p25_array_index_1081094_comb = p24_literal_1076351[p25_array_index_1081030_comb];
  assign p25_array_index_1081095_comb = p24_literal_1076353[p25_array_index_1081031_comb];
  assign p25_array_index_1081096_comb = p24_literal_1076355[p25_array_index_1081032_comb];
  assign p25_array_index_1081177_comb = p24_literal_1076347[p25_res7__545_comb];
  assign p25_array_index_1081178_comb = p24_literal_1076349[p25_res7__544_comb];
  assign p25_array_index_1081179_comb = p24_literal_1076351[p25_array_index_1081118_comb];
  assign p25_array_index_1081180_comb = p24_literal_1076353[p25_array_index_1081119_comb];
  assign p25_array_index_1081181_comb = p24_literal_1076355[p25_array_index_1081120_comb];
  assign p25_res7__131_comb = p24_literal_1076345[p25_res7__130_comb] ^ p25_array_index_1081092_comb ^ p25_array_index_1081093_comb ^ p25_array_index_1081094_comb ^ p25_array_index_1081095_comb ^ p25_array_index_1081096_comb ^ p25_array_index_1081033_comb ^ p24_literal_1076358[p25_array_index_1081034_comb] ^ p25_array_index_1081035_comb ^ p24_literal_1076355[p25_array_index_1081052_comb] ^ p24_literal_1076353[p25_array_index_1081037_comb] ^ p24_literal_1076351[p25_array_index_1081054_comb] ^ p24_literal_1076349[p25_array_index_1081039_comb] ^ p24_literal_1076347[p25_array_index_1081040_comb] ^ p24_literal_1076345[p25_array_index_1081041_comb] ^ p25_array_index_1081042_comb;
  assign p25_res7__547_comb = p24_literal_1076345[p25_res7__546_comb] ^ p25_array_index_1081177_comb ^ p25_array_index_1081178_comb ^ p25_array_index_1081179_comb ^ p25_array_index_1081180_comb ^ p25_array_index_1081181_comb ^ p25_array_index_1081121_comb ^ p24_literal_1076358[p25_array_index_1081122_comb] ^ p25_array_index_1081123_comb ^ p24_literal_1076355[p25_array_index_1081137_comb] ^ p24_literal_1076353[p25_array_index_1081124_comb] ^ p24_literal_1076351[p25_array_index_1081139_comb] ^ p24_literal_1076349[p25_array_index_1081125_comb] ^ p24_literal_1076347[p25_array_index_1081126_comb] ^ p24_literal_1076345[p25_array_index_1081127_comb] ^ p25_array_index_1081128_comb;
  assign p25_array_index_1081107_comb = p24_literal_1076349[p25_res7__129_comb];
  assign p25_array_index_1081108_comb = p24_literal_1076351[p25_res7__128_comb];
  assign p25_array_index_1081109_comb = p24_literal_1076353[p25_array_index_1081030_comb];
  assign p25_array_index_1081110_comb = p24_literal_1076355[p25_array_index_1081031_comb];
  assign p25_array_index_1081192_comb = p24_literal_1076349[p25_res7__545_comb];
  assign p25_array_index_1081193_comb = p24_literal_1076351[p25_res7__544_comb];
  assign p25_array_index_1081194_comb = p24_literal_1076353[p25_array_index_1081118_comb];
  assign p25_array_index_1081195_comb = p24_literal_1076355[p25_array_index_1081119_comb];
  assign p25_res7__132_comb = p24_literal_1076345[p25_res7__131_comb] ^ p24_literal_1076347[p25_res7__130_comb] ^ p25_array_index_1081107_comb ^ p25_array_index_1081108_comb ^ p25_array_index_1081109_comb ^ p25_array_index_1081110_comb ^ p25_array_index_1081032_comb ^ p24_literal_1076358[p25_array_index_1081033_comb] ^ p25_array_index_1081034_comb ^ p25_array_index_1081051_comb ^ p24_literal_1076353[p25_array_index_1081052_comb] ^ p24_literal_1076351[p25_array_index_1081037_comb] ^ p24_literal_1076349[p25_array_index_1081054_comb] ^ p24_literal_1076347[p25_array_index_1081039_comb] ^ p24_literal_1076345[p25_array_index_1081040_comb] ^ p25_array_index_1081041_comb;
  assign p25_res7__548_comb = p24_literal_1076345[p25_res7__547_comb] ^ p24_literal_1076347[p25_res7__546_comb] ^ p25_array_index_1081192_comb ^ p25_array_index_1081193_comb ^ p25_array_index_1081194_comb ^ p25_array_index_1081195_comb ^ p25_array_index_1081120_comb ^ p24_literal_1076358[p25_array_index_1081121_comb] ^ p25_array_index_1081122_comb ^ p25_array_index_1081136_comb ^ p24_literal_1076353[p25_array_index_1081137_comb] ^ p24_literal_1076351[p25_array_index_1081124_comb] ^ p24_literal_1076349[p25_array_index_1081139_comb] ^ p24_literal_1076347[p25_array_index_1081125_comb] ^ p24_literal_1076345[p25_array_index_1081126_comb] ^ p25_array_index_1081127_comb;

  // Registers for pipe stage 25:
  reg [127:0] p25_k3;
  reg [127:0] p25_k2;
  reg [7:0] p25_array_index_1081030;
  reg [7:0] p25_array_index_1081031;
  reg [7:0] p25_array_index_1081032;
  reg [7:0] p25_array_index_1081033;
  reg [7:0] p25_array_index_1081034;
  reg [7:0] p25_array_index_1081035;
  reg [7:0] p25_array_index_1081037;
  reg [7:0] p25_array_index_1081039;
  reg [7:0] p25_array_index_1081040;
  reg [7:0] p25_array_index_1081046;
  reg [7:0] p25_array_index_1081047;
  reg [7:0] p25_array_index_1081048;
  reg [7:0] p25_array_index_1081049;
  reg [7:0] p25_array_index_1081050;
  reg [7:0] p25_array_index_1081052;
  reg [7:0] p25_array_index_1081054;
  reg [7:0] p25_res7__128;
  reg [7:0] p25_array_index_1081063;
  reg [7:0] p25_array_index_1081064;
  reg [7:0] p25_array_index_1081065;
  reg [7:0] p25_array_index_1081066;
  reg [7:0] p25_array_index_1081067;
  reg [7:0] p25_array_index_1081068;
  reg [7:0] p25_res7__129;
  reg [7:0] p25_array_index_1081078;
  reg [7:0] p25_array_index_1081079;
  reg [7:0] p25_array_index_1081080;
  reg [7:0] p25_array_index_1081081;
  reg [7:0] p25_array_index_1081082;
  reg [7:0] p25_res7__130;
  reg [7:0] p25_array_index_1081092;
  reg [7:0] p25_array_index_1081093;
  reg [7:0] p25_array_index_1081094;
  reg [7:0] p25_array_index_1081095;
  reg [7:0] p25_array_index_1081096;
  reg [7:0] p25_res7__131;
  reg [7:0] p25_array_index_1081107;
  reg [7:0] p25_array_index_1081108;
  reg [7:0] p25_array_index_1081109;
  reg [7:0] p25_array_index_1081110;
  reg [7:0] p25_res7__132;
  reg [7:0] p25_array_index_1081118;
  reg [7:0] p25_array_index_1081119;
  reg [7:0] p25_array_index_1081120;
  reg [7:0] p25_array_index_1081121;
  reg [7:0] p25_array_index_1081122;
  reg [7:0] p25_array_index_1081123;
  reg [7:0] p25_array_index_1081124;
  reg [7:0] p25_array_index_1081125;
  reg [7:0] p25_array_index_1081126;
  reg [7:0] p25_array_index_1081131;
  reg [7:0] p25_array_index_1081132;
  reg [7:0] p25_array_index_1081133;
  reg [7:0] p25_array_index_1081134;
  reg [7:0] p25_array_index_1081135;
  reg [7:0] p25_array_index_1081137;
  reg [7:0] p25_array_index_1081139;
  reg [7:0] p25_res7__544;
  reg [7:0] p25_array_index_1081148;
  reg [7:0] p25_array_index_1081149;
  reg [7:0] p25_array_index_1081150;
  reg [7:0] p25_array_index_1081151;
  reg [7:0] p25_array_index_1081152;
  reg [7:0] p25_array_index_1081153;
  reg [7:0] p25_res7__545;
  reg [7:0] p25_array_index_1081163;
  reg [7:0] p25_array_index_1081164;
  reg [7:0] p25_array_index_1081165;
  reg [7:0] p25_array_index_1081166;
  reg [7:0] p25_array_index_1081167;
  reg [7:0] p25_res7__546;
  reg [7:0] p25_array_index_1081177;
  reg [7:0] p25_array_index_1081178;
  reg [7:0] p25_array_index_1081179;
  reg [7:0] p25_array_index_1081180;
  reg [7:0] p25_array_index_1081181;
  reg [7:0] p25_res7__547;
  reg [7:0] p25_array_index_1081192;
  reg [7:0] p25_array_index_1081193;
  reg [7:0] p25_array_index_1081194;
  reg [7:0] p25_array_index_1081195;
  reg [7:0] p25_res7__548;
  reg [7:0] p26_arr[256];
  reg [7:0] p26_literal_1076345[256];
  reg [7:0] p26_literal_1076347[256];
  reg [7:0] p26_literal_1076349[256];
  reg [7:0] p26_literal_1076351[256];
  reg [7:0] p26_literal_1076353[256];
  reg [7:0] p26_literal_1076355[256];
  reg [7:0] p26_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p25_k3 <= p24_k3;
    p25_k2 <= p24_k2;
    p25_array_index_1081030 <= p25_array_index_1081030_comb;
    p25_array_index_1081031 <= p25_array_index_1081031_comb;
    p25_array_index_1081032 <= p25_array_index_1081032_comb;
    p25_array_index_1081033 <= p25_array_index_1081033_comb;
    p25_array_index_1081034 <= p25_array_index_1081034_comb;
    p25_array_index_1081035 <= p25_array_index_1081035_comb;
    p25_array_index_1081037 <= p25_array_index_1081037_comb;
    p25_array_index_1081039 <= p25_array_index_1081039_comb;
    p25_array_index_1081040 <= p25_array_index_1081040_comb;
    p25_array_index_1081046 <= p25_array_index_1081046_comb;
    p25_array_index_1081047 <= p25_array_index_1081047_comb;
    p25_array_index_1081048 <= p25_array_index_1081048_comb;
    p25_array_index_1081049 <= p25_array_index_1081049_comb;
    p25_array_index_1081050 <= p25_array_index_1081050_comb;
    p25_array_index_1081052 <= p25_array_index_1081052_comb;
    p25_array_index_1081054 <= p25_array_index_1081054_comb;
    p25_res7__128 <= p25_res7__128_comb;
    p25_array_index_1081063 <= p25_array_index_1081063_comb;
    p25_array_index_1081064 <= p25_array_index_1081064_comb;
    p25_array_index_1081065 <= p25_array_index_1081065_comb;
    p25_array_index_1081066 <= p25_array_index_1081066_comb;
    p25_array_index_1081067 <= p25_array_index_1081067_comb;
    p25_array_index_1081068 <= p25_array_index_1081068_comb;
    p25_res7__129 <= p25_res7__129_comb;
    p25_array_index_1081078 <= p25_array_index_1081078_comb;
    p25_array_index_1081079 <= p25_array_index_1081079_comb;
    p25_array_index_1081080 <= p25_array_index_1081080_comb;
    p25_array_index_1081081 <= p25_array_index_1081081_comb;
    p25_array_index_1081082 <= p25_array_index_1081082_comb;
    p25_res7__130 <= p25_res7__130_comb;
    p25_array_index_1081092 <= p25_array_index_1081092_comb;
    p25_array_index_1081093 <= p25_array_index_1081093_comb;
    p25_array_index_1081094 <= p25_array_index_1081094_comb;
    p25_array_index_1081095 <= p25_array_index_1081095_comb;
    p25_array_index_1081096 <= p25_array_index_1081096_comb;
    p25_res7__131 <= p25_res7__131_comb;
    p25_array_index_1081107 <= p25_array_index_1081107_comb;
    p25_array_index_1081108 <= p25_array_index_1081108_comb;
    p25_array_index_1081109 <= p25_array_index_1081109_comb;
    p25_array_index_1081110 <= p25_array_index_1081110_comb;
    p25_res7__132 <= p25_res7__132_comb;
    p25_array_index_1081118 <= p25_array_index_1081118_comb;
    p25_array_index_1081119 <= p25_array_index_1081119_comb;
    p25_array_index_1081120 <= p25_array_index_1081120_comb;
    p25_array_index_1081121 <= p25_array_index_1081121_comb;
    p25_array_index_1081122 <= p25_array_index_1081122_comb;
    p25_array_index_1081123 <= p25_array_index_1081123_comb;
    p25_array_index_1081124 <= p25_array_index_1081124_comb;
    p25_array_index_1081125 <= p25_array_index_1081125_comb;
    p25_array_index_1081126 <= p25_array_index_1081126_comb;
    p25_array_index_1081131 <= p25_array_index_1081131_comb;
    p25_array_index_1081132 <= p25_array_index_1081132_comb;
    p25_array_index_1081133 <= p25_array_index_1081133_comb;
    p25_array_index_1081134 <= p25_array_index_1081134_comb;
    p25_array_index_1081135 <= p25_array_index_1081135_comb;
    p25_array_index_1081137 <= p25_array_index_1081137_comb;
    p25_array_index_1081139 <= p25_array_index_1081139_comb;
    p25_res7__544 <= p25_res7__544_comb;
    p25_array_index_1081148 <= p25_array_index_1081148_comb;
    p25_array_index_1081149 <= p25_array_index_1081149_comb;
    p25_array_index_1081150 <= p25_array_index_1081150_comb;
    p25_array_index_1081151 <= p25_array_index_1081151_comb;
    p25_array_index_1081152 <= p25_array_index_1081152_comb;
    p25_array_index_1081153 <= p25_array_index_1081153_comb;
    p25_res7__545 <= p25_res7__545_comb;
    p25_array_index_1081163 <= p25_array_index_1081163_comb;
    p25_array_index_1081164 <= p25_array_index_1081164_comb;
    p25_array_index_1081165 <= p25_array_index_1081165_comb;
    p25_array_index_1081166 <= p25_array_index_1081166_comb;
    p25_array_index_1081167 <= p25_array_index_1081167_comb;
    p25_res7__546 <= p25_res7__546_comb;
    p25_array_index_1081177 <= p25_array_index_1081177_comb;
    p25_array_index_1081178 <= p25_array_index_1081178_comb;
    p25_array_index_1081179 <= p25_array_index_1081179_comb;
    p25_array_index_1081180 <= p25_array_index_1081180_comb;
    p25_array_index_1081181 <= p25_array_index_1081181_comb;
    p25_res7__547 <= p25_res7__547_comb;
    p25_array_index_1081192 <= p25_array_index_1081192_comb;
    p25_array_index_1081193 <= p25_array_index_1081193_comb;
    p25_array_index_1081194 <= p25_array_index_1081194_comb;
    p25_array_index_1081195 <= p25_array_index_1081195_comb;
    p25_res7__548 <= p25_res7__548_comb;
    p26_arr <= p25_arr;
    p26_literal_1076345 <= p25_literal_1076345;
    p26_literal_1076347 <= p25_literal_1076347;
    p26_literal_1076349 <= p25_literal_1076349;
    p26_literal_1076351 <= p25_literal_1076351;
    p26_literal_1076353 <= p25_literal_1076353;
    p26_literal_1076355 <= p25_literal_1076355;
    p26_literal_1076358 <= p25_literal_1076358;
  end

  // ===== Pipe stage 26:
  wire [7:0] p26_array_index_1081389_comb;
  wire [7:0] p26_array_index_1081390_comb;
  wire [7:0] p26_array_index_1081391_comb;
  wire [7:0] p26_array_index_1081392_comb;
  wire [7:0] p26_array_index_1081457_comb;
  wire [7:0] p26_array_index_1081458_comb;
  wire [7:0] p26_array_index_1081459_comb;
  wire [7:0] p26_array_index_1081460_comb;
  wire [7:0] p26_res7__133_comb;
  wire [7:0] p26_res7__549_comb;
  wire [7:0] p26_array_index_1081403_comb;
  wire [7:0] p26_array_index_1081404_comb;
  wire [7:0] p26_array_index_1081405_comb;
  wire [7:0] p26_array_index_1081471_comb;
  wire [7:0] p26_array_index_1081472_comb;
  wire [7:0] p26_array_index_1081473_comb;
  wire [7:0] p26_res7__134_comb;
  wire [7:0] p26_res7__550_comb;
  wire [7:0] p26_array_index_1081415_comb;
  wire [7:0] p26_array_index_1081416_comb;
  wire [7:0] p26_array_index_1081417_comb;
  wire [7:0] p26_array_index_1081483_comb;
  wire [7:0] p26_array_index_1081484_comb;
  wire [7:0] p26_array_index_1081485_comb;
  wire [7:0] p26_res7__135_comb;
  wire [7:0] p26_res7__551_comb;
  wire [7:0] p26_array_index_1081428_comb;
  wire [7:0] p26_array_index_1081429_comb;
  wire [7:0] p26_array_index_1081496_comb;
  wire [7:0] p26_array_index_1081497_comb;
  wire [7:0] p26_res7__136_comb;
  wire [7:0] p26_res7__552_comb;
  wire [7:0] p26_array_index_1081439_comb;
  wire [7:0] p26_array_index_1081440_comb;
  wire [7:0] p26_array_index_1081507_comb;
  wire [7:0] p26_array_index_1081508_comb;
  wire [7:0] p26_res7__137_comb;
  wire [7:0] p26_res7__553_comb;
  wire [7:0] p26_array_index_1081446_comb;
  wire [7:0] p26_array_index_1081447_comb;
  wire [7:0] p26_array_index_1081448_comb;
  wire [7:0] p26_array_index_1081449_comb;
  wire [7:0] p26_array_index_1081450_comb;
  wire [7:0] p26_array_index_1081451_comb;
  wire [7:0] p26_array_index_1081452_comb;
  wire [7:0] p26_array_index_1081453_comb;
  wire [7:0] p26_array_index_1081454_comb;
  wire [7:0] p26_array_index_1081514_comb;
  wire [7:0] p26_array_index_1081515_comb;
  wire [7:0] p26_array_index_1081516_comb;
  wire [7:0] p26_array_index_1081517_comb;
  wire [7:0] p26_array_index_1081518_comb;
  wire [7:0] p26_array_index_1081519_comb;
  wire [7:0] p26_array_index_1081520_comb;
  wire [7:0] p26_array_index_1081521_comb;
  wire [7:0] p26_array_index_1081522_comb;
  assign p26_array_index_1081389_comb = p25_literal_1076349[p25_res7__130];
  assign p26_array_index_1081390_comb = p25_literal_1076351[p25_res7__129];
  assign p26_array_index_1081391_comb = p25_literal_1076353[p25_res7__128];
  assign p26_array_index_1081392_comb = p25_literal_1076355[p25_array_index_1081030];
  assign p26_array_index_1081457_comb = p25_literal_1076349[p25_res7__546];
  assign p26_array_index_1081458_comb = p25_literal_1076351[p25_res7__545];
  assign p26_array_index_1081459_comb = p25_literal_1076353[p25_res7__544];
  assign p26_array_index_1081460_comb = p25_literal_1076355[p25_array_index_1081118];
  assign p26_res7__133_comb = p25_literal_1076345[p25_res7__132] ^ p25_literal_1076347[p25_res7__131] ^ p26_array_index_1081389_comb ^ p26_array_index_1081390_comb ^ p26_array_index_1081391_comb ^ p26_array_index_1081392_comb ^ p25_array_index_1081031 ^ p25_literal_1076358[p25_array_index_1081032] ^ p25_array_index_1081033 ^ p25_array_index_1081068 ^ p25_literal_1076353[p25_array_index_1081035] ^ p25_literal_1076351[p25_array_index_1081052] ^ p25_literal_1076349[p25_array_index_1081037] ^ p25_literal_1076347[p25_array_index_1081054] ^ p25_literal_1076345[p25_array_index_1081039] ^ p25_array_index_1081040;
  assign p26_res7__549_comb = p25_literal_1076345[p25_res7__548] ^ p25_literal_1076347[p25_res7__547] ^ p26_array_index_1081457_comb ^ p26_array_index_1081458_comb ^ p26_array_index_1081459_comb ^ p26_array_index_1081460_comb ^ p25_array_index_1081119 ^ p25_literal_1076358[p25_array_index_1081120] ^ p25_array_index_1081121 ^ p25_array_index_1081153 ^ p25_literal_1076353[p25_array_index_1081123] ^ p25_literal_1076351[p25_array_index_1081137] ^ p25_literal_1076349[p25_array_index_1081124] ^ p25_literal_1076347[p25_array_index_1081139] ^ p25_literal_1076345[p25_array_index_1081125] ^ p25_array_index_1081126;
  assign p26_array_index_1081403_comb = p25_literal_1076351[p25_res7__130];
  assign p26_array_index_1081404_comb = p25_literal_1076353[p25_res7__129];
  assign p26_array_index_1081405_comb = p25_literal_1076355[p25_res7__128];
  assign p26_array_index_1081471_comb = p25_literal_1076351[p25_res7__546];
  assign p26_array_index_1081472_comb = p25_literal_1076353[p25_res7__545];
  assign p26_array_index_1081473_comb = p25_literal_1076355[p25_res7__544];
  assign p26_res7__134_comb = p25_literal_1076345[p26_res7__133_comb] ^ p25_literal_1076347[p25_res7__132] ^ p25_literal_1076349[p25_res7__131] ^ p26_array_index_1081403_comb ^ p26_array_index_1081404_comb ^ p26_array_index_1081405_comb ^ p25_array_index_1081030 ^ p25_literal_1076358[p25_array_index_1081031] ^ p25_array_index_1081032 ^ p25_array_index_1081082 ^ p25_array_index_1081050 ^ p25_literal_1076351[p25_array_index_1081035] ^ p25_literal_1076349[p25_array_index_1081052] ^ p25_literal_1076347[p25_array_index_1081037] ^ p25_literal_1076345[p25_array_index_1081054] ^ p25_array_index_1081039;
  assign p26_res7__550_comb = p25_literal_1076345[p26_res7__549_comb] ^ p25_literal_1076347[p25_res7__548] ^ p25_literal_1076349[p25_res7__547] ^ p26_array_index_1081471_comb ^ p26_array_index_1081472_comb ^ p26_array_index_1081473_comb ^ p25_array_index_1081118 ^ p25_literal_1076358[p25_array_index_1081119] ^ p25_array_index_1081120 ^ p25_array_index_1081167 ^ p25_array_index_1081135 ^ p25_literal_1076351[p25_array_index_1081123] ^ p25_literal_1076349[p25_array_index_1081137] ^ p25_literal_1076347[p25_array_index_1081124] ^ p25_literal_1076345[p25_array_index_1081139] ^ p25_array_index_1081125;
  assign p26_array_index_1081415_comb = p25_literal_1076351[p25_res7__131];
  assign p26_array_index_1081416_comb = p25_literal_1076353[p25_res7__130];
  assign p26_array_index_1081417_comb = p25_literal_1076355[p25_res7__129];
  assign p26_array_index_1081483_comb = p25_literal_1076351[p25_res7__547];
  assign p26_array_index_1081484_comb = p25_literal_1076353[p25_res7__546];
  assign p26_array_index_1081485_comb = p25_literal_1076355[p25_res7__545];
  assign p26_res7__135_comb = p25_literal_1076345[p26_res7__134_comb] ^ p25_literal_1076347[p26_res7__133_comb] ^ p25_literal_1076349[p25_res7__132] ^ p26_array_index_1081415_comb ^ p26_array_index_1081416_comb ^ p26_array_index_1081417_comb ^ p25_res7__128 ^ p25_literal_1076358[p25_array_index_1081030] ^ p25_array_index_1081031 ^ p25_array_index_1081096 ^ p25_array_index_1081067 ^ p25_literal_1076351[p25_array_index_1081034] ^ p25_literal_1076349[p25_array_index_1081035] ^ p25_literal_1076347[p25_array_index_1081052] ^ p25_literal_1076345[p25_array_index_1081037] ^ p25_array_index_1081054;
  assign p26_res7__551_comb = p25_literal_1076345[p26_res7__550_comb] ^ p25_literal_1076347[p26_res7__549_comb] ^ p25_literal_1076349[p25_res7__548] ^ p26_array_index_1081483_comb ^ p26_array_index_1081484_comb ^ p26_array_index_1081485_comb ^ p25_res7__544 ^ p25_literal_1076358[p25_array_index_1081118] ^ p25_array_index_1081119 ^ p25_array_index_1081181 ^ p25_array_index_1081152 ^ p25_literal_1076351[p25_array_index_1081122] ^ p25_literal_1076349[p25_array_index_1081123] ^ p25_literal_1076347[p25_array_index_1081137] ^ p25_literal_1076345[p25_array_index_1081124] ^ p25_array_index_1081139;
  assign p26_array_index_1081428_comb = p25_literal_1076353[p25_res7__131];
  assign p26_array_index_1081429_comb = p25_literal_1076355[p25_res7__130];
  assign p26_array_index_1081496_comb = p25_literal_1076353[p25_res7__547];
  assign p26_array_index_1081497_comb = p25_literal_1076355[p25_res7__546];
  assign p26_res7__136_comb = p25_literal_1076345[p26_res7__135_comb] ^ p25_literal_1076347[p26_res7__134_comb] ^ p25_literal_1076349[p26_res7__133_comb] ^ p25_literal_1076351[p25_res7__132] ^ p26_array_index_1081428_comb ^ p26_array_index_1081429_comb ^ p25_res7__129 ^ p25_literal_1076358[p25_res7__128] ^ p25_array_index_1081030 ^ p25_array_index_1081110 ^ p25_array_index_1081081 ^ p25_array_index_1081049 ^ p25_literal_1076349[p25_array_index_1081034] ^ p25_literal_1076347[p25_array_index_1081035] ^ p25_literal_1076345[p25_array_index_1081052] ^ p25_array_index_1081037;
  assign p26_res7__552_comb = p25_literal_1076345[p26_res7__551_comb] ^ p25_literal_1076347[p26_res7__550_comb] ^ p25_literal_1076349[p26_res7__549_comb] ^ p25_literal_1076351[p25_res7__548] ^ p26_array_index_1081496_comb ^ p26_array_index_1081497_comb ^ p25_res7__545 ^ p25_literal_1076358[p25_res7__544] ^ p25_array_index_1081118 ^ p25_array_index_1081195 ^ p25_array_index_1081166 ^ p25_array_index_1081134 ^ p25_literal_1076349[p25_array_index_1081122] ^ p25_literal_1076347[p25_array_index_1081123] ^ p25_literal_1076345[p25_array_index_1081137] ^ p25_array_index_1081124;
  assign p26_array_index_1081439_comb = p25_literal_1076353[p25_res7__132];
  assign p26_array_index_1081440_comb = p25_literal_1076355[p25_res7__131];
  assign p26_array_index_1081507_comb = p25_literal_1076353[p25_res7__548];
  assign p26_array_index_1081508_comb = p25_literal_1076355[p25_res7__547];
  assign p26_res7__137_comb = p25_literal_1076345[p26_res7__136_comb] ^ p25_literal_1076347[p26_res7__135_comb] ^ p25_literal_1076349[p26_res7__134_comb] ^ p25_literal_1076351[p26_res7__133_comb] ^ p26_array_index_1081439_comb ^ p26_array_index_1081440_comb ^ p25_res7__130 ^ p25_literal_1076358[p25_res7__129] ^ p25_res7__128 ^ p26_array_index_1081392_comb ^ p25_array_index_1081095 ^ p25_array_index_1081066 ^ p25_literal_1076349[p25_array_index_1081033] ^ p25_literal_1076347[p25_array_index_1081034] ^ p25_literal_1076345[p25_array_index_1081035] ^ p25_array_index_1081052;
  assign p26_res7__553_comb = p25_literal_1076345[p26_res7__552_comb] ^ p25_literal_1076347[p26_res7__551_comb] ^ p25_literal_1076349[p26_res7__550_comb] ^ p25_literal_1076351[p26_res7__549_comb] ^ p26_array_index_1081507_comb ^ p26_array_index_1081508_comb ^ p25_res7__546 ^ p25_literal_1076358[p25_res7__545] ^ p25_res7__544 ^ p26_array_index_1081460_comb ^ p25_array_index_1081180 ^ p25_array_index_1081151 ^ p25_literal_1076349[p25_array_index_1081121] ^ p25_literal_1076347[p25_array_index_1081122] ^ p25_literal_1076345[p25_array_index_1081123] ^ p25_array_index_1081137;
  assign p26_array_index_1081446_comb = p25_literal_1076345[p26_res7__137_comb];
  assign p26_array_index_1081447_comb = p25_literal_1076347[p26_res7__136_comb];
  assign p26_array_index_1081448_comb = p25_literal_1076349[p26_res7__135_comb];
  assign p26_array_index_1081449_comb = p25_literal_1076351[p26_res7__134_comb];
  assign p26_array_index_1081450_comb = p25_literal_1076353[p26_res7__133_comb];
  assign p26_array_index_1081451_comb = p25_literal_1076355[p25_res7__132];
  assign p26_array_index_1081452_comb = p25_literal_1076358[p25_res7__130];
  assign p26_array_index_1081453_comb = p25_literal_1076347[p25_array_index_1081033];
  assign p26_array_index_1081454_comb = p25_literal_1076345[p25_array_index_1081034];
  assign p26_array_index_1081514_comb = p25_literal_1076345[p26_res7__553_comb];
  assign p26_array_index_1081515_comb = p25_literal_1076347[p26_res7__552_comb];
  assign p26_array_index_1081516_comb = p25_literal_1076349[p26_res7__551_comb];
  assign p26_array_index_1081517_comb = p25_literal_1076351[p26_res7__550_comb];
  assign p26_array_index_1081518_comb = p25_literal_1076353[p26_res7__549_comb];
  assign p26_array_index_1081519_comb = p25_literal_1076355[p25_res7__548];
  assign p26_array_index_1081520_comb = p25_literal_1076358[p25_res7__546];
  assign p26_array_index_1081521_comb = p25_literal_1076347[p25_array_index_1081121];
  assign p26_array_index_1081522_comb = p25_literal_1076345[p25_array_index_1081122];

  // Registers for pipe stage 26:
  reg [127:0] p26_k3;
  reg [127:0] p26_k2;
  reg [7:0] p26_array_index_1081030;
  reg [7:0] p26_array_index_1081031;
  reg [7:0] p26_array_index_1081032;
  reg [7:0] p26_array_index_1081033;
  reg [7:0] p26_array_index_1081034;
  reg [7:0] p26_array_index_1081035;
  reg [7:0] p26_array_index_1081046;
  reg [7:0] p26_array_index_1081047;
  reg [7:0] p26_array_index_1081048;
  reg [7:0] p26_res7__128;
  reg [7:0] p26_array_index_1081063;
  reg [7:0] p26_array_index_1081064;
  reg [7:0] p26_array_index_1081065;
  reg [7:0] p26_res7__129;
  reg [7:0] p26_array_index_1081078;
  reg [7:0] p26_array_index_1081079;
  reg [7:0] p26_array_index_1081080;
  reg [7:0] p26_res7__130;
  reg [7:0] p26_array_index_1081092;
  reg [7:0] p26_array_index_1081093;
  reg [7:0] p26_array_index_1081094;
  reg [7:0] p26_res7__131;
  reg [7:0] p26_array_index_1081107;
  reg [7:0] p26_array_index_1081108;
  reg [7:0] p26_array_index_1081109;
  reg [7:0] p26_res7__132;
  reg [7:0] p26_array_index_1081389;
  reg [7:0] p26_array_index_1081390;
  reg [7:0] p26_array_index_1081391;
  reg [7:0] p26_res7__133;
  reg [7:0] p26_array_index_1081403;
  reg [7:0] p26_array_index_1081404;
  reg [7:0] p26_array_index_1081405;
  reg [7:0] p26_res7__134;
  reg [7:0] p26_array_index_1081415;
  reg [7:0] p26_array_index_1081416;
  reg [7:0] p26_array_index_1081417;
  reg [7:0] p26_res7__135;
  reg [7:0] p26_array_index_1081428;
  reg [7:0] p26_array_index_1081429;
  reg [7:0] p26_res7__136;
  reg [7:0] p26_array_index_1081439;
  reg [7:0] p26_array_index_1081440;
  reg [7:0] p26_res7__137;
  reg [7:0] p26_array_index_1081446;
  reg [7:0] p26_array_index_1081447;
  reg [7:0] p26_array_index_1081448;
  reg [7:0] p26_array_index_1081449;
  reg [7:0] p26_array_index_1081450;
  reg [7:0] p26_array_index_1081451;
  reg [7:0] p26_array_index_1081452;
  reg [7:0] p26_array_index_1081453;
  reg [7:0] p26_array_index_1081454;
  reg [7:0] p26_array_index_1081118;
  reg [7:0] p26_array_index_1081119;
  reg [7:0] p26_array_index_1081120;
  reg [7:0] p26_array_index_1081121;
  reg [7:0] p26_array_index_1081122;
  reg [7:0] p26_array_index_1081123;
  reg [7:0] p26_array_index_1081131;
  reg [7:0] p26_array_index_1081132;
  reg [7:0] p26_array_index_1081133;
  reg [7:0] p26_res7__544;
  reg [7:0] p26_array_index_1081148;
  reg [7:0] p26_array_index_1081149;
  reg [7:0] p26_array_index_1081150;
  reg [7:0] p26_res7__545;
  reg [7:0] p26_array_index_1081163;
  reg [7:0] p26_array_index_1081164;
  reg [7:0] p26_array_index_1081165;
  reg [7:0] p26_res7__546;
  reg [7:0] p26_array_index_1081177;
  reg [7:0] p26_array_index_1081178;
  reg [7:0] p26_array_index_1081179;
  reg [7:0] p26_res7__547;
  reg [7:0] p26_array_index_1081192;
  reg [7:0] p26_array_index_1081193;
  reg [7:0] p26_array_index_1081194;
  reg [7:0] p26_res7__548;
  reg [7:0] p26_array_index_1081457;
  reg [7:0] p26_array_index_1081458;
  reg [7:0] p26_array_index_1081459;
  reg [7:0] p26_res7__549;
  reg [7:0] p26_array_index_1081471;
  reg [7:0] p26_array_index_1081472;
  reg [7:0] p26_array_index_1081473;
  reg [7:0] p26_res7__550;
  reg [7:0] p26_array_index_1081483;
  reg [7:0] p26_array_index_1081484;
  reg [7:0] p26_array_index_1081485;
  reg [7:0] p26_res7__551;
  reg [7:0] p26_array_index_1081496;
  reg [7:0] p26_array_index_1081497;
  reg [7:0] p26_res7__552;
  reg [7:0] p26_array_index_1081507;
  reg [7:0] p26_array_index_1081508;
  reg [7:0] p26_res7__553;
  reg [7:0] p26_array_index_1081514;
  reg [7:0] p26_array_index_1081515;
  reg [7:0] p26_array_index_1081516;
  reg [7:0] p26_array_index_1081517;
  reg [7:0] p26_array_index_1081518;
  reg [7:0] p26_array_index_1081519;
  reg [7:0] p26_array_index_1081520;
  reg [7:0] p26_array_index_1081521;
  reg [7:0] p26_array_index_1081522;
  reg [7:0] p27_arr[256];
  reg [7:0] p27_literal_1076345[256];
  reg [7:0] p27_literal_1076347[256];
  reg [7:0] p27_literal_1076349[256];
  reg [7:0] p27_literal_1076351[256];
  reg [7:0] p27_literal_1076353[256];
  reg [7:0] p27_literal_1076355[256];
  reg [7:0] p27_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p26_k3 <= p25_k3;
    p26_k2 <= p25_k2;
    p26_array_index_1081030 <= p25_array_index_1081030;
    p26_array_index_1081031 <= p25_array_index_1081031;
    p26_array_index_1081032 <= p25_array_index_1081032;
    p26_array_index_1081033 <= p25_array_index_1081033;
    p26_array_index_1081034 <= p25_array_index_1081034;
    p26_array_index_1081035 <= p25_array_index_1081035;
    p26_array_index_1081046 <= p25_array_index_1081046;
    p26_array_index_1081047 <= p25_array_index_1081047;
    p26_array_index_1081048 <= p25_array_index_1081048;
    p26_res7__128 <= p25_res7__128;
    p26_array_index_1081063 <= p25_array_index_1081063;
    p26_array_index_1081064 <= p25_array_index_1081064;
    p26_array_index_1081065 <= p25_array_index_1081065;
    p26_res7__129 <= p25_res7__129;
    p26_array_index_1081078 <= p25_array_index_1081078;
    p26_array_index_1081079 <= p25_array_index_1081079;
    p26_array_index_1081080 <= p25_array_index_1081080;
    p26_res7__130 <= p25_res7__130;
    p26_array_index_1081092 <= p25_array_index_1081092;
    p26_array_index_1081093 <= p25_array_index_1081093;
    p26_array_index_1081094 <= p25_array_index_1081094;
    p26_res7__131 <= p25_res7__131;
    p26_array_index_1081107 <= p25_array_index_1081107;
    p26_array_index_1081108 <= p25_array_index_1081108;
    p26_array_index_1081109 <= p25_array_index_1081109;
    p26_res7__132 <= p25_res7__132;
    p26_array_index_1081389 <= p26_array_index_1081389_comb;
    p26_array_index_1081390 <= p26_array_index_1081390_comb;
    p26_array_index_1081391 <= p26_array_index_1081391_comb;
    p26_res7__133 <= p26_res7__133_comb;
    p26_array_index_1081403 <= p26_array_index_1081403_comb;
    p26_array_index_1081404 <= p26_array_index_1081404_comb;
    p26_array_index_1081405 <= p26_array_index_1081405_comb;
    p26_res7__134 <= p26_res7__134_comb;
    p26_array_index_1081415 <= p26_array_index_1081415_comb;
    p26_array_index_1081416 <= p26_array_index_1081416_comb;
    p26_array_index_1081417 <= p26_array_index_1081417_comb;
    p26_res7__135 <= p26_res7__135_comb;
    p26_array_index_1081428 <= p26_array_index_1081428_comb;
    p26_array_index_1081429 <= p26_array_index_1081429_comb;
    p26_res7__136 <= p26_res7__136_comb;
    p26_array_index_1081439 <= p26_array_index_1081439_comb;
    p26_array_index_1081440 <= p26_array_index_1081440_comb;
    p26_res7__137 <= p26_res7__137_comb;
    p26_array_index_1081446 <= p26_array_index_1081446_comb;
    p26_array_index_1081447 <= p26_array_index_1081447_comb;
    p26_array_index_1081448 <= p26_array_index_1081448_comb;
    p26_array_index_1081449 <= p26_array_index_1081449_comb;
    p26_array_index_1081450 <= p26_array_index_1081450_comb;
    p26_array_index_1081451 <= p26_array_index_1081451_comb;
    p26_array_index_1081452 <= p26_array_index_1081452_comb;
    p26_array_index_1081453 <= p26_array_index_1081453_comb;
    p26_array_index_1081454 <= p26_array_index_1081454_comb;
    p26_array_index_1081118 <= p25_array_index_1081118;
    p26_array_index_1081119 <= p25_array_index_1081119;
    p26_array_index_1081120 <= p25_array_index_1081120;
    p26_array_index_1081121 <= p25_array_index_1081121;
    p26_array_index_1081122 <= p25_array_index_1081122;
    p26_array_index_1081123 <= p25_array_index_1081123;
    p26_array_index_1081131 <= p25_array_index_1081131;
    p26_array_index_1081132 <= p25_array_index_1081132;
    p26_array_index_1081133 <= p25_array_index_1081133;
    p26_res7__544 <= p25_res7__544;
    p26_array_index_1081148 <= p25_array_index_1081148;
    p26_array_index_1081149 <= p25_array_index_1081149;
    p26_array_index_1081150 <= p25_array_index_1081150;
    p26_res7__545 <= p25_res7__545;
    p26_array_index_1081163 <= p25_array_index_1081163;
    p26_array_index_1081164 <= p25_array_index_1081164;
    p26_array_index_1081165 <= p25_array_index_1081165;
    p26_res7__546 <= p25_res7__546;
    p26_array_index_1081177 <= p25_array_index_1081177;
    p26_array_index_1081178 <= p25_array_index_1081178;
    p26_array_index_1081179 <= p25_array_index_1081179;
    p26_res7__547 <= p25_res7__547;
    p26_array_index_1081192 <= p25_array_index_1081192;
    p26_array_index_1081193 <= p25_array_index_1081193;
    p26_array_index_1081194 <= p25_array_index_1081194;
    p26_res7__548 <= p25_res7__548;
    p26_array_index_1081457 <= p26_array_index_1081457_comb;
    p26_array_index_1081458 <= p26_array_index_1081458_comb;
    p26_array_index_1081459 <= p26_array_index_1081459_comb;
    p26_res7__549 <= p26_res7__549_comb;
    p26_array_index_1081471 <= p26_array_index_1081471_comb;
    p26_array_index_1081472 <= p26_array_index_1081472_comb;
    p26_array_index_1081473 <= p26_array_index_1081473_comb;
    p26_res7__550 <= p26_res7__550_comb;
    p26_array_index_1081483 <= p26_array_index_1081483_comb;
    p26_array_index_1081484 <= p26_array_index_1081484_comb;
    p26_array_index_1081485 <= p26_array_index_1081485_comb;
    p26_res7__551 <= p26_res7__551_comb;
    p26_array_index_1081496 <= p26_array_index_1081496_comb;
    p26_array_index_1081497 <= p26_array_index_1081497_comb;
    p26_res7__552 <= p26_res7__552_comb;
    p26_array_index_1081507 <= p26_array_index_1081507_comb;
    p26_array_index_1081508 <= p26_array_index_1081508_comb;
    p26_res7__553 <= p26_res7__553_comb;
    p26_array_index_1081514 <= p26_array_index_1081514_comb;
    p26_array_index_1081515 <= p26_array_index_1081515_comb;
    p26_array_index_1081516 <= p26_array_index_1081516_comb;
    p26_array_index_1081517 <= p26_array_index_1081517_comb;
    p26_array_index_1081518 <= p26_array_index_1081518_comb;
    p26_array_index_1081519 <= p26_array_index_1081519_comb;
    p26_array_index_1081520 <= p26_array_index_1081520_comb;
    p26_array_index_1081521 <= p26_array_index_1081521_comb;
    p26_array_index_1081522 <= p26_array_index_1081522_comb;
    p27_arr <= p26_arr;
    p27_literal_1076345 <= p26_literal_1076345;
    p27_literal_1076347 <= p26_literal_1076347;
    p27_literal_1076349 <= p26_literal_1076349;
    p27_literal_1076351 <= p26_literal_1076351;
    p27_literal_1076353 <= p26_literal_1076353;
    p27_literal_1076355 <= p26_literal_1076355;
    p27_literal_1076358 <= p26_literal_1076358;
  end

  // ===== Pipe stage 27:
  wire [7:0] p27_res7__554_comb;
  wire [7:0] p27_res7__138_comb;
  wire [7:0] p27_array_index_1081808_comb;
  wire [7:0] p27_array_index_1081761_comb;
  wire [7:0] p27_res7__555_comb;
  wire [7:0] p27_res7__139_comb;
  wire [7:0] p27_res7__556_comb;
  wire [7:0] p27_res7__140_comb;
  wire [7:0] p27_res7__557_comb;
  wire [7:0] p27_res7__141_comb;
  wire [7:0] p27_res7__558_comb;
  wire [7:0] p27_res7__142_comb;
  wire [7:0] p27_res7__559_comb;
  wire [7:0] p27_res7__143_comb;
  wire [127:0] p27_res__34_comb;
  wire [127:0] p27_res__8_comb;
  wire [127:0] p27_addedKey__35_comb;
  wire [127:0] p27_xor_1081801_comb;
  wire [7:0] p27_bit_slice_1081849_comb;
  wire [7:0] p27_bit_slice_1081850_comb;
  wire [7:0] p27_bit_slice_1081851_comb;
  wire [7:0] p27_bit_slice_1081852_comb;
  wire [7:0] p27_bit_slice_1081853_comb;
  wire [7:0] p27_bit_slice_1081854_comb;
  wire [7:0] p27_bit_slice_1081855_comb;
  wire [7:0] p27_bit_slice_1081856_comb;
  wire [7:0] p27_bit_slice_1081857_comb;
  wire [7:0] p27_bit_slice_1081858_comb;
  wire [7:0] p27_bit_slice_1081859_comb;
  wire [7:0] p27_bit_slice_1081860_comb;
  wire [7:0] p27_bit_slice_1081861_comb;
  wire [7:0] p27_bit_slice_1081862_comb;
  wire [7:0] p27_bit_slice_1081863_comb;
  wire [7:0] p27_bit_slice_1081864_comb;
  assign p27_res7__554_comb = p26_array_index_1081514 ^ p26_array_index_1081515 ^ p26_array_index_1081516 ^ p26_array_index_1081517 ^ p26_array_index_1081518 ^ p26_array_index_1081519 ^ p26_res7__547 ^ p26_array_index_1081520 ^ p26_res7__545 ^ p26_array_index_1081473 ^ p26_array_index_1081194 ^ p26_array_index_1081165 ^ p26_array_index_1081133 ^ p26_array_index_1081521 ^ p26_array_index_1081522 ^ p26_array_index_1081123;
  assign p27_res7__138_comb = p26_array_index_1081446 ^ p26_array_index_1081447 ^ p26_array_index_1081448 ^ p26_array_index_1081449 ^ p26_array_index_1081450 ^ p26_array_index_1081451 ^ p26_res7__131 ^ p26_array_index_1081452 ^ p26_res7__129 ^ p26_array_index_1081405 ^ p26_array_index_1081109 ^ p26_array_index_1081080 ^ p26_array_index_1081048 ^ p26_array_index_1081453 ^ p26_array_index_1081454 ^ p26_array_index_1081035;
  assign p27_array_index_1081808_comb = p26_literal_1076355[p26_res7__549];
  assign p27_array_index_1081761_comb = p26_literal_1076355[p26_res7__133];
  assign p27_res7__555_comb = p26_literal_1076345[p27_res7__554_comb] ^ p26_literal_1076347[p26_res7__553] ^ p26_literal_1076349[p26_res7__552] ^ p26_literal_1076351[p26_res7__551] ^ p26_literal_1076353[p26_res7__550] ^ p27_array_index_1081808_comb ^ p26_res7__548 ^ p26_literal_1076358[p26_res7__547] ^ p26_res7__546 ^ p26_array_index_1081485 ^ p26_array_index_1081459 ^ p26_array_index_1081179 ^ p26_array_index_1081150 ^ p26_literal_1076347[p26_array_index_1081120] ^ p26_literal_1076345[p26_array_index_1081121] ^ p26_array_index_1081122;
  assign p27_res7__139_comb = p26_literal_1076345[p27_res7__138_comb] ^ p26_literal_1076347[p26_res7__137] ^ p26_literal_1076349[p26_res7__136] ^ p26_literal_1076351[p26_res7__135] ^ p26_literal_1076353[p26_res7__134] ^ p27_array_index_1081761_comb ^ p26_res7__132 ^ p26_literal_1076358[p26_res7__131] ^ p26_res7__130 ^ p26_array_index_1081417 ^ p26_array_index_1081391 ^ p26_array_index_1081094 ^ p26_array_index_1081065 ^ p26_literal_1076347[p26_array_index_1081032] ^ p26_literal_1076345[p26_array_index_1081033] ^ p26_array_index_1081034;
  assign p27_res7__556_comb = p26_literal_1076345[p27_res7__555_comb] ^ p26_literal_1076347[p27_res7__554_comb] ^ p26_literal_1076349[p26_res7__553] ^ p26_literal_1076351[p26_res7__552] ^ p26_literal_1076353[p26_res7__551] ^ p26_literal_1076355[p26_res7__550] ^ p26_res7__549 ^ p26_literal_1076358[p26_res7__548] ^ p26_res7__547 ^ p26_array_index_1081497 ^ p26_array_index_1081472 ^ p26_array_index_1081193 ^ p26_array_index_1081164 ^ p26_array_index_1081132 ^ p26_literal_1076345[p26_array_index_1081120] ^ p26_array_index_1081121;
  assign p27_res7__140_comb = p26_literal_1076345[p27_res7__139_comb] ^ p26_literal_1076347[p27_res7__138_comb] ^ p26_literal_1076349[p26_res7__137] ^ p26_literal_1076351[p26_res7__136] ^ p26_literal_1076353[p26_res7__135] ^ p26_literal_1076355[p26_res7__134] ^ p26_res7__133 ^ p26_literal_1076358[p26_res7__132] ^ p26_res7__131 ^ p26_array_index_1081429 ^ p26_array_index_1081404 ^ p26_array_index_1081108 ^ p26_array_index_1081079 ^ p26_array_index_1081047 ^ p26_literal_1076345[p26_array_index_1081032] ^ p26_array_index_1081033;
  assign p27_res7__557_comb = p26_literal_1076345[p27_res7__556_comb] ^ p26_literal_1076347[p27_res7__555_comb] ^ p26_literal_1076349[p27_res7__554_comb] ^ p26_literal_1076351[p26_res7__553] ^ p26_literal_1076353[p26_res7__552] ^ p26_literal_1076355[p26_res7__551] ^ p26_res7__550 ^ p26_literal_1076358[p26_res7__549] ^ p26_res7__548 ^ p26_array_index_1081508 ^ p26_array_index_1081484 ^ p26_array_index_1081458 ^ p26_array_index_1081178 ^ p26_array_index_1081149 ^ p26_literal_1076345[p26_array_index_1081119] ^ p26_array_index_1081120;
  assign p27_res7__141_comb = p26_literal_1076345[p27_res7__140_comb] ^ p26_literal_1076347[p27_res7__139_comb] ^ p26_literal_1076349[p27_res7__138_comb] ^ p26_literal_1076351[p26_res7__137] ^ p26_literal_1076353[p26_res7__136] ^ p26_literal_1076355[p26_res7__135] ^ p26_res7__134 ^ p26_literal_1076358[p26_res7__133] ^ p26_res7__132 ^ p26_array_index_1081440 ^ p26_array_index_1081416 ^ p26_array_index_1081390 ^ p26_array_index_1081093 ^ p26_array_index_1081064 ^ p26_literal_1076345[p26_array_index_1081031] ^ p26_array_index_1081032;
  assign p27_res7__558_comb = p26_literal_1076345[p27_res7__557_comb] ^ p26_literal_1076347[p27_res7__556_comb] ^ p26_literal_1076349[p27_res7__555_comb] ^ p26_literal_1076351[p27_res7__554_comb] ^ p26_literal_1076353[p26_res7__553] ^ p26_literal_1076355[p26_res7__552] ^ p26_res7__551 ^ p26_literal_1076358[p26_res7__550] ^ p26_res7__549 ^ p26_array_index_1081519 ^ p26_array_index_1081496 ^ p26_array_index_1081471 ^ p26_array_index_1081192 ^ p26_array_index_1081163 ^ p26_array_index_1081131 ^ p26_array_index_1081119;
  assign p27_res7__142_comb = p26_literal_1076345[p27_res7__141_comb] ^ p26_literal_1076347[p27_res7__140_comb] ^ p26_literal_1076349[p27_res7__139_comb] ^ p26_literal_1076351[p27_res7__138_comb] ^ p26_literal_1076353[p26_res7__137] ^ p26_literal_1076355[p26_res7__136] ^ p26_res7__135 ^ p26_literal_1076358[p26_res7__134] ^ p26_res7__133 ^ p26_array_index_1081451 ^ p26_array_index_1081428 ^ p26_array_index_1081403 ^ p26_array_index_1081107 ^ p26_array_index_1081078 ^ p26_array_index_1081046 ^ p26_array_index_1081031;
  assign p27_res7__559_comb = p26_literal_1076345[p27_res7__558_comb] ^ p26_literal_1076347[p27_res7__557_comb] ^ p26_literal_1076349[p27_res7__556_comb] ^ p26_literal_1076351[p27_res7__555_comb] ^ p26_literal_1076353[p27_res7__554_comb] ^ p26_literal_1076355[p26_res7__553] ^ p26_res7__552 ^ p26_literal_1076358[p26_res7__551] ^ p26_res7__550 ^ p27_array_index_1081808_comb ^ p26_array_index_1081507 ^ p26_array_index_1081483 ^ p26_array_index_1081457 ^ p26_array_index_1081177 ^ p26_array_index_1081148 ^ p26_array_index_1081118;
  assign p27_res7__143_comb = p26_literal_1076345[p27_res7__142_comb] ^ p26_literal_1076347[p27_res7__141_comb] ^ p26_literal_1076349[p27_res7__140_comb] ^ p26_literal_1076351[p27_res7__139_comb] ^ p26_literal_1076353[p27_res7__138_comb] ^ p26_literal_1076355[p26_res7__137] ^ p26_res7__136 ^ p26_literal_1076358[p26_res7__135] ^ p26_res7__134 ^ p27_array_index_1081761_comb ^ p26_array_index_1081439 ^ p26_array_index_1081415 ^ p26_array_index_1081389 ^ p26_array_index_1081092 ^ p26_array_index_1081063 ^ p26_array_index_1081030;
  assign p27_res__34_comb = {p27_res7__559_comb, p27_res7__558_comb, p27_res7__557_comb, p27_res7__556_comb, p27_res7__555_comb, p27_res7__554_comb, p26_res7__553, p26_res7__552, p26_res7__551, p26_res7__550, p26_res7__549, p26_res7__548, p26_res7__547, p26_res7__546, p26_res7__545, p26_res7__544};
  assign p27_res__8_comb = {p27_res7__143_comb, p27_res7__142_comb, p27_res7__141_comb, p27_res7__140_comb, p27_res7__139_comb, p27_res7__138_comb, p26_res7__137, p26_res7__136, p26_res7__135, p26_res7__134, p26_res7__133, p26_res7__132, p26_res7__131, p26_res7__130, p26_res7__129, p26_res7__128};
  assign p27_addedKey__35_comb = p26_k3 ^ p27_res__34_comb;
  assign p27_xor_1081801_comb = p27_res__8_comb ^ p26_k3;
  assign p27_bit_slice_1081849_comb = p27_addedKey__35_comb[127:120];
  assign p27_bit_slice_1081850_comb = p27_addedKey__35_comb[119:112];
  assign p27_bit_slice_1081851_comb = p27_addedKey__35_comb[111:104];
  assign p27_bit_slice_1081852_comb = p27_addedKey__35_comb[103:96];
  assign p27_bit_slice_1081853_comb = p27_addedKey__35_comb[95:88];
  assign p27_bit_slice_1081854_comb = p27_addedKey__35_comb[87:80];
  assign p27_bit_slice_1081855_comb = p27_addedKey__35_comb[71:64];
  assign p27_bit_slice_1081856_comb = p27_addedKey__35_comb[55:48];
  assign p27_bit_slice_1081857_comb = p27_addedKey__35_comb[47:40];
  assign p27_bit_slice_1081858_comb = p27_addedKey__35_comb[39:32];
  assign p27_bit_slice_1081859_comb = p27_addedKey__35_comb[31:24];
  assign p27_bit_slice_1081860_comb = p27_addedKey__35_comb[23:16];
  assign p27_bit_slice_1081861_comb = p27_addedKey__35_comb[15:8];
  assign p27_bit_slice_1081862_comb = p27_addedKey__35_comb[79:72];
  assign p27_bit_slice_1081863_comb = p27_addedKey__35_comb[63:56];
  assign p27_bit_slice_1081864_comb = p27_addedKey__35_comb[7:0];

  // Registers for pipe stage 27:
  reg [127:0] p27_k2;
  reg [127:0] p27_xor_1081801;
  reg [7:0] p27_bit_slice_1081849;
  reg [7:0] p27_bit_slice_1081850;
  reg [7:0] p27_bit_slice_1081851;
  reg [7:0] p27_bit_slice_1081852;
  reg [7:0] p27_bit_slice_1081853;
  reg [7:0] p27_bit_slice_1081854;
  reg [7:0] p27_bit_slice_1081855;
  reg [7:0] p27_bit_slice_1081856;
  reg [7:0] p27_bit_slice_1081857;
  reg [7:0] p27_bit_slice_1081858;
  reg [7:0] p27_bit_slice_1081859;
  reg [7:0] p27_bit_slice_1081860;
  reg [7:0] p27_bit_slice_1081861;
  reg [7:0] p27_bit_slice_1081862;
  reg [7:0] p27_bit_slice_1081863;
  reg [7:0] p27_bit_slice_1081864;
  reg [7:0] p28_arr[256];
  reg [7:0] p28_literal_1076345[256];
  reg [7:0] p28_literal_1076347[256];
  reg [7:0] p28_literal_1076349[256];
  reg [7:0] p28_literal_1076351[256];
  reg [7:0] p28_literal_1076353[256];
  reg [7:0] p28_literal_1076355[256];
  reg [7:0] p28_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p27_k2 <= p26_k2;
    p27_xor_1081801 <= p27_xor_1081801_comb;
    p27_bit_slice_1081849 <= p27_bit_slice_1081849_comb;
    p27_bit_slice_1081850 <= p27_bit_slice_1081850_comb;
    p27_bit_slice_1081851 <= p27_bit_slice_1081851_comb;
    p27_bit_slice_1081852 <= p27_bit_slice_1081852_comb;
    p27_bit_slice_1081853 <= p27_bit_slice_1081853_comb;
    p27_bit_slice_1081854 <= p27_bit_slice_1081854_comb;
    p27_bit_slice_1081855 <= p27_bit_slice_1081855_comb;
    p27_bit_slice_1081856 <= p27_bit_slice_1081856_comb;
    p27_bit_slice_1081857 <= p27_bit_slice_1081857_comb;
    p27_bit_slice_1081858 <= p27_bit_slice_1081858_comb;
    p27_bit_slice_1081859 <= p27_bit_slice_1081859_comb;
    p27_bit_slice_1081860 <= p27_bit_slice_1081860_comb;
    p27_bit_slice_1081861 <= p27_bit_slice_1081861_comb;
    p27_bit_slice_1081862 <= p27_bit_slice_1081862_comb;
    p27_bit_slice_1081863 <= p27_bit_slice_1081863_comb;
    p27_bit_slice_1081864 <= p27_bit_slice_1081864_comb;
    p28_arr <= p27_arr;
    p28_literal_1076345 <= p27_literal_1076345;
    p28_literal_1076347 <= p27_literal_1076347;
    p28_literal_1076349 <= p27_literal_1076349;
    p28_literal_1076351 <= p27_literal_1076351;
    p28_literal_1076353 <= p27_literal_1076353;
    p28_literal_1076355 <= p27_literal_1076355;
    p28_literal_1076358 <= p27_literal_1076358;
  end

  // ===== Pipe stage 28:
  wire [127:0] p28_addedKey__50_comb;
  wire [7:0] p28_array_index_1081932_comb;
  wire [7:0] p28_array_index_1081933_comb;
  wire [7:0] p28_array_index_1081934_comb;
  wire [7:0] p28_array_index_1081935_comb;
  wire [7:0] p28_array_index_1081936_comb;
  wire [7:0] p28_array_index_1081937_comb;
  wire [7:0] p28_array_index_1081939_comb;
  wire [7:0] p28_array_index_1081941_comb;
  wire [7:0] p28_array_index_1081942_comb;
  wire [7:0] p28_array_index_1081943_comb;
  wire [7:0] p28_array_index_1081944_comb;
  wire [7:0] p28_array_index_1081945_comb;
  wire [7:0] p28_array_index_1081946_comb;
  wire [7:0] p28_array_index_1082020_comb;
  wire [7:0] p28_array_index_1082021_comb;
  wire [7:0] p28_array_index_1082022_comb;
  wire [7:0] p28_array_index_1082023_comb;
  wire [7:0] p28_array_index_1082024_comb;
  wire [7:0] p28_array_index_1082025_comb;
  wire [7:0] p28_array_index_1082026_comb;
  wire [7:0] p28_array_index_1082027_comb;
  wire [7:0] p28_array_index_1082028_comb;
  wire [7:0] p28_array_index_1082029_comb;
  wire [7:0] p28_array_index_1082030_comb;
  wire [7:0] p28_array_index_1082031_comb;
  wire [7:0] p28_array_index_1082032_comb;
  wire [7:0] p28_array_index_1081948_comb;
  wire [7:0] p28_array_index_1081949_comb;
  wire [7:0] p28_array_index_1081950_comb;
  wire [7:0] p28_array_index_1081951_comb;
  wire [7:0] p28_array_index_1081952_comb;
  wire [7:0] p28_array_index_1081953_comb;
  wire [7:0] p28_array_index_1081954_comb;
  wire [7:0] p28_array_index_1081956_comb;
  wire [7:0] p28_array_index_1082033_comb;
  wire [7:0] p28_array_index_1082034_comb;
  wire [7:0] p28_array_index_1082035_comb;
  wire [7:0] p28_array_index_1082036_comb;
  wire [7:0] p28_array_index_1082037_comb;
  wire [7:0] p28_array_index_1082038_comb;
  wire [7:0] p28_array_index_1082039_comb;
  wire [7:0] p28_array_index_1082041_comb;
  wire [7:0] p28_res7__144_comb;
  wire [7:0] p28_res7__560_comb;
  wire [7:0] p28_array_index_1081965_comb;
  wire [7:0] p28_array_index_1081966_comb;
  wire [7:0] p28_array_index_1081967_comb;
  wire [7:0] p28_array_index_1081968_comb;
  wire [7:0] p28_array_index_1081969_comb;
  wire [7:0] p28_array_index_1081970_comb;
  wire [7:0] p28_array_index_1082050_comb;
  wire [7:0] p28_array_index_1082051_comb;
  wire [7:0] p28_array_index_1082052_comb;
  wire [7:0] p28_array_index_1082053_comb;
  wire [7:0] p28_array_index_1082054_comb;
  wire [7:0] p28_array_index_1082055_comb;
  wire [7:0] p28_res7__145_comb;
  wire [7:0] p28_res7__561_comb;
  wire [7:0] p28_array_index_1081980_comb;
  wire [7:0] p28_array_index_1081981_comb;
  wire [7:0] p28_array_index_1081982_comb;
  wire [7:0] p28_array_index_1081983_comb;
  wire [7:0] p28_array_index_1081984_comb;
  wire [7:0] p28_array_index_1082065_comb;
  wire [7:0] p28_array_index_1082066_comb;
  wire [7:0] p28_array_index_1082067_comb;
  wire [7:0] p28_array_index_1082068_comb;
  wire [7:0] p28_array_index_1082069_comb;
  wire [7:0] p28_res7__146_comb;
  wire [7:0] p28_res7__562_comb;
  wire [7:0] p28_array_index_1081994_comb;
  wire [7:0] p28_array_index_1081995_comb;
  wire [7:0] p28_array_index_1081996_comb;
  wire [7:0] p28_array_index_1081997_comb;
  wire [7:0] p28_array_index_1081998_comb;
  wire [7:0] p28_array_index_1082079_comb;
  wire [7:0] p28_array_index_1082080_comb;
  wire [7:0] p28_array_index_1082081_comb;
  wire [7:0] p28_array_index_1082082_comb;
  wire [7:0] p28_array_index_1082083_comb;
  wire [7:0] p28_res7__147_comb;
  wire [7:0] p28_res7__563_comb;
  wire [7:0] p28_array_index_1082009_comb;
  wire [7:0] p28_array_index_1082010_comb;
  wire [7:0] p28_array_index_1082011_comb;
  wire [7:0] p28_array_index_1082012_comb;
  wire [7:0] p28_array_index_1082094_comb;
  wire [7:0] p28_array_index_1082095_comb;
  wire [7:0] p28_array_index_1082096_comb;
  wire [7:0] p28_array_index_1082097_comb;
  wire [7:0] p28_res7__148_comb;
  wire [7:0] p28_res7__564_comb;
  assign p28_addedKey__50_comb = p27_xor_1081801 ^ 128'h2ade_daf2_3e95_a23a_17b5_18a0_5e61_c10a;
  assign p28_array_index_1081932_comb = p27_arr[p28_addedKey__50_comb[127:120]];
  assign p28_array_index_1081933_comb = p27_arr[p28_addedKey__50_comb[119:112]];
  assign p28_array_index_1081934_comb = p27_arr[p28_addedKey__50_comb[111:104]];
  assign p28_array_index_1081935_comb = p27_arr[p28_addedKey__50_comb[103:96]];
  assign p28_array_index_1081936_comb = p27_arr[p28_addedKey__50_comb[95:88]];
  assign p28_array_index_1081937_comb = p27_arr[p28_addedKey__50_comb[87:80]];
  assign p28_array_index_1081939_comb = p27_arr[p28_addedKey__50_comb[71:64]];
  assign p28_array_index_1081941_comb = p27_arr[p28_addedKey__50_comb[55:48]];
  assign p28_array_index_1081942_comb = p27_arr[p28_addedKey__50_comb[47:40]];
  assign p28_array_index_1081943_comb = p27_arr[p28_addedKey__50_comb[39:32]];
  assign p28_array_index_1081944_comb = p27_arr[p28_addedKey__50_comb[31:24]];
  assign p28_array_index_1081945_comb = p27_arr[p28_addedKey__50_comb[23:16]];
  assign p28_array_index_1081946_comb = p27_arr[p28_addedKey__50_comb[15:8]];
  assign p28_array_index_1082020_comb = p27_arr[p27_bit_slice_1081849];
  assign p28_array_index_1082021_comb = p27_arr[p27_bit_slice_1081850];
  assign p28_array_index_1082022_comb = p27_arr[p27_bit_slice_1081851];
  assign p28_array_index_1082023_comb = p27_arr[p27_bit_slice_1081852];
  assign p28_array_index_1082024_comb = p27_arr[p27_bit_slice_1081853];
  assign p28_array_index_1082025_comb = p27_arr[p27_bit_slice_1081854];
  assign p28_array_index_1082026_comb = p27_arr[p27_bit_slice_1081855];
  assign p28_array_index_1082027_comb = p27_arr[p27_bit_slice_1081856];
  assign p28_array_index_1082028_comb = p27_arr[p27_bit_slice_1081857];
  assign p28_array_index_1082029_comb = p27_arr[p27_bit_slice_1081858];
  assign p28_array_index_1082030_comb = p27_arr[p27_bit_slice_1081859];
  assign p28_array_index_1082031_comb = p27_arr[p27_bit_slice_1081860];
  assign p28_array_index_1082032_comb = p27_arr[p27_bit_slice_1081861];
  assign p28_array_index_1081948_comb = p27_literal_1076345[p28_array_index_1081932_comb];
  assign p28_array_index_1081949_comb = p27_literal_1076347[p28_array_index_1081933_comb];
  assign p28_array_index_1081950_comb = p27_literal_1076349[p28_array_index_1081934_comb];
  assign p28_array_index_1081951_comb = p27_literal_1076351[p28_array_index_1081935_comb];
  assign p28_array_index_1081952_comb = p27_literal_1076353[p28_array_index_1081936_comb];
  assign p28_array_index_1081953_comb = p27_literal_1076355[p28_array_index_1081937_comb];
  assign p28_array_index_1081954_comb = p27_arr[p28_addedKey__50_comb[79:72]];
  assign p28_array_index_1081956_comb = p27_arr[p28_addedKey__50_comb[63:56]];
  assign p28_array_index_1082033_comb = p27_literal_1076345[p28_array_index_1082020_comb];
  assign p28_array_index_1082034_comb = p27_literal_1076347[p28_array_index_1082021_comb];
  assign p28_array_index_1082035_comb = p27_literal_1076349[p28_array_index_1082022_comb];
  assign p28_array_index_1082036_comb = p27_literal_1076351[p28_array_index_1082023_comb];
  assign p28_array_index_1082037_comb = p27_literal_1076353[p28_array_index_1082024_comb];
  assign p28_array_index_1082038_comb = p27_literal_1076355[p28_array_index_1082025_comb];
  assign p28_array_index_1082039_comb = p27_arr[p27_bit_slice_1081862];
  assign p28_array_index_1082041_comb = p27_arr[p27_bit_slice_1081863];
  assign p28_res7__144_comb = p28_array_index_1081948_comb ^ p28_array_index_1081949_comb ^ p28_array_index_1081950_comb ^ p28_array_index_1081951_comb ^ p28_array_index_1081952_comb ^ p28_array_index_1081953_comb ^ p28_array_index_1081954_comb ^ p27_literal_1076358[p28_array_index_1081939_comb] ^ p28_array_index_1081956_comb ^ p27_literal_1076355[p28_array_index_1081941_comb] ^ p27_literal_1076353[p28_array_index_1081942_comb] ^ p27_literal_1076351[p28_array_index_1081943_comb] ^ p27_literal_1076349[p28_array_index_1081944_comb] ^ p27_literal_1076347[p28_array_index_1081945_comb] ^ p27_literal_1076345[p28_array_index_1081946_comb] ^ p27_arr[p28_addedKey__50_comb[7:0]];
  assign p28_res7__560_comb = p28_array_index_1082033_comb ^ p28_array_index_1082034_comb ^ p28_array_index_1082035_comb ^ p28_array_index_1082036_comb ^ p28_array_index_1082037_comb ^ p28_array_index_1082038_comb ^ p28_array_index_1082039_comb ^ p27_literal_1076358[p28_array_index_1082026_comb] ^ p28_array_index_1082041_comb ^ p27_literal_1076355[p28_array_index_1082027_comb] ^ p27_literal_1076353[p28_array_index_1082028_comb] ^ p27_literal_1076351[p28_array_index_1082029_comb] ^ p27_literal_1076349[p28_array_index_1082030_comb] ^ p27_literal_1076347[p28_array_index_1082031_comb] ^ p27_literal_1076345[p28_array_index_1082032_comb] ^ p27_arr[p27_bit_slice_1081864];
  assign p28_array_index_1081965_comb = p27_literal_1076345[p28_res7__144_comb];
  assign p28_array_index_1081966_comb = p27_literal_1076347[p28_array_index_1081932_comb];
  assign p28_array_index_1081967_comb = p27_literal_1076349[p28_array_index_1081933_comb];
  assign p28_array_index_1081968_comb = p27_literal_1076351[p28_array_index_1081934_comb];
  assign p28_array_index_1081969_comb = p27_literal_1076353[p28_array_index_1081935_comb];
  assign p28_array_index_1081970_comb = p27_literal_1076355[p28_array_index_1081936_comb];
  assign p28_array_index_1082050_comb = p27_literal_1076345[p28_res7__560_comb];
  assign p28_array_index_1082051_comb = p27_literal_1076347[p28_array_index_1082020_comb];
  assign p28_array_index_1082052_comb = p27_literal_1076349[p28_array_index_1082021_comb];
  assign p28_array_index_1082053_comb = p27_literal_1076351[p28_array_index_1082022_comb];
  assign p28_array_index_1082054_comb = p27_literal_1076353[p28_array_index_1082023_comb];
  assign p28_array_index_1082055_comb = p27_literal_1076355[p28_array_index_1082024_comb];
  assign p28_res7__145_comb = p28_array_index_1081965_comb ^ p28_array_index_1081966_comb ^ p28_array_index_1081967_comb ^ p28_array_index_1081968_comb ^ p28_array_index_1081969_comb ^ p28_array_index_1081970_comb ^ p28_array_index_1081937_comb ^ p27_literal_1076358[p28_array_index_1081954_comb] ^ p28_array_index_1081939_comb ^ p27_literal_1076355[p28_array_index_1081956_comb] ^ p27_literal_1076353[p28_array_index_1081941_comb] ^ p27_literal_1076351[p28_array_index_1081942_comb] ^ p27_literal_1076349[p28_array_index_1081943_comb] ^ p27_literal_1076347[p28_array_index_1081944_comb] ^ p27_literal_1076345[p28_array_index_1081945_comb] ^ p28_array_index_1081946_comb;
  assign p28_res7__561_comb = p28_array_index_1082050_comb ^ p28_array_index_1082051_comb ^ p28_array_index_1082052_comb ^ p28_array_index_1082053_comb ^ p28_array_index_1082054_comb ^ p28_array_index_1082055_comb ^ p28_array_index_1082025_comb ^ p27_literal_1076358[p28_array_index_1082039_comb] ^ p28_array_index_1082026_comb ^ p27_literal_1076355[p28_array_index_1082041_comb] ^ p27_literal_1076353[p28_array_index_1082027_comb] ^ p27_literal_1076351[p28_array_index_1082028_comb] ^ p27_literal_1076349[p28_array_index_1082029_comb] ^ p27_literal_1076347[p28_array_index_1082030_comb] ^ p27_literal_1076345[p28_array_index_1082031_comb] ^ p28_array_index_1082032_comb;
  assign p28_array_index_1081980_comb = p27_literal_1076347[p28_res7__144_comb];
  assign p28_array_index_1081981_comb = p27_literal_1076349[p28_array_index_1081932_comb];
  assign p28_array_index_1081982_comb = p27_literal_1076351[p28_array_index_1081933_comb];
  assign p28_array_index_1081983_comb = p27_literal_1076353[p28_array_index_1081934_comb];
  assign p28_array_index_1081984_comb = p27_literal_1076355[p28_array_index_1081935_comb];
  assign p28_array_index_1082065_comb = p27_literal_1076347[p28_res7__560_comb];
  assign p28_array_index_1082066_comb = p27_literal_1076349[p28_array_index_1082020_comb];
  assign p28_array_index_1082067_comb = p27_literal_1076351[p28_array_index_1082021_comb];
  assign p28_array_index_1082068_comb = p27_literal_1076353[p28_array_index_1082022_comb];
  assign p28_array_index_1082069_comb = p27_literal_1076355[p28_array_index_1082023_comb];
  assign p28_res7__146_comb = p27_literal_1076345[p28_res7__145_comb] ^ p28_array_index_1081980_comb ^ p28_array_index_1081981_comb ^ p28_array_index_1081982_comb ^ p28_array_index_1081983_comb ^ p28_array_index_1081984_comb ^ p28_array_index_1081936_comb ^ p27_literal_1076358[p28_array_index_1081937_comb] ^ p28_array_index_1081954_comb ^ p27_literal_1076355[p28_array_index_1081939_comb] ^ p27_literal_1076353[p28_array_index_1081956_comb] ^ p27_literal_1076351[p28_array_index_1081941_comb] ^ p27_literal_1076349[p28_array_index_1081942_comb] ^ p27_literal_1076347[p28_array_index_1081943_comb] ^ p27_literal_1076345[p28_array_index_1081944_comb] ^ p28_array_index_1081945_comb;
  assign p28_res7__562_comb = p27_literal_1076345[p28_res7__561_comb] ^ p28_array_index_1082065_comb ^ p28_array_index_1082066_comb ^ p28_array_index_1082067_comb ^ p28_array_index_1082068_comb ^ p28_array_index_1082069_comb ^ p28_array_index_1082024_comb ^ p27_literal_1076358[p28_array_index_1082025_comb] ^ p28_array_index_1082039_comb ^ p27_literal_1076355[p28_array_index_1082026_comb] ^ p27_literal_1076353[p28_array_index_1082041_comb] ^ p27_literal_1076351[p28_array_index_1082027_comb] ^ p27_literal_1076349[p28_array_index_1082028_comb] ^ p27_literal_1076347[p28_array_index_1082029_comb] ^ p27_literal_1076345[p28_array_index_1082030_comb] ^ p28_array_index_1082031_comb;
  assign p28_array_index_1081994_comb = p27_literal_1076347[p28_res7__145_comb];
  assign p28_array_index_1081995_comb = p27_literal_1076349[p28_res7__144_comb];
  assign p28_array_index_1081996_comb = p27_literal_1076351[p28_array_index_1081932_comb];
  assign p28_array_index_1081997_comb = p27_literal_1076353[p28_array_index_1081933_comb];
  assign p28_array_index_1081998_comb = p27_literal_1076355[p28_array_index_1081934_comb];
  assign p28_array_index_1082079_comb = p27_literal_1076347[p28_res7__561_comb];
  assign p28_array_index_1082080_comb = p27_literal_1076349[p28_res7__560_comb];
  assign p28_array_index_1082081_comb = p27_literal_1076351[p28_array_index_1082020_comb];
  assign p28_array_index_1082082_comb = p27_literal_1076353[p28_array_index_1082021_comb];
  assign p28_array_index_1082083_comb = p27_literal_1076355[p28_array_index_1082022_comb];
  assign p28_res7__147_comb = p27_literal_1076345[p28_res7__146_comb] ^ p28_array_index_1081994_comb ^ p28_array_index_1081995_comb ^ p28_array_index_1081996_comb ^ p28_array_index_1081997_comb ^ p28_array_index_1081998_comb ^ p28_array_index_1081935_comb ^ p27_literal_1076358[p28_array_index_1081936_comb] ^ p28_array_index_1081937_comb ^ p27_literal_1076355[p28_array_index_1081954_comb] ^ p27_literal_1076353[p28_array_index_1081939_comb] ^ p27_literal_1076351[p28_array_index_1081956_comb] ^ p27_literal_1076349[p28_array_index_1081941_comb] ^ p27_literal_1076347[p28_array_index_1081942_comb] ^ p27_literal_1076345[p28_array_index_1081943_comb] ^ p28_array_index_1081944_comb;
  assign p28_res7__563_comb = p27_literal_1076345[p28_res7__562_comb] ^ p28_array_index_1082079_comb ^ p28_array_index_1082080_comb ^ p28_array_index_1082081_comb ^ p28_array_index_1082082_comb ^ p28_array_index_1082083_comb ^ p28_array_index_1082023_comb ^ p27_literal_1076358[p28_array_index_1082024_comb] ^ p28_array_index_1082025_comb ^ p27_literal_1076355[p28_array_index_1082039_comb] ^ p27_literal_1076353[p28_array_index_1082026_comb] ^ p27_literal_1076351[p28_array_index_1082041_comb] ^ p27_literal_1076349[p28_array_index_1082027_comb] ^ p27_literal_1076347[p28_array_index_1082028_comb] ^ p27_literal_1076345[p28_array_index_1082029_comb] ^ p28_array_index_1082030_comb;
  assign p28_array_index_1082009_comb = p27_literal_1076349[p28_res7__145_comb];
  assign p28_array_index_1082010_comb = p27_literal_1076351[p28_res7__144_comb];
  assign p28_array_index_1082011_comb = p27_literal_1076353[p28_array_index_1081932_comb];
  assign p28_array_index_1082012_comb = p27_literal_1076355[p28_array_index_1081933_comb];
  assign p28_array_index_1082094_comb = p27_literal_1076349[p28_res7__561_comb];
  assign p28_array_index_1082095_comb = p27_literal_1076351[p28_res7__560_comb];
  assign p28_array_index_1082096_comb = p27_literal_1076353[p28_array_index_1082020_comb];
  assign p28_array_index_1082097_comb = p27_literal_1076355[p28_array_index_1082021_comb];
  assign p28_res7__148_comb = p27_literal_1076345[p28_res7__147_comb] ^ p27_literal_1076347[p28_res7__146_comb] ^ p28_array_index_1082009_comb ^ p28_array_index_1082010_comb ^ p28_array_index_1082011_comb ^ p28_array_index_1082012_comb ^ p28_array_index_1081934_comb ^ p27_literal_1076358[p28_array_index_1081935_comb] ^ p28_array_index_1081936_comb ^ p28_array_index_1081953_comb ^ p27_literal_1076353[p28_array_index_1081954_comb] ^ p27_literal_1076351[p28_array_index_1081939_comb] ^ p27_literal_1076349[p28_array_index_1081956_comb] ^ p27_literal_1076347[p28_array_index_1081941_comb] ^ p27_literal_1076345[p28_array_index_1081942_comb] ^ p28_array_index_1081943_comb;
  assign p28_res7__564_comb = p27_literal_1076345[p28_res7__563_comb] ^ p27_literal_1076347[p28_res7__562_comb] ^ p28_array_index_1082094_comb ^ p28_array_index_1082095_comb ^ p28_array_index_1082096_comb ^ p28_array_index_1082097_comb ^ p28_array_index_1082022_comb ^ p27_literal_1076358[p28_array_index_1082023_comb] ^ p28_array_index_1082024_comb ^ p28_array_index_1082038_comb ^ p27_literal_1076353[p28_array_index_1082039_comb] ^ p27_literal_1076351[p28_array_index_1082026_comb] ^ p27_literal_1076349[p28_array_index_1082041_comb] ^ p27_literal_1076347[p28_array_index_1082027_comb] ^ p27_literal_1076345[p28_array_index_1082028_comb] ^ p28_array_index_1082029_comb;

  // Registers for pipe stage 28:
  reg [127:0] p28_k2;
  reg [127:0] p28_xor_1081801;
  reg [7:0] p28_array_index_1081932;
  reg [7:0] p28_array_index_1081933;
  reg [7:0] p28_array_index_1081934;
  reg [7:0] p28_array_index_1081935;
  reg [7:0] p28_array_index_1081936;
  reg [7:0] p28_array_index_1081937;
  reg [7:0] p28_array_index_1081939;
  reg [7:0] p28_array_index_1081941;
  reg [7:0] p28_array_index_1081942;
  reg [7:0] p28_array_index_1081948;
  reg [7:0] p28_array_index_1081949;
  reg [7:0] p28_array_index_1081950;
  reg [7:0] p28_array_index_1081951;
  reg [7:0] p28_array_index_1081952;
  reg [7:0] p28_array_index_1081954;
  reg [7:0] p28_array_index_1081956;
  reg [7:0] p28_res7__144;
  reg [7:0] p28_array_index_1081965;
  reg [7:0] p28_array_index_1081966;
  reg [7:0] p28_array_index_1081967;
  reg [7:0] p28_array_index_1081968;
  reg [7:0] p28_array_index_1081969;
  reg [7:0] p28_array_index_1081970;
  reg [7:0] p28_res7__145;
  reg [7:0] p28_array_index_1081980;
  reg [7:0] p28_array_index_1081981;
  reg [7:0] p28_array_index_1081982;
  reg [7:0] p28_array_index_1081983;
  reg [7:0] p28_array_index_1081984;
  reg [7:0] p28_res7__146;
  reg [7:0] p28_array_index_1081994;
  reg [7:0] p28_array_index_1081995;
  reg [7:0] p28_array_index_1081996;
  reg [7:0] p28_array_index_1081997;
  reg [7:0] p28_array_index_1081998;
  reg [7:0] p28_res7__147;
  reg [7:0] p28_array_index_1082009;
  reg [7:0] p28_array_index_1082010;
  reg [7:0] p28_array_index_1082011;
  reg [7:0] p28_array_index_1082012;
  reg [7:0] p28_res7__148;
  reg [7:0] p28_array_index_1082020;
  reg [7:0] p28_array_index_1082021;
  reg [7:0] p28_array_index_1082022;
  reg [7:0] p28_array_index_1082023;
  reg [7:0] p28_array_index_1082024;
  reg [7:0] p28_array_index_1082025;
  reg [7:0] p28_array_index_1082026;
  reg [7:0] p28_array_index_1082027;
  reg [7:0] p28_array_index_1082028;
  reg [7:0] p28_array_index_1082033;
  reg [7:0] p28_array_index_1082034;
  reg [7:0] p28_array_index_1082035;
  reg [7:0] p28_array_index_1082036;
  reg [7:0] p28_array_index_1082037;
  reg [7:0] p28_array_index_1082039;
  reg [7:0] p28_array_index_1082041;
  reg [7:0] p28_res7__560;
  reg [7:0] p28_array_index_1082050;
  reg [7:0] p28_array_index_1082051;
  reg [7:0] p28_array_index_1082052;
  reg [7:0] p28_array_index_1082053;
  reg [7:0] p28_array_index_1082054;
  reg [7:0] p28_array_index_1082055;
  reg [7:0] p28_res7__561;
  reg [7:0] p28_array_index_1082065;
  reg [7:0] p28_array_index_1082066;
  reg [7:0] p28_array_index_1082067;
  reg [7:0] p28_array_index_1082068;
  reg [7:0] p28_array_index_1082069;
  reg [7:0] p28_res7__562;
  reg [7:0] p28_array_index_1082079;
  reg [7:0] p28_array_index_1082080;
  reg [7:0] p28_array_index_1082081;
  reg [7:0] p28_array_index_1082082;
  reg [7:0] p28_array_index_1082083;
  reg [7:0] p28_res7__563;
  reg [7:0] p28_array_index_1082094;
  reg [7:0] p28_array_index_1082095;
  reg [7:0] p28_array_index_1082096;
  reg [7:0] p28_array_index_1082097;
  reg [7:0] p28_res7__564;
  reg [7:0] p29_arr[256];
  reg [7:0] p29_literal_1076345[256];
  reg [7:0] p29_literal_1076347[256];
  reg [7:0] p29_literal_1076349[256];
  reg [7:0] p29_literal_1076351[256];
  reg [7:0] p29_literal_1076353[256];
  reg [7:0] p29_literal_1076355[256];
  reg [7:0] p29_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p28_k2 <= p27_k2;
    p28_xor_1081801 <= p27_xor_1081801;
    p28_array_index_1081932 <= p28_array_index_1081932_comb;
    p28_array_index_1081933 <= p28_array_index_1081933_comb;
    p28_array_index_1081934 <= p28_array_index_1081934_comb;
    p28_array_index_1081935 <= p28_array_index_1081935_comb;
    p28_array_index_1081936 <= p28_array_index_1081936_comb;
    p28_array_index_1081937 <= p28_array_index_1081937_comb;
    p28_array_index_1081939 <= p28_array_index_1081939_comb;
    p28_array_index_1081941 <= p28_array_index_1081941_comb;
    p28_array_index_1081942 <= p28_array_index_1081942_comb;
    p28_array_index_1081948 <= p28_array_index_1081948_comb;
    p28_array_index_1081949 <= p28_array_index_1081949_comb;
    p28_array_index_1081950 <= p28_array_index_1081950_comb;
    p28_array_index_1081951 <= p28_array_index_1081951_comb;
    p28_array_index_1081952 <= p28_array_index_1081952_comb;
    p28_array_index_1081954 <= p28_array_index_1081954_comb;
    p28_array_index_1081956 <= p28_array_index_1081956_comb;
    p28_res7__144 <= p28_res7__144_comb;
    p28_array_index_1081965 <= p28_array_index_1081965_comb;
    p28_array_index_1081966 <= p28_array_index_1081966_comb;
    p28_array_index_1081967 <= p28_array_index_1081967_comb;
    p28_array_index_1081968 <= p28_array_index_1081968_comb;
    p28_array_index_1081969 <= p28_array_index_1081969_comb;
    p28_array_index_1081970 <= p28_array_index_1081970_comb;
    p28_res7__145 <= p28_res7__145_comb;
    p28_array_index_1081980 <= p28_array_index_1081980_comb;
    p28_array_index_1081981 <= p28_array_index_1081981_comb;
    p28_array_index_1081982 <= p28_array_index_1081982_comb;
    p28_array_index_1081983 <= p28_array_index_1081983_comb;
    p28_array_index_1081984 <= p28_array_index_1081984_comb;
    p28_res7__146 <= p28_res7__146_comb;
    p28_array_index_1081994 <= p28_array_index_1081994_comb;
    p28_array_index_1081995 <= p28_array_index_1081995_comb;
    p28_array_index_1081996 <= p28_array_index_1081996_comb;
    p28_array_index_1081997 <= p28_array_index_1081997_comb;
    p28_array_index_1081998 <= p28_array_index_1081998_comb;
    p28_res7__147 <= p28_res7__147_comb;
    p28_array_index_1082009 <= p28_array_index_1082009_comb;
    p28_array_index_1082010 <= p28_array_index_1082010_comb;
    p28_array_index_1082011 <= p28_array_index_1082011_comb;
    p28_array_index_1082012 <= p28_array_index_1082012_comb;
    p28_res7__148 <= p28_res7__148_comb;
    p28_array_index_1082020 <= p28_array_index_1082020_comb;
    p28_array_index_1082021 <= p28_array_index_1082021_comb;
    p28_array_index_1082022 <= p28_array_index_1082022_comb;
    p28_array_index_1082023 <= p28_array_index_1082023_comb;
    p28_array_index_1082024 <= p28_array_index_1082024_comb;
    p28_array_index_1082025 <= p28_array_index_1082025_comb;
    p28_array_index_1082026 <= p28_array_index_1082026_comb;
    p28_array_index_1082027 <= p28_array_index_1082027_comb;
    p28_array_index_1082028 <= p28_array_index_1082028_comb;
    p28_array_index_1082033 <= p28_array_index_1082033_comb;
    p28_array_index_1082034 <= p28_array_index_1082034_comb;
    p28_array_index_1082035 <= p28_array_index_1082035_comb;
    p28_array_index_1082036 <= p28_array_index_1082036_comb;
    p28_array_index_1082037 <= p28_array_index_1082037_comb;
    p28_array_index_1082039 <= p28_array_index_1082039_comb;
    p28_array_index_1082041 <= p28_array_index_1082041_comb;
    p28_res7__560 <= p28_res7__560_comb;
    p28_array_index_1082050 <= p28_array_index_1082050_comb;
    p28_array_index_1082051 <= p28_array_index_1082051_comb;
    p28_array_index_1082052 <= p28_array_index_1082052_comb;
    p28_array_index_1082053 <= p28_array_index_1082053_comb;
    p28_array_index_1082054 <= p28_array_index_1082054_comb;
    p28_array_index_1082055 <= p28_array_index_1082055_comb;
    p28_res7__561 <= p28_res7__561_comb;
    p28_array_index_1082065 <= p28_array_index_1082065_comb;
    p28_array_index_1082066 <= p28_array_index_1082066_comb;
    p28_array_index_1082067 <= p28_array_index_1082067_comb;
    p28_array_index_1082068 <= p28_array_index_1082068_comb;
    p28_array_index_1082069 <= p28_array_index_1082069_comb;
    p28_res7__562 <= p28_res7__562_comb;
    p28_array_index_1082079 <= p28_array_index_1082079_comb;
    p28_array_index_1082080 <= p28_array_index_1082080_comb;
    p28_array_index_1082081 <= p28_array_index_1082081_comb;
    p28_array_index_1082082 <= p28_array_index_1082082_comb;
    p28_array_index_1082083 <= p28_array_index_1082083_comb;
    p28_res7__563 <= p28_res7__563_comb;
    p28_array_index_1082094 <= p28_array_index_1082094_comb;
    p28_array_index_1082095 <= p28_array_index_1082095_comb;
    p28_array_index_1082096 <= p28_array_index_1082096_comb;
    p28_array_index_1082097 <= p28_array_index_1082097_comb;
    p28_res7__564 <= p28_res7__564_comb;
    p29_arr <= p28_arr;
    p29_literal_1076345 <= p28_literal_1076345;
    p29_literal_1076347 <= p28_literal_1076347;
    p29_literal_1076349 <= p28_literal_1076349;
    p29_literal_1076351 <= p28_literal_1076351;
    p29_literal_1076353 <= p28_literal_1076353;
    p29_literal_1076355 <= p28_literal_1076355;
    p29_literal_1076358 <= p28_literal_1076358;
  end

  // ===== Pipe stage 29:
  wire [7:0] p29_array_index_1082291_comb;
  wire [7:0] p29_array_index_1082292_comb;
  wire [7:0] p29_array_index_1082293_comb;
  wire [7:0] p29_array_index_1082294_comb;
  wire [7:0] p29_res7__149_comb;
  wire [7:0] p29_array_index_1082359_comb;
  wire [7:0] p29_array_index_1082360_comb;
  wire [7:0] p29_array_index_1082361_comb;
  wire [7:0] p29_array_index_1082362_comb;
  wire [7:0] p29_array_index_1082305_comb;
  wire [7:0] p29_array_index_1082306_comb;
  wire [7:0] p29_array_index_1082307_comb;
  wire [7:0] p29_res7__565_comb;
  wire [7:0] p29_res7__150_comb;
  wire [7:0] p29_array_index_1082373_comb;
  wire [7:0] p29_array_index_1082374_comb;
  wire [7:0] p29_array_index_1082375_comb;
  wire [7:0] p29_array_index_1082317_comb;
  wire [7:0] p29_array_index_1082318_comb;
  wire [7:0] p29_array_index_1082319_comb;
  wire [7:0] p29_res7__566_comb;
  wire [7:0] p29_res7__151_comb;
  wire [7:0] p29_array_index_1082385_comb;
  wire [7:0] p29_array_index_1082386_comb;
  wire [7:0] p29_array_index_1082387_comb;
  wire [7:0] p29_array_index_1082330_comb;
  wire [7:0] p29_array_index_1082331_comb;
  wire [7:0] p29_res7__567_comb;
  wire [7:0] p29_res7__152_comb;
  wire [7:0] p29_array_index_1082398_comb;
  wire [7:0] p29_array_index_1082399_comb;
  wire [7:0] p29_array_index_1082341_comb;
  wire [7:0] p29_array_index_1082342_comb;
  wire [7:0] p29_res7__568_comb;
  wire [7:0] p29_res7__153_comb;
  wire [7:0] p29_array_index_1082409_comb;
  wire [7:0] p29_array_index_1082410_comb;
  wire [7:0] p29_array_index_1082348_comb;
  wire [7:0] p29_array_index_1082349_comb;
  wire [7:0] p29_array_index_1082350_comb;
  wire [7:0] p29_array_index_1082351_comb;
  wire [7:0] p29_array_index_1082352_comb;
  wire [7:0] p29_array_index_1082353_comb;
  wire [7:0] p29_array_index_1082354_comb;
  wire [7:0] p29_array_index_1082355_comb;
  wire [7:0] p29_array_index_1082356_comb;
  wire [7:0] p29_res7__569_comb;
  assign p29_array_index_1082291_comb = p28_literal_1076349[p28_res7__146];
  assign p29_array_index_1082292_comb = p28_literal_1076351[p28_res7__145];
  assign p29_array_index_1082293_comb = p28_literal_1076353[p28_res7__144];
  assign p29_array_index_1082294_comb = p28_literal_1076355[p28_array_index_1081932];
  assign p29_res7__149_comb = p28_literal_1076345[p28_res7__148] ^ p28_literal_1076347[p28_res7__147] ^ p29_array_index_1082291_comb ^ p29_array_index_1082292_comb ^ p29_array_index_1082293_comb ^ p29_array_index_1082294_comb ^ p28_array_index_1081933 ^ p28_literal_1076358[p28_array_index_1081934] ^ p28_array_index_1081935 ^ p28_array_index_1081970 ^ p28_literal_1076353[p28_array_index_1081937] ^ p28_literal_1076351[p28_array_index_1081954] ^ p28_literal_1076349[p28_array_index_1081939] ^ p28_literal_1076347[p28_array_index_1081956] ^ p28_literal_1076345[p28_array_index_1081941] ^ p28_array_index_1081942;
  assign p29_array_index_1082359_comb = p28_literal_1076349[p28_res7__562];
  assign p29_array_index_1082360_comb = p28_literal_1076351[p28_res7__561];
  assign p29_array_index_1082361_comb = p28_literal_1076353[p28_res7__560];
  assign p29_array_index_1082362_comb = p28_literal_1076355[p28_array_index_1082020];
  assign p29_array_index_1082305_comb = p28_literal_1076351[p28_res7__146];
  assign p29_array_index_1082306_comb = p28_literal_1076353[p28_res7__145];
  assign p29_array_index_1082307_comb = p28_literal_1076355[p28_res7__144];
  assign p29_res7__565_comb = p28_literal_1076345[p28_res7__564] ^ p28_literal_1076347[p28_res7__563] ^ p29_array_index_1082359_comb ^ p29_array_index_1082360_comb ^ p29_array_index_1082361_comb ^ p29_array_index_1082362_comb ^ p28_array_index_1082021 ^ p28_literal_1076358[p28_array_index_1082022] ^ p28_array_index_1082023 ^ p28_array_index_1082055 ^ p28_literal_1076353[p28_array_index_1082025] ^ p28_literal_1076351[p28_array_index_1082039] ^ p28_literal_1076349[p28_array_index_1082026] ^ p28_literal_1076347[p28_array_index_1082041] ^ p28_literal_1076345[p28_array_index_1082027] ^ p28_array_index_1082028;
  assign p29_res7__150_comb = p28_literal_1076345[p29_res7__149_comb] ^ p28_literal_1076347[p28_res7__148] ^ p28_literal_1076349[p28_res7__147] ^ p29_array_index_1082305_comb ^ p29_array_index_1082306_comb ^ p29_array_index_1082307_comb ^ p28_array_index_1081932 ^ p28_literal_1076358[p28_array_index_1081933] ^ p28_array_index_1081934 ^ p28_array_index_1081984 ^ p28_array_index_1081952 ^ p28_literal_1076351[p28_array_index_1081937] ^ p28_literal_1076349[p28_array_index_1081954] ^ p28_literal_1076347[p28_array_index_1081939] ^ p28_literal_1076345[p28_array_index_1081956] ^ p28_array_index_1081941;
  assign p29_array_index_1082373_comb = p28_literal_1076351[p28_res7__562];
  assign p29_array_index_1082374_comb = p28_literal_1076353[p28_res7__561];
  assign p29_array_index_1082375_comb = p28_literal_1076355[p28_res7__560];
  assign p29_array_index_1082317_comb = p28_literal_1076351[p28_res7__147];
  assign p29_array_index_1082318_comb = p28_literal_1076353[p28_res7__146];
  assign p29_array_index_1082319_comb = p28_literal_1076355[p28_res7__145];
  assign p29_res7__566_comb = p28_literal_1076345[p29_res7__565_comb] ^ p28_literal_1076347[p28_res7__564] ^ p28_literal_1076349[p28_res7__563] ^ p29_array_index_1082373_comb ^ p29_array_index_1082374_comb ^ p29_array_index_1082375_comb ^ p28_array_index_1082020 ^ p28_literal_1076358[p28_array_index_1082021] ^ p28_array_index_1082022 ^ p28_array_index_1082069 ^ p28_array_index_1082037 ^ p28_literal_1076351[p28_array_index_1082025] ^ p28_literal_1076349[p28_array_index_1082039] ^ p28_literal_1076347[p28_array_index_1082026] ^ p28_literal_1076345[p28_array_index_1082041] ^ p28_array_index_1082027;
  assign p29_res7__151_comb = p28_literal_1076345[p29_res7__150_comb] ^ p28_literal_1076347[p29_res7__149_comb] ^ p28_literal_1076349[p28_res7__148] ^ p29_array_index_1082317_comb ^ p29_array_index_1082318_comb ^ p29_array_index_1082319_comb ^ p28_res7__144 ^ p28_literal_1076358[p28_array_index_1081932] ^ p28_array_index_1081933 ^ p28_array_index_1081998 ^ p28_array_index_1081969 ^ p28_literal_1076351[p28_array_index_1081936] ^ p28_literal_1076349[p28_array_index_1081937] ^ p28_literal_1076347[p28_array_index_1081954] ^ p28_literal_1076345[p28_array_index_1081939] ^ p28_array_index_1081956;
  assign p29_array_index_1082385_comb = p28_literal_1076351[p28_res7__563];
  assign p29_array_index_1082386_comb = p28_literal_1076353[p28_res7__562];
  assign p29_array_index_1082387_comb = p28_literal_1076355[p28_res7__561];
  assign p29_array_index_1082330_comb = p28_literal_1076353[p28_res7__147];
  assign p29_array_index_1082331_comb = p28_literal_1076355[p28_res7__146];
  assign p29_res7__567_comb = p28_literal_1076345[p29_res7__566_comb] ^ p28_literal_1076347[p29_res7__565_comb] ^ p28_literal_1076349[p28_res7__564] ^ p29_array_index_1082385_comb ^ p29_array_index_1082386_comb ^ p29_array_index_1082387_comb ^ p28_res7__560 ^ p28_literal_1076358[p28_array_index_1082020] ^ p28_array_index_1082021 ^ p28_array_index_1082083 ^ p28_array_index_1082054 ^ p28_literal_1076351[p28_array_index_1082024] ^ p28_literal_1076349[p28_array_index_1082025] ^ p28_literal_1076347[p28_array_index_1082039] ^ p28_literal_1076345[p28_array_index_1082026] ^ p28_array_index_1082041;
  assign p29_res7__152_comb = p28_literal_1076345[p29_res7__151_comb] ^ p28_literal_1076347[p29_res7__150_comb] ^ p28_literal_1076349[p29_res7__149_comb] ^ p28_literal_1076351[p28_res7__148] ^ p29_array_index_1082330_comb ^ p29_array_index_1082331_comb ^ p28_res7__145 ^ p28_literal_1076358[p28_res7__144] ^ p28_array_index_1081932 ^ p28_array_index_1082012 ^ p28_array_index_1081983 ^ p28_array_index_1081951 ^ p28_literal_1076349[p28_array_index_1081936] ^ p28_literal_1076347[p28_array_index_1081937] ^ p28_literal_1076345[p28_array_index_1081954] ^ p28_array_index_1081939;
  assign p29_array_index_1082398_comb = p28_literal_1076353[p28_res7__563];
  assign p29_array_index_1082399_comb = p28_literal_1076355[p28_res7__562];
  assign p29_array_index_1082341_comb = p28_literal_1076353[p28_res7__148];
  assign p29_array_index_1082342_comb = p28_literal_1076355[p28_res7__147];
  assign p29_res7__568_comb = p28_literal_1076345[p29_res7__567_comb] ^ p28_literal_1076347[p29_res7__566_comb] ^ p28_literal_1076349[p29_res7__565_comb] ^ p28_literal_1076351[p28_res7__564] ^ p29_array_index_1082398_comb ^ p29_array_index_1082399_comb ^ p28_res7__561 ^ p28_literal_1076358[p28_res7__560] ^ p28_array_index_1082020 ^ p28_array_index_1082097 ^ p28_array_index_1082068 ^ p28_array_index_1082036 ^ p28_literal_1076349[p28_array_index_1082024] ^ p28_literal_1076347[p28_array_index_1082025] ^ p28_literal_1076345[p28_array_index_1082039] ^ p28_array_index_1082026;
  assign p29_res7__153_comb = p28_literal_1076345[p29_res7__152_comb] ^ p28_literal_1076347[p29_res7__151_comb] ^ p28_literal_1076349[p29_res7__150_comb] ^ p28_literal_1076351[p29_res7__149_comb] ^ p29_array_index_1082341_comb ^ p29_array_index_1082342_comb ^ p28_res7__146 ^ p28_literal_1076358[p28_res7__145] ^ p28_res7__144 ^ p29_array_index_1082294_comb ^ p28_array_index_1081997 ^ p28_array_index_1081968 ^ p28_literal_1076349[p28_array_index_1081935] ^ p28_literal_1076347[p28_array_index_1081936] ^ p28_literal_1076345[p28_array_index_1081937] ^ p28_array_index_1081954;
  assign p29_array_index_1082409_comb = p28_literal_1076353[p28_res7__564];
  assign p29_array_index_1082410_comb = p28_literal_1076355[p28_res7__563];
  assign p29_array_index_1082348_comb = p28_literal_1076345[p29_res7__153_comb];
  assign p29_array_index_1082349_comb = p28_literal_1076347[p29_res7__152_comb];
  assign p29_array_index_1082350_comb = p28_literal_1076349[p29_res7__151_comb];
  assign p29_array_index_1082351_comb = p28_literal_1076351[p29_res7__150_comb];
  assign p29_array_index_1082352_comb = p28_literal_1076353[p29_res7__149_comb];
  assign p29_array_index_1082353_comb = p28_literal_1076355[p28_res7__148];
  assign p29_array_index_1082354_comb = p28_literal_1076358[p28_res7__146];
  assign p29_array_index_1082355_comb = p28_literal_1076347[p28_array_index_1081935];
  assign p29_array_index_1082356_comb = p28_literal_1076345[p28_array_index_1081936];
  assign p29_res7__569_comb = p28_literal_1076345[p29_res7__568_comb] ^ p28_literal_1076347[p29_res7__567_comb] ^ p28_literal_1076349[p29_res7__566_comb] ^ p28_literal_1076351[p29_res7__565_comb] ^ p29_array_index_1082409_comb ^ p29_array_index_1082410_comb ^ p28_res7__562 ^ p28_literal_1076358[p28_res7__561] ^ p28_res7__560 ^ p29_array_index_1082362_comb ^ p28_array_index_1082082 ^ p28_array_index_1082053 ^ p28_literal_1076349[p28_array_index_1082023] ^ p28_literal_1076347[p28_array_index_1082024] ^ p28_literal_1076345[p28_array_index_1082025] ^ p28_array_index_1082039;

  // Registers for pipe stage 29:
  reg [127:0] p29_k2;
  reg [127:0] p29_xor_1081801;
  reg [7:0] p29_array_index_1081932;
  reg [7:0] p29_array_index_1081933;
  reg [7:0] p29_array_index_1081934;
  reg [7:0] p29_array_index_1081935;
  reg [7:0] p29_array_index_1081936;
  reg [7:0] p29_array_index_1081937;
  reg [7:0] p29_array_index_1081948;
  reg [7:0] p29_array_index_1081949;
  reg [7:0] p29_array_index_1081950;
  reg [7:0] p29_res7__144;
  reg [7:0] p29_array_index_1081965;
  reg [7:0] p29_array_index_1081966;
  reg [7:0] p29_array_index_1081967;
  reg [7:0] p29_res7__145;
  reg [7:0] p29_array_index_1081980;
  reg [7:0] p29_array_index_1081981;
  reg [7:0] p29_array_index_1081982;
  reg [7:0] p29_res7__146;
  reg [7:0] p29_array_index_1081994;
  reg [7:0] p29_array_index_1081995;
  reg [7:0] p29_array_index_1081996;
  reg [7:0] p29_res7__147;
  reg [7:0] p29_array_index_1082009;
  reg [7:0] p29_array_index_1082010;
  reg [7:0] p29_array_index_1082011;
  reg [7:0] p29_res7__148;
  reg [7:0] p29_array_index_1082291;
  reg [7:0] p29_array_index_1082292;
  reg [7:0] p29_array_index_1082293;
  reg [7:0] p29_res7__149;
  reg [7:0] p29_array_index_1082305;
  reg [7:0] p29_array_index_1082306;
  reg [7:0] p29_array_index_1082307;
  reg [7:0] p29_res7__150;
  reg [7:0] p29_array_index_1082317;
  reg [7:0] p29_array_index_1082318;
  reg [7:0] p29_array_index_1082319;
  reg [7:0] p29_res7__151;
  reg [7:0] p29_array_index_1082330;
  reg [7:0] p29_array_index_1082331;
  reg [7:0] p29_res7__152;
  reg [7:0] p29_array_index_1082341;
  reg [7:0] p29_array_index_1082342;
  reg [7:0] p29_res7__153;
  reg [7:0] p29_array_index_1082348;
  reg [7:0] p29_array_index_1082349;
  reg [7:0] p29_array_index_1082350;
  reg [7:0] p29_array_index_1082351;
  reg [7:0] p29_array_index_1082352;
  reg [7:0] p29_array_index_1082353;
  reg [7:0] p29_array_index_1082354;
  reg [7:0] p29_array_index_1082355;
  reg [7:0] p29_array_index_1082356;
  reg [7:0] p29_array_index_1082020;
  reg [7:0] p29_array_index_1082021;
  reg [7:0] p29_array_index_1082022;
  reg [7:0] p29_array_index_1082023;
  reg [7:0] p29_array_index_1082024;
  reg [7:0] p29_array_index_1082025;
  reg [7:0] p29_array_index_1082033;
  reg [7:0] p29_array_index_1082034;
  reg [7:0] p29_array_index_1082035;
  reg [7:0] p29_res7__560;
  reg [7:0] p29_array_index_1082050;
  reg [7:0] p29_array_index_1082051;
  reg [7:0] p29_array_index_1082052;
  reg [7:0] p29_res7__561;
  reg [7:0] p29_array_index_1082065;
  reg [7:0] p29_array_index_1082066;
  reg [7:0] p29_array_index_1082067;
  reg [7:0] p29_res7__562;
  reg [7:0] p29_array_index_1082079;
  reg [7:0] p29_array_index_1082080;
  reg [7:0] p29_array_index_1082081;
  reg [7:0] p29_res7__563;
  reg [7:0] p29_array_index_1082094;
  reg [7:0] p29_array_index_1082095;
  reg [7:0] p29_array_index_1082096;
  reg [7:0] p29_res7__564;
  reg [7:0] p29_array_index_1082359;
  reg [7:0] p29_array_index_1082360;
  reg [7:0] p29_array_index_1082361;
  reg [7:0] p29_res7__565;
  reg [7:0] p29_array_index_1082373;
  reg [7:0] p29_array_index_1082374;
  reg [7:0] p29_array_index_1082375;
  reg [7:0] p29_res7__566;
  reg [7:0] p29_array_index_1082385;
  reg [7:0] p29_array_index_1082386;
  reg [7:0] p29_array_index_1082387;
  reg [7:0] p29_res7__567;
  reg [7:0] p29_array_index_1082398;
  reg [7:0] p29_array_index_1082399;
  reg [7:0] p29_res7__568;
  reg [7:0] p29_array_index_1082409;
  reg [7:0] p29_array_index_1082410;
  reg [7:0] p29_res7__569;
  reg [7:0] p30_arr[256];
  reg [7:0] p30_literal_1076345[256];
  reg [7:0] p30_literal_1076347[256];
  reg [7:0] p30_literal_1076349[256];
  reg [7:0] p30_literal_1076351[256];
  reg [7:0] p30_literal_1076353[256];
  reg [7:0] p30_literal_1076355[256];
  reg [7:0] p30_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p29_k2 <= p28_k2;
    p29_xor_1081801 <= p28_xor_1081801;
    p29_array_index_1081932 <= p28_array_index_1081932;
    p29_array_index_1081933 <= p28_array_index_1081933;
    p29_array_index_1081934 <= p28_array_index_1081934;
    p29_array_index_1081935 <= p28_array_index_1081935;
    p29_array_index_1081936 <= p28_array_index_1081936;
    p29_array_index_1081937 <= p28_array_index_1081937;
    p29_array_index_1081948 <= p28_array_index_1081948;
    p29_array_index_1081949 <= p28_array_index_1081949;
    p29_array_index_1081950 <= p28_array_index_1081950;
    p29_res7__144 <= p28_res7__144;
    p29_array_index_1081965 <= p28_array_index_1081965;
    p29_array_index_1081966 <= p28_array_index_1081966;
    p29_array_index_1081967 <= p28_array_index_1081967;
    p29_res7__145 <= p28_res7__145;
    p29_array_index_1081980 <= p28_array_index_1081980;
    p29_array_index_1081981 <= p28_array_index_1081981;
    p29_array_index_1081982 <= p28_array_index_1081982;
    p29_res7__146 <= p28_res7__146;
    p29_array_index_1081994 <= p28_array_index_1081994;
    p29_array_index_1081995 <= p28_array_index_1081995;
    p29_array_index_1081996 <= p28_array_index_1081996;
    p29_res7__147 <= p28_res7__147;
    p29_array_index_1082009 <= p28_array_index_1082009;
    p29_array_index_1082010 <= p28_array_index_1082010;
    p29_array_index_1082011 <= p28_array_index_1082011;
    p29_res7__148 <= p28_res7__148;
    p29_array_index_1082291 <= p29_array_index_1082291_comb;
    p29_array_index_1082292 <= p29_array_index_1082292_comb;
    p29_array_index_1082293 <= p29_array_index_1082293_comb;
    p29_res7__149 <= p29_res7__149_comb;
    p29_array_index_1082305 <= p29_array_index_1082305_comb;
    p29_array_index_1082306 <= p29_array_index_1082306_comb;
    p29_array_index_1082307 <= p29_array_index_1082307_comb;
    p29_res7__150 <= p29_res7__150_comb;
    p29_array_index_1082317 <= p29_array_index_1082317_comb;
    p29_array_index_1082318 <= p29_array_index_1082318_comb;
    p29_array_index_1082319 <= p29_array_index_1082319_comb;
    p29_res7__151 <= p29_res7__151_comb;
    p29_array_index_1082330 <= p29_array_index_1082330_comb;
    p29_array_index_1082331 <= p29_array_index_1082331_comb;
    p29_res7__152 <= p29_res7__152_comb;
    p29_array_index_1082341 <= p29_array_index_1082341_comb;
    p29_array_index_1082342 <= p29_array_index_1082342_comb;
    p29_res7__153 <= p29_res7__153_comb;
    p29_array_index_1082348 <= p29_array_index_1082348_comb;
    p29_array_index_1082349 <= p29_array_index_1082349_comb;
    p29_array_index_1082350 <= p29_array_index_1082350_comb;
    p29_array_index_1082351 <= p29_array_index_1082351_comb;
    p29_array_index_1082352 <= p29_array_index_1082352_comb;
    p29_array_index_1082353 <= p29_array_index_1082353_comb;
    p29_array_index_1082354 <= p29_array_index_1082354_comb;
    p29_array_index_1082355 <= p29_array_index_1082355_comb;
    p29_array_index_1082356 <= p29_array_index_1082356_comb;
    p29_array_index_1082020 <= p28_array_index_1082020;
    p29_array_index_1082021 <= p28_array_index_1082021;
    p29_array_index_1082022 <= p28_array_index_1082022;
    p29_array_index_1082023 <= p28_array_index_1082023;
    p29_array_index_1082024 <= p28_array_index_1082024;
    p29_array_index_1082025 <= p28_array_index_1082025;
    p29_array_index_1082033 <= p28_array_index_1082033;
    p29_array_index_1082034 <= p28_array_index_1082034;
    p29_array_index_1082035 <= p28_array_index_1082035;
    p29_res7__560 <= p28_res7__560;
    p29_array_index_1082050 <= p28_array_index_1082050;
    p29_array_index_1082051 <= p28_array_index_1082051;
    p29_array_index_1082052 <= p28_array_index_1082052;
    p29_res7__561 <= p28_res7__561;
    p29_array_index_1082065 <= p28_array_index_1082065;
    p29_array_index_1082066 <= p28_array_index_1082066;
    p29_array_index_1082067 <= p28_array_index_1082067;
    p29_res7__562 <= p28_res7__562;
    p29_array_index_1082079 <= p28_array_index_1082079;
    p29_array_index_1082080 <= p28_array_index_1082080;
    p29_array_index_1082081 <= p28_array_index_1082081;
    p29_res7__563 <= p28_res7__563;
    p29_array_index_1082094 <= p28_array_index_1082094;
    p29_array_index_1082095 <= p28_array_index_1082095;
    p29_array_index_1082096 <= p28_array_index_1082096;
    p29_res7__564 <= p28_res7__564;
    p29_array_index_1082359 <= p29_array_index_1082359_comb;
    p29_array_index_1082360 <= p29_array_index_1082360_comb;
    p29_array_index_1082361 <= p29_array_index_1082361_comb;
    p29_res7__565 <= p29_res7__565_comb;
    p29_array_index_1082373 <= p29_array_index_1082373_comb;
    p29_array_index_1082374 <= p29_array_index_1082374_comb;
    p29_array_index_1082375 <= p29_array_index_1082375_comb;
    p29_res7__566 <= p29_res7__566_comb;
    p29_array_index_1082385 <= p29_array_index_1082385_comb;
    p29_array_index_1082386 <= p29_array_index_1082386_comb;
    p29_array_index_1082387 <= p29_array_index_1082387_comb;
    p29_res7__567 <= p29_res7__567_comb;
    p29_array_index_1082398 <= p29_array_index_1082398_comb;
    p29_array_index_1082399 <= p29_array_index_1082399_comb;
    p29_res7__568 <= p29_res7__568_comb;
    p29_array_index_1082409 <= p29_array_index_1082409_comb;
    p29_array_index_1082410 <= p29_array_index_1082410_comb;
    p29_res7__569 <= p29_res7__569_comb;
    p30_arr <= p29_arr;
    p30_literal_1076345 <= p29_literal_1076345;
    p30_literal_1076347 <= p29_literal_1076347;
    p30_literal_1076349 <= p29_literal_1076349;
    p30_literal_1076351 <= p29_literal_1076351;
    p30_literal_1076353 <= p29_literal_1076353;
    p30_literal_1076355 <= p29_literal_1076355;
    p30_literal_1076358 <= p29_literal_1076358;
  end

  // ===== Pipe stage 30:
  wire [7:0] p30_res7__154_comb;
  wire [7:0] p30_array_index_1082636_comb;
  wire [7:0] p30_res7__155_comb;
  wire [7:0] p30_array_index_1082682_comb;
  wire [7:0] p30_res7__156_comb;
  wire [7:0] p30_res7__570_comb;
  wire [7:0] p30_array_index_1082692_comb;
  wire [7:0] p30_res7__157_comb;
  wire [7:0] p30_res7__571_comb;
  wire [7:0] p30_res7__158_comb;
  wire [7:0] p30_res7__572_comb;
  wire [7:0] p30_res7__159_comb;
  wire [7:0] p30_res7__573_comb;
  wire [127:0] p30_res__9_comb;
  wire [127:0] p30_xor_1082676_comb;
  wire [7:0] p30_res7__574_comb;
  assign p30_res7__154_comb = p29_array_index_1082348 ^ p29_array_index_1082349 ^ p29_array_index_1082350 ^ p29_array_index_1082351 ^ p29_array_index_1082352 ^ p29_array_index_1082353 ^ p29_res7__147 ^ p29_array_index_1082354 ^ p29_res7__145 ^ p29_array_index_1082307 ^ p29_array_index_1082011 ^ p29_array_index_1081982 ^ p29_array_index_1081950 ^ p29_array_index_1082355 ^ p29_array_index_1082356 ^ p29_array_index_1081937;
  assign p30_array_index_1082636_comb = p29_literal_1076355[p29_res7__149];
  assign p30_res7__155_comb = p29_literal_1076345[p30_res7__154_comb] ^ p29_literal_1076347[p29_res7__153] ^ p29_literal_1076349[p29_res7__152] ^ p29_literal_1076351[p29_res7__151] ^ p29_literal_1076353[p29_res7__150] ^ p30_array_index_1082636_comb ^ p29_res7__148 ^ p29_literal_1076358[p29_res7__147] ^ p29_res7__146 ^ p29_array_index_1082319 ^ p29_array_index_1082293 ^ p29_array_index_1081996 ^ p29_array_index_1081967 ^ p29_literal_1076347[p29_array_index_1081934] ^ p29_literal_1076345[p29_array_index_1081935] ^ p29_array_index_1081936;
  assign p30_array_index_1082682_comb = p29_literal_1076355[p29_res7__564];
  assign p30_res7__156_comb = p29_literal_1076345[p30_res7__155_comb] ^ p29_literal_1076347[p30_res7__154_comb] ^ p29_literal_1076349[p29_res7__153] ^ p29_literal_1076351[p29_res7__152] ^ p29_literal_1076353[p29_res7__151] ^ p29_literal_1076355[p29_res7__150] ^ p29_res7__149 ^ p29_literal_1076358[p29_res7__148] ^ p29_res7__147 ^ p29_array_index_1082331 ^ p29_array_index_1082306 ^ p29_array_index_1082010 ^ p29_array_index_1081981 ^ p29_array_index_1081949 ^ p29_literal_1076345[p29_array_index_1081934] ^ p29_array_index_1081935;
  assign p30_res7__570_comb = p29_literal_1076345[p29_res7__569] ^ p29_literal_1076347[p29_res7__568] ^ p29_literal_1076349[p29_res7__567] ^ p29_literal_1076351[p29_res7__566] ^ p29_literal_1076353[p29_res7__565] ^ p30_array_index_1082682_comb ^ p29_res7__563 ^ p29_literal_1076358[p29_res7__562] ^ p29_res7__561 ^ p29_array_index_1082375 ^ p29_array_index_1082096 ^ p29_array_index_1082067 ^ p29_array_index_1082035 ^ p29_literal_1076347[p29_array_index_1082023] ^ p29_literal_1076345[p29_array_index_1082024] ^ p29_array_index_1082025;
  assign p30_array_index_1082692_comb = p29_literal_1076355[p29_res7__565];
  assign p30_res7__157_comb = p29_literal_1076345[p30_res7__156_comb] ^ p29_literal_1076347[p30_res7__155_comb] ^ p29_literal_1076349[p30_res7__154_comb] ^ p29_literal_1076351[p29_res7__153] ^ p29_literal_1076353[p29_res7__152] ^ p29_literal_1076355[p29_res7__151] ^ p29_res7__150 ^ p29_literal_1076358[p29_res7__149] ^ p29_res7__148 ^ p29_array_index_1082342 ^ p29_array_index_1082318 ^ p29_array_index_1082292 ^ p29_array_index_1081995 ^ p29_array_index_1081966 ^ p29_literal_1076345[p29_array_index_1081933] ^ p29_array_index_1081934;
  assign p30_res7__571_comb = p29_literal_1076345[p30_res7__570_comb] ^ p29_literal_1076347[p29_res7__569] ^ p29_literal_1076349[p29_res7__568] ^ p29_literal_1076351[p29_res7__567] ^ p29_literal_1076353[p29_res7__566] ^ p30_array_index_1082692_comb ^ p29_res7__564 ^ p29_literal_1076358[p29_res7__563] ^ p29_res7__562 ^ p29_array_index_1082387 ^ p29_array_index_1082361 ^ p29_array_index_1082081 ^ p29_array_index_1082052 ^ p29_literal_1076347[p29_array_index_1082022] ^ p29_literal_1076345[p29_array_index_1082023] ^ p29_array_index_1082024;
  assign p30_res7__158_comb = p29_literal_1076345[p30_res7__157_comb] ^ p29_literal_1076347[p30_res7__156_comb] ^ p29_literal_1076349[p30_res7__155_comb] ^ p29_literal_1076351[p30_res7__154_comb] ^ p29_literal_1076353[p29_res7__153] ^ p29_literal_1076355[p29_res7__152] ^ p29_res7__151 ^ p29_literal_1076358[p29_res7__150] ^ p29_res7__149 ^ p29_array_index_1082353 ^ p29_array_index_1082330 ^ p29_array_index_1082305 ^ p29_array_index_1082009 ^ p29_array_index_1081980 ^ p29_array_index_1081948 ^ p29_array_index_1081933;
  assign p30_res7__572_comb = p29_literal_1076345[p30_res7__571_comb] ^ p29_literal_1076347[p30_res7__570_comb] ^ p29_literal_1076349[p29_res7__569] ^ p29_literal_1076351[p29_res7__568] ^ p29_literal_1076353[p29_res7__567] ^ p29_literal_1076355[p29_res7__566] ^ p29_res7__565 ^ p29_literal_1076358[p29_res7__564] ^ p29_res7__563 ^ p29_array_index_1082399 ^ p29_array_index_1082374 ^ p29_array_index_1082095 ^ p29_array_index_1082066 ^ p29_array_index_1082034 ^ p29_literal_1076345[p29_array_index_1082022] ^ p29_array_index_1082023;
  assign p30_res7__159_comb = p29_literal_1076345[p30_res7__158_comb] ^ p29_literal_1076347[p30_res7__157_comb] ^ p29_literal_1076349[p30_res7__156_comb] ^ p29_literal_1076351[p30_res7__155_comb] ^ p29_literal_1076353[p30_res7__154_comb] ^ p29_literal_1076355[p29_res7__153] ^ p29_res7__152 ^ p29_literal_1076358[p29_res7__151] ^ p29_res7__150 ^ p30_array_index_1082636_comb ^ p29_array_index_1082341 ^ p29_array_index_1082317 ^ p29_array_index_1082291 ^ p29_array_index_1081994 ^ p29_array_index_1081965 ^ p29_array_index_1081932;
  assign p30_res7__573_comb = p29_literal_1076345[p30_res7__572_comb] ^ p29_literal_1076347[p30_res7__571_comb] ^ p29_literal_1076349[p30_res7__570_comb] ^ p29_literal_1076351[p29_res7__569] ^ p29_literal_1076353[p29_res7__568] ^ p29_literal_1076355[p29_res7__567] ^ p29_res7__566 ^ p29_literal_1076358[p29_res7__565] ^ p29_res7__564 ^ p29_array_index_1082410 ^ p29_array_index_1082386 ^ p29_array_index_1082360 ^ p29_array_index_1082080 ^ p29_array_index_1082051 ^ p29_literal_1076345[p29_array_index_1082021] ^ p29_array_index_1082022;
  assign p30_res__9_comb = {p30_res7__159_comb, p30_res7__158_comb, p30_res7__157_comb, p30_res7__156_comb, p30_res7__155_comb, p30_res7__154_comb, p29_res7__153, p29_res7__152, p29_res7__151, p29_res7__150, p29_res7__149, p29_res7__148, p29_res7__147, p29_res7__146, p29_res7__145, p29_res7__144};
  assign p30_xor_1082676_comb = p30_res__9_comb ^ p29_k2;
  assign p30_res7__574_comb = p29_literal_1076345[p30_res7__573_comb] ^ p29_literal_1076347[p30_res7__572_comb] ^ p29_literal_1076349[p30_res7__571_comb] ^ p29_literal_1076351[p30_res7__570_comb] ^ p29_literal_1076353[p29_res7__569] ^ p29_literal_1076355[p29_res7__568] ^ p29_res7__567 ^ p29_literal_1076358[p29_res7__566] ^ p29_res7__565 ^ p30_array_index_1082682_comb ^ p29_array_index_1082398 ^ p29_array_index_1082373 ^ p29_array_index_1082094 ^ p29_array_index_1082065 ^ p29_array_index_1082033 ^ p29_array_index_1082021;

  // Registers for pipe stage 30:
  reg [127:0] p30_xor_1081801;
  reg [127:0] p30_xor_1082676;
  reg [7:0] p30_array_index_1082020;
  reg [7:0] p30_res7__560;
  reg [7:0] p30_array_index_1082050;
  reg [7:0] p30_res7__561;
  reg [7:0] p30_res7__562;
  reg [7:0] p30_array_index_1082079;
  reg [7:0] p30_res7__563;
  reg [7:0] p30_res7__564;
  reg [7:0] p30_array_index_1082359;
  reg [7:0] p30_res7__565;
  reg [7:0] p30_res7__566;
  reg [7:0] p30_array_index_1082385;
  reg [7:0] p30_res7__567;
  reg [7:0] p30_res7__568;
  reg [7:0] p30_array_index_1082409;
  reg [7:0] p30_res7__569;
  reg [7:0] p30_res7__570;
  reg [7:0] p30_array_index_1082692;
  reg [7:0] p30_res7__571;
  reg [7:0] p30_res7__572;
  reg [7:0] p30_res7__573;
  reg [7:0] p30_res7__574;
  reg [7:0] p31_arr[256];
  reg [7:0] p31_literal_1076345[256];
  reg [7:0] p31_literal_1076347[256];
  reg [7:0] p31_literal_1076349[256];
  reg [7:0] p31_literal_1076351[256];
  reg [7:0] p31_literal_1076353[256];
  reg [7:0] p31_literal_1076355[256];
  reg [7:0] p31_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p30_xor_1081801 <= p29_xor_1081801;
    p30_xor_1082676 <= p30_xor_1082676_comb;
    p30_array_index_1082020 <= p29_array_index_1082020;
    p30_res7__560 <= p29_res7__560;
    p30_array_index_1082050 <= p29_array_index_1082050;
    p30_res7__561 <= p29_res7__561;
    p30_res7__562 <= p29_res7__562;
    p30_array_index_1082079 <= p29_array_index_1082079;
    p30_res7__563 <= p29_res7__563;
    p30_res7__564 <= p29_res7__564;
    p30_array_index_1082359 <= p29_array_index_1082359;
    p30_res7__565 <= p29_res7__565;
    p30_res7__566 <= p29_res7__566;
    p30_array_index_1082385 <= p29_array_index_1082385;
    p30_res7__567 <= p29_res7__567;
    p30_res7__568 <= p29_res7__568;
    p30_array_index_1082409 <= p29_array_index_1082409;
    p30_res7__569 <= p29_res7__569;
    p30_res7__570 <= p30_res7__570_comb;
    p30_array_index_1082692 <= p30_array_index_1082692_comb;
    p30_res7__571 <= p30_res7__571_comb;
    p30_res7__572 <= p30_res7__572_comb;
    p30_res7__573 <= p30_res7__573_comb;
    p30_res7__574 <= p30_res7__574_comb;
    p31_arr <= p30_arr;
    p31_literal_1076345 <= p30_literal_1076345;
    p31_literal_1076347 <= p30_literal_1076347;
    p31_literal_1076349 <= p30_literal_1076349;
    p31_literal_1076351 <= p30_literal_1076351;
    p31_literal_1076353 <= p30_literal_1076353;
    p31_literal_1076355 <= p30_literal_1076355;
    p31_literal_1076358 <= p30_literal_1076358;
  end

  // ===== Pipe stage 31:
  wire [127:0] p31_addedKey__51_comb;
  wire [7:0] p31_array_index_1082802_comb;
  wire [7:0] p31_array_index_1082803_comb;
  wire [7:0] p31_array_index_1082804_comb;
  wire [7:0] p31_array_index_1082805_comb;
  wire [7:0] p31_array_index_1082806_comb;
  wire [7:0] p31_array_index_1082807_comb;
  wire [7:0] p31_array_index_1082809_comb;
  wire [7:0] p31_array_index_1082811_comb;
  wire [7:0] p31_array_index_1082812_comb;
  wire [7:0] p31_array_index_1082813_comb;
  wire [7:0] p31_array_index_1082814_comb;
  wire [7:0] p31_array_index_1082815_comb;
  wire [7:0] p31_array_index_1082816_comb;
  wire [7:0] p31_array_index_1082818_comb;
  wire [7:0] p31_array_index_1082819_comb;
  wire [7:0] p31_array_index_1082820_comb;
  wire [7:0] p31_array_index_1082821_comb;
  wire [7:0] p31_array_index_1082822_comb;
  wire [7:0] p31_array_index_1082823_comb;
  wire [7:0] p31_array_index_1082824_comb;
  wire [7:0] p31_array_index_1082826_comb;
  wire [7:0] p31_res7__160_comb;
  wire [7:0] p31_array_index_1082835_comb;
  wire [7:0] p31_array_index_1082836_comb;
  wire [7:0] p31_array_index_1082837_comb;
  wire [7:0] p31_array_index_1082838_comb;
  wire [7:0] p31_array_index_1082839_comb;
  wire [7:0] p31_array_index_1082840_comb;
  wire [7:0] p31_res7__161_comb;
  wire [7:0] p31_array_index_1082850_comb;
  wire [7:0] p31_array_index_1082851_comb;
  wire [7:0] p31_array_index_1082852_comb;
  wire [7:0] p31_array_index_1082853_comb;
  wire [7:0] p31_array_index_1082854_comb;
  wire [7:0] p31_res7__162_comb;
  wire [7:0] p31_array_index_1082864_comb;
  wire [7:0] p31_array_index_1082865_comb;
  wire [7:0] p31_array_index_1082866_comb;
  wire [7:0] p31_array_index_1082867_comb;
  wire [7:0] p31_array_index_1082868_comb;
  wire [7:0] p31_res7__163_comb;
  wire [7:0] p31_array_index_1082879_comb;
  wire [7:0] p31_array_index_1082880_comb;
  wire [7:0] p31_array_index_1082881_comb;
  wire [7:0] p31_array_index_1082882_comb;
  wire [7:0] p31_res7__575_comb;
  wire [7:0] p31_res7__164_comb;
  wire [127:0] p31_res__35_comb;
  assign p31_addedKey__51_comb = p30_xor_1082676 ^ 128'h447c_ac80_52dd_d882_4a92_a5b0_83e5_550b;
  assign p31_array_index_1082802_comb = p30_arr[p31_addedKey__51_comb[127:120]];
  assign p31_array_index_1082803_comb = p30_arr[p31_addedKey__51_comb[119:112]];
  assign p31_array_index_1082804_comb = p30_arr[p31_addedKey__51_comb[111:104]];
  assign p31_array_index_1082805_comb = p30_arr[p31_addedKey__51_comb[103:96]];
  assign p31_array_index_1082806_comb = p30_arr[p31_addedKey__51_comb[95:88]];
  assign p31_array_index_1082807_comb = p30_arr[p31_addedKey__51_comb[87:80]];
  assign p31_array_index_1082809_comb = p30_arr[p31_addedKey__51_comb[71:64]];
  assign p31_array_index_1082811_comb = p30_arr[p31_addedKey__51_comb[55:48]];
  assign p31_array_index_1082812_comb = p30_arr[p31_addedKey__51_comb[47:40]];
  assign p31_array_index_1082813_comb = p30_arr[p31_addedKey__51_comb[39:32]];
  assign p31_array_index_1082814_comb = p30_arr[p31_addedKey__51_comb[31:24]];
  assign p31_array_index_1082815_comb = p30_arr[p31_addedKey__51_comb[23:16]];
  assign p31_array_index_1082816_comb = p30_arr[p31_addedKey__51_comb[15:8]];
  assign p31_array_index_1082818_comb = p30_literal_1076345[p31_array_index_1082802_comb];
  assign p31_array_index_1082819_comb = p30_literal_1076347[p31_array_index_1082803_comb];
  assign p31_array_index_1082820_comb = p30_literal_1076349[p31_array_index_1082804_comb];
  assign p31_array_index_1082821_comb = p30_literal_1076351[p31_array_index_1082805_comb];
  assign p31_array_index_1082822_comb = p30_literal_1076353[p31_array_index_1082806_comb];
  assign p31_array_index_1082823_comb = p30_literal_1076355[p31_array_index_1082807_comb];
  assign p31_array_index_1082824_comb = p30_arr[p31_addedKey__51_comb[79:72]];
  assign p31_array_index_1082826_comb = p30_arr[p31_addedKey__51_comb[63:56]];
  assign p31_res7__160_comb = p31_array_index_1082818_comb ^ p31_array_index_1082819_comb ^ p31_array_index_1082820_comb ^ p31_array_index_1082821_comb ^ p31_array_index_1082822_comb ^ p31_array_index_1082823_comb ^ p31_array_index_1082824_comb ^ p30_literal_1076358[p31_array_index_1082809_comb] ^ p31_array_index_1082826_comb ^ p30_literal_1076355[p31_array_index_1082811_comb] ^ p30_literal_1076353[p31_array_index_1082812_comb] ^ p30_literal_1076351[p31_array_index_1082813_comb] ^ p30_literal_1076349[p31_array_index_1082814_comb] ^ p30_literal_1076347[p31_array_index_1082815_comb] ^ p30_literal_1076345[p31_array_index_1082816_comb] ^ p30_arr[p31_addedKey__51_comb[7:0]];
  assign p31_array_index_1082835_comb = p30_literal_1076345[p31_res7__160_comb];
  assign p31_array_index_1082836_comb = p30_literal_1076347[p31_array_index_1082802_comb];
  assign p31_array_index_1082837_comb = p30_literal_1076349[p31_array_index_1082803_comb];
  assign p31_array_index_1082838_comb = p30_literal_1076351[p31_array_index_1082804_comb];
  assign p31_array_index_1082839_comb = p30_literal_1076353[p31_array_index_1082805_comb];
  assign p31_array_index_1082840_comb = p30_literal_1076355[p31_array_index_1082806_comb];
  assign p31_res7__161_comb = p31_array_index_1082835_comb ^ p31_array_index_1082836_comb ^ p31_array_index_1082837_comb ^ p31_array_index_1082838_comb ^ p31_array_index_1082839_comb ^ p31_array_index_1082840_comb ^ p31_array_index_1082807_comb ^ p30_literal_1076358[p31_array_index_1082824_comb] ^ p31_array_index_1082809_comb ^ p30_literal_1076355[p31_array_index_1082826_comb] ^ p30_literal_1076353[p31_array_index_1082811_comb] ^ p30_literal_1076351[p31_array_index_1082812_comb] ^ p30_literal_1076349[p31_array_index_1082813_comb] ^ p30_literal_1076347[p31_array_index_1082814_comb] ^ p30_literal_1076345[p31_array_index_1082815_comb] ^ p31_array_index_1082816_comb;
  assign p31_array_index_1082850_comb = p30_literal_1076347[p31_res7__160_comb];
  assign p31_array_index_1082851_comb = p30_literal_1076349[p31_array_index_1082802_comb];
  assign p31_array_index_1082852_comb = p30_literal_1076351[p31_array_index_1082803_comb];
  assign p31_array_index_1082853_comb = p30_literal_1076353[p31_array_index_1082804_comb];
  assign p31_array_index_1082854_comb = p30_literal_1076355[p31_array_index_1082805_comb];
  assign p31_res7__162_comb = p30_literal_1076345[p31_res7__161_comb] ^ p31_array_index_1082850_comb ^ p31_array_index_1082851_comb ^ p31_array_index_1082852_comb ^ p31_array_index_1082853_comb ^ p31_array_index_1082854_comb ^ p31_array_index_1082806_comb ^ p30_literal_1076358[p31_array_index_1082807_comb] ^ p31_array_index_1082824_comb ^ p30_literal_1076355[p31_array_index_1082809_comb] ^ p30_literal_1076353[p31_array_index_1082826_comb] ^ p30_literal_1076351[p31_array_index_1082811_comb] ^ p30_literal_1076349[p31_array_index_1082812_comb] ^ p30_literal_1076347[p31_array_index_1082813_comb] ^ p30_literal_1076345[p31_array_index_1082814_comb] ^ p31_array_index_1082815_comb;
  assign p31_array_index_1082864_comb = p30_literal_1076347[p31_res7__161_comb];
  assign p31_array_index_1082865_comb = p30_literal_1076349[p31_res7__160_comb];
  assign p31_array_index_1082866_comb = p30_literal_1076351[p31_array_index_1082802_comb];
  assign p31_array_index_1082867_comb = p30_literal_1076353[p31_array_index_1082803_comb];
  assign p31_array_index_1082868_comb = p30_literal_1076355[p31_array_index_1082804_comb];
  assign p31_res7__163_comb = p30_literal_1076345[p31_res7__162_comb] ^ p31_array_index_1082864_comb ^ p31_array_index_1082865_comb ^ p31_array_index_1082866_comb ^ p31_array_index_1082867_comb ^ p31_array_index_1082868_comb ^ p31_array_index_1082805_comb ^ p30_literal_1076358[p31_array_index_1082806_comb] ^ p31_array_index_1082807_comb ^ p30_literal_1076355[p31_array_index_1082824_comb] ^ p30_literal_1076353[p31_array_index_1082809_comb] ^ p30_literal_1076351[p31_array_index_1082826_comb] ^ p30_literal_1076349[p31_array_index_1082811_comb] ^ p30_literal_1076347[p31_array_index_1082812_comb] ^ p30_literal_1076345[p31_array_index_1082813_comb] ^ p31_array_index_1082814_comb;
  assign p31_array_index_1082879_comb = p30_literal_1076349[p31_res7__161_comb];
  assign p31_array_index_1082880_comb = p30_literal_1076351[p31_res7__160_comb];
  assign p31_array_index_1082881_comb = p30_literal_1076353[p31_array_index_1082802_comb];
  assign p31_array_index_1082882_comb = p30_literal_1076355[p31_array_index_1082803_comb];
  assign p31_res7__575_comb = p30_literal_1076345[p30_res7__574] ^ p30_literal_1076347[p30_res7__573] ^ p30_literal_1076349[p30_res7__572] ^ p30_literal_1076351[p30_res7__571] ^ p30_literal_1076353[p30_res7__570] ^ p30_literal_1076355[p30_res7__569] ^ p30_res7__568 ^ p30_literal_1076358[p30_res7__567] ^ p30_res7__566 ^ p30_array_index_1082692 ^ p30_array_index_1082409 ^ p30_array_index_1082385 ^ p30_array_index_1082359 ^ p30_array_index_1082079 ^ p30_array_index_1082050 ^ p30_array_index_1082020;
  assign p31_res7__164_comb = p30_literal_1076345[p31_res7__163_comb] ^ p30_literal_1076347[p31_res7__162_comb] ^ p31_array_index_1082879_comb ^ p31_array_index_1082880_comb ^ p31_array_index_1082881_comb ^ p31_array_index_1082882_comb ^ p31_array_index_1082804_comb ^ p30_literal_1076358[p31_array_index_1082805_comb] ^ p31_array_index_1082806_comb ^ p31_array_index_1082823_comb ^ p30_literal_1076353[p31_array_index_1082824_comb] ^ p30_literal_1076351[p31_array_index_1082809_comb] ^ p30_literal_1076349[p31_array_index_1082826_comb] ^ p30_literal_1076347[p31_array_index_1082811_comb] ^ p30_literal_1076345[p31_array_index_1082812_comb] ^ p31_array_index_1082813_comb;
  assign p31_res__35_comb = {p31_res7__575_comb, p30_res7__574, p30_res7__573, p30_res7__572, p30_res7__571, p30_res7__570, p30_res7__569, p30_res7__568, p30_res7__567, p30_res7__566, p30_res7__565, p30_res7__564, p30_res7__563, p30_res7__562, p30_res7__561, p30_res7__560};

  // Registers for pipe stage 31:
  reg [127:0] p31_xor_1081801;
  reg [127:0] p31_xor_1082676;
  reg [7:0] p31_array_index_1082802;
  reg [7:0] p31_array_index_1082803;
  reg [7:0] p31_array_index_1082804;
  reg [7:0] p31_array_index_1082805;
  reg [7:0] p31_array_index_1082806;
  reg [7:0] p31_array_index_1082807;
  reg [7:0] p31_array_index_1082809;
  reg [7:0] p31_array_index_1082811;
  reg [7:0] p31_array_index_1082812;
  reg [7:0] p31_array_index_1082818;
  reg [7:0] p31_array_index_1082819;
  reg [7:0] p31_array_index_1082820;
  reg [7:0] p31_array_index_1082821;
  reg [7:0] p31_array_index_1082822;
  reg [7:0] p31_array_index_1082824;
  reg [7:0] p31_array_index_1082826;
  reg [7:0] p31_res7__160;
  reg [7:0] p31_array_index_1082835;
  reg [7:0] p31_array_index_1082836;
  reg [7:0] p31_array_index_1082837;
  reg [7:0] p31_array_index_1082838;
  reg [7:0] p31_array_index_1082839;
  reg [7:0] p31_array_index_1082840;
  reg [7:0] p31_res7__161;
  reg [7:0] p31_array_index_1082850;
  reg [7:0] p31_array_index_1082851;
  reg [7:0] p31_array_index_1082852;
  reg [7:0] p31_array_index_1082853;
  reg [7:0] p31_array_index_1082854;
  reg [7:0] p31_res7__162;
  reg [7:0] p31_array_index_1082864;
  reg [7:0] p31_array_index_1082865;
  reg [7:0] p31_array_index_1082866;
  reg [7:0] p31_array_index_1082867;
  reg [7:0] p31_array_index_1082868;
  reg [7:0] p31_res7__163;
  reg [7:0] p31_array_index_1082879;
  reg [7:0] p31_array_index_1082880;
  reg [7:0] p31_array_index_1082881;
  reg [7:0] p31_array_index_1082882;
  reg [7:0] p31_res7__164;
  reg [127:0] p31_res__35;
  reg [7:0] p32_arr[256];
  reg [7:0] p32_literal_1076345[256];
  reg [7:0] p32_literal_1076347[256];
  reg [7:0] p32_literal_1076349[256];
  reg [7:0] p32_literal_1076351[256];
  reg [7:0] p32_literal_1076353[256];
  reg [7:0] p32_literal_1076355[256];
  reg [7:0] p32_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p31_xor_1081801 <= p30_xor_1081801;
    p31_xor_1082676 <= p30_xor_1082676;
    p31_array_index_1082802 <= p31_array_index_1082802_comb;
    p31_array_index_1082803 <= p31_array_index_1082803_comb;
    p31_array_index_1082804 <= p31_array_index_1082804_comb;
    p31_array_index_1082805 <= p31_array_index_1082805_comb;
    p31_array_index_1082806 <= p31_array_index_1082806_comb;
    p31_array_index_1082807 <= p31_array_index_1082807_comb;
    p31_array_index_1082809 <= p31_array_index_1082809_comb;
    p31_array_index_1082811 <= p31_array_index_1082811_comb;
    p31_array_index_1082812 <= p31_array_index_1082812_comb;
    p31_array_index_1082818 <= p31_array_index_1082818_comb;
    p31_array_index_1082819 <= p31_array_index_1082819_comb;
    p31_array_index_1082820 <= p31_array_index_1082820_comb;
    p31_array_index_1082821 <= p31_array_index_1082821_comb;
    p31_array_index_1082822 <= p31_array_index_1082822_comb;
    p31_array_index_1082824 <= p31_array_index_1082824_comb;
    p31_array_index_1082826 <= p31_array_index_1082826_comb;
    p31_res7__160 <= p31_res7__160_comb;
    p31_array_index_1082835 <= p31_array_index_1082835_comb;
    p31_array_index_1082836 <= p31_array_index_1082836_comb;
    p31_array_index_1082837 <= p31_array_index_1082837_comb;
    p31_array_index_1082838 <= p31_array_index_1082838_comb;
    p31_array_index_1082839 <= p31_array_index_1082839_comb;
    p31_array_index_1082840 <= p31_array_index_1082840_comb;
    p31_res7__161 <= p31_res7__161_comb;
    p31_array_index_1082850 <= p31_array_index_1082850_comb;
    p31_array_index_1082851 <= p31_array_index_1082851_comb;
    p31_array_index_1082852 <= p31_array_index_1082852_comb;
    p31_array_index_1082853 <= p31_array_index_1082853_comb;
    p31_array_index_1082854 <= p31_array_index_1082854_comb;
    p31_res7__162 <= p31_res7__162_comb;
    p31_array_index_1082864 <= p31_array_index_1082864_comb;
    p31_array_index_1082865 <= p31_array_index_1082865_comb;
    p31_array_index_1082866 <= p31_array_index_1082866_comb;
    p31_array_index_1082867 <= p31_array_index_1082867_comb;
    p31_array_index_1082868 <= p31_array_index_1082868_comb;
    p31_res7__163 <= p31_res7__163_comb;
    p31_array_index_1082879 <= p31_array_index_1082879_comb;
    p31_array_index_1082880 <= p31_array_index_1082880_comb;
    p31_array_index_1082881 <= p31_array_index_1082881_comb;
    p31_array_index_1082882 <= p31_array_index_1082882_comb;
    p31_res7__164 <= p31_res7__164_comb;
    p31_res__35 <= p31_res__35_comb;
    p32_arr <= p31_arr;
    p32_literal_1076345 <= p31_literal_1076345;
    p32_literal_1076347 <= p31_literal_1076347;
    p32_literal_1076349 <= p31_literal_1076349;
    p32_literal_1076351 <= p31_literal_1076351;
    p32_literal_1076353 <= p31_literal_1076353;
    p32_literal_1076355 <= p31_literal_1076355;
    p32_literal_1076358 <= p31_literal_1076358;
  end

  // ===== Pipe stage 32:
  wire [7:0] p32_array_index_1083005_comb;
  wire [7:0] p32_array_index_1083006_comb;
  wire [7:0] p32_array_index_1083007_comb;
  wire [7:0] p32_array_index_1083008_comb;
  wire [7:0] p32_res7__165_comb;
  wire [7:0] p32_array_index_1083019_comb;
  wire [7:0] p32_array_index_1083020_comb;
  wire [7:0] p32_array_index_1083021_comb;
  wire [7:0] p32_res7__166_comb;
  wire [7:0] p32_array_index_1083031_comb;
  wire [7:0] p32_array_index_1083032_comb;
  wire [7:0] p32_array_index_1083033_comb;
  wire [7:0] p32_res7__167_comb;
  wire [7:0] p32_array_index_1083044_comb;
  wire [7:0] p32_array_index_1083045_comb;
  wire [7:0] p32_res7__168_comb;
  wire [7:0] p32_array_index_1083055_comb;
  wire [7:0] p32_array_index_1083056_comb;
  wire [7:0] p32_res7__169_comb;
  wire [7:0] p32_array_index_1083062_comb;
  wire [7:0] p32_array_index_1083063_comb;
  wire [7:0] p32_array_index_1083064_comb;
  wire [7:0] p32_array_index_1083065_comb;
  wire [7:0] p32_array_index_1083066_comb;
  wire [7:0] p32_array_index_1083067_comb;
  wire [7:0] p32_array_index_1083068_comb;
  wire [7:0] p32_array_index_1083069_comb;
  wire [7:0] p32_array_index_1083070_comb;
  assign p32_array_index_1083005_comb = p31_literal_1076349[p31_res7__162];
  assign p32_array_index_1083006_comb = p31_literal_1076351[p31_res7__161];
  assign p32_array_index_1083007_comb = p31_literal_1076353[p31_res7__160];
  assign p32_array_index_1083008_comb = p31_literal_1076355[p31_array_index_1082802];
  assign p32_res7__165_comb = p31_literal_1076345[p31_res7__164] ^ p31_literal_1076347[p31_res7__163] ^ p32_array_index_1083005_comb ^ p32_array_index_1083006_comb ^ p32_array_index_1083007_comb ^ p32_array_index_1083008_comb ^ p31_array_index_1082803 ^ p31_literal_1076358[p31_array_index_1082804] ^ p31_array_index_1082805 ^ p31_array_index_1082840 ^ p31_literal_1076353[p31_array_index_1082807] ^ p31_literal_1076351[p31_array_index_1082824] ^ p31_literal_1076349[p31_array_index_1082809] ^ p31_literal_1076347[p31_array_index_1082826] ^ p31_literal_1076345[p31_array_index_1082811] ^ p31_array_index_1082812;
  assign p32_array_index_1083019_comb = p31_literal_1076351[p31_res7__162];
  assign p32_array_index_1083020_comb = p31_literal_1076353[p31_res7__161];
  assign p32_array_index_1083021_comb = p31_literal_1076355[p31_res7__160];
  assign p32_res7__166_comb = p31_literal_1076345[p32_res7__165_comb] ^ p31_literal_1076347[p31_res7__164] ^ p31_literal_1076349[p31_res7__163] ^ p32_array_index_1083019_comb ^ p32_array_index_1083020_comb ^ p32_array_index_1083021_comb ^ p31_array_index_1082802 ^ p31_literal_1076358[p31_array_index_1082803] ^ p31_array_index_1082804 ^ p31_array_index_1082854 ^ p31_array_index_1082822 ^ p31_literal_1076351[p31_array_index_1082807] ^ p31_literal_1076349[p31_array_index_1082824] ^ p31_literal_1076347[p31_array_index_1082809] ^ p31_literal_1076345[p31_array_index_1082826] ^ p31_array_index_1082811;
  assign p32_array_index_1083031_comb = p31_literal_1076351[p31_res7__163];
  assign p32_array_index_1083032_comb = p31_literal_1076353[p31_res7__162];
  assign p32_array_index_1083033_comb = p31_literal_1076355[p31_res7__161];
  assign p32_res7__167_comb = p31_literal_1076345[p32_res7__166_comb] ^ p31_literal_1076347[p32_res7__165_comb] ^ p31_literal_1076349[p31_res7__164] ^ p32_array_index_1083031_comb ^ p32_array_index_1083032_comb ^ p32_array_index_1083033_comb ^ p31_res7__160 ^ p31_literal_1076358[p31_array_index_1082802] ^ p31_array_index_1082803 ^ p31_array_index_1082868 ^ p31_array_index_1082839 ^ p31_literal_1076351[p31_array_index_1082806] ^ p31_literal_1076349[p31_array_index_1082807] ^ p31_literal_1076347[p31_array_index_1082824] ^ p31_literal_1076345[p31_array_index_1082809] ^ p31_array_index_1082826;
  assign p32_array_index_1083044_comb = p31_literal_1076353[p31_res7__163];
  assign p32_array_index_1083045_comb = p31_literal_1076355[p31_res7__162];
  assign p32_res7__168_comb = p31_literal_1076345[p32_res7__167_comb] ^ p31_literal_1076347[p32_res7__166_comb] ^ p31_literal_1076349[p32_res7__165_comb] ^ p31_literal_1076351[p31_res7__164] ^ p32_array_index_1083044_comb ^ p32_array_index_1083045_comb ^ p31_res7__161 ^ p31_literal_1076358[p31_res7__160] ^ p31_array_index_1082802 ^ p31_array_index_1082882 ^ p31_array_index_1082853 ^ p31_array_index_1082821 ^ p31_literal_1076349[p31_array_index_1082806] ^ p31_literal_1076347[p31_array_index_1082807] ^ p31_literal_1076345[p31_array_index_1082824] ^ p31_array_index_1082809;
  assign p32_array_index_1083055_comb = p31_literal_1076353[p31_res7__164];
  assign p32_array_index_1083056_comb = p31_literal_1076355[p31_res7__163];
  assign p32_res7__169_comb = p31_literal_1076345[p32_res7__168_comb] ^ p31_literal_1076347[p32_res7__167_comb] ^ p31_literal_1076349[p32_res7__166_comb] ^ p31_literal_1076351[p32_res7__165_comb] ^ p32_array_index_1083055_comb ^ p32_array_index_1083056_comb ^ p31_res7__162 ^ p31_literal_1076358[p31_res7__161] ^ p31_res7__160 ^ p32_array_index_1083008_comb ^ p31_array_index_1082867 ^ p31_array_index_1082838 ^ p31_literal_1076349[p31_array_index_1082805] ^ p31_literal_1076347[p31_array_index_1082806] ^ p31_literal_1076345[p31_array_index_1082807] ^ p31_array_index_1082824;
  assign p32_array_index_1083062_comb = p31_literal_1076345[p32_res7__169_comb];
  assign p32_array_index_1083063_comb = p31_literal_1076347[p32_res7__168_comb];
  assign p32_array_index_1083064_comb = p31_literal_1076349[p32_res7__167_comb];
  assign p32_array_index_1083065_comb = p31_literal_1076351[p32_res7__166_comb];
  assign p32_array_index_1083066_comb = p31_literal_1076353[p32_res7__165_comb];
  assign p32_array_index_1083067_comb = p31_literal_1076355[p31_res7__164];
  assign p32_array_index_1083068_comb = p31_literal_1076358[p31_res7__162];
  assign p32_array_index_1083069_comb = p31_literal_1076347[p31_array_index_1082805];
  assign p32_array_index_1083070_comb = p31_literal_1076345[p31_array_index_1082806];

  // Registers for pipe stage 32:
  reg [127:0] p32_xor_1081801;
  reg [127:0] p32_xor_1082676;
  reg [7:0] p32_array_index_1082802;
  reg [7:0] p32_array_index_1082803;
  reg [7:0] p32_array_index_1082804;
  reg [7:0] p32_array_index_1082805;
  reg [7:0] p32_array_index_1082806;
  reg [7:0] p32_array_index_1082807;
  reg [7:0] p32_array_index_1082818;
  reg [7:0] p32_array_index_1082819;
  reg [7:0] p32_array_index_1082820;
  reg [7:0] p32_res7__160;
  reg [7:0] p32_array_index_1082835;
  reg [7:0] p32_array_index_1082836;
  reg [7:0] p32_array_index_1082837;
  reg [7:0] p32_res7__161;
  reg [7:0] p32_array_index_1082850;
  reg [7:0] p32_array_index_1082851;
  reg [7:0] p32_array_index_1082852;
  reg [7:0] p32_res7__162;
  reg [7:0] p32_array_index_1082864;
  reg [7:0] p32_array_index_1082865;
  reg [7:0] p32_array_index_1082866;
  reg [7:0] p32_res7__163;
  reg [7:0] p32_array_index_1082879;
  reg [7:0] p32_array_index_1082880;
  reg [7:0] p32_array_index_1082881;
  reg [7:0] p32_res7__164;
  reg [7:0] p32_array_index_1083005;
  reg [7:0] p32_array_index_1083006;
  reg [7:0] p32_array_index_1083007;
  reg [7:0] p32_res7__165;
  reg [7:0] p32_array_index_1083019;
  reg [7:0] p32_array_index_1083020;
  reg [7:0] p32_array_index_1083021;
  reg [7:0] p32_res7__166;
  reg [7:0] p32_array_index_1083031;
  reg [7:0] p32_array_index_1083032;
  reg [7:0] p32_array_index_1083033;
  reg [7:0] p32_res7__167;
  reg [7:0] p32_array_index_1083044;
  reg [7:0] p32_array_index_1083045;
  reg [7:0] p32_res7__168;
  reg [7:0] p32_array_index_1083055;
  reg [7:0] p32_array_index_1083056;
  reg [7:0] p32_res7__169;
  reg [7:0] p32_array_index_1083062;
  reg [7:0] p32_array_index_1083063;
  reg [7:0] p32_array_index_1083064;
  reg [7:0] p32_array_index_1083065;
  reg [7:0] p32_array_index_1083066;
  reg [7:0] p32_array_index_1083067;
  reg [7:0] p32_array_index_1083068;
  reg [7:0] p32_array_index_1083069;
  reg [7:0] p32_array_index_1083070;
  reg [127:0] p32_res__35;
  reg [7:0] p33_arr[256];
  reg [7:0] p33_literal_1076345[256];
  reg [7:0] p33_literal_1076347[256];
  reg [7:0] p33_literal_1076349[256];
  reg [7:0] p33_literal_1076351[256];
  reg [7:0] p33_literal_1076353[256];
  reg [7:0] p33_literal_1076355[256];
  reg [7:0] p33_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p32_xor_1081801 <= p31_xor_1081801;
    p32_xor_1082676 <= p31_xor_1082676;
    p32_array_index_1082802 <= p31_array_index_1082802;
    p32_array_index_1082803 <= p31_array_index_1082803;
    p32_array_index_1082804 <= p31_array_index_1082804;
    p32_array_index_1082805 <= p31_array_index_1082805;
    p32_array_index_1082806 <= p31_array_index_1082806;
    p32_array_index_1082807 <= p31_array_index_1082807;
    p32_array_index_1082818 <= p31_array_index_1082818;
    p32_array_index_1082819 <= p31_array_index_1082819;
    p32_array_index_1082820 <= p31_array_index_1082820;
    p32_res7__160 <= p31_res7__160;
    p32_array_index_1082835 <= p31_array_index_1082835;
    p32_array_index_1082836 <= p31_array_index_1082836;
    p32_array_index_1082837 <= p31_array_index_1082837;
    p32_res7__161 <= p31_res7__161;
    p32_array_index_1082850 <= p31_array_index_1082850;
    p32_array_index_1082851 <= p31_array_index_1082851;
    p32_array_index_1082852 <= p31_array_index_1082852;
    p32_res7__162 <= p31_res7__162;
    p32_array_index_1082864 <= p31_array_index_1082864;
    p32_array_index_1082865 <= p31_array_index_1082865;
    p32_array_index_1082866 <= p31_array_index_1082866;
    p32_res7__163 <= p31_res7__163;
    p32_array_index_1082879 <= p31_array_index_1082879;
    p32_array_index_1082880 <= p31_array_index_1082880;
    p32_array_index_1082881 <= p31_array_index_1082881;
    p32_res7__164 <= p31_res7__164;
    p32_array_index_1083005 <= p32_array_index_1083005_comb;
    p32_array_index_1083006 <= p32_array_index_1083006_comb;
    p32_array_index_1083007 <= p32_array_index_1083007_comb;
    p32_res7__165 <= p32_res7__165_comb;
    p32_array_index_1083019 <= p32_array_index_1083019_comb;
    p32_array_index_1083020 <= p32_array_index_1083020_comb;
    p32_array_index_1083021 <= p32_array_index_1083021_comb;
    p32_res7__166 <= p32_res7__166_comb;
    p32_array_index_1083031 <= p32_array_index_1083031_comb;
    p32_array_index_1083032 <= p32_array_index_1083032_comb;
    p32_array_index_1083033 <= p32_array_index_1083033_comb;
    p32_res7__167 <= p32_res7__167_comb;
    p32_array_index_1083044 <= p32_array_index_1083044_comb;
    p32_array_index_1083045 <= p32_array_index_1083045_comb;
    p32_res7__168 <= p32_res7__168_comb;
    p32_array_index_1083055 <= p32_array_index_1083055_comb;
    p32_array_index_1083056 <= p32_array_index_1083056_comb;
    p32_res7__169 <= p32_res7__169_comb;
    p32_array_index_1083062 <= p32_array_index_1083062_comb;
    p32_array_index_1083063 <= p32_array_index_1083063_comb;
    p32_array_index_1083064 <= p32_array_index_1083064_comb;
    p32_array_index_1083065 <= p32_array_index_1083065_comb;
    p32_array_index_1083066 <= p32_array_index_1083066_comb;
    p32_array_index_1083067 <= p32_array_index_1083067_comb;
    p32_array_index_1083068 <= p32_array_index_1083068_comb;
    p32_array_index_1083069 <= p32_array_index_1083069_comb;
    p32_array_index_1083070 <= p32_array_index_1083070_comb;
    p32_res__35 <= p31_res__35;
    p33_arr <= p32_arr;
    p33_literal_1076345 <= p32_literal_1076345;
    p33_literal_1076347 <= p32_literal_1076347;
    p33_literal_1076349 <= p32_literal_1076349;
    p33_literal_1076351 <= p32_literal_1076351;
    p33_literal_1076353 <= p32_literal_1076353;
    p33_literal_1076355 <= p32_literal_1076355;
    p33_literal_1076358 <= p32_literal_1076358;
  end

  // ===== Pipe stage 33:
  wire [7:0] p33_res7__170_comb;
  wire [7:0] p33_array_index_1083205_comb;
  wire [7:0] p33_res7__171_comb;
  wire [7:0] p33_res7__172_comb;
  wire [7:0] p33_res7__173_comb;
  wire [7:0] p33_res7__174_comb;
  wire [7:0] p33_res7__175_comb;
  wire [127:0] p33_res__10_comb;
  wire [127:0] p33_xor_1083245_comb;
  assign p33_res7__170_comb = p32_array_index_1083062 ^ p32_array_index_1083063 ^ p32_array_index_1083064 ^ p32_array_index_1083065 ^ p32_array_index_1083066 ^ p32_array_index_1083067 ^ p32_res7__163 ^ p32_array_index_1083068 ^ p32_res7__161 ^ p32_array_index_1083021 ^ p32_array_index_1082881 ^ p32_array_index_1082852 ^ p32_array_index_1082820 ^ p32_array_index_1083069 ^ p32_array_index_1083070 ^ p32_array_index_1082807;
  assign p33_array_index_1083205_comb = p32_literal_1076355[p32_res7__165];
  assign p33_res7__171_comb = p32_literal_1076345[p33_res7__170_comb] ^ p32_literal_1076347[p32_res7__169] ^ p32_literal_1076349[p32_res7__168] ^ p32_literal_1076351[p32_res7__167] ^ p32_literal_1076353[p32_res7__166] ^ p33_array_index_1083205_comb ^ p32_res7__164 ^ p32_literal_1076358[p32_res7__163] ^ p32_res7__162 ^ p32_array_index_1083033 ^ p32_array_index_1083007 ^ p32_array_index_1082866 ^ p32_array_index_1082837 ^ p32_literal_1076347[p32_array_index_1082804] ^ p32_literal_1076345[p32_array_index_1082805] ^ p32_array_index_1082806;
  assign p33_res7__172_comb = p32_literal_1076345[p33_res7__171_comb] ^ p32_literal_1076347[p33_res7__170_comb] ^ p32_literal_1076349[p32_res7__169] ^ p32_literal_1076351[p32_res7__168] ^ p32_literal_1076353[p32_res7__167] ^ p32_literal_1076355[p32_res7__166] ^ p32_res7__165 ^ p32_literal_1076358[p32_res7__164] ^ p32_res7__163 ^ p32_array_index_1083045 ^ p32_array_index_1083020 ^ p32_array_index_1082880 ^ p32_array_index_1082851 ^ p32_array_index_1082819 ^ p32_literal_1076345[p32_array_index_1082804] ^ p32_array_index_1082805;
  assign p33_res7__173_comb = p32_literal_1076345[p33_res7__172_comb] ^ p32_literal_1076347[p33_res7__171_comb] ^ p32_literal_1076349[p33_res7__170_comb] ^ p32_literal_1076351[p32_res7__169] ^ p32_literal_1076353[p32_res7__168] ^ p32_literal_1076355[p32_res7__167] ^ p32_res7__166 ^ p32_literal_1076358[p32_res7__165] ^ p32_res7__164 ^ p32_array_index_1083056 ^ p32_array_index_1083032 ^ p32_array_index_1083006 ^ p32_array_index_1082865 ^ p32_array_index_1082836 ^ p32_literal_1076345[p32_array_index_1082803] ^ p32_array_index_1082804;
  assign p33_res7__174_comb = p32_literal_1076345[p33_res7__173_comb] ^ p32_literal_1076347[p33_res7__172_comb] ^ p32_literal_1076349[p33_res7__171_comb] ^ p32_literal_1076351[p33_res7__170_comb] ^ p32_literal_1076353[p32_res7__169] ^ p32_literal_1076355[p32_res7__168] ^ p32_res7__167 ^ p32_literal_1076358[p32_res7__166] ^ p32_res7__165 ^ p32_array_index_1083067 ^ p32_array_index_1083044 ^ p32_array_index_1083019 ^ p32_array_index_1082879 ^ p32_array_index_1082850 ^ p32_array_index_1082818 ^ p32_array_index_1082803;
  assign p33_res7__175_comb = p32_literal_1076345[p33_res7__174_comb] ^ p32_literal_1076347[p33_res7__173_comb] ^ p32_literal_1076349[p33_res7__172_comb] ^ p32_literal_1076351[p33_res7__171_comb] ^ p32_literal_1076353[p33_res7__170_comb] ^ p32_literal_1076355[p32_res7__169] ^ p32_res7__168 ^ p32_literal_1076358[p32_res7__167] ^ p32_res7__166 ^ p33_array_index_1083205_comb ^ p32_array_index_1083055 ^ p32_array_index_1083031 ^ p32_array_index_1083005 ^ p32_array_index_1082864 ^ p32_array_index_1082835 ^ p32_array_index_1082802;
  assign p33_res__10_comb = {p33_res7__175_comb, p33_res7__174_comb, p33_res7__173_comb, p33_res7__172_comb, p33_res7__171_comb, p33_res7__170_comb, p32_res7__169, p32_res7__168, p32_res7__167, p32_res7__166, p32_res7__165, p32_res7__164, p32_res7__163, p32_res7__162, p32_res7__161, p32_res7__160};
  assign p33_xor_1083245_comb = p33_res__10_comb ^ p32_xor_1081801;

  // Registers for pipe stage 33:
  reg [127:0] p33_xor_1082676;
  reg [127:0] p33_xor_1083245;
  reg [127:0] p33_res__35;
  reg [7:0] p34_arr[256];
  reg [7:0] p34_literal_1076345[256];
  reg [7:0] p34_literal_1076347[256];
  reg [7:0] p34_literal_1076349[256];
  reg [7:0] p34_literal_1076351[256];
  reg [7:0] p34_literal_1076353[256];
  reg [7:0] p34_literal_1076355[256];
  reg [7:0] p34_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p33_xor_1082676 <= p32_xor_1082676;
    p33_xor_1083245 <= p33_xor_1083245_comb;
    p33_res__35 <= p32_res__35;
    p34_arr <= p33_arr;
    p34_literal_1076345 <= p33_literal_1076345;
    p34_literal_1076347 <= p33_literal_1076347;
    p34_literal_1076349 <= p33_literal_1076349;
    p34_literal_1076351 <= p33_literal_1076351;
    p34_literal_1076353 <= p33_literal_1076353;
    p34_literal_1076355 <= p33_literal_1076355;
    p34_literal_1076358 <= p33_literal_1076358;
  end

  // ===== Pipe stage 34:
  wire [127:0] p34_addedKey__52_comb;
  wire [7:0] p34_array_index_1083283_comb;
  wire [7:0] p34_array_index_1083284_comb;
  wire [7:0] p34_array_index_1083285_comb;
  wire [7:0] p34_array_index_1083286_comb;
  wire [7:0] p34_array_index_1083287_comb;
  wire [7:0] p34_array_index_1083288_comb;
  wire [7:0] p34_array_index_1083290_comb;
  wire [7:0] p34_array_index_1083292_comb;
  wire [7:0] p34_array_index_1083293_comb;
  wire [7:0] p34_array_index_1083294_comb;
  wire [7:0] p34_array_index_1083295_comb;
  wire [7:0] p34_array_index_1083296_comb;
  wire [7:0] p34_array_index_1083297_comb;
  wire [7:0] p34_array_index_1083299_comb;
  wire [7:0] p34_array_index_1083300_comb;
  wire [7:0] p34_array_index_1083301_comb;
  wire [7:0] p34_array_index_1083302_comb;
  wire [7:0] p34_array_index_1083303_comb;
  wire [7:0] p34_array_index_1083304_comb;
  wire [7:0] p34_array_index_1083305_comb;
  wire [7:0] p34_array_index_1083307_comb;
  wire [7:0] p34_res7__176_comb;
  wire [7:0] p34_array_index_1083316_comb;
  wire [7:0] p34_array_index_1083317_comb;
  wire [7:0] p34_array_index_1083318_comb;
  wire [7:0] p34_array_index_1083319_comb;
  wire [7:0] p34_array_index_1083320_comb;
  wire [7:0] p34_array_index_1083321_comb;
  wire [7:0] p34_res7__177_comb;
  wire [7:0] p34_array_index_1083331_comb;
  wire [7:0] p34_array_index_1083332_comb;
  wire [7:0] p34_array_index_1083333_comb;
  wire [7:0] p34_array_index_1083334_comb;
  wire [7:0] p34_array_index_1083335_comb;
  wire [7:0] p34_res7__178_comb;
  wire [7:0] p34_array_index_1083345_comb;
  wire [7:0] p34_array_index_1083346_comb;
  wire [7:0] p34_array_index_1083347_comb;
  wire [7:0] p34_array_index_1083348_comb;
  wire [7:0] p34_array_index_1083349_comb;
  wire [7:0] p34_res7__179_comb;
  wire [7:0] p34_array_index_1083360_comb;
  wire [7:0] p34_array_index_1083361_comb;
  wire [7:0] p34_array_index_1083362_comb;
  wire [7:0] p34_array_index_1083363_comb;
  wire [7:0] p34_res7__180_comb;
  assign p34_addedKey__52_comb = p33_xor_1083245 ^ 128'h8d94_2d1d_95e6_7d2c_1a67_10c0_d5ff_3f0c;
  assign p34_array_index_1083283_comb = p33_arr[p34_addedKey__52_comb[127:120]];
  assign p34_array_index_1083284_comb = p33_arr[p34_addedKey__52_comb[119:112]];
  assign p34_array_index_1083285_comb = p33_arr[p34_addedKey__52_comb[111:104]];
  assign p34_array_index_1083286_comb = p33_arr[p34_addedKey__52_comb[103:96]];
  assign p34_array_index_1083287_comb = p33_arr[p34_addedKey__52_comb[95:88]];
  assign p34_array_index_1083288_comb = p33_arr[p34_addedKey__52_comb[87:80]];
  assign p34_array_index_1083290_comb = p33_arr[p34_addedKey__52_comb[71:64]];
  assign p34_array_index_1083292_comb = p33_arr[p34_addedKey__52_comb[55:48]];
  assign p34_array_index_1083293_comb = p33_arr[p34_addedKey__52_comb[47:40]];
  assign p34_array_index_1083294_comb = p33_arr[p34_addedKey__52_comb[39:32]];
  assign p34_array_index_1083295_comb = p33_arr[p34_addedKey__52_comb[31:24]];
  assign p34_array_index_1083296_comb = p33_arr[p34_addedKey__52_comb[23:16]];
  assign p34_array_index_1083297_comb = p33_arr[p34_addedKey__52_comb[15:8]];
  assign p34_array_index_1083299_comb = p33_literal_1076345[p34_array_index_1083283_comb];
  assign p34_array_index_1083300_comb = p33_literal_1076347[p34_array_index_1083284_comb];
  assign p34_array_index_1083301_comb = p33_literal_1076349[p34_array_index_1083285_comb];
  assign p34_array_index_1083302_comb = p33_literal_1076351[p34_array_index_1083286_comb];
  assign p34_array_index_1083303_comb = p33_literal_1076353[p34_array_index_1083287_comb];
  assign p34_array_index_1083304_comb = p33_literal_1076355[p34_array_index_1083288_comb];
  assign p34_array_index_1083305_comb = p33_arr[p34_addedKey__52_comb[79:72]];
  assign p34_array_index_1083307_comb = p33_arr[p34_addedKey__52_comb[63:56]];
  assign p34_res7__176_comb = p34_array_index_1083299_comb ^ p34_array_index_1083300_comb ^ p34_array_index_1083301_comb ^ p34_array_index_1083302_comb ^ p34_array_index_1083303_comb ^ p34_array_index_1083304_comb ^ p34_array_index_1083305_comb ^ p33_literal_1076358[p34_array_index_1083290_comb] ^ p34_array_index_1083307_comb ^ p33_literal_1076355[p34_array_index_1083292_comb] ^ p33_literal_1076353[p34_array_index_1083293_comb] ^ p33_literal_1076351[p34_array_index_1083294_comb] ^ p33_literal_1076349[p34_array_index_1083295_comb] ^ p33_literal_1076347[p34_array_index_1083296_comb] ^ p33_literal_1076345[p34_array_index_1083297_comb] ^ p33_arr[p34_addedKey__52_comb[7:0]];
  assign p34_array_index_1083316_comb = p33_literal_1076345[p34_res7__176_comb];
  assign p34_array_index_1083317_comb = p33_literal_1076347[p34_array_index_1083283_comb];
  assign p34_array_index_1083318_comb = p33_literal_1076349[p34_array_index_1083284_comb];
  assign p34_array_index_1083319_comb = p33_literal_1076351[p34_array_index_1083285_comb];
  assign p34_array_index_1083320_comb = p33_literal_1076353[p34_array_index_1083286_comb];
  assign p34_array_index_1083321_comb = p33_literal_1076355[p34_array_index_1083287_comb];
  assign p34_res7__177_comb = p34_array_index_1083316_comb ^ p34_array_index_1083317_comb ^ p34_array_index_1083318_comb ^ p34_array_index_1083319_comb ^ p34_array_index_1083320_comb ^ p34_array_index_1083321_comb ^ p34_array_index_1083288_comb ^ p33_literal_1076358[p34_array_index_1083305_comb] ^ p34_array_index_1083290_comb ^ p33_literal_1076355[p34_array_index_1083307_comb] ^ p33_literal_1076353[p34_array_index_1083292_comb] ^ p33_literal_1076351[p34_array_index_1083293_comb] ^ p33_literal_1076349[p34_array_index_1083294_comb] ^ p33_literal_1076347[p34_array_index_1083295_comb] ^ p33_literal_1076345[p34_array_index_1083296_comb] ^ p34_array_index_1083297_comb;
  assign p34_array_index_1083331_comb = p33_literal_1076347[p34_res7__176_comb];
  assign p34_array_index_1083332_comb = p33_literal_1076349[p34_array_index_1083283_comb];
  assign p34_array_index_1083333_comb = p33_literal_1076351[p34_array_index_1083284_comb];
  assign p34_array_index_1083334_comb = p33_literal_1076353[p34_array_index_1083285_comb];
  assign p34_array_index_1083335_comb = p33_literal_1076355[p34_array_index_1083286_comb];
  assign p34_res7__178_comb = p33_literal_1076345[p34_res7__177_comb] ^ p34_array_index_1083331_comb ^ p34_array_index_1083332_comb ^ p34_array_index_1083333_comb ^ p34_array_index_1083334_comb ^ p34_array_index_1083335_comb ^ p34_array_index_1083287_comb ^ p33_literal_1076358[p34_array_index_1083288_comb] ^ p34_array_index_1083305_comb ^ p33_literal_1076355[p34_array_index_1083290_comb] ^ p33_literal_1076353[p34_array_index_1083307_comb] ^ p33_literal_1076351[p34_array_index_1083292_comb] ^ p33_literal_1076349[p34_array_index_1083293_comb] ^ p33_literal_1076347[p34_array_index_1083294_comb] ^ p33_literal_1076345[p34_array_index_1083295_comb] ^ p34_array_index_1083296_comb;
  assign p34_array_index_1083345_comb = p33_literal_1076347[p34_res7__177_comb];
  assign p34_array_index_1083346_comb = p33_literal_1076349[p34_res7__176_comb];
  assign p34_array_index_1083347_comb = p33_literal_1076351[p34_array_index_1083283_comb];
  assign p34_array_index_1083348_comb = p33_literal_1076353[p34_array_index_1083284_comb];
  assign p34_array_index_1083349_comb = p33_literal_1076355[p34_array_index_1083285_comb];
  assign p34_res7__179_comb = p33_literal_1076345[p34_res7__178_comb] ^ p34_array_index_1083345_comb ^ p34_array_index_1083346_comb ^ p34_array_index_1083347_comb ^ p34_array_index_1083348_comb ^ p34_array_index_1083349_comb ^ p34_array_index_1083286_comb ^ p33_literal_1076358[p34_array_index_1083287_comb] ^ p34_array_index_1083288_comb ^ p33_literal_1076355[p34_array_index_1083305_comb] ^ p33_literal_1076353[p34_array_index_1083290_comb] ^ p33_literal_1076351[p34_array_index_1083307_comb] ^ p33_literal_1076349[p34_array_index_1083292_comb] ^ p33_literal_1076347[p34_array_index_1083293_comb] ^ p33_literal_1076345[p34_array_index_1083294_comb] ^ p34_array_index_1083295_comb;
  assign p34_array_index_1083360_comb = p33_literal_1076349[p34_res7__177_comb];
  assign p34_array_index_1083361_comb = p33_literal_1076351[p34_res7__176_comb];
  assign p34_array_index_1083362_comb = p33_literal_1076353[p34_array_index_1083283_comb];
  assign p34_array_index_1083363_comb = p33_literal_1076355[p34_array_index_1083284_comb];
  assign p34_res7__180_comb = p33_literal_1076345[p34_res7__179_comb] ^ p33_literal_1076347[p34_res7__178_comb] ^ p34_array_index_1083360_comb ^ p34_array_index_1083361_comb ^ p34_array_index_1083362_comb ^ p34_array_index_1083363_comb ^ p34_array_index_1083285_comb ^ p33_literal_1076358[p34_array_index_1083286_comb] ^ p34_array_index_1083287_comb ^ p34_array_index_1083304_comb ^ p33_literal_1076353[p34_array_index_1083305_comb] ^ p33_literal_1076351[p34_array_index_1083290_comb] ^ p33_literal_1076349[p34_array_index_1083307_comb] ^ p33_literal_1076347[p34_array_index_1083292_comb] ^ p33_literal_1076345[p34_array_index_1083293_comb] ^ p34_array_index_1083294_comb;

  // Registers for pipe stage 34:
  reg [127:0] p34_xor_1082676;
  reg [127:0] p34_xor_1083245;
  reg [7:0] p34_array_index_1083283;
  reg [7:0] p34_array_index_1083284;
  reg [7:0] p34_array_index_1083285;
  reg [7:0] p34_array_index_1083286;
  reg [7:0] p34_array_index_1083287;
  reg [7:0] p34_array_index_1083288;
  reg [7:0] p34_array_index_1083290;
  reg [7:0] p34_array_index_1083292;
  reg [7:0] p34_array_index_1083293;
  reg [7:0] p34_array_index_1083299;
  reg [7:0] p34_array_index_1083300;
  reg [7:0] p34_array_index_1083301;
  reg [7:0] p34_array_index_1083302;
  reg [7:0] p34_array_index_1083303;
  reg [7:0] p34_array_index_1083305;
  reg [7:0] p34_array_index_1083307;
  reg [7:0] p34_res7__176;
  reg [7:0] p34_array_index_1083316;
  reg [7:0] p34_array_index_1083317;
  reg [7:0] p34_array_index_1083318;
  reg [7:0] p34_array_index_1083319;
  reg [7:0] p34_array_index_1083320;
  reg [7:0] p34_array_index_1083321;
  reg [7:0] p34_res7__177;
  reg [7:0] p34_array_index_1083331;
  reg [7:0] p34_array_index_1083332;
  reg [7:0] p34_array_index_1083333;
  reg [7:0] p34_array_index_1083334;
  reg [7:0] p34_array_index_1083335;
  reg [7:0] p34_res7__178;
  reg [7:0] p34_array_index_1083345;
  reg [7:0] p34_array_index_1083346;
  reg [7:0] p34_array_index_1083347;
  reg [7:0] p34_array_index_1083348;
  reg [7:0] p34_array_index_1083349;
  reg [7:0] p34_res7__179;
  reg [7:0] p34_array_index_1083360;
  reg [7:0] p34_array_index_1083361;
  reg [7:0] p34_array_index_1083362;
  reg [7:0] p34_array_index_1083363;
  reg [7:0] p34_res7__180;
  reg [127:0] p34_res__35;
  reg [7:0] p35_arr[256];
  reg [7:0] p35_literal_1076345[256];
  reg [7:0] p35_literal_1076347[256];
  reg [7:0] p35_literal_1076349[256];
  reg [7:0] p35_literal_1076351[256];
  reg [7:0] p35_literal_1076353[256];
  reg [7:0] p35_literal_1076355[256];
  reg [7:0] p35_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p34_xor_1082676 <= p33_xor_1082676;
    p34_xor_1083245 <= p33_xor_1083245;
    p34_array_index_1083283 <= p34_array_index_1083283_comb;
    p34_array_index_1083284 <= p34_array_index_1083284_comb;
    p34_array_index_1083285 <= p34_array_index_1083285_comb;
    p34_array_index_1083286 <= p34_array_index_1083286_comb;
    p34_array_index_1083287 <= p34_array_index_1083287_comb;
    p34_array_index_1083288 <= p34_array_index_1083288_comb;
    p34_array_index_1083290 <= p34_array_index_1083290_comb;
    p34_array_index_1083292 <= p34_array_index_1083292_comb;
    p34_array_index_1083293 <= p34_array_index_1083293_comb;
    p34_array_index_1083299 <= p34_array_index_1083299_comb;
    p34_array_index_1083300 <= p34_array_index_1083300_comb;
    p34_array_index_1083301 <= p34_array_index_1083301_comb;
    p34_array_index_1083302 <= p34_array_index_1083302_comb;
    p34_array_index_1083303 <= p34_array_index_1083303_comb;
    p34_array_index_1083305 <= p34_array_index_1083305_comb;
    p34_array_index_1083307 <= p34_array_index_1083307_comb;
    p34_res7__176 <= p34_res7__176_comb;
    p34_array_index_1083316 <= p34_array_index_1083316_comb;
    p34_array_index_1083317 <= p34_array_index_1083317_comb;
    p34_array_index_1083318 <= p34_array_index_1083318_comb;
    p34_array_index_1083319 <= p34_array_index_1083319_comb;
    p34_array_index_1083320 <= p34_array_index_1083320_comb;
    p34_array_index_1083321 <= p34_array_index_1083321_comb;
    p34_res7__177 <= p34_res7__177_comb;
    p34_array_index_1083331 <= p34_array_index_1083331_comb;
    p34_array_index_1083332 <= p34_array_index_1083332_comb;
    p34_array_index_1083333 <= p34_array_index_1083333_comb;
    p34_array_index_1083334 <= p34_array_index_1083334_comb;
    p34_array_index_1083335 <= p34_array_index_1083335_comb;
    p34_res7__178 <= p34_res7__178_comb;
    p34_array_index_1083345 <= p34_array_index_1083345_comb;
    p34_array_index_1083346 <= p34_array_index_1083346_comb;
    p34_array_index_1083347 <= p34_array_index_1083347_comb;
    p34_array_index_1083348 <= p34_array_index_1083348_comb;
    p34_array_index_1083349 <= p34_array_index_1083349_comb;
    p34_res7__179 <= p34_res7__179_comb;
    p34_array_index_1083360 <= p34_array_index_1083360_comb;
    p34_array_index_1083361 <= p34_array_index_1083361_comb;
    p34_array_index_1083362 <= p34_array_index_1083362_comb;
    p34_array_index_1083363 <= p34_array_index_1083363_comb;
    p34_res7__180 <= p34_res7__180_comb;
    p34_res__35 <= p33_res__35;
    p35_arr <= p34_arr;
    p35_literal_1076345 <= p34_literal_1076345;
    p35_literal_1076347 <= p34_literal_1076347;
    p35_literal_1076349 <= p34_literal_1076349;
    p35_literal_1076351 <= p34_literal_1076351;
    p35_literal_1076353 <= p34_literal_1076353;
    p35_literal_1076355 <= p34_literal_1076355;
    p35_literal_1076358 <= p34_literal_1076358;
  end

  // ===== Pipe stage 35:
  wire [7:0] p35_array_index_1083477_comb;
  wire [7:0] p35_array_index_1083478_comb;
  wire [7:0] p35_array_index_1083479_comb;
  wire [7:0] p35_array_index_1083480_comb;
  wire [7:0] p35_res7__181_comb;
  wire [7:0] p35_array_index_1083491_comb;
  wire [7:0] p35_array_index_1083492_comb;
  wire [7:0] p35_array_index_1083493_comb;
  wire [7:0] p35_res7__182_comb;
  wire [7:0] p35_array_index_1083503_comb;
  wire [7:0] p35_array_index_1083504_comb;
  wire [7:0] p35_array_index_1083505_comb;
  wire [7:0] p35_res7__183_comb;
  wire [7:0] p35_array_index_1083516_comb;
  wire [7:0] p35_array_index_1083517_comb;
  wire [7:0] p35_res7__184_comb;
  wire [7:0] p35_array_index_1083527_comb;
  wire [7:0] p35_array_index_1083528_comb;
  wire [7:0] p35_res7__185_comb;
  wire [7:0] p35_array_index_1083534_comb;
  wire [7:0] p35_array_index_1083535_comb;
  wire [7:0] p35_array_index_1083536_comb;
  wire [7:0] p35_array_index_1083537_comb;
  wire [7:0] p35_array_index_1083538_comb;
  wire [7:0] p35_array_index_1083539_comb;
  wire [7:0] p35_array_index_1083540_comb;
  wire [7:0] p35_array_index_1083541_comb;
  wire [7:0] p35_array_index_1083542_comb;
  assign p35_array_index_1083477_comb = p34_literal_1076349[p34_res7__178];
  assign p35_array_index_1083478_comb = p34_literal_1076351[p34_res7__177];
  assign p35_array_index_1083479_comb = p34_literal_1076353[p34_res7__176];
  assign p35_array_index_1083480_comb = p34_literal_1076355[p34_array_index_1083283];
  assign p35_res7__181_comb = p34_literal_1076345[p34_res7__180] ^ p34_literal_1076347[p34_res7__179] ^ p35_array_index_1083477_comb ^ p35_array_index_1083478_comb ^ p35_array_index_1083479_comb ^ p35_array_index_1083480_comb ^ p34_array_index_1083284 ^ p34_literal_1076358[p34_array_index_1083285] ^ p34_array_index_1083286 ^ p34_array_index_1083321 ^ p34_literal_1076353[p34_array_index_1083288] ^ p34_literal_1076351[p34_array_index_1083305] ^ p34_literal_1076349[p34_array_index_1083290] ^ p34_literal_1076347[p34_array_index_1083307] ^ p34_literal_1076345[p34_array_index_1083292] ^ p34_array_index_1083293;
  assign p35_array_index_1083491_comb = p34_literal_1076351[p34_res7__178];
  assign p35_array_index_1083492_comb = p34_literal_1076353[p34_res7__177];
  assign p35_array_index_1083493_comb = p34_literal_1076355[p34_res7__176];
  assign p35_res7__182_comb = p34_literal_1076345[p35_res7__181_comb] ^ p34_literal_1076347[p34_res7__180] ^ p34_literal_1076349[p34_res7__179] ^ p35_array_index_1083491_comb ^ p35_array_index_1083492_comb ^ p35_array_index_1083493_comb ^ p34_array_index_1083283 ^ p34_literal_1076358[p34_array_index_1083284] ^ p34_array_index_1083285 ^ p34_array_index_1083335 ^ p34_array_index_1083303 ^ p34_literal_1076351[p34_array_index_1083288] ^ p34_literal_1076349[p34_array_index_1083305] ^ p34_literal_1076347[p34_array_index_1083290] ^ p34_literal_1076345[p34_array_index_1083307] ^ p34_array_index_1083292;
  assign p35_array_index_1083503_comb = p34_literal_1076351[p34_res7__179];
  assign p35_array_index_1083504_comb = p34_literal_1076353[p34_res7__178];
  assign p35_array_index_1083505_comb = p34_literal_1076355[p34_res7__177];
  assign p35_res7__183_comb = p34_literal_1076345[p35_res7__182_comb] ^ p34_literal_1076347[p35_res7__181_comb] ^ p34_literal_1076349[p34_res7__180] ^ p35_array_index_1083503_comb ^ p35_array_index_1083504_comb ^ p35_array_index_1083505_comb ^ p34_res7__176 ^ p34_literal_1076358[p34_array_index_1083283] ^ p34_array_index_1083284 ^ p34_array_index_1083349 ^ p34_array_index_1083320 ^ p34_literal_1076351[p34_array_index_1083287] ^ p34_literal_1076349[p34_array_index_1083288] ^ p34_literal_1076347[p34_array_index_1083305] ^ p34_literal_1076345[p34_array_index_1083290] ^ p34_array_index_1083307;
  assign p35_array_index_1083516_comb = p34_literal_1076353[p34_res7__179];
  assign p35_array_index_1083517_comb = p34_literal_1076355[p34_res7__178];
  assign p35_res7__184_comb = p34_literal_1076345[p35_res7__183_comb] ^ p34_literal_1076347[p35_res7__182_comb] ^ p34_literal_1076349[p35_res7__181_comb] ^ p34_literal_1076351[p34_res7__180] ^ p35_array_index_1083516_comb ^ p35_array_index_1083517_comb ^ p34_res7__177 ^ p34_literal_1076358[p34_res7__176] ^ p34_array_index_1083283 ^ p34_array_index_1083363 ^ p34_array_index_1083334 ^ p34_array_index_1083302 ^ p34_literal_1076349[p34_array_index_1083287] ^ p34_literal_1076347[p34_array_index_1083288] ^ p34_literal_1076345[p34_array_index_1083305] ^ p34_array_index_1083290;
  assign p35_array_index_1083527_comb = p34_literal_1076353[p34_res7__180];
  assign p35_array_index_1083528_comb = p34_literal_1076355[p34_res7__179];
  assign p35_res7__185_comb = p34_literal_1076345[p35_res7__184_comb] ^ p34_literal_1076347[p35_res7__183_comb] ^ p34_literal_1076349[p35_res7__182_comb] ^ p34_literal_1076351[p35_res7__181_comb] ^ p35_array_index_1083527_comb ^ p35_array_index_1083528_comb ^ p34_res7__178 ^ p34_literal_1076358[p34_res7__177] ^ p34_res7__176 ^ p35_array_index_1083480_comb ^ p34_array_index_1083348 ^ p34_array_index_1083319 ^ p34_literal_1076349[p34_array_index_1083286] ^ p34_literal_1076347[p34_array_index_1083287] ^ p34_literal_1076345[p34_array_index_1083288] ^ p34_array_index_1083305;
  assign p35_array_index_1083534_comb = p34_literal_1076345[p35_res7__185_comb];
  assign p35_array_index_1083535_comb = p34_literal_1076347[p35_res7__184_comb];
  assign p35_array_index_1083536_comb = p34_literal_1076349[p35_res7__183_comb];
  assign p35_array_index_1083537_comb = p34_literal_1076351[p35_res7__182_comb];
  assign p35_array_index_1083538_comb = p34_literal_1076353[p35_res7__181_comb];
  assign p35_array_index_1083539_comb = p34_literal_1076355[p34_res7__180];
  assign p35_array_index_1083540_comb = p34_literal_1076358[p34_res7__178];
  assign p35_array_index_1083541_comb = p34_literal_1076347[p34_array_index_1083286];
  assign p35_array_index_1083542_comb = p34_literal_1076345[p34_array_index_1083287];

  // Registers for pipe stage 35:
  reg [127:0] p35_xor_1082676;
  reg [127:0] p35_xor_1083245;
  reg [7:0] p35_array_index_1083283;
  reg [7:0] p35_array_index_1083284;
  reg [7:0] p35_array_index_1083285;
  reg [7:0] p35_array_index_1083286;
  reg [7:0] p35_array_index_1083287;
  reg [7:0] p35_array_index_1083288;
  reg [7:0] p35_array_index_1083299;
  reg [7:0] p35_array_index_1083300;
  reg [7:0] p35_array_index_1083301;
  reg [7:0] p35_res7__176;
  reg [7:0] p35_array_index_1083316;
  reg [7:0] p35_array_index_1083317;
  reg [7:0] p35_array_index_1083318;
  reg [7:0] p35_res7__177;
  reg [7:0] p35_array_index_1083331;
  reg [7:0] p35_array_index_1083332;
  reg [7:0] p35_array_index_1083333;
  reg [7:0] p35_res7__178;
  reg [7:0] p35_array_index_1083345;
  reg [7:0] p35_array_index_1083346;
  reg [7:0] p35_array_index_1083347;
  reg [7:0] p35_res7__179;
  reg [7:0] p35_array_index_1083360;
  reg [7:0] p35_array_index_1083361;
  reg [7:0] p35_array_index_1083362;
  reg [7:0] p35_res7__180;
  reg [7:0] p35_array_index_1083477;
  reg [7:0] p35_array_index_1083478;
  reg [7:0] p35_array_index_1083479;
  reg [7:0] p35_res7__181;
  reg [7:0] p35_array_index_1083491;
  reg [7:0] p35_array_index_1083492;
  reg [7:0] p35_array_index_1083493;
  reg [7:0] p35_res7__182;
  reg [7:0] p35_array_index_1083503;
  reg [7:0] p35_array_index_1083504;
  reg [7:0] p35_array_index_1083505;
  reg [7:0] p35_res7__183;
  reg [7:0] p35_array_index_1083516;
  reg [7:0] p35_array_index_1083517;
  reg [7:0] p35_res7__184;
  reg [7:0] p35_array_index_1083527;
  reg [7:0] p35_array_index_1083528;
  reg [7:0] p35_res7__185;
  reg [7:0] p35_array_index_1083534;
  reg [7:0] p35_array_index_1083535;
  reg [7:0] p35_array_index_1083536;
  reg [7:0] p35_array_index_1083537;
  reg [7:0] p35_array_index_1083538;
  reg [7:0] p35_array_index_1083539;
  reg [7:0] p35_array_index_1083540;
  reg [7:0] p35_array_index_1083541;
  reg [7:0] p35_array_index_1083542;
  reg [127:0] p35_res__35;
  reg [7:0] p36_arr[256];
  reg [7:0] p36_literal_1076345[256];
  reg [7:0] p36_literal_1076347[256];
  reg [7:0] p36_literal_1076349[256];
  reg [7:0] p36_literal_1076351[256];
  reg [7:0] p36_literal_1076353[256];
  reg [7:0] p36_literal_1076355[256];
  reg [7:0] p36_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p35_xor_1082676 <= p34_xor_1082676;
    p35_xor_1083245 <= p34_xor_1083245;
    p35_array_index_1083283 <= p34_array_index_1083283;
    p35_array_index_1083284 <= p34_array_index_1083284;
    p35_array_index_1083285 <= p34_array_index_1083285;
    p35_array_index_1083286 <= p34_array_index_1083286;
    p35_array_index_1083287 <= p34_array_index_1083287;
    p35_array_index_1083288 <= p34_array_index_1083288;
    p35_array_index_1083299 <= p34_array_index_1083299;
    p35_array_index_1083300 <= p34_array_index_1083300;
    p35_array_index_1083301 <= p34_array_index_1083301;
    p35_res7__176 <= p34_res7__176;
    p35_array_index_1083316 <= p34_array_index_1083316;
    p35_array_index_1083317 <= p34_array_index_1083317;
    p35_array_index_1083318 <= p34_array_index_1083318;
    p35_res7__177 <= p34_res7__177;
    p35_array_index_1083331 <= p34_array_index_1083331;
    p35_array_index_1083332 <= p34_array_index_1083332;
    p35_array_index_1083333 <= p34_array_index_1083333;
    p35_res7__178 <= p34_res7__178;
    p35_array_index_1083345 <= p34_array_index_1083345;
    p35_array_index_1083346 <= p34_array_index_1083346;
    p35_array_index_1083347 <= p34_array_index_1083347;
    p35_res7__179 <= p34_res7__179;
    p35_array_index_1083360 <= p34_array_index_1083360;
    p35_array_index_1083361 <= p34_array_index_1083361;
    p35_array_index_1083362 <= p34_array_index_1083362;
    p35_res7__180 <= p34_res7__180;
    p35_array_index_1083477 <= p35_array_index_1083477_comb;
    p35_array_index_1083478 <= p35_array_index_1083478_comb;
    p35_array_index_1083479 <= p35_array_index_1083479_comb;
    p35_res7__181 <= p35_res7__181_comb;
    p35_array_index_1083491 <= p35_array_index_1083491_comb;
    p35_array_index_1083492 <= p35_array_index_1083492_comb;
    p35_array_index_1083493 <= p35_array_index_1083493_comb;
    p35_res7__182 <= p35_res7__182_comb;
    p35_array_index_1083503 <= p35_array_index_1083503_comb;
    p35_array_index_1083504 <= p35_array_index_1083504_comb;
    p35_array_index_1083505 <= p35_array_index_1083505_comb;
    p35_res7__183 <= p35_res7__183_comb;
    p35_array_index_1083516 <= p35_array_index_1083516_comb;
    p35_array_index_1083517 <= p35_array_index_1083517_comb;
    p35_res7__184 <= p35_res7__184_comb;
    p35_array_index_1083527 <= p35_array_index_1083527_comb;
    p35_array_index_1083528 <= p35_array_index_1083528_comb;
    p35_res7__185 <= p35_res7__185_comb;
    p35_array_index_1083534 <= p35_array_index_1083534_comb;
    p35_array_index_1083535 <= p35_array_index_1083535_comb;
    p35_array_index_1083536 <= p35_array_index_1083536_comb;
    p35_array_index_1083537 <= p35_array_index_1083537_comb;
    p35_array_index_1083538 <= p35_array_index_1083538_comb;
    p35_array_index_1083539 <= p35_array_index_1083539_comb;
    p35_array_index_1083540 <= p35_array_index_1083540_comb;
    p35_array_index_1083541 <= p35_array_index_1083541_comb;
    p35_array_index_1083542 <= p35_array_index_1083542_comb;
    p35_res__35 <= p34_res__35;
    p36_arr <= p35_arr;
    p36_literal_1076345 <= p35_literal_1076345;
    p36_literal_1076347 <= p35_literal_1076347;
    p36_literal_1076349 <= p35_literal_1076349;
    p36_literal_1076351 <= p35_literal_1076351;
    p36_literal_1076353 <= p35_literal_1076353;
    p36_literal_1076355 <= p35_literal_1076355;
    p36_literal_1076358 <= p35_literal_1076358;
  end

  // ===== Pipe stage 36:
  wire [7:0] p36_res7__186_comb;
  wire [7:0] p36_array_index_1083677_comb;
  wire [7:0] p36_res7__187_comb;
  wire [7:0] p36_res7__188_comb;
  wire [7:0] p36_res7__189_comb;
  wire [7:0] p36_res7__190_comb;
  wire [7:0] p36_res7__191_comb;
  wire [127:0] p36_res__11_comb;
  wire [127:0] p36_xor_1083717_comb;
  assign p36_res7__186_comb = p35_array_index_1083534 ^ p35_array_index_1083535 ^ p35_array_index_1083536 ^ p35_array_index_1083537 ^ p35_array_index_1083538 ^ p35_array_index_1083539 ^ p35_res7__179 ^ p35_array_index_1083540 ^ p35_res7__177 ^ p35_array_index_1083493 ^ p35_array_index_1083362 ^ p35_array_index_1083333 ^ p35_array_index_1083301 ^ p35_array_index_1083541 ^ p35_array_index_1083542 ^ p35_array_index_1083288;
  assign p36_array_index_1083677_comb = p35_literal_1076355[p35_res7__181];
  assign p36_res7__187_comb = p35_literal_1076345[p36_res7__186_comb] ^ p35_literal_1076347[p35_res7__185] ^ p35_literal_1076349[p35_res7__184] ^ p35_literal_1076351[p35_res7__183] ^ p35_literal_1076353[p35_res7__182] ^ p36_array_index_1083677_comb ^ p35_res7__180 ^ p35_literal_1076358[p35_res7__179] ^ p35_res7__178 ^ p35_array_index_1083505 ^ p35_array_index_1083479 ^ p35_array_index_1083347 ^ p35_array_index_1083318 ^ p35_literal_1076347[p35_array_index_1083285] ^ p35_literal_1076345[p35_array_index_1083286] ^ p35_array_index_1083287;
  assign p36_res7__188_comb = p35_literal_1076345[p36_res7__187_comb] ^ p35_literal_1076347[p36_res7__186_comb] ^ p35_literal_1076349[p35_res7__185] ^ p35_literal_1076351[p35_res7__184] ^ p35_literal_1076353[p35_res7__183] ^ p35_literal_1076355[p35_res7__182] ^ p35_res7__181 ^ p35_literal_1076358[p35_res7__180] ^ p35_res7__179 ^ p35_array_index_1083517 ^ p35_array_index_1083492 ^ p35_array_index_1083361 ^ p35_array_index_1083332 ^ p35_array_index_1083300 ^ p35_literal_1076345[p35_array_index_1083285] ^ p35_array_index_1083286;
  assign p36_res7__189_comb = p35_literal_1076345[p36_res7__188_comb] ^ p35_literal_1076347[p36_res7__187_comb] ^ p35_literal_1076349[p36_res7__186_comb] ^ p35_literal_1076351[p35_res7__185] ^ p35_literal_1076353[p35_res7__184] ^ p35_literal_1076355[p35_res7__183] ^ p35_res7__182 ^ p35_literal_1076358[p35_res7__181] ^ p35_res7__180 ^ p35_array_index_1083528 ^ p35_array_index_1083504 ^ p35_array_index_1083478 ^ p35_array_index_1083346 ^ p35_array_index_1083317 ^ p35_literal_1076345[p35_array_index_1083284] ^ p35_array_index_1083285;
  assign p36_res7__190_comb = p35_literal_1076345[p36_res7__189_comb] ^ p35_literal_1076347[p36_res7__188_comb] ^ p35_literal_1076349[p36_res7__187_comb] ^ p35_literal_1076351[p36_res7__186_comb] ^ p35_literal_1076353[p35_res7__185] ^ p35_literal_1076355[p35_res7__184] ^ p35_res7__183 ^ p35_literal_1076358[p35_res7__182] ^ p35_res7__181 ^ p35_array_index_1083539 ^ p35_array_index_1083516 ^ p35_array_index_1083491 ^ p35_array_index_1083360 ^ p35_array_index_1083331 ^ p35_array_index_1083299 ^ p35_array_index_1083284;
  assign p36_res7__191_comb = p35_literal_1076345[p36_res7__190_comb] ^ p35_literal_1076347[p36_res7__189_comb] ^ p35_literal_1076349[p36_res7__188_comb] ^ p35_literal_1076351[p36_res7__187_comb] ^ p35_literal_1076353[p36_res7__186_comb] ^ p35_literal_1076355[p35_res7__185] ^ p35_res7__184 ^ p35_literal_1076358[p35_res7__183] ^ p35_res7__182 ^ p36_array_index_1083677_comb ^ p35_array_index_1083527 ^ p35_array_index_1083503 ^ p35_array_index_1083477 ^ p35_array_index_1083345 ^ p35_array_index_1083316 ^ p35_array_index_1083283;
  assign p36_res__11_comb = {p36_res7__191_comb, p36_res7__190_comb, p36_res7__189_comb, p36_res7__188_comb, p36_res7__187_comb, p36_res7__186_comb, p35_res7__185, p35_res7__184, p35_res7__183, p35_res7__182, p35_res7__181, p35_res7__180, p35_res7__179, p35_res7__178, p35_res7__177, p35_res7__176};
  assign p36_xor_1083717_comb = p36_res__11_comb ^ p35_xor_1082676;

  // Registers for pipe stage 36:
  reg [127:0] p36_xor_1083245;
  reg [127:0] p36_xor_1083717;
  reg [127:0] p36_res__35;
  reg [7:0] p37_arr[256];
  reg [7:0] p37_literal_1076345[256];
  reg [7:0] p37_literal_1076347[256];
  reg [7:0] p37_literal_1076349[256];
  reg [7:0] p37_literal_1076351[256];
  reg [7:0] p37_literal_1076353[256];
  reg [7:0] p37_literal_1076355[256];
  reg [7:0] p37_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p36_xor_1083245 <= p35_xor_1083245;
    p36_xor_1083717 <= p36_xor_1083717_comb;
    p36_res__35 <= p35_res__35;
    p37_arr <= p36_arr;
    p37_literal_1076345 <= p36_literal_1076345;
    p37_literal_1076347 <= p36_literal_1076347;
    p37_literal_1076349 <= p36_literal_1076349;
    p37_literal_1076351 <= p36_literal_1076351;
    p37_literal_1076353 <= p36_literal_1076353;
    p37_literal_1076355 <= p36_literal_1076355;
    p37_literal_1076358 <= p36_literal_1076358;
  end

  // ===== Pipe stage 37:
  wire [127:0] p37_addedKey__53_comb;
  wire [7:0] p37_array_index_1083755_comb;
  wire [7:0] p37_array_index_1083756_comb;
  wire [7:0] p37_array_index_1083757_comb;
  wire [7:0] p37_array_index_1083758_comb;
  wire [7:0] p37_array_index_1083759_comb;
  wire [7:0] p37_array_index_1083760_comb;
  wire [7:0] p37_array_index_1083762_comb;
  wire [7:0] p37_array_index_1083764_comb;
  wire [7:0] p37_array_index_1083765_comb;
  wire [7:0] p37_array_index_1083766_comb;
  wire [7:0] p37_array_index_1083767_comb;
  wire [7:0] p37_array_index_1083768_comb;
  wire [7:0] p37_array_index_1083769_comb;
  wire [7:0] p37_array_index_1083771_comb;
  wire [7:0] p37_array_index_1083772_comb;
  wire [7:0] p37_array_index_1083773_comb;
  wire [7:0] p37_array_index_1083774_comb;
  wire [7:0] p37_array_index_1083775_comb;
  wire [7:0] p37_array_index_1083776_comb;
  wire [7:0] p37_array_index_1083777_comb;
  wire [7:0] p37_array_index_1083779_comb;
  wire [7:0] p37_res7__192_comb;
  wire [7:0] p37_array_index_1083788_comb;
  wire [7:0] p37_array_index_1083789_comb;
  wire [7:0] p37_array_index_1083790_comb;
  wire [7:0] p37_array_index_1083791_comb;
  wire [7:0] p37_array_index_1083792_comb;
  wire [7:0] p37_array_index_1083793_comb;
  wire [7:0] p37_res7__193_comb;
  wire [7:0] p37_array_index_1083803_comb;
  wire [7:0] p37_array_index_1083804_comb;
  wire [7:0] p37_array_index_1083805_comb;
  wire [7:0] p37_array_index_1083806_comb;
  wire [7:0] p37_array_index_1083807_comb;
  wire [7:0] p37_res7__194_comb;
  wire [7:0] p37_array_index_1083817_comb;
  wire [7:0] p37_array_index_1083818_comb;
  wire [7:0] p37_array_index_1083819_comb;
  wire [7:0] p37_array_index_1083820_comb;
  wire [7:0] p37_array_index_1083821_comb;
  wire [7:0] p37_res7__195_comb;
  wire [7:0] p37_array_index_1083832_comb;
  wire [7:0] p37_array_index_1083833_comb;
  wire [7:0] p37_array_index_1083834_comb;
  wire [7:0] p37_array_index_1083835_comb;
  wire [7:0] p37_res7__196_comb;
  assign p37_addedKey__53_comb = p36_xor_1083717 ^ 128'he336_5b6f_f9ae_0794_4740_add0_087b_ab0d;
  assign p37_array_index_1083755_comb = p36_arr[p37_addedKey__53_comb[127:120]];
  assign p37_array_index_1083756_comb = p36_arr[p37_addedKey__53_comb[119:112]];
  assign p37_array_index_1083757_comb = p36_arr[p37_addedKey__53_comb[111:104]];
  assign p37_array_index_1083758_comb = p36_arr[p37_addedKey__53_comb[103:96]];
  assign p37_array_index_1083759_comb = p36_arr[p37_addedKey__53_comb[95:88]];
  assign p37_array_index_1083760_comb = p36_arr[p37_addedKey__53_comb[87:80]];
  assign p37_array_index_1083762_comb = p36_arr[p37_addedKey__53_comb[71:64]];
  assign p37_array_index_1083764_comb = p36_arr[p37_addedKey__53_comb[55:48]];
  assign p37_array_index_1083765_comb = p36_arr[p37_addedKey__53_comb[47:40]];
  assign p37_array_index_1083766_comb = p36_arr[p37_addedKey__53_comb[39:32]];
  assign p37_array_index_1083767_comb = p36_arr[p37_addedKey__53_comb[31:24]];
  assign p37_array_index_1083768_comb = p36_arr[p37_addedKey__53_comb[23:16]];
  assign p37_array_index_1083769_comb = p36_arr[p37_addedKey__53_comb[15:8]];
  assign p37_array_index_1083771_comb = p36_literal_1076345[p37_array_index_1083755_comb];
  assign p37_array_index_1083772_comb = p36_literal_1076347[p37_array_index_1083756_comb];
  assign p37_array_index_1083773_comb = p36_literal_1076349[p37_array_index_1083757_comb];
  assign p37_array_index_1083774_comb = p36_literal_1076351[p37_array_index_1083758_comb];
  assign p37_array_index_1083775_comb = p36_literal_1076353[p37_array_index_1083759_comb];
  assign p37_array_index_1083776_comb = p36_literal_1076355[p37_array_index_1083760_comb];
  assign p37_array_index_1083777_comb = p36_arr[p37_addedKey__53_comb[79:72]];
  assign p37_array_index_1083779_comb = p36_arr[p37_addedKey__53_comb[63:56]];
  assign p37_res7__192_comb = p37_array_index_1083771_comb ^ p37_array_index_1083772_comb ^ p37_array_index_1083773_comb ^ p37_array_index_1083774_comb ^ p37_array_index_1083775_comb ^ p37_array_index_1083776_comb ^ p37_array_index_1083777_comb ^ p36_literal_1076358[p37_array_index_1083762_comb] ^ p37_array_index_1083779_comb ^ p36_literal_1076355[p37_array_index_1083764_comb] ^ p36_literal_1076353[p37_array_index_1083765_comb] ^ p36_literal_1076351[p37_array_index_1083766_comb] ^ p36_literal_1076349[p37_array_index_1083767_comb] ^ p36_literal_1076347[p37_array_index_1083768_comb] ^ p36_literal_1076345[p37_array_index_1083769_comb] ^ p36_arr[p37_addedKey__53_comb[7:0]];
  assign p37_array_index_1083788_comb = p36_literal_1076345[p37_res7__192_comb];
  assign p37_array_index_1083789_comb = p36_literal_1076347[p37_array_index_1083755_comb];
  assign p37_array_index_1083790_comb = p36_literal_1076349[p37_array_index_1083756_comb];
  assign p37_array_index_1083791_comb = p36_literal_1076351[p37_array_index_1083757_comb];
  assign p37_array_index_1083792_comb = p36_literal_1076353[p37_array_index_1083758_comb];
  assign p37_array_index_1083793_comb = p36_literal_1076355[p37_array_index_1083759_comb];
  assign p37_res7__193_comb = p37_array_index_1083788_comb ^ p37_array_index_1083789_comb ^ p37_array_index_1083790_comb ^ p37_array_index_1083791_comb ^ p37_array_index_1083792_comb ^ p37_array_index_1083793_comb ^ p37_array_index_1083760_comb ^ p36_literal_1076358[p37_array_index_1083777_comb] ^ p37_array_index_1083762_comb ^ p36_literal_1076355[p37_array_index_1083779_comb] ^ p36_literal_1076353[p37_array_index_1083764_comb] ^ p36_literal_1076351[p37_array_index_1083765_comb] ^ p36_literal_1076349[p37_array_index_1083766_comb] ^ p36_literal_1076347[p37_array_index_1083767_comb] ^ p36_literal_1076345[p37_array_index_1083768_comb] ^ p37_array_index_1083769_comb;
  assign p37_array_index_1083803_comb = p36_literal_1076347[p37_res7__192_comb];
  assign p37_array_index_1083804_comb = p36_literal_1076349[p37_array_index_1083755_comb];
  assign p37_array_index_1083805_comb = p36_literal_1076351[p37_array_index_1083756_comb];
  assign p37_array_index_1083806_comb = p36_literal_1076353[p37_array_index_1083757_comb];
  assign p37_array_index_1083807_comb = p36_literal_1076355[p37_array_index_1083758_comb];
  assign p37_res7__194_comb = p36_literal_1076345[p37_res7__193_comb] ^ p37_array_index_1083803_comb ^ p37_array_index_1083804_comb ^ p37_array_index_1083805_comb ^ p37_array_index_1083806_comb ^ p37_array_index_1083807_comb ^ p37_array_index_1083759_comb ^ p36_literal_1076358[p37_array_index_1083760_comb] ^ p37_array_index_1083777_comb ^ p36_literal_1076355[p37_array_index_1083762_comb] ^ p36_literal_1076353[p37_array_index_1083779_comb] ^ p36_literal_1076351[p37_array_index_1083764_comb] ^ p36_literal_1076349[p37_array_index_1083765_comb] ^ p36_literal_1076347[p37_array_index_1083766_comb] ^ p36_literal_1076345[p37_array_index_1083767_comb] ^ p37_array_index_1083768_comb;
  assign p37_array_index_1083817_comb = p36_literal_1076347[p37_res7__193_comb];
  assign p37_array_index_1083818_comb = p36_literal_1076349[p37_res7__192_comb];
  assign p37_array_index_1083819_comb = p36_literal_1076351[p37_array_index_1083755_comb];
  assign p37_array_index_1083820_comb = p36_literal_1076353[p37_array_index_1083756_comb];
  assign p37_array_index_1083821_comb = p36_literal_1076355[p37_array_index_1083757_comb];
  assign p37_res7__195_comb = p36_literal_1076345[p37_res7__194_comb] ^ p37_array_index_1083817_comb ^ p37_array_index_1083818_comb ^ p37_array_index_1083819_comb ^ p37_array_index_1083820_comb ^ p37_array_index_1083821_comb ^ p37_array_index_1083758_comb ^ p36_literal_1076358[p37_array_index_1083759_comb] ^ p37_array_index_1083760_comb ^ p36_literal_1076355[p37_array_index_1083777_comb] ^ p36_literal_1076353[p37_array_index_1083762_comb] ^ p36_literal_1076351[p37_array_index_1083779_comb] ^ p36_literal_1076349[p37_array_index_1083764_comb] ^ p36_literal_1076347[p37_array_index_1083765_comb] ^ p36_literal_1076345[p37_array_index_1083766_comb] ^ p37_array_index_1083767_comb;
  assign p37_array_index_1083832_comb = p36_literal_1076349[p37_res7__193_comb];
  assign p37_array_index_1083833_comb = p36_literal_1076351[p37_res7__192_comb];
  assign p37_array_index_1083834_comb = p36_literal_1076353[p37_array_index_1083755_comb];
  assign p37_array_index_1083835_comb = p36_literal_1076355[p37_array_index_1083756_comb];
  assign p37_res7__196_comb = p36_literal_1076345[p37_res7__195_comb] ^ p36_literal_1076347[p37_res7__194_comb] ^ p37_array_index_1083832_comb ^ p37_array_index_1083833_comb ^ p37_array_index_1083834_comb ^ p37_array_index_1083835_comb ^ p37_array_index_1083757_comb ^ p36_literal_1076358[p37_array_index_1083758_comb] ^ p37_array_index_1083759_comb ^ p37_array_index_1083776_comb ^ p36_literal_1076353[p37_array_index_1083777_comb] ^ p36_literal_1076351[p37_array_index_1083762_comb] ^ p36_literal_1076349[p37_array_index_1083779_comb] ^ p36_literal_1076347[p37_array_index_1083764_comb] ^ p36_literal_1076345[p37_array_index_1083765_comb] ^ p37_array_index_1083766_comb;

  // Registers for pipe stage 37:
  reg [127:0] p37_xor_1083245;
  reg [127:0] p37_xor_1083717;
  reg [7:0] p37_array_index_1083755;
  reg [7:0] p37_array_index_1083756;
  reg [7:0] p37_array_index_1083757;
  reg [7:0] p37_array_index_1083758;
  reg [7:0] p37_array_index_1083759;
  reg [7:0] p37_array_index_1083760;
  reg [7:0] p37_array_index_1083762;
  reg [7:0] p37_array_index_1083764;
  reg [7:0] p37_array_index_1083765;
  reg [7:0] p37_array_index_1083771;
  reg [7:0] p37_array_index_1083772;
  reg [7:0] p37_array_index_1083773;
  reg [7:0] p37_array_index_1083774;
  reg [7:0] p37_array_index_1083775;
  reg [7:0] p37_array_index_1083777;
  reg [7:0] p37_array_index_1083779;
  reg [7:0] p37_res7__192;
  reg [7:0] p37_array_index_1083788;
  reg [7:0] p37_array_index_1083789;
  reg [7:0] p37_array_index_1083790;
  reg [7:0] p37_array_index_1083791;
  reg [7:0] p37_array_index_1083792;
  reg [7:0] p37_array_index_1083793;
  reg [7:0] p37_res7__193;
  reg [7:0] p37_array_index_1083803;
  reg [7:0] p37_array_index_1083804;
  reg [7:0] p37_array_index_1083805;
  reg [7:0] p37_array_index_1083806;
  reg [7:0] p37_array_index_1083807;
  reg [7:0] p37_res7__194;
  reg [7:0] p37_array_index_1083817;
  reg [7:0] p37_array_index_1083818;
  reg [7:0] p37_array_index_1083819;
  reg [7:0] p37_array_index_1083820;
  reg [7:0] p37_array_index_1083821;
  reg [7:0] p37_res7__195;
  reg [7:0] p37_array_index_1083832;
  reg [7:0] p37_array_index_1083833;
  reg [7:0] p37_array_index_1083834;
  reg [7:0] p37_array_index_1083835;
  reg [7:0] p37_res7__196;
  reg [127:0] p37_res__35;
  reg [7:0] p38_arr[256];
  reg [7:0] p38_literal_1076345[256];
  reg [7:0] p38_literal_1076347[256];
  reg [7:0] p38_literal_1076349[256];
  reg [7:0] p38_literal_1076351[256];
  reg [7:0] p38_literal_1076353[256];
  reg [7:0] p38_literal_1076355[256];
  reg [7:0] p38_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p37_xor_1083245 <= p36_xor_1083245;
    p37_xor_1083717 <= p36_xor_1083717;
    p37_array_index_1083755 <= p37_array_index_1083755_comb;
    p37_array_index_1083756 <= p37_array_index_1083756_comb;
    p37_array_index_1083757 <= p37_array_index_1083757_comb;
    p37_array_index_1083758 <= p37_array_index_1083758_comb;
    p37_array_index_1083759 <= p37_array_index_1083759_comb;
    p37_array_index_1083760 <= p37_array_index_1083760_comb;
    p37_array_index_1083762 <= p37_array_index_1083762_comb;
    p37_array_index_1083764 <= p37_array_index_1083764_comb;
    p37_array_index_1083765 <= p37_array_index_1083765_comb;
    p37_array_index_1083771 <= p37_array_index_1083771_comb;
    p37_array_index_1083772 <= p37_array_index_1083772_comb;
    p37_array_index_1083773 <= p37_array_index_1083773_comb;
    p37_array_index_1083774 <= p37_array_index_1083774_comb;
    p37_array_index_1083775 <= p37_array_index_1083775_comb;
    p37_array_index_1083777 <= p37_array_index_1083777_comb;
    p37_array_index_1083779 <= p37_array_index_1083779_comb;
    p37_res7__192 <= p37_res7__192_comb;
    p37_array_index_1083788 <= p37_array_index_1083788_comb;
    p37_array_index_1083789 <= p37_array_index_1083789_comb;
    p37_array_index_1083790 <= p37_array_index_1083790_comb;
    p37_array_index_1083791 <= p37_array_index_1083791_comb;
    p37_array_index_1083792 <= p37_array_index_1083792_comb;
    p37_array_index_1083793 <= p37_array_index_1083793_comb;
    p37_res7__193 <= p37_res7__193_comb;
    p37_array_index_1083803 <= p37_array_index_1083803_comb;
    p37_array_index_1083804 <= p37_array_index_1083804_comb;
    p37_array_index_1083805 <= p37_array_index_1083805_comb;
    p37_array_index_1083806 <= p37_array_index_1083806_comb;
    p37_array_index_1083807 <= p37_array_index_1083807_comb;
    p37_res7__194 <= p37_res7__194_comb;
    p37_array_index_1083817 <= p37_array_index_1083817_comb;
    p37_array_index_1083818 <= p37_array_index_1083818_comb;
    p37_array_index_1083819 <= p37_array_index_1083819_comb;
    p37_array_index_1083820 <= p37_array_index_1083820_comb;
    p37_array_index_1083821 <= p37_array_index_1083821_comb;
    p37_res7__195 <= p37_res7__195_comb;
    p37_array_index_1083832 <= p37_array_index_1083832_comb;
    p37_array_index_1083833 <= p37_array_index_1083833_comb;
    p37_array_index_1083834 <= p37_array_index_1083834_comb;
    p37_array_index_1083835 <= p37_array_index_1083835_comb;
    p37_res7__196 <= p37_res7__196_comb;
    p37_res__35 <= p36_res__35;
    p38_arr <= p37_arr;
    p38_literal_1076345 <= p37_literal_1076345;
    p38_literal_1076347 <= p37_literal_1076347;
    p38_literal_1076349 <= p37_literal_1076349;
    p38_literal_1076351 <= p37_literal_1076351;
    p38_literal_1076353 <= p37_literal_1076353;
    p38_literal_1076355 <= p37_literal_1076355;
    p38_literal_1076358 <= p37_literal_1076358;
  end

  // ===== Pipe stage 38:
  wire [7:0] p38_array_index_1083949_comb;
  wire [7:0] p38_array_index_1083950_comb;
  wire [7:0] p38_array_index_1083951_comb;
  wire [7:0] p38_array_index_1083952_comb;
  wire [7:0] p38_res7__197_comb;
  wire [7:0] p38_array_index_1083963_comb;
  wire [7:0] p38_array_index_1083964_comb;
  wire [7:0] p38_array_index_1083965_comb;
  wire [7:0] p38_res7__198_comb;
  wire [7:0] p38_array_index_1083975_comb;
  wire [7:0] p38_array_index_1083976_comb;
  wire [7:0] p38_array_index_1083977_comb;
  wire [7:0] p38_res7__199_comb;
  wire [7:0] p38_array_index_1083988_comb;
  wire [7:0] p38_array_index_1083989_comb;
  wire [7:0] p38_res7__200_comb;
  wire [7:0] p38_array_index_1083999_comb;
  wire [7:0] p38_array_index_1084000_comb;
  wire [7:0] p38_res7__201_comb;
  wire [7:0] p38_array_index_1084006_comb;
  wire [7:0] p38_array_index_1084007_comb;
  wire [7:0] p38_array_index_1084008_comb;
  wire [7:0] p38_array_index_1084009_comb;
  wire [7:0] p38_array_index_1084010_comb;
  wire [7:0] p38_array_index_1084011_comb;
  wire [7:0] p38_array_index_1084012_comb;
  wire [7:0] p38_array_index_1084013_comb;
  wire [7:0] p38_array_index_1084014_comb;
  assign p38_array_index_1083949_comb = p37_literal_1076349[p37_res7__194];
  assign p38_array_index_1083950_comb = p37_literal_1076351[p37_res7__193];
  assign p38_array_index_1083951_comb = p37_literal_1076353[p37_res7__192];
  assign p38_array_index_1083952_comb = p37_literal_1076355[p37_array_index_1083755];
  assign p38_res7__197_comb = p37_literal_1076345[p37_res7__196] ^ p37_literal_1076347[p37_res7__195] ^ p38_array_index_1083949_comb ^ p38_array_index_1083950_comb ^ p38_array_index_1083951_comb ^ p38_array_index_1083952_comb ^ p37_array_index_1083756 ^ p37_literal_1076358[p37_array_index_1083757] ^ p37_array_index_1083758 ^ p37_array_index_1083793 ^ p37_literal_1076353[p37_array_index_1083760] ^ p37_literal_1076351[p37_array_index_1083777] ^ p37_literal_1076349[p37_array_index_1083762] ^ p37_literal_1076347[p37_array_index_1083779] ^ p37_literal_1076345[p37_array_index_1083764] ^ p37_array_index_1083765;
  assign p38_array_index_1083963_comb = p37_literal_1076351[p37_res7__194];
  assign p38_array_index_1083964_comb = p37_literal_1076353[p37_res7__193];
  assign p38_array_index_1083965_comb = p37_literal_1076355[p37_res7__192];
  assign p38_res7__198_comb = p37_literal_1076345[p38_res7__197_comb] ^ p37_literal_1076347[p37_res7__196] ^ p37_literal_1076349[p37_res7__195] ^ p38_array_index_1083963_comb ^ p38_array_index_1083964_comb ^ p38_array_index_1083965_comb ^ p37_array_index_1083755 ^ p37_literal_1076358[p37_array_index_1083756] ^ p37_array_index_1083757 ^ p37_array_index_1083807 ^ p37_array_index_1083775 ^ p37_literal_1076351[p37_array_index_1083760] ^ p37_literal_1076349[p37_array_index_1083777] ^ p37_literal_1076347[p37_array_index_1083762] ^ p37_literal_1076345[p37_array_index_1083779] ^ p37_array_index_1083764;
  assign p38_array_index_1083975_comb = p37_literal_1076351[p37_res7__195];
  assign p38_array_index_1083976_comb = p37_literal_1076353[p37_res7__194];
  assign p38_array_index_1083977_comb = p37_literal_1076355[p37_res7__193];
  assign p38_res7__199_comb = p37_literal_1076345[p38_res7__198_comb] ^ p37_literal_1076347[p38_res7__197_comb] ^ p37_literal_1076349[p37_res7__196] ^ p38_array_index_1083975_comb ^ p38_array_index_1083976_comb ^ p38_array_index_1083977_comb ^ p37_res7__192 ^ p37_literal_1076358[p37_array_index_1083755] ^ p37_array_index_1083756 ^ p37_array_index_1083821 ^ p37_array_index_1083792 ^ p37_literal_1076351[p37_array_index_1083759] ^ p37_literal_1076349[p37_array_index_1083760] ^ p37_literal_1076347[p37_array_index_1083777] ^ p37_literal_1076345[p37_array_index_1083762] ^ p37_array_index_1083779;
  assign p38_array_index_1083988_comb = p37_literal_1076353[p37_res7__195];
  assign p38_array_index_1083989_comb = p37_literal_1076355[p37_res7__194];
  assign p38_res7__200_comb = p37_literal_1076345[p38_res7__199_comb] ^ p37_literal_1076347[p38_res7__198_comb] ^ p37_literal_1076349[p38_res7__197_comb] ^ p37_literal_1076351[p37_res7__196] ^ p38_array_index_1083988_comb ^ p38_array_index_1083989_comb ^ p37_res7__193 ^ p37_literal_1076358[p37_res7__192] ^ p37_array_index_1083755 ^ p37_array_index_1083835 ^ p37_array_index_1083806 ^ p37_array_index_1083774 ^ p37_literal_1076349[p37_array_index_1083759] ^ p37_literal_1076347[p37_array_index_1083760] ^ p37_literal_1076345[p37_array_index_1083777] ^ p37_array_index_1083762;
  assign p38_array_index_1083999_comb = p37_literal_1076353[p37_res7__196];
  assign p38_array_index_1084000_comb = p37_literal_1076355[p37_res7__195];
  assign p38_res7__201_comb = p37_literal_1076345[p38_res7__200_comb] ^ p37_literal_1076347[p38_res7__199_comb] ^ p37_literal_1076349[p38_res7__198_comb] ^ p37_literal_1076351[p38_res7__197_comb] ^ p38_array_index_1083999_comb ^ p38_array_index_1084000_comb ^ p37_res7__194 ^ p37_literal_1076358[p37_res7__193] ^ p37_res7__192 ^ p38_array_index_1083952_comb ^ p37_array_index_1083820 ^ p37_array_index_1083791 ^ p37_literal_1076349[p37_array_index_1083758] ^ p37_literal_1076347[p37_array_index_1083759] ^ p37_literal_1076345[p37_array_index_1083760] ^ p37_array_index_1083777;
  assign p38_array_index_1084006_comb = p37_literal_1076345[p38_res7__201_comb];
  assign p38_array_index_1084007_comb = p37_literal_1076347[p38_res7__200_comb];
  assign p38_array_index_1084008_comb = p37_literal_1076349[p38_res7__199_comb];
  assign p38_array_index_1084009_comb = p37_literal_1076351[p38_res7__198_comb];
  assign p38_array_index_1084010_comb = p37_literal_1076353[p38_res7__197_comb];
  assign p38_array_index_1084011_comb = p37_literal_1076355[p37_res7__196];
  assign p38_array_index_1084012_comb = p37_literal_1076358[p37_res7__194];
  assign p38_array_index_1084013_comb = p37_literal_1076347[p37_array_index_1083758];
  assign p38_array_index_1084014_comb = p37_literal_1076345[p37_array_index_1083759];

  // Registers for pipe stage 38:
  reg [127:0] p38_xor_1083245;
  reg [127:0] p38_xor_1083717;
  reg [7:0] p38_array_index_1083755;
  reg [7:0] p38_array_index_1083756;
  reg [7:0] p38_array_index_1083757;
  reg [7:0] p38_array_index_1083758;
  reg [7:0] p38_array_index_1083759;
  reg [7:0] p38_array_index_1083760;
  reg [7:0] p38_array_index_1083771;
  reg [7:0] p38_array_index_1083772;
  reg [7:0] p38_array_index_1083773;
  reg [7:0] p38_res7__192;
  reg [7:0] p38_array_index_1083788;
  reg [7:0] p38_array_index_1083789;
  reg [7:0] p38_array_index_1083790;
  reg [7:0] p38_res7__193;
  reg [7:0] p38_array_index_1083803;
  reg [7:0] p38_array_index_1083804;
  reg [7:0] p38_array_index_1083805;
  reg [7:0] p38_res7__194;
  reg [7:0] p38_array_index_1083817;
  reg [7:0] p38_array_index_1083818;
  reg [7:0] p38_array_index_1083819;
  reg [7:0] p38_res7__195;
  reg [7:0] p38_array_index_1083832;
  reg [7:0] p38_array_index_1083833;
  reg [7:0] p38_array_index_1083834;
  reg [7:0] p38_res7__196;
  reg [7:0] p38_array_index_1083949;
  reg [7:0] p38_array_index_1083950;
  reg [7:0] p38_array_index_1083951;
  reg [7:0] p38_res7__197;
  reg [7:0] p38_array_index_1083963;
  reg [7:0] p38_array_index_1083964;
  reg [7:0] p38_array_index_1083965;
  reg [7:0] p38_res7__198;
  reg [7:0] p38_array_index_1083975;
  reg [7:0] p38_array_index_1083976;
  reg [7:0] p38_array_index_1083977;
  reg [7:0] p38_res7__199;
  reg [7:0] p38_array_index_1083988;
  reg [7:0] p38_array_index_1083989;
  reg [7:0] p38_res7__200;
  reg [7:0] p38_array_index_1083999;
  reg [7:0] p38_array_index_1084000;
  reg [7:0] p38_res7__201;
  reg [7:0] p38_array_index_1084006;
  reg [7:0] p38_array_index_1084007;
  reg [7:0] p38_array_index_1084008;
  reg [7:0] p38_array_index_1084009;
  reg [7:0] p38_array_index_1084010;
  reg [7:0] p38_array_index_1084011;
  reg [7:0] p38_array_index_1084012;
  reg [7:0] p38_array_index_1084013;
  reg [7:0] p38_array_index_1084014;
  reg [127:0] p38_res__35;
  reg [7:0] p39_arr[256];
  reg [7:0] p39_literal_1076345[256];
  reg [7:0] p39_literal_1076347[256];
  reg [7:0] p39_literal_1076349[256];
  reg [7:0] p39_literal_1076351[256];
  reg [7:0] p39_literal_1076353[256];
  reg [7:0] p39_literal_1076355[256];
  reg [7:0] p39_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p38_xor_1083245 <= p37_xor_1083245;
    p38_xor_1083717 <= p37_xor_1083717;
    p38_array_index_1083755 <= p37_array_index_1083755;
    p38_array_index_1083756 <= p37_array_index_1083756;
    p38_array_index_1083757 <= p37_array_index_1083757;
    p38_array_index_1083758 <= p37_array_index_1083758;
    p38_array_index_1083759 <= p37_array_index_1083759;
    p38_array_index_1083760 <= p37_array_index_1083760;
    p38_array_index_1083771 <= p37_array_index_1083771;
    p38_array_index_1083772 <= p37_array_index_1083772;
    p38_array_index_1083773 <= p37_array_index_1083773;
    p38_res7__192 <= p37_res7__192;
    p38_array_index_1083788 <= p37_array_index_1083788;
    p38_array_index_1083789 <= p37_array_index_1083789;
    p38_array_index_1083790 <= p37_array_index_1083790;
    p38_res7__193 <= p37_res7__193;
    p38_array_index_1083803 <= p37_array_index_1083803;
    p38_array_index_1083804 <= p37_array_index_1083804;
    p38_array_index_1083805 <= p37_array_index_1083805;
    p38_res7__194 <= p37_res7__194;
    p38_array_index_1083817 <= p37_array_index_1083817;
    p38_array_index_1083818 <= p37_array_index_1083818;
    p38_array_index_1083819 <= p37_array_index_1083819;
    p38_res7__195 <= p37_res7__195;
    p38_array_index_1083832 <= p37_array_index_1083832;
    p38_array_index_1083833 <= p37_array_index_1083833;
    p38_array_index_1083834 <= p37_array_index_1083834;
    p38_res7__196 <= p37_res7__196;
    p38_array_index_1083949 <= p38_array_index_1083949_comb;
    p38_array_index_1083950 <= p38_array_index_1083950_comb;
    p38_array_index_1083951 <= p38_array_index_1083951_comb;
    p38_res7__197 <= p38_res7__197_comb;
    p38_array_index_1083963 <= p38_array_index_1083963_comb;
    p38_array_index_1083964 <= p38_array_index_1083964_comb;
    p38_array_index_1083965 <= p38_array_index_1083965_comb;
    p38_res7__198 <= p38_res7__198_comb;
    p38_array_index_1083975 <= p38_array_index_1083975_comb;
    p38_array_index_1083976 <= p38_array_index_1083976_comb;
    p38_array_index_1083977 <= p38_array_index_1083977_comb;
    p38_res7__199 <= p38_res7__199_comb;
    p38_array_index_1083988 <= p38_array_index_1083988_comb;
    p38_array_index_1083989 <= p38_array_index_1083989_comb;
    p38_res7__200 <= p38_res7__200_comb;
    p38_array_index_1083999 <= p38_array_index_1083999_comb;
    p38_array_index_1084000 <= p38_array_index_1084000_comb;
    p38_res7__201 <= p38_res7__201_comb;
    p38_array_index_1084006 <= p38_array_index_1084006_comb;
    p38_array_index_1084007 <= p38_array_index_1084007_comb;
    p38_array_index_1084008 <= p38_array_index_1084008_comb;
    p38_array_index_1084009 <= p38_array_index_1084009_comb;
    p38_array_index_1084010 <= p38_array_index_1084010_comb;
    p38_array_index_1084011 <= p38_array_index_1084011_comb;
    p38_array_index_1084012 <= p38_array_index_1084012_comb;
    p38_array_index_1084013 <= p38_array_index_1084013_comb;
    p38_array_index_1084014 <= p38_array_index_1084014_comb;
    p38_res__35 <= p37_res__35;
    p39_arr <= p38_arr;
    p39_literal_1076345 <= p38_literal_1076345;
    p39_literal_1076347 <= p38_literal_1076347;
    p39_literal_1076349 <= p38_literal_1076349;
    p39_literal_1076351 <= p38_literal_1076351;
    p39_literal_1076353 <= p38_literal_1076353;
    p39_literal_1076355 <= p38_literal_1076355;
    p39_literal_1076358 <= p38_literal_1076358;
  end

  // ===== Pipe stage 39:
  wire [7:0] p39_res7__202_comb;
  wire [7:0] p39_array_index_1084149_comb;
  wire [7:0] p39_res7__203_comb;
  wire [7:0] p39_res7__204_comb;
  wire [7:0] p39_res7__205_comb;
  wire [7:0] p39_res7__206_comb;
  wire [7:0] p39_res7__207_comb;
  wire [127:0] p39_res__12_comb;
  wire [127:0] p39_xor_1084189_comb;
  assign p39_res7__202_comb = p38_array_index_1084006 ^ p38_array_index_1084007 ^ p38_array_index_1084008 ^ p38_array_index_1084009 ^ p38_array_index_1084010 ^ p38_array_index_1084011 ^ p38_res7__195 ^ p38_array_index_1084012 ^ p38_res7__193 ^ p38_array_index_1083965 ^ p38_array_index_1083834 ^ p38_array_index_1083805 ^ p38_array_index_1083773 ^ p38_array_index_1084013 ^ p38_array_index_1084014 ^ p38_array_index_1083760;
  assign p39_array_index_1084149_comb = p38_literal_1076355[p38_res7__197];
  assign p39_res7__203_comb = p38_literal_1076345[p39_res7__202_comb] ^ p38_literal_1076347[p38_res7__201] ^ p38_literal_1076349[p38_res7__200] ^ p38_literal_1076351[p38_res7__199] ^ p38_literal_1076353[p38_res7__198] ^ p39_array_index_1084149_comb ^ p38_res7__196 ^ p38_literal_1076358[p38_res7__195] ^ p38_res7__194 ^ p38_array_index_1083977 ^ p38_array_index_1083951 ^ p38_array_index_1083819 ^ p38_array_index_1083790 ^ p38_literal_1076347[p38_array_index_1083757] ^ p38_literal_1076345[p38_array_index_1083758] ^ p38_array_index_1083759;
  assign p39_res7__204_comb = p38_literal_1076345[p39_res7__203_comb] ^ p38_literal_1076347[p39_res7__202_comb] ^ p38_literal_1076349[p38_res7__201] ^ p38_literal_1076351[p38_res7__200] ^ p38_literal_1076353[p38_res7__199] ^ p38_literal_1076355[p38_res7__198] ^ p38_res7__197 ^ p38_literal_1076358[p38_res7__196] ^ p38_res7__195 ^ p38_array_index_1083989 ^ p38_array_index_1083964 ^ p38_array_index_1083833 ^ p38_array_index_1083804 ^ p38_array_index_1083772 ^ p38_literal_1076345[p38_array_index_1083757] ^ p38_array_index_1083758;
  assign p39_res7__205_comb = p38_literal_1076345[p39_res7__204_comb] ^ p38_literal_1076347[p39_res7__203_comb] ^ p38_literal_1076349[p39_res7__202_comb] ^ p38_literal_1076351[p38_res7__201] ^ p38_literal_1076353[p38_res7__200] ^ p38_literal_1076355[p38_res7__199] ^ p38_res7__198 ^ p38_literal_1076358[p38_res7__197] ^ p38_res7__196 ^ p38_array_index_1084000 ^ p38_array_index_1083976 ^ p38_array_index_1083950 ^ p38_array_index_1083818 ^ p38_array_index_1083789 ^ p38_literal_1076345[p38_array_index_1083756] ^ p38_array_index_1083757;
  assign p39_res7__206_comb = p38_literal_1076345[p39_res7__205_comb] ^ p38_literal_1076347[p39_res7__204_comb] ^ p38_literal_1076349[p39_res7__203_comb] ^ p38_literal_1076351[p39_res7__202_comb] ^ p38_literal_1076353[p38_res7__201] ^ p38_literal_1076355[p38_res7__200] ^ p38_res7__199 ^ p38_literal_1076358[p38_res7__198] ^ p38_res7__197 ^ p38_array_index_1084011 ^ p38_array_index_1083988 ^ p38_array_index_1083963 ^ p38_array_index_1083832 ^ p38_array_index_1083803 ^ p38_array_index_1083771 ^ p38_array_index_1083756;
  assign p39_res7__207_comb = p38_literal_1076345[p39_res7__206_comb] ^ p38_literal_1076347[p39_res7__205_comb] ^ p38_literal_1076349[p39_res7__204_comb] ^ p38_literal_1076351[p39_res7__203_comb] ^ p38_literal_1076353[p39_res7__202_comb] ^ p38_literal_1076355[p38_res7__201] ^ p38_res7__200 ^ p38_literal_1076358[p38_res7__199] ^ p38_res7__198 ^ p39_array_index_1084149_comb ^ p38_array_index_1083999 ^ p38_array_index_1083975 ^ p38_array_index_1083949 ^ p38_array_index_1083817 ^ p38_array_index_1083788 ^ p38_array_index_1083755;
  assign p39_res__12_comb = {p39_res7__207_comb, p39_res7__206_comb, p39_res7__205_comb, p39_res7__204_comb, p39_res7__203_comb, p39_res7__202_comb, p38_res7__201, p38_res7__200, p38_res7__199, p38_res7__198, p38_res7__197, p38_res7__196, p38_res7__195, p38_res7__194, p38_res7__193, p38_res7__192};
  assign p39_xor_1084189_comb = p39_res__12_comb ^ p38_xor_1083245;

  // Registers for pipe stage 39:
  reg [127:0] p39_xor_1083717;
  reg [127:0] p39_xor_1084189;
  reg [127:0] p39_res__35;
  reg [7:0] p40_arr[256];
  reg [7:0] p40_literal_1076345[256];
  reg [7:0] p40_literal_1076347[256];
  reg [7:0] p40_literal_1076349[256];
  reg [7:0] p40_literal_1076351[256];
  reg [7:0] p40_literal_1076353[256];
  reg [7:0] p40_literal_1076355[256];
  reg [7:0] p40_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p39_xor_1083717 <= p38_xor_1083717;
    p39_xor_1084189 <= p39_xor_1084189_comb;
    p39_res__35 <= p38_res__35;
    p40_arr <= p39_arr;
    p40_literal_1076345 <= p39_literal_1076345;
    p40_literal_1076347 <= p39_literal_1076347;
    p40_literal_1076349 <= p39_literal_1076349;
    p40_literal_1076351 <= p39_literal_1076351;
    p40_literal_1076353 <= p39_literal_1076353;
    p40_literal_1076355 <= p39_literal_1076355;
    p40_literal_1076358 <= p39_literal_1076358;
  end

  // ===== Pipe stage 40:
  wire [127:0] p40_addedKey__54_comb;
  wire [7:0] p40_array_index_1084227_comb;
  wire [7:0] p40_array_index_1084228_comb;
  wire [7:0] p40_array_index_1084229_comb;
  wire [7:0] p40_array_index_1084230_comb;
  wire [7:0] p40_array_index_1084231_comb;
  wire [7:0] p40_array_index_1084232_comb;
  wire [7:0] p40_array_index_1084234_comb;
  wire [7:0] p40_array_index_1084236_comb;
  wire [7:0] p40_array_index_1084237_comb;
  wire [7:0] p40_array_index_1084238_comb;
  wire [7:0] p40_array_index_1084239_comb;
  wire [7:0] p40_array_index_1084240_comb;
  wire [7:0] p40_array_index_1084241_comb;
  wire [7:0] p40_array_index_1084243_comb;
  wire [7:0] p40_array_index_1084244_comb;
  wire [7:0] p40_array_index_1084245_comb;
  wire [7:0] p40_array_index_1084246_comb;
  wire [7:0] p40_array_index_1084247_comb;
  wire [7:0] p40_array_index_1084248_comb;
  wire [7:0] p40_array_index_1084249_comb;
  wire [7:0] p40_array_index_1084251_comb;
  wire [7:0] p40_res7__208_comb;
  wire [7:0] p40_array_index_1084260_comb;
  wire [7:0] p40_array_index_1084261_comb;
  wire [7:0] p40_array_index_1084262_comb;
  wire [7:0] p40_array_index_1084263_comb;
  wire [7:0] p40_array_index_1084264_comb;
  wire [7:0] p40_array_index_1084265_comb;
  wire [7:0] p40_res7__209_comb;
  wire [7:0] p40_array_index_1084275_comb;
  wire [7:0] p40_array_index_1084276_comb;
  wire [7:0] p40_array_index_1084277_comb;
  wire [7:0] p40_array_index_1084278_comb;
  wire [7:0] p40_array_index_1084279_comb;
  wire [7:0] p40_res7__210_comb;
  wire [7:0] p40_array_index_1084289_comb;
  wire [7:0] p40_array_index_1084290_comb;
  wire [7:0] p40_array_index_1084291_comb;
  wire [7:0] p40_array_index_1084292_comb;
  wire [7:0] p40_array_index_1084293_comb;
  wire [7:0] p40_res7__211_comb;
  wire [7:0] p40_array_index_1084304_comb;
  wire [7:0] p40_array_index_1084305_comb;
  wire [7:0] p40_array_index_1084306_comb;
  wire [7:0] p40_array_index_1084307_comb;
  wire [7:0] p40_res7__212_comb;
  assign p40_addedKey__54_comb = p39_xor_1084189 ^ 128'h5113_c1f9_4d76_899f_a029_a9e0_ac34_d40e;
  assign p40_array_index_1084227_comb = p39_arr[p40_addedKey__54_comb[127:120]];
  assign p40_array_index_1084228_comb = p39_arr[p40_addedKey__54_comb[119:112]];
  assign p40_array_index_1084229_comb = p39_arr[p40_addedKey__54_comb[111:104]];
  assign p40_array_index_1084230_comb = p39_arr[p40_addedKey__54_comb[103:96]];
  assign p40_array_index_1084231_comb = p39_arr[p40_addedKey__54_comb[95:88]];
  assign p40_array_index_1084232_comb = p39_arr[p40_addedKey__54_comb[87:80]];
  assign p40_array_index_1084234_comb = p39_arr[p40_addedKey__54_comb[71:64]];
  assign p40_array_index_1084236_comb = p39_arr[p40_addedKey__54_comb[55:48]];
  assign p40_array_index_1084237_comb = p39_arr[p40_addedKey__54_comb[47:40]];
  assign p40_array_index_1084238_comb = p39_arr[p40_addedKey__54_comb[39:32]];
  assign p40_array_index_1084239_comb = p39_arr[p40_addedKey__54_comb[31:24]];
  assign p40_array_index_1084240_comb = p39_arr[p40_addedKey__54_comb[23:16]];
  assign p40_array_index_1084241_comb = p39_arr[p40_addedKey__54_comb[15:8]];
  assign p40_array_index_1084243_comb = p39_literal_1076345[p40_array_index_1084227_comb];
  assign p40_array_index_1084244_comb = p39_literal_1076347[p40_array_index_1084228_comb];
  assign p40_array_index_1084245_comb = p39_literal_1076349[p40_array_index_1084229_comb];
  assign p40_array_index_1084246_comb = p39_literal_1076351[p40_array_index_1084230_comb];
  assign p40_array_index_1084247_comb = p39_literal_1076353[p40_array_index_1084231_comb];
  assign p40_array_index_1084248_comb = p39_literal_1076355[p40_array_index_1084232_comb];
  assign p40_array_index_1084249_comb = p39_arr[p40_addedKey__54_comb[79:72]];
  assign p40_array_index_1084251_comb = p39_arr[p40_addedKey__54_comb[63:56]];
  assign p40_res7__208_comb = p40_array_index_1084243_comb ^ p40_array_index_1084244_comb ^ p40_array_index_1084245_comb ^ p40_array_index_1084246_comb ^ p40_array_index_1084247_comb ^ p40_array_index_1084248_comb ^ p40_array_index_1084249_comb ^ p39_literal_1076358[p40_array_index_1084234_comb] ^ p40_array_index_1084251_comb ^ p39_literal_1076355[p40_array_index_1084236_comb] ^ p39_literal_1076353[p40_array_index_1084237_comb] ^ p39_literal_1076351[p40_array_index_1084238_comb] ^ p39_literal_1076349[p40_array_index_1084239_comb] ^ p39_literal_1076347[p40_array_index_1084240_comb] ^ p39_literal_1076345[p40_array_index_1084241_comb] ^ p39_arr[p40_addedKey__54_comb[7:0]];
  assign p40_array_index_1084260_comb = p39_literal_1076345[p40_res7__208_comb];
  assign p40_array_index_1084261_comb = p39_literal_1076347[p40_array_index_1084227_comb];
  assign p40_array_index_1084262_comb = p39_literal_1076349[p40_array_index_1084228_comb];
  assign p40_array_index_1084263_comb = p39_literal_1076351[p40_array_index_1084229_comb];
  assign p40_array_index_1084264_comb = p39_literal_1076353[p40_array_index_1084230_comb];
  assign p40_array_index_1084265_comb = p39_literal_1076355[p40_array_index_1084231_comb];
  assign p40_res7__209_comb = p40_array_index_1084260_comb ^ p40_array_index_1084261_comb ^ p40_array_index_1084262_comb ^ p40_array_index_1084263_comb ^ p40_array_index_1084264_comb ^ p40_array_index_1084265_comb ^ p40_array_index_1084232_comb ^ p39_literal_1076358[p40_array_index_1084249_comb] ^ p40_array_index_1084234_comb ^ p39_literal_1076355[p40_array_index_1084251_comb] ^ p39_literal_1076353[p40_array_index_1084236_comb] ^ p39_literal_1076351[p40_array_index_1084237_comb] ^ p39_literal_1076349[p40_array_index_1084238_comb] ^ p39_literal_1076347[p40_array_index_1084239_comb] ^ p39_literal_1076345[p40_array_index_1084240_comb] ^ p40_array_index_1084241_comb;
  assign p40_array_index_1084275_comb = p39_literal_1076347[p40_res7__208_comb];
  assign p40_array_index_1084276_comb = p39_literal_1076349[p40_array_index_1084227_comb];
  assign p40_array_index_1084277_comb = p39_literal_1076351[p40_array_index_1084228_comb];
  assign p40_array_index_1084278_comb = p39_literal_1076353[p40_array_index_1084229_comb];
  assign p40_array_index_1084279_comb = p39_literal_1076355[p40_array_index_1084230_comb];
  assign p40_res7__210_comb = p39_literal_1076345[p40_res7__209_comb] ^ p40_array_index_1084275_comb ^ p40_array_index_1084276_comb ^ p40_array_index_1084277_comb ^ p40_array_index_1084278_comb ^ p40_array_index_1084279_comb ^ p40_array_index_1084231_comb ^ p39_literal_1076358[p40_array_index_1084232_comb] ^ p40_array_index_1084249_comb ^ p39_literal_1076355[p40_array_index_1084234_comb] ^ p39_literal_1076353[p40_array_index_1084251_comb] ^ p39_literal_1076351[p40_array_index_1084236_comb] ^ p39_literal_1076349[p40_array_index_1084237_comb] ^ p39_literal_1076347[p40_array_index_1084238_comb] ^ p39_literal_1076345[p40_array_index_1084239_comb] ^ p40_array_index_1084240_comb;
  assign p40_array_index_1084289_comb = p39_literal_1076347[p40_res7__209_comb];
  assign p40_array_index_1084290_comb = p39_literal_1076349[p40_res7__208_comb];
  assign p40_array_index_1084291_comb = p39_literal_1076351[p40_array_index_1084227_comb];
  assign p40_array_index_1084292_comb = p39_literal_1076353[p40_array_index_1084228_comb];
  assign p40_array_index_1084293_comb = p39_literal_1076355[p40_array_index_1084229_comb];
  assign p40_res7__211_comb = p39_literal_1076345[p40_res7__210_comb] ^ p40_array_index_1084289_comb ^ p40_array_index_1084290_comb ^ p40_array_index_1084291_comb ^ p40_array_index_1084292_comb ^ p40_array_index_1084293_comb ^ p40_array_index_1084230_comb ^ p39_literal_1076358[p40_array_index_1084231_comb] ^ p40_array_index_1084232_comb ^ p39_literal_1076355[p40_array_index_1084249_comb] ^ p39_literal_1076353[p40_array_index_1084234_comb] ^ p39_literal_1076351[p40_array_index_1084251_comb] ^ p39_literal_1076349[p40_array_index_1084236_comb] ^ p39_literal_1076347[p40_array_index_1084237_comb] ^ p39_literal_1076345[p40_array_index_1084238_comb] ^ p40_array_index_1084239_comb;
  assign p40_array_index_1084304_comb = p39_literal_1076349[p40_res7__209_comb];
  assign p40_array_index_1084305_comb = p39_literal_1076351[p40_res7__208_comb];
  assign p40_array_index_1084306_comb = p39_literal_1076353[p40_array_index_1084227_comb];
  assign p40_array_index_1084307_comb = p39_literal_1076355[p40_array_index_1084228_comb];
  assign p40_res7__212_comb = p39_literal_1076345[p40_res7__211_comb] ^ p39_literal_1076347[p40_res7__210_comb] ^ p40_array_index_1084304_comb ^ p40_array_index_1084305_comb ^ p40_array_index_1084306_comb ^ p40_array_index_1084307_comb ^ p40_array_index_1084229_comb ^ p39_literal_1076358[p40_array_index_1084230_comb] ^ p40_array_index_1084231_comb ^ p40_array_index_1084248_comb ^ p39_literal_1076353[p40_array_index_1084249_comb] ^ p39_literal_1076351[p40_array_index_1084234_comb] ^ p39_literal_1076349[p40_array_index_1084251_comb] ^ p39_literal_1076347[p40_array_index_1084236_comb] ^ p39_literal_1076345[p40_array_index_1084237_comb] ^ p40_array_index_1084238_comb;

  // Registers for pipe stage 40:
  reg [127:0] p40_xor_1083717;
  reg [127:0] p40_xor_1084189;
  reg [7:0] p40_array_index_1084227;
  reg [7:0] p40_array_index_1084228;
  reg [7:0] p40_array_index_1084229;
  reg [7:0] p40_array_index_1084230;
  reg [7:0] p40_array_index_1084231;
  reg [7:0] p40_array_index_1084232;
  reg [7:0] p40_array_index_1084234;
  reg [7:0] p40_array_index_1084236;
  reg [7:0] p40_array_index_1084237;
  reg [7:0] p40_array_index_1084243;
  reg [7:0] p40_array_index_1084244;
  reg [7:0] p40_array_index_1084245;
  reg [7:0] p40_array_index_1084246;
  reg [7:0] p40_array_index_1084247;
  reg [7:0] p40_array_index_1084249;
  reg [7:0] p40_array_index_1084251;
  reg [7:0] p40_res7__208;
  reg [7:0] p40_array_index_1084260;
  reg [7:0] p40_array_index_1084261;
  reg [7:0] p40_array_index_1084262;
  reg [7:0] p40_array_index_1084263;
  reg [7:0] p40_array_index_1084264;
  reg [7:0] p40_array_index_1084265;
  reg [7:0] p40_res7__209;
  reg [7:0] p40_array_index_1084275;
  reg [7:0] p40_array_index_1084276;
  reg [7:0] p40_array_index_1084277;
  reg [7:0] p40_array_index_1084278;
  reg [7:0] p40_array_index_1084279;
  reg [7:0] p40_res7__210;
  reg [7:0] p40_array_index_1084289;
  reg [7:0] p40_array_index_1084290;
  reg [7:0] p40_array_index_1084291;
  reg [7:0] p40_array_index_1084292;
  reg [7:0] p40_array_index_1084293;
  reg [7:0] p40_res7__211;
  reg [7:0] p40_array_index_1084304;
  reg [7:0] p40_array_index_1084305;
  reg [7:0] p40_array_index_1084306;
  reg [7:0] p40_array_index_1084307;
  reg [7:0] p40_res7__212;
  reg [127:0] p40_res__35;
  reg [7:0] p41_arr[256];
  reg [7:0] p41_literal_1076345[256];
  reg [7:0] p41_literal_1076347[256];
  reg [7:0] p41_literal_1076349[256];
  reg [7:0] p41_literal_1076351[256];
  reg [7:0] p41_literal_1076353[256];
  reg [7:0] p41_literal_1076355[256];
  reg [7:0] p41_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p40_xor_1083717 <= p39_xor_1083717;
    p40_xor_1084189 <= p39_xor_1084189;
    p40_array_index_1084227 <= p40_array_index_1084227_comb;
    p40_array_index_1084228 <= p40_array_index_1084228_comb;
    p40_array_index_1084229 <= p40_array_index_1084229_comb;
    p40_array_index_1084230 <= p40_array_index_1084230_comb;
    p40_array_index_1084231 <= p40_array_index_1084231_comb;
    p40_array_index_1084232 <= p40_array_index_1084232_comb;
    p40_array_index_1084234 <= p40_array_index_1084234_comb;
    p40_array_index_1084236 <= p40_array_index_1084236_comb;
    p40_array_index_1084237 <= p40_array_index_1084237_comb;
    p40_array_index_1084243 <= p40_array_index_1084243_comb;
    p40_array_index_1084244 <= p40_array_index_1084244_comb;
    p40_array_index_1084245 <= p40_array_index_1084245_comb;
    p40_array_index_1084246 <= p40_array_index_1084246_comb;
    p40_array_index_1084247 <= p40_array_index_1084247_comb;
    p40_array_index_1084249 <= p40_array_index_1084249_comb;
    p40_array_index_1084251 <= p40_array_index_1084251_comb;
    p40_res7__208 <= p40_res7__208_comb;
    p40_array_index_1084260 <= p40_array_index_1084260_comb;
    p40_array_index_1084261 <= p40_array_index_1084261_comb;
    p40_array_index_1084262 <= p40_array_index_1084262_comb;
    p40_array_index_1084263 <= p40_array_index_1084263_comb;
    p40_array_index_1084264 <= p40_array_index_1084264_comb;
    p40_array_index_1084265 <= p40_array_index_1084265_comb;
    p40_res7__209 <= p40_res7__209_comb;
    p40_array_index_1084275 <= p40_array_index_1084275_comb;
    p40_array_index_1084276 <= p40_array_index_1084276_comb;
    p40_array_index_1084277 <= p40_array_index_1084277_comb;
    p40_array_index_1084278 <= p40_array_index_1084278_comb;
    p40_array_index_1084279 <= p40_array_index_1084279_comb;
    p40_res7__210 <= p40_res7__210_comb;
    p40_array_index_1084289 <= p40_array_index_1084289_comb;
    p40_array_index_1084290 <= p40_array_index_1084290_comb;
    p40_array_index_1084291 <= p40_array_index_1084291_comb;
    p40_array_index_1084292 <= p40_array_index_1084292_comb;
    p40_array_index_1084293 <= p40_array_index_1084293_comb;
    p40_res7__211 <= p40_res7__211_comb;
    p40_array_index_1084304 <= p40_array_index_1084304_comb;
    p40_array_index_1084305 <= p40_array_index_1084305_comb;
    p40_array_index_1084306 <= p40_array_index_1084306_comb;
    p40_array_index_1084307 <= p40_array_index_1084307_comb;
    p40_res7__212 <= p40_res7__212_comb;
    p40_res__35 <= p39_res__35;
    p41_arr <= p40_arr;
    p41_literal_1076345 <= p40_literal_1076345;
    p41_literal_1076347 <= p40_literal_1076347;
    p41_literal_1076349 <= p40_literal_1076349;
    p41_literal_1076351 <= p40_literal_1076351;
    p41_literal_1076353 <= p40_literal_1076353;
    p41_literal_1076355 <= p40_literal_1076355;
    p41_literal_1076358 <= p40_literal_1076358;
  end

  // ===== Pipe stage 41:
  wire [7:0] p41_array_index_1084421_comb;
  wire [7:0] p41_array_index_1084422_comb;
  wire [7:0] p41_array_index_1084423_comb;
  wire [7:0] p41_array_index_1084424_comb;
  wire [7:0] p41_res7__213_comb;
  wire [7:0] p41_array_index_1084435_comb;
  wire [7:0] p41_array_index_1084436_comb;
  wire [7:0] p41_array_index_1084437_comb;
  wire [7:0] p41_res7__214_comb;
  wire [7:0] p41_array_index_1084447_comb;
  wire [7:0] p41_array_index_1084448_comb;
  wire [7:0] p41_array_index_1084449_comb;
  wire [7:0] p41_res7__215_comb;
  wire [7:0] p41_array_index_1084460_comb;
  wire [7:0] p41_array_index_1084461_comb;
  wire [7:0] p41_res7__216_comb;
  wire [7:0] p41_array_index_1084471_comb;
  wire [7:0] p41_array_index_1084472_comb;
  wire [7:0] p41_res7__217_comb;
  wire [7:0] p41_array_index_1084478_comb;
  wire [7:0] p41_array_index_1084479_comb;
  wire [7:0] p41_array_index_1084480_comb;
  wire [7:0] p41_array_index_1084481_comb;
  wire [7:0] p41_array_index_1084482_comb;
  wire [7:0] p41_array_index_1084483_comb;
  wire [7:0] p41_array_index_1084484_comb;
  wire [7:0] p41_array_index_1084485_comb;
  wire [7:0] p41_array_index_1084486_comb;
  assign p41_array_index_1084421_comb = p40_literal_1076349[p40_res7__210];
  assign p41_array_index_1084422_comb = p40_literal_1076351[p40_res7__209];
  assign p41_array_index_1084423_comb = p40_literal_1076353[p40_res7__208];
  assign p41_array_index_1084424_comb = p40_literal_1076355[p40_array_index_1084227];
  assign p41_res7__213_comb = p40_literal_1076345[p40_res7__212] ^ p40_literal_1076347[p40_res7__211] ^ p41_array_index_1084421_comb ^ p41_array_index_1084422_comb ^ p41_array_index_1084423_comb ^ p41_array_index_1084424_comb ^ p40_array_index_1084228 ^ p40_literal_1076358[p40_array_index_1084229] ^ p40_array_index_1084230 ^ p40_array_index_1084265 ^ p40_literal_1076353[p40_array_index_1084232] ^ p40_literal_1076351[p40_array_index_1084249] ^ p40_literal_1076349[p40_array_index_1084234] ^ p40_literal_1076347[p40_array_index_1084251] ^ p40_literal_1076345[p40_array_index_1084236] ^ p40_array_index_1084237;
  assign p41_array_index_1084435_comb = p40_literal_1076351[p40_res7__210];
  assign p41_array_index_1084436_comb = p40_literal_1076353[p40_res7__209];
  assign p41_array_index_1084437_comb = p40_literal_1076355[p40_res7__208];
  assign p41_res7__214_comb = p40_literal_1076345[p41_res7__213_comb] ^ p40_literal_1076347[p40_res7__212] ^ p40_literal_1076349[p40_res7__211] ^ p41_array_index_1084435_comb ^ p41_array_index_1084436_comb ^ p41_array_index_1084437_comb ^ p40_array_index_1084227 ^ p40_literal_1076358[p40_array_index_1084228] ^ p40_array_index_1084229 ^ p40_array_index_1084279 ^ p40_array_index_1084247 ^ p40_literal_1076351[p40_array_index_1084232] ^ p40_literal_1076349[p40_array_index_1084249] ^ p40_literal_1076347[p40_array_index_1084234] ^ p40_literal_1076345[p40_array_index_1084251] ^ p40_array_index_1084236;
  assign p41_array_index_1084447_comb = p40_literal_1076351[p40_res7__211];
  assign p41_array_index_1084448_comb = p40_literal_1076353[p40_res7__210];
  assign p41_array_index_1084449_comb = p40_literal_1076355[p40_res7__209];
  assign p41_res7__215_comb = p40_literal_1076345[p41_res7__214_comb] ^ p40_literal_1076347[p41_res7__213_comb] ^ p40_literal_1076349[p40_res7__212] ^ p41_array_index_1084447_comb ^ p41_array_index_1084448_comb ^ p41_array_index_1084449_comb ^ p40_res7__208 ^ p40_literal_1076358[p40_array_index_1084227] ^ p40_array_index_1084228 ^ p40_array_index_1084293 ^ p40_array_index_1084264 ^ p40_literal_1076351[p40_array_index_1084231] ^ p40_literal_1076349[p40_array_index_1084232] ^ p40_literal_1076347[p40_array_index_1084249] ^ p40_literal_1076345[p40_array_index_1084234] ^ p40_array_index_1084251;
  assign p41_array_index_1084460_comb = p40_literal_1076353[p40_res7__211];
  assign p41_array_index_1084461_comb = p40_literal_1076355[p40_res7__210];
  assign p41_res7__216_comb = p40_literal_1076345[p41_res7__215_comb] ^ p40_literal_1076347[p41_res7__214_comb] ^ p40_literal_1076349[p41_res7__213_comb] ^ p40_literal_1076351[p40_res7__212] ^ p41_array_index_1084460_comb ^ p41_array_index_1084461_comb ^ p40_res7__209 ^ p40_literal_1076358[p40_res7__208] ^ p40_array_index_1084227 ^ p40_array_index_1084307 ^ p40_array_index_1084278 ^ p40_array_index_1084246 ^ p40_literal_1076349[p40_array_index_1084231] ^ p40_literal_1076347[p40_array_index_1084232] ^ p40_literal_1076345[p40_array_index_1084249] ^ p40_array_index_1084234;
  assign p41_array_index_1084471_comb = p40_literal_1076353[p40_res7__212];
  assign p41_array_index_1084472_comb = p40_literal_1076355[p40_res7__211];
  assign p41_res7__217_comb = p40_literal_1076345[p41_res7__216_comb] ^ p40_literal_1076347[p41_res7__215_comb] ^ p40_literal_1076349[p41_res7__214_comb] ^ p40_literal_1076351[p41_res7__213_comb] ^ p41_array_index_1084471_comb ^ p41_array_index_1084472_comb ^ p40_res7__210 ^ p40_literal_1076358[p40_res7__209] ^ p40_res7__208 ^ p41_array_index_1084424_comb ^ p40_array_index_1084292 ^ p40_array_index_1084263 ^ p40_literal_1076349[p40_array_index_1084230] ^ p40_literal_1076347[p40_array_index_1084231] ^ p40_literal_1076345[p40_array_index_1084232] ^ p40_array_index_1084249;
  assign p41_array_index_1084478_comb = p40_literal_1076345[p41_res7__217_comb];
  assign p41_array_index_1084479_comb = p40_literal_1076347[p41_res7__216_comb];
  assign p41_array_index_1084480_comb = p40_literal_1076349[p41_res7__215_comb];
  assign p41_array_index_1084481_comb = p40_literal_1076351[p41_res7__214_comb];
  assign p41_array_index_1084482_comb = p40_literal_1076353[p41_res7__213_comb];
  assign p41_array_index_1084483_comb = p40_literal_1076355[p40_res7__212];
  assign p41_array_index_1084484_comb = p40_literal_1076358[p40_res7__210];
  assign p41_array_index_1084485_comb = p40_literal_1076347[p40_array_index_1084230];
  assign p41_array_index_1084486_comb = p40_literal_1076345[p40_array_index_1084231];

  // Registers for pipe stage 41:
  reg [127:0] p41_xor_1083717;
  reg [127:0] p41_xor_1084189;
  reg [7:0] p41_array_index_1084227;
  reg [7:0] p41_array_index_1084228;
  reg [7:0] p41_array_index_1084229;
  reg [7:0] p41_array_index_1084230;
  reg [7:0] p41_array_index_1084231;
  reg [7:0] p41_array_index_1084232;
  reg [7:0] p41_array_index_1084243;
  reg [7:0] p41_array_index_1084244;
  reg [7:0] p41_array_index_1084245;
  reg [7:0] p41_res7__208;
  reg [7:0] p41_array_index_1084260;
  reg [7:0] p41_array_index_1084261;
  reg [7:0] p41_array_index_1084262;
  reg [7:0] p41_res7__209;
  reg [7:0] p41_array_index_1084275;
  reg [7:0] p41_array_index_1084276;
  reg [7:0] p41_array_index_1084277;
  reg [7:0] p41_res7__210;
  reg [7:0] p41_array_index_1084289;
  reg [7:0] p41_array_index_1084290;
  reg [7:0] p41_array_index_1084291;
  reg [7:0] p41_res7__211;
  reg [7:0] p41_array_index_1084304;
  reg [7:0] p41_array_index_1084305;
  reg [7:0] p41_array_index_1084306;
  reg [7:0] p41_res7__212;
  reg [7:0] p41_array_index_1084421;
  reg [7:0] p41_array_index_1084422;
  reg [7:0] p41_array_index_1084423;
  reg [7:0] p41_res7__213;
  reg [7:0] p41_array_index_1084435;
  reg [7:0] p41_array_index_1084436;
  reg [7:0] p41_array_index_1084437;
  reg [7:0] p41_res7__214;
  reg [7:0] p41_array_index_1084447;
  reg [7:0] p41_array_index_1084448;
  reg [7:0] p41_array_index_1084449;
  reg [7:0] p41_res7__215;
  reg [7:0] p41_array_index_1084460;
  reg [7:0] p41_array_index_1084461;
  reg [7:0] p41_res7__216;
  reg [7:0] p41_array_index_1084471;
  reg [7:0] p41_array_index_1084472;
  reg [7:0] p41_res7__217;
  reg [7:0] p41_array_index_1084478;
  reg [7:0] p41_array_index_1084479;
  reg [7:0] p41_array_index_1084480;
  reg [7:0] p41_array_index_1084481;
  reg [7:0] p41_array_index_1084482;
  reg [7:0] p41_array_index_1084483;
  reg [7:0] p41_array_index_1084484;
  reg [7:0] p41_array_index_1084485;
  reg [7:0] p41_array_index_1084486;
  reg [127:0] p41_res__35;
  reg [7:0] p42_arr[256];
  reg [7:0] p42_literal_1076345[256];
  reg [7:0] p42_literal_1076347[256];
  reg [7:0] p42_literal_1076349[256];
  reg [7:0] p42_literal_1076351[256];
  reg [7:0] p42_literal_1076353[256];
  reg [7:0] p42_literal_1076355[256];
  reg [7:0] p42_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p41_xor_1083717 <= p40_xor_1083717;
    p41_xor_1084189 <= p40_xor_1084189;
    p41_array_index_1084227 <= p40_array_index_1084227;
    p41_array_index_1084228 <= p40_array_index_1084228;
    p41_array_index_1084229 <= p40_array_index_1084229;
    p41_array_index_1084230 <= p40_array_index_1084230;
    p41_array_index_1084231 <= p40_array_index_1084231;
    p41_array_index_1084232 <= p40_array_index_1084232;
    p41_array_index_1084243 <= p40_array_index_1084243;
    p41_array_index_1084244 <= p40_array_index_1084244;
    p41_array_index_1084245 <= p40_array_index_1084245;
    p41_res7__208 <= p40_res7__208;
    p41_array_index_1084260 <= p40_array_index_1084260;
    p41_array_index_1084261 <= p40_array_index_1084261;
    p41_array_index_1084262 <= p40_array_index_1084262;
    p41_res7__209 <= p40_res7__209;
    p41_array_index_1084275 <= p40_array_index_1084275;
    p41_array_index_1084276 <= p40_array_index_1084276;
    p41_array_index_1084277 <= p40_array_index_1084277;
    p41_res7__210 <= p40_res7__210;
    p41_array_index_1084289 <= p40_array_index_1084289;
    p41_array_index_1084290 <= p40_array_index_1084290;
    p41_array_index_1084291 <= p40_array_index_1084291;
    p41_res7__211 <= p40_res7__211;
    p41_array_index_1084304 <= p40_array_index_1084304;
    p41_array_index_1084305 <= p40_array_index_1084305;
    p41_array_index_1084306 <= p40_array_index_1084306;
    p41_res7__212 <= p40_res7__212;
    p41_array_index_1084421 <= p41_array_index_1084421_comb;
    p41_array_index_1084422 <= p41_array_index_1084422_comb;
    p41_array_index_1084423 <= p41_array_index_1084423_comb;
    p41_res7__213 <= p41_res7__213_comb;
    p41_array_index_1084435 <= p41_array_index_1084435_comb;
    p41_array_index_1084436 <= p41_array_index_1084436_comb;
    p41_array_index_1084437 <= p41_array_index_1084437_comb;
    p41_res7__214 <= p41_res7__214_comb;
    p41_array_index_1084447 <= p41_array_index_1084447_comb;
    p41_array_index_1084448 <= p41_array_index_1084448_comb;
    p41_array_index_1084449 <= p41_array_index_1084449_comb;
    p41_res7__215 <= p41_res7__215_comb;
    p41_array_index_1084460 <= p41_array_index_1084460_comb;
    p41_array_index_1084461 <= p41_array_index_1084461_comb;
    p41_res7__216 <= p41_res7__216_comb;
    p41_array_index_1084471 <= p41_array_index_1084471_comb;
    p41_array_index_1084472 <= p41_array_index_1084472_comb;
    p41_res7__217 <= p41_res7__217_comb;
    p41_array_index_1084478 <= p41_array_index_1084478_comb;
    p41_array_index_1084479 <= p41_array_index_1084479_comb;
    p41_array_index_1084480 <= p41_array_index_1084480_comb;
    p41_array_index_1084481 <= p41_array_index_1084481_comb;
    p41_array_index_1084482 <= p41_array_index_1084482_comb;
    p41_array_index_1084483 <= p41_array_index_1084483_comb;
    p41_array_index_1084484 <= p41_array_index_1084484_comb;
    p41_array_index_1084485 <= p41_array_index_1084485_comb;
    p41_array_index_1084486 <= p41_array_index_1084486_comb;
    p41_res__35 <= p40_res__35;
    p42_arr <= p41_arr;
    p42_literal_1076345 <= p41_literal_1076345;
    p42_literal_1076347 <= p41_literal_1076347;
    p42_literal_1076349 <= p41_literal_1076349;
    p42_literal_1076351 <= p41_literal_1076351;
    p42_literal_1076353 <= p41_literal_1076353;
    p42_literal_1076355 <= p41_literal_1076355;
    p42_literal_1076358 <= p41_literal_1076358;
  end

  // ===== Pipe stage 42:
  wire [7:0] p42_res7__218_comb;
  wire [7:0] p42_array_index_1084621_comb;
  wire [7:0] p42_res7__219_comb;
  wire [7:0] p42_res7__220_comb;
  wire [7:0] p42_res7__221_comb;
  wire [7:0] p42_res7__222_comb;
  wire [7:0] p42_res7__223_comb;
  wire [127:0] p42_res__13_comb;
  wire [127:0] p42_xor_1084661_comb;
  assign p42_res7__218_comb = p41_array_index_1084478 ^ p41_array_index_1084479 ^ p41_array_index_1084480 ^ p41_array_index_1084481 ^ p41_array_index_1084482 ^ p41_array_index_1084483 ^ p41_res7__211 ^ p41_array_index_1084484 ^ p41_res7__209 ^ p41_array_index_1084437 ^ p41_array_index_1084306 ^ p41_array_index_1084277 ^ p41_array_index_1084245 ^ p41_array_index_1084485 ^ p41_array_index_1084486 ^ p41_array_index_1084232;
  assign p42_array_index_1084621_comb = p41_literal_1076355[p41_res7__213];
  assign p42_res7__219_comb = p41_literal_1076345[p42_res7__218_comb] ^ p41_literal_1076347[p41_res7__217] ^ p41_literal_1076349[p41_res7__216] ^ p41_literal_1076351[p41_res7__215] ^ p41_literal_1076353[p41_res7__214] ^ p42_array_index_1084621_comb ^ p41_res7__212 ^ p41_literal_1076358[p41_res7__211] ^ p41_res7__210 ^ p41_array_index_1084449 ^ p41_array_index_1084423 ^ p41_array_index_1084291 ^ p41_array_index_1084262 ^ p41_literal_1076347[p41_array_index_1084229] ^ p41_literal_1076345[p41_array_index_1084230] ^ p41_array_index_1084231;
  assign p42_res7__220_comb = p41_literal_1076345[p42_res7__219_comb] ^ p41_literal_1076347[p42_res7__218_comb] ^ p41_literal_1076349[p41_res7__217] ^ p41_literal_1076351[p41_res7__216] ^ p41_literal_1076353[p41_res7__215] ^ p41_literal_1076355[p41_res7__214] ^ p41_res7__213 ^ p41_literal_1076358[p41_res7__212] ^ p41_res7__211 ^ p41_array_index_1084461 ^ p41_array_index_1084436 ^ p41_array_index_1084305 ^ p41_array_index_1084276 ^ p41_array_index_1084244 ^ p41_literal_1076345[p41_array_index_1084229] ^ p41_array_index_1084230;
  assign p42_res7__221_comb = p41_literal_1076345[p42_res7__220_comb] ^ p41_literal_1076347[p42_res7__219_comb] ^ p41_literal_1076349[p42_res7__218_comb] ^ p41_literal_1076351[p41_res7__217] ^ p41_literal_1076353[p41_res7__216] ^ p41_literal_1076355[p41_res7__215] ^ p41_res7__214 ^ p41_literal_1076358[p41_res7__213] ^ p41_res7__212 ^ p41_array_index_1084472 ^ p41_array_index_1084448 ^ p41_array_index_1084422 ^ p41_array_index_1084290 ^ p41_array_index_1084261 ^ p41_literal_1076345[p41_array_index_1084228] ^ p41_array_index_1084229;
  assign p42_res7__222_comb = p41_literal_1076345[p42_res7__221_comb] ^ p41_literal_1076347[p42_res7__220_comb] ^ p41_literal_1076349[p42_res7__219_comb] ^ p41_literal_1076351[p42_res7__218_comb] ^ p41_literal_1076353[p41_res7__217] ^ p41_literal_1076355[p41_res7__216] ^ p41_res7__215 ^ p41_literal_1076358[p41_res7__214] ^ p41_res7__213 ^ p41_array_index_1084483 ^ p41_array_index_1084460 ^ p41_array_index_1084435 ^ p41_array_index_1084304 ^ p41_array_index_1084275 ^ p41_array_index_1084243 ^ p41_array_index_1084228;
  assign p42_res7__223_comb = p41_literal_1076345[p42_res7__222_comb] ^ p41_literal_1076347[p42_res7__221_comb] ^ p41_literal_1076349[p42_res7__220_comb] ^ p41_literal_1076351[p42_res7__219_comb] ^ p41_literal_1076353[p42_res7__218_comb] ^ p41_literal_1076355[p41_res7__217] ^ p41_res7__216 ^ p41_literal_1076358[p41_res7__215] ^ p41_res7__214 ^ p42_array_index_1084621_comb ^ p41_array_index_1084471 ^ p41_array_index_1084447 ^ p41_array_index_1084421 ^ p41_array_index_1084289 ^ p41_array_index_1084260 ^ p41_array_index_1084227;
  assign p42_res__13_comb = {p42_res7__223_comb, p42_res7__222_comb, p42_res7__221_comb, p42_res7__220_comb, p42_res7__219_comb, p42_res7__218_comb, p41_res7__217, p41_res7__216, p41_res7__215, p41_res7__214, p41_res7__213, p41_res7__212, p41_res7__211, p41_res7__210, p41_res7__209, p41_res7__208};
  assign p42_xor_1084661_comb = p42_res__13_comb ^ p41_xor_1083717;

  // Registers for pipe stage 42:
  reg [127:0] p42_xor_1084189;
  reg [127:0] p42_xor_1084661;
  reg [127:0] p42_res__35;
  reg [7:0] p43_arr[256];
  reg [7:0] p43_literal_1076345[256];
  reg [7:0] p43_literal_1076347[256];
  reg [7:0] p43_literal_1076349[256];
  reg [7:0] p43_literal_1076351[256];
  reg [7:0] p43_literal_1076353[256];
  reg [7:0] p43_literal_1076355[256];
  reg [7:0] p43_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p42_xor_1084189 <= p41_xor_1084189;
    p42_xor_1084661 <= p42_xor_1084661_comb;
    p42_res__35 <= p41_res__35;
    p43_arr <= p42_arr;
    p43_literal_1076345 <= p42_literal_1076345;
    p43_literal_1076347 <= p42_literal_1076347;
    p43_literal_1076349 <= p42_literal_1076349;
    p43_literal_1076351 <= p42_literal_1076351;
    p43_literal_1076353 <= p42_literal_1076353;
    p43_literal_1076355 <= p42_literal_1076355;
    p43_literal_1076358 <= p42_literal_1076358;
  end

  // ===== Pipe stage 43:
  wire [127:0] p43_addedKey__55_comb;
  wire [7:0] p43_array_index_1084699_comb;
  wire [7:0] p43_array_index_1084700_comb;
  wire [7:0] p43_array_index_1084701_comb;
  wire [7:0] p43_array_index_1084702_comb;
  wire [7:0] p43_array_index_1084703_comb;
  wire [7:0] p43_array_index_1084704_comb;
  wire [7:0] p43_array_index_1084706_comb;
  wire [7:0] p43_array_index_1084708_comb;
  wire [7:0] p43_array_index_1084709_comb;
  wire [7:0] p43_array_index_1084710_comb;
  wire [7:0] p43_array_index_1084711_comb;
  wire [7:0] p43_array_index_1084712_comb;
  wire [7:0] p43_array_index_1084713_comb;
  wire [7:0] p43_array_index_1084715_comb;
  wire [7:0] p43_array_index_1084716_comb;
  wire [7:0] p43_array_index_1084717_comb;
  wire [7:0] p43_array_index_1084718_comb;
  wire [7:0] p43_array_index_1084719_comb;
  wire [7:0] p43_array_index_1084720_comb;
  wire [7:0] p43_array_index_1084721_comb;
  wire [7:0] p43_array_index_1084723_comb;
  wire [7:0] p43_res7__224_comb;
  wire [7:0] p43_array_index_1084732_comb;
  wire [7:0] p43_array_index_1084733_comb;
  wire [7:0] p43_array_index_1084734_comb;
  wire [7:0] p43_array_index_1084735_comb;
  wire [7:0] p43_array_index_1084736_comb;
  wire [7:0] p43_array_index_1084737_comb;
  wire [7:0] p43_res7__225_comb;
  wire [7:0] p43_array_index_1084747_comb;
  wire [7:0] p43_array_index_1084748_comb;
  wire [7:0] p43_array_index_1084749_comb;
  wire [7:0] p43_array_index_1084750_comb;
  wire [7:0] p43_array_index_1084751_comb;
  wire [7:0] p43_res7__226_comb;
  wire [7:0] p43_array_index_1084761_comb;
  wire [7:0] p43_array_index_1084762_comb;
  wire [7:0] p43_array_index_1084763_comb;
  wire [7:0] p43_array_index_1084764_comb;
  wire [7:0] p43_array_index_1084765_comb;
  wire [7:0] p43_res7__227_comb;
  wire [7:0] p43_array_index_1084776_comb;
  wire [7:0] p43_array_index_1084777_comb;
  wire [7:0] p43_array_index_1084778_comb;
  wire [7:0] p43_array_index_1084779_comb;
  wire [7:0] p43_res7__228_comb;
  assign p43_addedKey__55_comb = p42_xor_1084661 ^ 128'h3fb1_b78b_213e_f327_fd0e_14f0_71b0_400f;
  assign p43_array_index_1084699_comb = p42_arr[p43_addedKey__55_comb[127:120]];
  assign p43_array_index_1084700_comb = p42_arr[p43_addedKey__55_comb[119:112]];
  assign p43_array_index_1084701_comb = p42_arr[p43_addedKey__55_comb[111:104]];
  assign p43_array_index_1084702_comb = p42_arr[p43_addedKey__55_comb[103:96]];
  assign p43_array_index_1084703_comb = p42_arr[p43_addedKey__55_comb[95:88]];
  assign p43_array_index_1084704_comb = p42_arr[p43_addedKey__55_comb[87:80]];
  assign p43_array_index_1084706_comb = p42_arr[p43_addedKey__55_comb[71:64]];
  assign p43_array_index_1084708_comb = p42_arr[p43_addedKey__55_comb[55:48]];
  assign p43_array_index_1084709_comb = p42_arr[p43_addedKey__55_comb[47:40]];
  assign p43_array_index_1084710_comb = p42_arr[p43_addedKey__55_comb[39:32]];
  assign p43_array_index_1084711_comb = p42_arr[p43_addedKey__55_comb[31:24]];
  assign p43_array_index_1084712_comb = p42_arr[p43_addedKey__55_comb[23:16]];
  assign p43_array_index_1084713_comb = p42_arr[p43_addedKey__55_comb[15:8]];
  assign p43_array_index_1084715_comb = p42_literal_1076345[p43_array_index_1084699_comb];
  assign p43_array_index_1084716_comb = p42_literal_1076347[p43_array_index_1084700_comb];
  assign p43_array_index_1084717_comb = p42_literal_1076349[p43_array_index_1084701_comb];
  assign p43_array_index_1084718_comb = p42_literal_1076351[p43_array_index_1084702_comb];
  assign p43_array_index_1084719_comb = p42_literal_1076353[p43_array_index_1084703_comb];
  assign p43_array_index_1084720_comb = p42_literal_1076355[p43_array_index_1084704_comb];
  assign p43_array_index_1084721_comb = p42_arr[p43_addedKey__55_comb[79:72]];
  assign p43_array_index_1084723_comb = p42_arr[p43_addedKey__55_comb[63:56]];
  assign p43_res7__224_comb = p43_array_index_1084715_comb ^ p43_array_index_1084716_comb ^ p43_array_index_1084717_comb ^ p43_array_index_1084718_comb ^ p43_array_index_1084719_comb ^ p43_array_index_1084720_comb ^ p43_array_index_1084721_comb ^ p42_literal_1076358[p43_array_index_1084706_comb] ^ p43_array_index_1084723_comb ^ p42_literal_1076355[p43_array_index_1084708_comb] ^ p42_literal_1076353[p43_array_index_1084709_comb] ^ p42_literal_1076351[p43_array_index_1084710_comb] ^ p42_literal_1076349[p43_array_index_1084711_comb] ^ p42_literal_1076347[p43_array_index_1084712_comb] ^ p42_literal_1076345[p43_array_index_1084713_comb] ^ p42_arr[p43_addedKey__55_comb[7:0]];
  assign p43_array_index_1084732_comb = p42_literal_1076345[p43_res7__224_comb];
  assign p43_array_index_1084733_comb = p42_literal_1076347[p43_array_index_1084699_comb];
  assign p43_array_index_1084734_comb = p42_literal_1076349[p43_array_index_1084700_comb];
  assign p43_array_index_1084735_comb = p42_literal_1076351[p43_array_index_1084701_comb];
  assign p43_array_index_1084736_comb = p42_literal_1076353[p43_array_index_1084702_comb];
  assign p43_array_index_1084737_comb = p42_literal_1076355[p43_array_index_1084703_comb];
  assign p43_res7__225_comb = p43_array_index_1084732_comb ^ p43_array_index_1084733_comb ^ p43_array_index_1084734_comb ^ p43_array_index_1084735_comb ^ p43_array_index_1084736_comb ^ p43_array_index_1084737_comb ^ p43_array_index_1084704_comb ^ p42_literal_1076358[p43_array_index_1084721_comb] ^ p43_array_index_1084706_comb ^ p42_literal_1076355[p43_array_index_1084723_comb] ^ p42_literal_1076353[p43_array_index_1084708_comb] ^ p42_literal_1076351[p43_array_index_1084709_comb] ^ p42_literal_1076349[p43_array_index_1084710_comb] ^ p42_literal_1076347[p43_array_index_1084711_comb] ^ p42_literal_1076345[p43_array_index_1084712_comb] ^ p43_array_index_1084713_comb;
  assign p43_array_index_1084747_comb = p42_literal_1076347[p43_res7__224_comb];
  assign p43_array_index_1084748_comb = p42_literal_1076349[p43_array_index_1084699_comb];
  assign p43_array_index_1084749_comb = p42_literal_1076351[p43_array_index_1084700_comb];
  assign p43_array_index_1084750_comb = p42_literal_1076353[p43_array_index_1084701_comb];
  assign p43_array_index_1084751_comb = p42_literal_1076355[p43_array_index_1084702_comb];
  assign p43_res7__226_comb = p42_literal_1076345[p43_res7__225_comb] ^ p43_array_index_1084747_comb ^ p43_array_index_1084748_comb ^ p43_array_index_1084749_comb ^ p43_array_index_1084750_comb ^ p43_array_index_1084751_comb ^ p43_array_index_1084703_comb ^ p42_literal_1076358[p43_array_index_1084704_comb] ^ p43_array_index_1084721_comb ^ p42_literal_1076355[p43_array_index_1084706_comb] ^ p42_literal_1076353[p43_array_index_1084723_comb] ^ p42_literal_1076351[p43_array_index_1084708_comb] ^ p42_literal_1076349[p43_array_index_1084709_comb] ^ p42_literal_1076347[p43_array_index_1084710_comb] ^ p42_literal_1076345[p43_array_index_1084711_comb] ^ p43_array_index_1084712_comb;
  assign p43_array_index_1084761_comb = p42_literal_1076347[p43_res7__225_comb];
  assign p43_array_index_1084762_comb = p42_literal_1076349[p43_res7__224_comb];
  assign p43_array_index_1084763_comb = p42_literal_1076351[p43_array_index_1084699_comb];
  assign p43_array_index_1084764_comb = p42_literal_1076353[p43_array_index_1084700_comb];
  assign p43_array_index_1084765_comb = p42_literal_1076355[p43_array_index_1084701_comb];
  assign p43_res7__227_comb = p42_literal_1076345[p43_res7__226_comb] ^ p43_array_index_1084761_comb ^ p43_array_index_1084762_comb ^ p43_array_index_1084763_comb ^ p43_array_index_1084764_comb ^ p43_array_index_1084765_comb ^ p43_array_index_1084702_comb ^ p42_literal_1076358[p43_array_index_1084703_comb] ^ p43_array_index_1084704_comb ^ p42_literal_1076355[p43_array_index_1084721_comb] ^ p42_literal_1076353[p43_array_index_1084706_comb] ^ p42_literal_1076351[p43_array_index_1084723_comb] ^ p42_literal_1076349[p43_array_index_1084708_comb] ^ p42_literal_1076347[p43_array_index_1084709_comb] ^ p42_literal_1076345[p43_array_index_1084710_comb] ^ p43_array_index_1084711_comb;
  assign p43_array_index_1084776_comb = p42_literal_1076349[p43_res7__225_comb];
  assign p43_array_index_1084777_comb = p42_literal_1076351[p43_res7__224_comb];
  assign p43_array_index_1084778_comb = p42_literal_1076353[p43_array_index_1084699_comb];
  assign p43_array_index_1084779_comb = p42_literal_1076355[p43_array_index_1084700_comb];
  assign p43_res7__228_comb = p42_literal_1076345[p43_res7__227_comb] ^ p42_literal_1076347[p43_res7__226_comb] ^ p43_array_index_1084776_comb ^ p43_array_index_1084777_comb ^ p43_array_index_1084778_comb ^ p43_array_index_1084779_comb ^ p43_array_index_1084701_comb ^ p42_literal_1076358[p43_array_index_1084702_comb] ^ p43_array_index_1084703_comb ^ p43_array_index_1084720_comb ^ p42_literal_1076353[p43_array_index_1084721_comb] ^ p42_literal_1076351[p43_array_index_1084706_comb] ^ p42_literal_1076349[p43_array_index_1084723_comb] ^ p42_literal_1076347[p43_array_index_1084708_comb] ^ p42_literal_1076345[p43_array_index_1084709_comb] ^ p43_array_index_1084710_comb;

  // Registers for pipe stage 43:
  reg [127:0] p43_xor_1084189;
  reg [127:0] p43_xor_1084661;
  reg [7:0] p43_array_index_1084699;
  reg [7:0] p43_array_index_1084700;
  reg [7:0] p43_array_index_1084701;
  reg [7:0] p43_array_index_1084702;
  reg [7:0] p43_array_index_1084703;
  reg [7:0] p43_array_index_1084704;
  reg [7:0] p43_array_index_1084706;
  reg [7:0] p43_array_index_1084708;
  reg [7:0] p43_array_index_1084709;
  reg [7:0] p43_array_index_1084715;
  reg [7:0] p43_array_index_1084716;
  reg [7:0] p43_array_index_1084717;
  reg [7:0] p43_array_index_1084718;
  reg [7:0] p43_array_index_1084719;
  reg [7:0] p43_array_index_1084721;
  reg [7:0] p43_array_index_1084723;
  reg [7:0] p43_res7__224;
  reg [7:0] p43_array_index_1084732;
  reg [7:0] p43_array_index_1084733;
  reg [7:0] p43_array_index_1084734;
  reg [7:0] p43_array_index_1084735;
  reg [7:0] p43_array_index_1084736;
  reg [7:0] p43_array_index_1084737;
  reg [7:0] p43_res7__225;
  reg [7:0] p43_array_index_1084747;
  reg [7:0] p43_array_index_1084748;
  reg [7:0] p43_array_index_1084749;
  reg [7:0] p43_array_index_1084750;
  reg [7:0] p43_array_index_1084751;
  reg [7:0] p43_res7__226;
  reg [7:0] p43_array_index_1084761;
  reg [7:0] p43_array_index_1084762;
  reg [7:0] p43_array_index_1084763;
  reg [7:0] p43_array_index_1084764;
  reg [7:0] p43_array_index_1084765;
  reg [7:0] p43_res7__227;
  reg [7:0] p43_array_index_1084776;
  reg [7:0] p43_array_index_1084777;
  reg [7:0] p43_array_index_1084778;
  reg [7:0] p43_array_index_1084779;
  reg [7:0] p43_res7__228;
  reg [127:0] p43_res__35;
  reg [7:0] p44_arr[256];
  reg [7:0] p44_literal_1076345[256];
  reg [7:0] p44_literal_1076347[256];
  reg [7:0] p44_literal_1076349[256];
  reg [7:0] p44_literal_1076351[256];
  reg [7:0] p44_literal_1076353[256];
  reg [7:0] p44_literal_1076355[256];
  reg [7:0] p44_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p43_xor_1084189 <= p42_xor_1084189;
    p43_xor_1084661 <= p42_xor_1084661;
    p43_array_index_1084699 <= p43_array_index_1084699_comb;
    p43_array_index_1084700 <= p43_array_index_1084700_comb;
    p43_array_index_1084701 <= p43_array_index_1084701_comb;
    p43_array_index_1084702 <= p43_array_index_1084702_comb;
    p43_array_index_1084703 <= p43_array_index_1084703_comb;
    p43_array_index_1084704 <= p43_array_index_1084704_comb;
    p43_array_index_1084706 <= p43_array_index_1084706_comb;
    p43_array_index_1084708 <= p43_array_index_1084708_comb;
    p43_array_index_1084709 <= p43_array_index_1084709_comb;
    p43_array_index_1084715 <= p43_array_index_1084715_comb;
    p43_array_index_1084716 <= p43_array_index_1084716_comb;
    p43_array_index_1084717 <= p43_array_index_1084717_comb;
    p43_array_index_1084718 <= p43_array_index_1084718_comb;
    p43_array_index_1084719 <= p43_array_index_1084719_comb;
    p43_array_index_1084721 <= p43_array_index_1084721_comb;
    p43_array_index_1084723 <= p43_array_index_1084723_comb;
    p43_res7__224 <= p43_res7__224_comb;
    p43_array_index_1084732 <= p43_array_index_1084732_comb;
    p43_array_index_1084733 <= p43_array_index_1084733_comb;
    p43_array_index_1084734 <= p43_array_index_1084734_comb;
    p43_array_index_1084735 <= p43_array_index_1084735_comb;
    p43_array_index_1084736 <= p43_array_index_1084736_comb;
    p43_array_index_1084737 <= p43_array_index_1084737_comb;
    p43_res7__225 <= p43_res7__225_comb;
    p43_array_index_1084747 <= p43_array_index_1084747_comb;
    p43_array_index_1084748 <= p43_array_index_1084748_comb;
    p43_array_index_1084749 <= p43_array_index_1084749_comb;
    p43_array_index_1084750 <= p43_array_index_1084750_comb;
    p43_array_index_1084751 <= p43_array_index_1084751_comb;
    p43_res7__226 <= p43_res7__226_comb;
    p43_array_index_1084761 <= p43_array_index_1084761_comb;
    p43_array_index_1084762 <= p43_array_index_1084762_comb;
    p43_array_index_1084763 <= p43_array_index_1084763_comb;
    p43_array_index_1084764 <= p43_array_index_1084764_comb;
    p43_array_index_1084765 <= p43_array_index_1084765_comb;
    p43_res7__227 <= p43_res7__227_comb;
    p43_array_index_1084776 <= p43_array_index_1084776_comb;
    p43_array_index_1084777 <= p43_array_index_1084777_comb;
    p43_array_index_1084778 <= p43_array_index_1084778_comb;
    p43_array_index_1084779 <= p43_array_index_1084779_comb;
    p43_res7__228 <= p43_res7__228_comb;
    p43_res__35 <= p42_res__35;
    p44_arr <= p43_arr;
    p44_literal_1076345 <= p43_literal_1076345;
    p44_literal_1076347 <= p43_literal_1076347;
    p44_literal_1076349 <= p43_literal_1076349;
    p44_literal_1076351 <= p43_literal_1076351;
    p44_literal_1076353 <= p43_literal_1076353;
    p44_literal_1076355 <= p43_literal_1076355;
    p44_literal_1076358 <= p43_literal_1076358;
  end

  // ===== Pipe stage 44:
  wire [7:0] p44_array_index_1084893_comb;
  wire [7:0] p44_array_index_1084894_comb;
  wire [7:0] p44_array_index_1084895_comb;
  wire [7:0] p44_array_index_1084896_comb;
  wire [7:0] p44_res7__229_comb;
  wire [7:0] p44_array_index_1084907_comb;
  wire [7:0] p44_array_index_1084908_comb;
  wire [7:0] p44_array_index_1084909_comb;
  wire [7:0] p44_res7__230_comb;
  wire [7:0] p44_array_index_1084919_comb;
  wire [7:0] p44_array_index_1084920_comb;
  wire [7:0] p44_array_index_1084921_comb;
  wire [7:0] p44_res7__231_comb;
  wire [7:0] p44_array_index_1084932_comb;
  wire [7:0] p44_array_index_1084933_comb;
  wire [7:0] p44_res7__232_comb;
  wire [7:0] p44_array_index_1084943_comb;
  wire [7:0] p44_array_index_1084944_comb;
  wire [7:0] p44_res7__233_comb;
  wire [7:0] p44_array_index_1084950_comb;
  wire [7:0] p44_array_index_1084951_comb;
  wire [7:0] p44_array_index_1084952_comb;
  wire [7:0] p44_array_index_1084953_comb;
  wire [7:0] p44_array_index_1084954_comb;
  wire [7:0] p44_array_index_1084955_comb;
  wire [7:0] p44_array_index_1084956_comb;
  wire [7:0] p44_array_index_1084957_comb;
  wire [7:0] p44_array_index_1084958_comb;
  assign p44_array_index_1084893_comb = p43_literal_1076349[p43_res7__226];
  assign p44_array_index_1084894_comb = p43_literal_1076351[p43_res7__225];
  assign p44_array_index_1084895_comb = p43_literal_1076353[p43_res7__224];
  assign p44_array_index_1084896_comb = p43_literal_1076355[p43_array_index_1084699];
  assign p44_res7__229_comb = p43_literal_1076345[p43_res7__228] ^ p43_literal_1076347[p43_res7__227] ^ p44_array_index_1084893_comb ^ p44_array_index_1084894_comb ^ p44_array_index_1084895_comb ^ p44_array_index_1084896_comb ^ p43_array_index_1084700 ^ p43_literal_1076358[p43_array_index_1084701] ^ p43_array_index_1084702 ^ p43_array_index_1084737 ^ p43_literal_1076353[p43_array_index_1084704] ^ p43_literal_1076351[p43_array_index_1084721] ^ p43_literal_1076349[p43_array_index_1084706] ^ p43_literal_1076347[p43_array_index_1084723] ^ p43_literal_1076345[p43_array_index_1084708] ^ p43_array_index_1084709;
  assign p44_array_index_1084907_comb = p43_literal_1076351[p43_res7__226];
  assign p44_array_index_1084908_comb = p43_literal_1076353[p43_res7__225];
  assign p44_array_index_1084909_comb = p43_literal_1076355[p43_res7__224];
  assign p44_res7__230_comb = p43_literal_1076345[p44_res7__229_comb] ^ p43_literal_1076347[p43_res7__228] ^ p43_literal_1076349[p43_res7__227] ^ p44_array_index_1084907_comb ^ p44_array_index_1084908_comb ^ p44_array_index_1084909_comb ^ p43_array_index_1084699 ^ p43_literal_1076358[p43_array_index_1084700] ^ p43_array_index_1084701 ^ p43_array_index_1084751 ^ p43_array_index_1084719 ^ p43_literal_1076351[p43_array_index_1084704] ^ p43_literal_1076349[p43_array_index_1084721] ^ p43_literal_1076347[p43_array_index_1084706] ^ p43_literal_1076345[p43_array_index_1084723] ^ p43_array_index_1084708;
  assign p44_array_index_1084919_comb = p43_literal_1076351[p43_res7__227];
  assign p44_array_index_1084920_comb = p43_literal_1076353[p43_res7__226];
  assign p44_array_index_1084921_comb = p43_literal_1076355[p43_res7__225];
  assign p44_res7__231_comb = p43_literal_1076345[p44_res7__230_comb] ^ p43_literal_1076347[p44_res7__229_comb] ^ p43_literal_1076349[p43_res7__228] ^ p44_array_index_1084919_comb ^ p44_array_index_1084920_comb ^ p44_array_index_1084921_comb ^ p43_res7__224 ^ p43_literal_1076358[p43_array_index_1084699] ^ p43_array_index_1084700 ^ p43_array_index_1084765 ^ p43_array_index_1084736 ^ p43_literal_1076351[p43_array_index_1084703] ^ p43_literal_1076349[p43_array_index_1084704] ^ p43_literal_1076347[p43_array_index_1084721] ^ p43_literal_1076345[p43_array_index_1084706] ^ p43_array_index_1084723;
  assign p44_array_index_1084932_comb = p43_literal_1076353[p43_res7__227];
  assign p44_array_index_1084933_comb = p43_literal_1076355[p43_res7__226];
  assign p44_res7__232_comb = p43_literal_1076345[p44_res7__231_comb] ^ p43_literal_1076347[p44_res7__230_comb] ^ p43_literal_1076349[p44_res7__229_comb] ^ p43_literal_1076351[p43_res7__228] ^ p44_array_index_1084932_comb ^ p44_array_index_1084933_comb ^ p43_res7__225 ^ p43_literal_1076358[p43_res7__224] ^ p43_array_index_1084699 ^ p43_array_index_1084779 ^ p43_array_index_1084750 ^ p43_array_index_1084718 ^ p43_literal_1076349[p43_array_index_1084703] ^ p43_literal_1076347[p43_array_index_1084704] ^ p43_literal_1076345[p43_array_index_1084721] ^ p43_array_index_1084706;
  assign p44_array_index_1084943_comb = p43_literal_1076353[p43_res7__228];
  assign p44_array_index_1084944_comb = p43_literal_1076355[p43_res7__227];
  assign p44_res7__233_comb = p43_literal_1076345[p44_res7__232_comb] ^ p43_literal_1076347[p44_res7__231_comb] ^ p43_literal_1076349[p44_res7__230_comb] ^ p43_literal_1076351[p44_res7__229_comb] ^ p44_array_index_1084943_comb ^ p44_array_index_1084944_comb ^ p43_res7__226 ^ p43_literal_1076358[p43_res7__225] ^ p43_res7__224 ^ p44_array_index_1084896_comb ^ p43_array_index_1084764 ^ p43_array_index_1084735 ^ p43_literal_1076349[p43_array_index_1084702] ^ p43_literal_1076347[p43_array_index_1084703] ^ p43_literal_1076345[p43_array_index_1084704] ^ p43_array_index_1084721;
  assign p44_array_index_1084950_comb = p43_literal_1076345[p44_res7__233_comb];
  assign p44_array_index_1084951_comb = p43_literal_1076347[p44_res7__232_comb];
  assign p44_array_index_1084952_comb = p43_literal_1076349[p44_res7__231_comb];
  assign p44_array_index_1084953_comb = p43_literal_1076351[p44_res7__230_comb];
  assign p44_array_index_1084954_comb = p43_literal_1076353[p44_res7__229_comb];
  assign p44_array_index_1084955_comb = p43_literal_1076355[p43_res7__228];
  assign p44_array_index_1084956_comb = p43_literal_1076358[p43_res7__226];
  assign p44_array_index_1084957_comb = p43_literal_1076347[p43_array_index_1084702];
  assign p44_array_index_1084958_comb = p43_literal_1076345[p43_array_index_1084703];

  // Registers for pipe stage 44:
  reg [127:0] p44_xor_1084189;
  reg [127:0] p44_xor_1084661;
  reg [7:0] p44_array_index_1084699;
  reg [7:0] p44_array_index_1084700;
  reg [7:0] p44_array_index_1084701;
  reg [7:0] p44_array_index_1084702;
  reg [7:0] p44_array_index_1084703;
  reg [7:0] p44_array_index_1084704;
  reg [7:0] p44_array_index_1084715;
  reg [7:0] p44_array_index_1084716;
  reg [7:0] p44_array_index_1084717;
  reg [7:0] p44_res7__224;
  reg [7:0] p44_array_index_1084732;
  reg [7:0] p44_array_index_1084733;
  reg [7:0] p44_array_index_1084734;
  reg [7:0] p44_res7__225;
  reg [7:0] p44_array_index_1084747;
  reg [7:0] p44_array_index_1084748;
  reg [7:0] p44_array_index_1084749;
  reg [7:0] p44_res7__226;
  reg [7:0] p44_array_index_1084761;
  reg [7:0] p44_array_index_1084762;
  reg [7:0] p44_array_index_1084763;
  reg [7:0] p44_res7__227;
  reg [7:0] p44_array_index_1084776;
  reg [7:0] p44_array_index_1084777;
  reg [7:0] p44_array_index_1084778;
  reg [7:0] p44_res7__228;
  reg [7:0] p44_array_index_1084893;
  reg [7:0] p44_array_index_1084894;
  reg [7:0] p44_array_index_1084895;
  reg [7:0] p44_res7__229;
  reg [7:0] p44_array_index_1084907;
  reg [7:0] p44_array_index_1084908;
  reg [7:0] p44_array_index_1084909;
  reg [7:0] p44_res7__230;
  reg [7:0] p44_array_index_1084919;
  reg [7:0] p44_array_index_1084920;
  reg [7:0] p44_array_index_1084921;
  reg [7:0] p44_res7__231;
  reg [7:0] p44_array_index_1084932;
  reg [7:0] p44_array_index_1084933;
  reg [7:0] p44_res7__232;
  reg [7:0] p44_array_index_1084943;
  reg [7:0] p44_array_index_1084944;
  reg [7:0] p44_res7__233;
  reg [7:0] p44_array_index_1084950;
  reg [7:0] p44_array_index_1084951;
  reg [7:0] p44_array_index_1084952;
  reg [7:0] p44_array_index_1084953;
  reg [7:0] p44_array_index_1084954;
  reg [7:0] p44_array_index_1084955;
  reg [7:0] p44_array_index_1084956;
  reg [7:0] p44_array_index_1084957;
  reg [7:0] p44_array_index_1084958;
  reg [127:0] p44_res__35;
  reg [7:0] p45_arr[256];
  reg [7:0] p45_literal_1076345[256];
  reg [7:0] p45_literal_1076347[256];
  reg [7:0] p45_literal_1076349[256];
  reg [7:0] p45_literal_1076351[256];
  reg [7:0] p45_literal_1076353[256];
  reg [7:0] p45_literal_1076355[256];
  reg [7:0] p45_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p44_xor_1084189 <= p43_xor_1084189;
    p44_xor_1084661 <= p43_xor_1084661;
    p44_array_index_1084699 <= p43_array_index_1084699;
    p44_array_index_1084700 <= p43_array_index_1084700;
    p44_array_index_1084701 <= p43_array_index_1084701;
    p44_array_index_1084702 <= p43_array_index_1084702;
    p44_array_index_1084703 <= p43_array_index_1084703;
    p44_array_index_1084704 <= p43_array_index_1084704;
    p44_array_index_1084715 <= p43_array_index_1084715;
    p44_array_index_1084716 <= p43_array_index_1084716;
    p44_array_index_1084717 <= p43_array_index_1084717;
    p44_res7__224 <= p43_res7__224;
    p44_array_index_1084732 <= p43_array_index_1084732;
    p44_array_index_1084733 <= p43_array_index_1084733;
    p44_array_index_1084734 <= p43_array_index_1084734;
    p44_res7__225 <= p43_res7__225;
    p44_array_index_1084747 <= p43_array_index_1084747;
    p44_array_index_1084748 <= p43_array_index_1084748;
    p44_array_index_1084749 <= p43_array_index_1084749;
    p44_res7__226 <= p43_res7__226;
    p44_array_index_1084761 <= p43_array_index_1084761;
    p44_array_index_1084762 <= p43_array_index_1084762;
    p44_array_index_1084763 <= p43_array_index_1084763;
    p44_res7__227 <= p43_res7__227;
    p44_array_index_1084776 <= p43_array_index_1084776;
    p44_array_index_1084777 <= p43_array_index_1084777;
    p44_array_index_1084778 <= p43_array_index_1084778;
    p44_res7__228 <= p43_res7__228;
    p44_array_index_1084893 <= p44_array_index_1084893_comb;
    p44_array_index_1084894 <= p44_array_index_1084894_comb;
    p44_array_index_1084895 <= p44_array_index_1084895_comb;
    p44_res7__229 <= p44_res7__229_comb;
    p44_array_index_1084907 <= p44_array_index_1084907_comb;
    p44_array_index_1084908 <= p44_array_index_1084908_comb;
    p44_array_index_1084909 <= p44_array_index_1084909_comb;
    p44_res7__230 <= p44_res7__230_comb;
    p44_array_index_1084919 <= p44_array_index_1084919_comb;
    p44_array_index_1084920 <= p44_array_index_1084920_comb;
    p44_array_index_1084921 <= p44_array_index_1084921_comb;
    p44_res7__231 <= p44_res7__231_comb;
    p44_array_index_1084932 <= p44_array_index_1084932_comb;
    p44_array_index_1084933 <= p44_array_index_1084933_comb;
    p44_res7__232 <= p44_res7__232_comb;
    p44_array_index_1084943 <= p44_array_index_1084943_comb;
    p44_array_index_1084944 <= p44_array_index_1084944_comb;
    p44_res7__233 <= p44_res7__233_comb;
    p44_array_index_1084950 <= p44_array_index_1084950_comb;
    p44_array_index_1084951 <= p44_array_index_1084951_comb;
    p44_array_index_1084952 <= p44_array_index_1084952_comb;
    p44_array_index_1084953 <= p44_array_index_1084953_comb;
    p44_array_index_1084954 <= p44_array_index_1084954_comb;
    p44_array_index_1084955 <= p44_array_index_1084955_comb;
    p44_array_index_1084956 <= p44_array_index_1084956_comb;
    p44_array_index_1084957 <= p44_array_index_1084957_comb;
    p44_array_index_1084958 <= p44_array_index_1084958_comb;
    p44_res__35 <= p43_res__35;
    p45_arr <= p44_arr;
    p45_literal_1076345 <= p44_literal_1076345;
    p45_literal_1076347 <= p44_literal_1076347;
    p45_literal_1076349 <= p44_literal_1076349;
    p45_literal_1076351 <= p44_literal_1076351;
    p45_literal_1076353 <= p44_literal_1076353;
    p45_literal_1076355 <= p44_literal_1076355;
    p45_literal_1076358 <= p44_literal_1076358;
  end

  // ===== Pipe stage 45:
  wire [7:0] p45_res7__234_comb;
  wire [7:0] p45_array_index_1085093_comb;
  wire [7:0] p45_res7__235_comb;
  wire [7:0] p45_res7__236_comb;
  wire [7:0] p45_res7__237_comb;
  wire [7:0] p45_res7__238_comb;
  wire [7:0] p45_res7__239_comb;
  wire [127:0] p45_res__14_comb;
  wire [127:0] p45_k5_comb;
  assign p45_res7__234_comb = p44_array_index_1084950 ^ p44_array_index_1084951 ^ p44_array_index_1084952 ^ p44_array_index_1084953 ^ p44_array_index_1084954 ^ p44_array_index_1084955 ^ p44_res7__227 ^ p44_array_index_1084956 ^ p44_res7__225 ^ p44_array_index_1084909 ^ p44_array_index_1084778 ^ p44_array_index_1084749 ^ p44_array_index_1084717 ^ p44_array_index_1084957 ^ p44_array_index_1084958 ^ p44_array_index_1084704;
  assign p45_array_index_1085093_comb = p44_literal_1076355[p44_res7__229];
  assign p45_res7__235_comb = p44_literal_1076345[p45_res7__234_comb] ^ p44_literal_1076347[p44_res7__233] ^ p44_literal_1076349[p44_res7__232] ^ p44_literal_1076351[p44_res7__231] ^ p44_literal_1076353[p44_res7__230] ^ p45_array_index_1085093_comb ^ p44_res7__228 ^ p44_literal_1076358[p44_res7__227] ^ p44_res7__226 ^ p44_array_index_1084921 ^ p44_array_index_1084895 ^ p44_array_index_1084763 ^ p44_array_index_1084734 ^ p44_literal_1076347[p44_array_index_1084701] ^ p44_literal_1076345[p44_array_index_1084702] ^ p44_array_index_1084703;
  assign p45_res7__236_comb = p44_literal_1076345[p45_res7__235_comb] ^ p44_literal_1076347[p45_res7__234_comb] ^ p44_literal_1076349[p44_res7__233] ^ p44_literal_1076351[p44_res7__232] ^ p44_literal_1076353[p44_res7__231] ^ p44_literal_1076355[p44_res7__230] ^ p44_res7__229 ^ p44_literal_1076358[p44_res7__228] ^ p44_res7__227 ^ p44_array_index_1084933 ^ p44_array_index_1084908 ^ p44_array_index_1084777 ^ p44_array_index_1084748 ^ p44_array_index_1084716 ^ p44_literal_1076345[p44_array_index_1084701] ^ p44_array_index_1084702;
  assign p45_res7__237_comb = p44_literal_1076345[p45_res7__236_comb] ^ p44_literal_1076347[p45_res7__235_comb] ^ p44_literal_1076349[p45_res7__234_comb] ^ p44_literal_1076351[p44_res7__233] ^ p44_literal_1076353[p44_res7__232] ^ p44_literal_1076355[p44_res7__231] ^ p44_res7__230 ^ p44_literal_1076358[p44_res7__229] ^ p44_res7__228 ^ p44_array_index_1084944 ^ p44_array_index_1084920 ^ p44_array_index_1084894 ^ p44_array_index_1084762 ^ p44_array_index_1084733 ^ p44_literal_1076345[p44_array_index_1084700] ^ p44_array_index_1084701;
  assign p45_res7__238_comb = p44_literal_1076345[p45_res7__237_comb] ^ p44_literal_1076347[p45_res7__236_comb] ^ p44_literal_1076349[p45_res7__235_comb] ^ p44_literal_1076351[p45_res7__234_comb] ^ p44_literal_1076353[p44_res7__233] ^ p44_literal_1076355[p44_res7__232] ^ p44_res7__231 ^ p44_literal_1076358[p44_res7__230] ^ p44_res7__229 ^ p44_array_index_1084955 ^ p44_array_index_1084932 ^ p44_array_index_1084907 ^ p44_array_index_1084776 ^ p44_array_index_1084747 ^ p44_array_index_1084715 ^ p44_array_index_1084700;
  assign p45_res7__239_comb = p44_literal_1076345[p45_res7__238_comb] ^ p44_literal_1076347[p45_res7__237_comb] ^ p44_literal_1076349[p45_res7__236_comb] ^ p44_literal_1076351[p45_res7__235_comb] ^ p44_literal_1076353[p45_res7__234_comb] ^ p44_literal_1076355[p44_res7__233] ^ p44_res7__232 ^ p44_literal_1076358[p44_res7__231] ^ p44_res7__230 ^ p45_array_index_1085093_comb ^ p44_array_index_1084943 ^ p44_array_index_1084919 ^ p44_array_index_1084893 ^ p44_array_index_1084761 ^ p44_array_index_1084732 ^ p44_array_index_1084699;
  assign p45_res__14_comb = {p45_res7__239_comb, p45_res7__238_comb, p45_res7__237_comb, p45_res7__236_comb, p45_res7__235_comb, p45_res7__234_comb, p44_res7__233, p44_res7__232, p44_res7__231, p44_res7__230, p44_res7__229, p44_res7__228, p44_res7__227, p44_res7__226, p44_res7__225, p44_res7__224};
  assign p45_k5_comb = p45_res__14_comb ^ p44_xor_1084189;

  // Registers for pipe stage 45:
  reg [127:0] p45_xor_1084661;
  reg [127:0] p45_k5;
  reg [127:0] p45_res__35;
  reg [7:0] p46_arr[256];
  reg [7:0] p46_literal_1076345[256];
  reg [7:0] p46_literal_1076347[256];
  reg [7:0] p46_literal_1076349[256];
  reg [7:0] p46_literal_1076351[256];
  reg [7:0] p46_literal_1076353[256];
  reg [7:0] p46_literal_1076355[256];
  reg [7:0] p46_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p45_xor_1084661 <= p44_xor_1084661;
    p45_k5 <= p45_k5_comb;
    p45_res__35 <= p44_res__35;
    p46_arr <= p45_arr;
    p46_literal_1076345 <= p45_literal_1076345;
    p46_literal_1076347 <= p45_literal_1076347;
    p46_literal_1076349 <= p45_literal_1076349;
    p46_literal_1076351 <= p45_literal_1076351;
    p46_literal_1076353 <= p45_literal_1076353;
    p46_literal_1076355 <= p45_literal_1076355;
    p46_literal_1076358 <= p45_literal_1076358;
  end

  // ===== Pipe stage 46:
  wire [127:0] p46_addedKey__56_comb;
  wire [7:0] p46_array_index_1085171_comb;
  wire [7:0] p46_array_index_1085172_comb;
  wire [7:0] p46_array_index_1085173_comb;
  wire [7:0] p46_array_index_1085174_comb;
  wire [7:0] p46_array_index_1085175_comb;
  wire [7:0] p46_array_index_1085176_comb;
  wire [7:0] p46_array_index_1085178_comb;
  wire [7:0] p46_array_index_1085180_comb;
  wire [7:0] p46_array_index_1085181_comb;
  wire [7:0] p46_array_index_1085182_comb;
  wire [7:0] p46_array_index_1085183_comb;
  wire [7:0] p46_array_index_1085184_comb;
  wire [7:0] p46_array_index_1085185_comb;
  wire [7:0] p46_array_index_1085187_comb;
  wire [7:0] p46_array_index_1085188_comb;
  wire [7:0] p46_array_index_1085189_comb;
  wire [7:0] p46_array_index_1085190_comb;
  wire [7:0] p46_array_index_1085191_comb;
  wire [7:0] p46_array_index_1085192_comb;
  wire [7:0] p46_array_index_1085193_comb;
  wire [7:0] p46_array_index_1085195_comb;
  wire [7:0] p46_res7__240_comb;
  wire [7:0] p46_array_index_1085204_comb;
  wire [7:0] p46_array_index_1085205_comb;
  wire [7:0] p46_array_index_1085206_comb;
  wire [7:0] p46_array_index_1085207_comb;
  wire [7:0] p46_array_index_1085208_comb;
  wire [7:0] p46_array_index_1085209_comb;
  wire [7:0] p46_res7__241_comb;
  wire [7:0] p46_array_index_1085219_comb;
  wire [7:0] p46_array_index_1085220_comb;
  wire [7:0] p46_array_index_1085221_comb;
  wire [7:0] p46_array_index_1085222_comb;
  wire [7:0] p46_array_index_1085223_comb;
  wire [7:0] p46_res7__242_comb;
  wire [7:0] p46_array_index_1085233_comb;
  wire [7:0] p46_array_index_1085234_comb;
  wire [7:0] p46_array_index_1085235_comb;
  wire [7:0] p46_array_index_1085236_comb;
  wire [7:0] p46_array_index_1085237_comb;
  wire [7:0] p46_res7__243_comb;
  wire [7:0] p46_array_index_1085248_comb;
  wire [7:0] p46_array_index_1085249_comb;
  wire [7:0] p46_array_index_1085250_comb;
  wire [7:0] p46_array_index_1085251_comb;
  wire [7:0] p46_res7__244_comb;
  assign p46_addedKey__56_comb = p45_k5 ^ 128'h2fb2_6c2c_0f0a_acd1_9935_81c3_4e97_5410;
  assign p46_array_index_1085171_comb = p45_arr[p46_addedKey__56_comb[127:120]];
  assign p46_array_index_1085172_comb = p45_arr[p46_addedKey__56_comb[119:112]];
  assign p46_array_index_1085173_comb = p45_arr[p46_addedKey__56_comb[111:104]];
  assign p46_array_index_1085174_comb = p45_arr[p46_addedKey__56_comb[103:96]];
  assign p46_array_index_1085175_comb = p45_arr[p46_addedKey__56_comb[95:88]];
  assign p46_array_index_1085176_comb = p45_arr[p46_addedKey__56_comb[87:80]];
  assign p46_array_index_1085178_comb = p45_arr[p46_addedKey__56_comb[71:64]];
  assign p46_array_index_1085180_comb = p45_arr[p46_addedKey__56_comb[55:48]];
  assign p46_array_index_1085181_comb = p45_arr[p46_addedKey__56_comb[47:40]];
  assign p46_array_index_1085182_comb = p45_arr[p46_addedKey__56_comb[39:32]];
  assign p46_array_index_1085183_comb = p45_arr[p46_addedKey__56_comb[31:24]];
  assign p46_array_index_1085184_comb = p45_arr[p46_addedKey__56_comb[23:16]];
  assign p46_array_index_1085185_comb = p45_arr[p46_addedKey__56_comb[15:8]];
  assign p46_array_index_1085187_comb = p45_literal_1076345[p46_array_index_1085171_comb];
  assign p46_array_index_1085188_comb = p45_literal_1076347[p46_array_index_1085172_comb];
  assign p46_array_index_1085189_comb = p45_literal_1076349[p46_array_index_1085173_comb];
  assign p46_array_index_1085190_comb = p45_literal_1076351[p46_array_index_1085174_comb];
  assign p46_array_index_1085191_comb = p45_literal_1076353[p46_array_index_1085175_comb];
  assign p46_array_index_1085192_comb = p45_literal_1076355[p46_array_index_1085176_comb];
  assign p46_array_index_1085193_comb = p45_arr[p46_addedKey__56_comb[79:72]];
  assign p46_array_index_1085195_comb = p45_arr[p46_addedKey__56_comb[63:56]];
  assign p46_res7__240_comb = p46_array_index_1085187_comb ^ p46_array_index_1085188_comb ^ p46_array_index_1085189_comb ^ p46_array_index_1085190_comb ^ p46_array_index_1085191_comb ^ p46_array_index_1085192_comb ^ p46_array_index_1085193_comb ^ p45_literal_1076358[p46_array_index_1085178_comb] ^ p46_array_index_1085195_comb ^ p45_literal_1076355[p46_array_index_1085180_comb] ^ p45_literal_1076353[p46_array_index_1085181_comb] ^ p45_literal_1076351[p46_array_index_1085182_comb] ^ p45_literal_1076349[p46_array_index_1085183_comb] ^ p45_literal_1076347[p46_array_index_1085184_comb] ^ p45_literal_1076345[p46_array_index_1085185_comb] ^ p45_arr[p46_addedKey__56_comb[7:0]];
  assign p46_array_index_1085204_comb = p45_literal_1076345[p46_res7__240_comb];
  assign p46_array_index_1085205_comb = p45_literal_1076347[p46_array_index_1085171_comb];
  assign p46_array_index_1085206_comb = p45_literal_1076349[p46_array_index_1085172_comb];
  assign p46_array_index_1085207_comb = p45_literal_1076351[p46_array_index_1085173_comb];
  assign p46_array_index_1085208_comb = p45_literal_1076353[p46_array_index_1085174_comb];
  assign p46_array_index_1085209_comb = p45_literal_1076355[p46_array_index_1085175_comb];
  assign p46_res7__241_comb = p46_array_index_1085204_comb ^ p46_array_index_1085205_comb ^ p46_array_index_1085206_comb ^ p46_array_index_1085207_comb ^ p46_array_index_1085208_comb ^ p46_array_index_1085209_comb ^ p46_array_index_1085176_comb ^ p45_literal_1076358[p46_array_index_1085193_comb] ^ p46_array_index_1085178_comb ^ p45_literal_1076355[p46_array_index_1085195_comb] ^ p45_literal_1076353[p46_array_index_1085180_comb] ^ p45_literal_1076351[p46_array_index_1085181_comb] ^ p45_literal_1076349[p46_array_index_1085182_comb] ^ p45_literal_1076347[p46_array_index_1085183_comb] ^ p45_literal_1076345[p46_array_index_1085184_comb] ^ p46_array_index_1085185_comb;
  assign p46_array_index_1085219_comb = p45_literal_1076347[p46_res7__240_comb];
  assign p46_array_index_1085220_comb = p45_literal_1076349[p46_array_index_1085171_comb];
  assign p46_array_index_1085221_comb = p45_literal_1076351[p46_array_index_1085172_comb];
  assign p46_array_index_1085222_comb = p45_literal_1076353[p46_array_index_1085173_comb];
  assign p46_array_index_1085223_comb = p45_literal_1076355[p46_array_index_1085174_comb];
  assign p46_res7__242_comb = p45_literal_1076345[p46_res7__241_comb] ^ p46_array_index_1085219_comb ^ p46_array_index_1085220_comb ^ p46_array_index_1085221_comb ^ p46_array_index_1085222_comb ^ p46_array_index_1085223_comb ^ p46_array_index_1085175_comb ^ p45_literal_1076358[p46_array_index_1085176_comb] ^ p46_array_index_1085193_comb ^ p45_literal_1076355[p46_array_index_1085178_comb] ^ p45_literal_1076353[p46_array_index_1085195_comb] ^ p45_literal_1076351[p46_array_index_1085180_comb] ^ p45_literal_1076349[p46_array_index_1085181_comb] ^ p45_literal_1076347[p46_array_index_1085182_comb] ^ p45_literal_1076345[p46_array_index_1085183_comb] ^ p46_array_index_1085184_comb;
  assign p46_array_index_1085233_comb = p45_literal_1076347[p46_res7__241_comb];
  assign p46_array_index_1085234_comb = p45_literal_1076349[p46_res7__240_comb];
  assign p46_array_index_1085235_comb = p45_literal_1076351[p46_array_index_1085171_comb];
  assign p46_array_index_1085236_comb = p45_literal_1076353[p46_array_index_1085172_comb];
  assign p46_array_index_1085237_comb = p45_literal_1076355[p46_array_index_1085173_comb];
  assign p46_res7__243_comb = p45_literal_1076345[p46_res7__242_comb] ^ p46_array_index_1085233_comb ^ p46_array_index_1085234_comb ^ p46_array_index_1085235_comb ^ p46_array_index_1085236_comb ^ p46_array_index_1085237_comb ^ p46_array_index_1085174_comb ^ p45_literal_1076358[p46_array_index_1085175_comb] ^ p46_array_index_1085176_comb ^ p45_literal_1076355[p46_array_index_1085193_comb] ^ p45_literal_1076353[p46_array_index_1085178_comb] ^ p45_literal_1076351[p46_array_index_1085195_comb] ^ p45_literal_1076349[p46_array_index_1085180_comb] ^ p45_literal_1076347[p46_array_index_1085181_comb] ^ p45_literal_1076345[p46_array_index_1085182_comb] ^ p46_array_index_1085183_comb;
  assign p46_array_index_1085248_comb = p45_literal_1076349[p46_res7__241_comb];
  assign p46_array_index_1085249_comb = p45_literal_1076351[p46_res7__240_comb];
  assign p46_array_index_1085250_comb = p45_literal_1076353[p46_array_index_1085171_comb];
  assign p46_array_index_1085251_comb = p45_literal_1076355[p46_array_index_1085172_comb];
  assign p46_res7__244_comb = p45_literal_1076345[p46_res7__243_comb] ^ p45_literal_1076347[p46_res7__242_comb] ^ p46_array_index_1085248_comb ^ p46_array_index_1085249_comb ^ p46_array_index_1085250_comb ^ p46_array_index_1085251_comb ^ p46_array_index_1085173_comb ^ p45_literal_1076358[p46_array_index_1085174_comb] ^ p46_array_index_1085175_comb ^ p46_array_index_1085192_comb ^ p45_literal_1076353[p46_array_index_1085193_comb] ^ p45_literal_1076351[p46_array_index_1085178_comb] ^ p45_literal_1076349[p46_array_index_1085195_comb] ^ p45_literal_1076347[p46_array_index_1085180_comb] ^ p45_literal_1076345[p46_array_index_1085181_comb] ^ p46_array_index_1085182_comb;

  // Registers for pipe stage 46:
  reg [127:0] p46_xor_1084661;
  reg [127:0] p46_k5;
  reg [7:0] p46_array_index_1085171;
  reg [7:0] p46_array_index_1085172;
  reg [7:0] p46_array_index_1085173;
  reg [7:0] p46_array_index_1085174;
  reg [7:0] p46_array_index_1085175;
  reg [7:0] p46_array_index_1085176;
  reg [7:0] p46_array_index_1085178;
  reg [7:0] p46_array_index_1085180;
  reg [7:0] p46_array_index_1085181;
  reg [7:0] p46_array_index_1085187;
  reg [7:0] p46_array_index_1085188;
  reg [7:0] p46_array_index_1085189;
  reg [7:0] p46_array_index_1085190;
  reg [7:0] p46_array_index_1085191;
  reg [7:0] p46_array_index_1085193;
  reg [7:0] p46_array_index_1085195;
  reg [7:0] p46_res7__240;
  reg [7:0] p46_array_index_1085204;
  reg [7:0] p46_array_index_1085205;
  reg [7:0] p46_array_index_1085206;
  reg [7:0] p46_array_index_1085207;
  reg [7:0] p46_array_index_1085208;
  reg [7:0] p46_array_index_1085209;
  reg [7:0] p46_res7__241;
  reg [7:0] p46_array_index_1085219;
  reg [7:0] p46_array_index_1085220;
  reg [7:0] p46_array_index_1085221;
  reg [7:0] p46_array_index_1085222;
  reg [7:0] p46_array_index_1085223;
  reg [7:0] p46_res7__242;
  reg [7:0] p46_array_index_1085233;
  reg [7:0] p46_array_index_1085234;
  reg [7:0] p46_array_index_1085235;
  reg [7:0] p46_array_index_1085236;
  reg [7:0] p46_array_index_1085237;
  reg [7:0] p46_res7__243;
  reg [7:0] p46_array_index_1085248;
  reg [7:0] p46_array_index_1085249;
  reg [7:0] p46_array_index_1085250;
  reg [7:0] p46_array_index_1085251;
  reg [7:0] p46_res7__244;
  reg [127:0] p46_res__35;
  reg [7:0] p47_arr[256];
  reg [7:0] p47_literal_1076345[256];
  reg [7:0] p47_literal_1076347[256];
  reg [7:0] p47_literal_1076349[256];
  reg [7:0] p47_literal_1076351[256];
  reg [7:0] p47_literal_1076353[256];
  reg [7:0] p47_literal_1076355[256];
  reg [7:0] p47_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p46_xor_1084661 <= p45_xor_1084661;
    p46_k5 <= p45_k5;
    p46_array_index_1085171 <= p46_array_index_1085171_comb;
    p46_array_index_1085172 <= p46_array_index_1085172_comb;
    p46_array_index_1085173 <= p46_array_index_1085173_comb;
    p46_array_index_1085174 <= p46_array_index_1085174_comb;
    p46_array_index_1085175 <= p46_array_index_1085175_comb;
    p46_array_index_1085176 <= p46_array_index_1085176_comb;
    p46_array_index_1085178 <= p46_array_index_1085178_comb;
    p46_array_index_1085180 <= p46_array_index_1085180_comb;
    p46_array_index_1085181 <= p46_array_index_1085181_comb;
    p46_array_index_1085187 <= p46_array_index_1085187_comb;
    p46_array_index_1085188 <= p46_array_index_1085188_comb;
    p46_array_index_1085189 <= p46_array_index_1085189_comb;
    p46_array_index_1085190 <= p46_array_index_1085190_comb;
    p46_array_index_1085191 <= p46_array_index_1085191_comb;
    p46_array_index_1085193 <= p46_array_index_1085193_comb;
    p46_array_index_1085195 <= p46_array_index_1085195_comb;
    p46_res7__240 <= p46_res7__240_comb;
    p46_array_index_1085204 <= p46_array_index_1085204_comb;
    p46_array_index_1085205 <= p46_array_index_1085205_comb;
    p46_array_index_1085206 <= p46_array_index_1085206_comb;
    p46_array_index_1085207 <= p46_array_index_1085207_comb;
    p46_array_index_1085208 <= p46_array_index_1085208_comb;
    p46_array_index_1085209 <= p46_array_index_1085209_comb;
    p46_res7__241 <= p46_res7__241_comb;
    p46_array_index_1085219 <= p46_array_index_1085219_comb;
    p46_array_index_1085220 <= p46_array_index_1085220_comb;
    p46_array_index_1085221 <= p46_array_index_1085221_comb;
    p46_array_index_1085222 <= p46_array_index_1085222_comb;
    p46_array_index_1085223 <= p46_array_index_1085223_comb;
    p46_res7__242 <= p46_res7__242_comb;
    p46_array_index_1085233 <= p46_array_index_1085233_comb;
    p46_array_index_1085234 <= p46_array_index_1085234_comb;
    p46_array_index_1085235 <= p46_array_index_1085235_comb;
    p46_array_index_1085236 <= p46_array_index_1085236_comb;
    p46_array_index_1085237 <= p46_array_index_1085237_comb;
    p46_res7__243 <= p46_res7__243_comb;
    p46_array_index_1085248 <= p46_array_index_1085248_comb;
    p46_array_index_1085249 <= p46_array_index_1085249_comb;
    p46_array_index_1085250 <= p46_array_index_1085250_comb;
    p46_array_index_1085251 <= p46_array_index_1085251_comb;
    p46_res7__244 <= p46_res7__244_comb;
    p46_res__35 <= p45_res__35;
    p47_arr <= p46_arr;
    p47_literal_1076345 <= p46_literal_1076345;
    p47_literal_1076347 <= p46_literal_1076347;
    p47_literal_1076349 <= p46_literal_1076349;
    p47_literal_1076351 <= p46_literal_1076351;
    p47_literal_1076353 <= p46_literal_1076353;
    p47_literal_1076355 <= p46_literal_1076355;
    p47_literal_1076358 <= p46_literal_1076358;
  end

  // ===== Pipe stage 47:
  wire [7:0] p47_array_index_1085365_comb;
  wire [7:0] p47_array_index_1085366_comb;
  wire [7:0] p47_array_index_1085367_comb;
  wire [7:0] p47_array_index_1085368_comb;
  wire [7:0] p47_res7__245_comb;
  wire [7:0] p47_array_index_1085379_comb;
  wire [7:0] p47_array_index_1085380_comb;
  wire [7:0] p47_array_index_1085381_comb;
  wire [7:0] p47_res7__246_comb;
  wire [7:0] p47_array_index_1085391_comb;
  wire [7:0] p47_array_index_1085392_comb;
  wire [7:0] p47_array_index_1085393_comb;
  wire [7:0] p47_res7__247_comb;
  wire [7:0] p47_array_index_1085404_comb;
  wire [7:0] p47_array_index_1085405_comb;
  wire [7:0] p47_res7__248_comb;
  wire [7:0] p47_array_index_1085415_comb;
  wire [7:0] p47_array_index_1085416_comb;
  wire [7:0] p47_res7__249_comb;
  wire [7:0] p47_array_index_1085422_comb;
  wire [7:0] p47_array_index_1085423_comb;
  wire [7:0] p47_array_index_1085424_comb;
  wire [7:0] p47_array_index_1085425_comb;
  wire [7:0] p47_array_index_1085426_comb;
  wire [7:0] p47_array_index_1085427_comb;
  wire [7:0] p47_array_index_1085428_comb;
  wire [7:0] p47_array_index_1085429_comb;
  wire [7:0] p47_array_index_1085430_comb;
  assign p47_array_index_1085365_comb = p46_literal_1076349[p46_res7__242];
  assign p47_array_index_1085366_comb = p46_literal_1076351[p46_res7__241];
  assign p47_array_index_1085367_comb = p46_literal_1076353[p46_res7__240];
  assign p47_array_index_1085368_comb = p46_literal_1076355[p46_array_index_1085171];
  assign p47_res7__245_comb = p46_literal_1076345[p46_res7__244] ^ p46_literal_1076347[p46_res7__243] ^ p47_array_index_1085365_comb ^ p47_array_index_1085366_comb ^ p47_array_index_1085367_comb ^ p47_array_index_1085368_comb ^ p46_array_index_1085172 ^ p46_literal_1076358[p46_array_index_1085173] ^ p46_array_index_1085174 ^ p46_array_index_1085209 ^ p46_literal_1076353[p46_array_index_1085176] ^ p46_literal_1076351[p46_array_index_1085193] ^ p46_literal_1076349[p46_array_index_1085178] ^ p46_literal_1076347[p46_array_index_1085195] ^ p46_literal_1076345[p46_array_index_1085180] ^ p46_array_index_1085181;
  assign p47_array_index_1085379_comb = p46_literal_1076351[p46_res7__242];
  assign p47_array_index_1085380_comb = p46_literal_1076353[p46_res7__241];
  assign p47_array_index_1085381_comb = p46_literal_1076355[p46_res7__240];
  assign p47_res7__246_comb = p46_literal_1076345[p47_res7__245_comb] ^ p46_literal_1076347[p46_res7__244] ^ p46_literal_1076349[p46_res7__243] ^ p47_array_index_1085379_comb ^ p47_array_index_1085380_comb ^ p47_array_index_1085381_comb ^ p46_array_index_1085171 ^ p46_literal_1076358[p46_array_index_1085172] ^ p46_array_index_1085173 ^ p46_array_index_1085223 ^ p46_array_index_1085191 ^ p46_literal_1076351[p46_array_index_1085176] ^ p46_literal_1076349[p46_array_index_1085193] ^ p46_literal_1076347[p46_array_index_1085178] ^ p46_literal_1076345[p46_array_index_1085195] ^ p46_array_index_1085180;
  assign p47_array_index_1085391_comb = p46_literal_1076351[p46_res7__243];
  assign p47_array_index_1085392_comb = p46_literal_1076353[p46_res7__242];
  assign p47_array_index_1085393_comb = p46_literal_1076355[p46_res7__241];
  assign p47_res7__247_comb = p46_literal_1076345[p47_res7__246_comb] ^ p46_literal_1076347[p47_res7__245_comb] ^ p46_literal_1076349[p46_res7__244] ^ p47_array_index_1085391_comb ^ p47_array_index_1085392_comb ^ p47_array_index_1085393_comb ^ p46_res7__240 ^ p46_literal_1076358[p46_array_index_1085171] ^ p46_array_index_1085172 ^ p46_array_index_1085237 ^ p46_array_index_1085208 ^ p46_literal_1076351[p46_array_index_1085175] ^ p46_literal_1076349[p46_array_index_1085176] ^ p46_literal_1076347[p46_array_index_1085193] ^ p46_literal_1076345[p46_array_index_1085178] ^ p46_array_index_1085195;
  assign p47_array_index_1085404_comb = p46_literal_1076353[p46_res7__243];
  assign p47_array_index_1085405_comb = p46_literal_1076355[p46_res7__242];
  assign p47_res7__248_comb = p46_literal_1076345[p47_res7__247_comb] ^ p46_literal_1076347[p47_res7__246_comb] ^ p46_literal_1076349[p47_res7__245_comb] ^ p46_literal_1076351[p46_res7__244] ^ p47_array_index_1085404_comb ^ p47_array_index_1085405_comb ^ p46_res7__241 ^ p46_literal_1076358[p46_res7__240] ^ p46_array_index_1085171 ^ p46_array_index_1085251 ^ p46_array_index_1085222 ^ p46_array_index_1085190 ^ p46_literal_1076349[p46_array_index_1085175] ^ p46_literal_1076347[p46_array_index_1085176] ^ p46_literal_1076345[p46_array_index_1085193] ^ p46_array_index_1085178;
  assign p47_array_index_1085415_comb = p46_literal_1076353[p46_res7__244];
  assign p47_array_index_1085416_comb = p46_literal_1076355[p46_res7__243];
  assign p47_res7__249_comb = p46_literal_1076345[p47_res7__248_comb] ^ p46_literal_1076347[p47_res7__247_comb] ^ p46_literal_1076349[p47_res7__246_comb] ^ p46_literal_1076351[p47_res7__245_comb] ^ p47_array_index_1085415_comb ^ p47_array_index_1085416_comb ^ p46_res7__242 ^ p46_literal_1076358[p46_res7__241] ^ p46_res7__240 ^ p47_array_index_1085368_comb ^ p46_array_index_1085236 ^ p46_array_index_1085207 ^ p46_literal_1076349[p46_array_index_1085174] ^ p46_literal_1076347[p46_array_index_1085175] ^ p46_literal_1076345[p46_array_index_1085176] ^ p46_array_index_1085193;
  assign p47_array_index_1085422_comb = p46_literal_1076345[p47_res7__249_comb];
  assign p47_array_index_1085423_comb = p46_literal_1076347[p47_res7__248_comb];
  assign p47_array_index_1085424_comb = p46_literal_1076349[p47_res7__247_comb];
  assign p47_array_index_1085425_comb = p46_literal_1076351[p47_res7__246_comb];
  assign p47_array_index_1085426_comb = p46_literal_1076353[p47_res7__245_comb];
  assign p47_array_index_1085427_comb = p46_literal_1076355[p46_res7__244];
  assign p47_array_index_1085428_comb = p46_literal_1076358[p46_res7__242];
  assign p47_array_index_1085429_comb = p46_literal_1076347[p46_array_index_1085174];
  assign p47_array_index_1085430_comb = p46_literal_1076345[p46_array_index_1085175];

  // Registers for pipe stage 47:
  reg [127:0] p47_xor_1084661;
  reg [127:0] p47_k5;
  reg [7:0] p47_array_index_1085171;
  reg [7:0] p47_array_index_1085172;
  reg [7:0] p47_array_index_1085173;
  reg [7:0] p47_array_index_1085174;
  reg [7:0] p47_array_index_1085175;
  reg [7:0] p47_array_index_1085176;
  reg [7:0] p47_array_index_1085187;
  reg [7:0] p47_array_index_1085188;
  reg [7:0] p47_array_index_1085189;
  reg [7:0] p47_res7__240;
  reg [7:0] p47_array_index_1085204;
  reg [7:0] p47_array_index_1085205;
  reg [7:0] p47_array_index_1085206;
  reg [7:0] p47_res7__241;
  reg [7:0] p47_array_index_1085219;
  reg [7:0] p47_array_index_1085220;
  reg [7:0] p47_array_index_1085221;
  reg [7:0] p47_res7__242;
  reg [7:0] p47_array_index_1085233;
  reg [7:0] p47_array_index_1085234;
  reg [7:0] p47_array_index_1085235;
  reg [7:0] p47_res7__243;
  reg [7:0] p47_array_index_1085248;
  reg [7:0] p47_array_index_1085249;
  reg [7:0] p47_array_index_1085250;
  reg [7:0] p47_res7__244;
  reg [7:0] p47_array_index_1085365;
  reg [7:0] p47_array_index_1085366;
  reg [7:0] p47_array_index_1085367;
  reg [7:0] p47_res7__245;
  reg [7:0] p47_array_index_1085379;
  reg [7:0] p47_array_index_1085380;
  reg [7:0] p47_array_index_1085381;
  reg [7:0] p47_res7__246;
  reg [7:0] p47_array_index_1085391;
  reg [7:0] p47_array_index_1085392;
  reg [7:0] p47_array_index_1085393;
  reg [7:0] p47_res7__247;
  reg [7:0] p47_array_index_1085404;
  reg [7:0] p47_array_index_1085405;
  reg [7:0] p47_res7__248;
  reg [7:0] p47_array_index_1085415;
  reg [7:0] p47_array_index_1085416;
  reg [7:0] p47_res7__249;
  reg [7:0] p47_array_index_1085422;
  reg [7:0] p47_array_index_1085423;
  reg [7:0] p47_array_index_1085424;
  reg [7:0] p47_array_index_1085425;
  reg [7:0] p47_array_index_1085426;
  reg [7:0] p47_array_index_1085427;
  reg [7:0] p47_array_index_1085428;
  reg [7:0] p47_array_index_1085429;
  reg [7:0] p47_array_index_1085430;
  reg [127:0] p47_res__35;
  reg [7:0] p48_arr[256];
  reg [7:0] p48_literal_1076345[256];
  reg [7:0] p48_literal_1076347[256];
  reg [7:0] p48_literal_1076349[256];
  reg [7:0] p48_literal_1076351[256];
  reg [7:0] p48_literal_1076353[256];
  reg [7:0] p48_literal_1076355[256];
  reg [7:0] p48_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p47_xor_1084661 <= p46_xor_1084661;
    p47_k5 <= p46_k5;
    p47_array_index_1085171 <= p46_array_index_1085171;
    p47_array_index_1085172 <= p46_array_index_1085172;
    p47_array_index_1085173 <= p46_array_index_1085173;
    p47_array_index_1085174 <= p46_array_index_1085174;
    p47_array_index_1085175 <= p46_array_index_1085175;
    p47_array_index_1085176 <= p46_array_index_1085176;
    p47_array_index_1085187 <= p46_array_index_1085187;
    p47_array_index_1085188 <= p46_array_index_1085188;
    p47_array_index_1085189 <= p46_array_index_1085189;
    p47_res7__240 <= p46_res7__240;
    p47_array_index_1085204 <= p46_array_index_1085204;
    p47_array_index_1085205 <= p46_array_index_1085205;
    p47_array_index_1085206 <= p46_array_index_1085206;
    p47_res7__241 <= p46_res7__241;
    p47_array_index_1085219 <= p46_array_index_1085219;
    p47_array_index_1085220 <= p46_array_index_1085220;
    p47_array_index_1085221 <= p46_array_index_1085221;
    p47_res7__242 <= p46_res7__242;
    p47_array_index_1085233 <= p46_array_index_1085233;
    p47_array_index_1085234 <= p46_array_index_1085234;
    p47_array_index_1085235 <= p46_array_index_1085235;
    p47_res7__243 <= p46_res7__243;
    p47_array_index_1085248 <= p46_array_index_1085248;
    p47_array_index_1085249 <= p46_array_index_1085249;
    p47_array_index_1085250 <= p46_array_index_1085250;
    p47_res7__244 <= p46_res7__244;
    p47_array_index_1085365 <= p47_array_index_1085365_comb;
    p47_array_index_1085366 <= p47_array_index_1085366_comb;
    p47_array_index_1085367 <= p47_array_index_1085367_comb;
    p47_res7__245 <= p47_res7__245_comb;
    p47_array_index_1085379 <= p47_array_index_1085379_comb;
    p47_array_index_1085380 <= p47_array_index_1085380_comb;
    p47_array_index_1085381 <= p47_array_index_1085381_comb;
    p47_res7__246 <= p47_res7__246_comb;
    p47_array_index_1085391 <= p47_array_index_1085391_comb;
    p47_array_index_1085392 <= p47_array_index_1085392_comb;
    p47_array_index_1085393 <= p47_array_index_1085393_comb;
    p47_res7__247 <= p47_res7__247_comb;
    p47_array_index_1085404 <= p47_array_index_1085404_comb;
    p47_array_index_1085405 <= p47_array_index_1085405_comb;
    p47_res7__248 <= p47_res7__248_comb;
    p47_array_index_1085415 <= p47_array_index_1085415_comb;
    p47_array_index_1085416 <= p47_array_index_1085416_comb;
    p47_res7__249 <= p47_res7__249_comb;
    p47_array_index_1085422 <= p47_array_index_1085422_comb;
    p47_array_index_1085423 <= p47_array_index_1085423_comb;
    p47_array_index_1085424 <= p47_array_index_1085424_comb;
    p47_array_index_1085425 <= p47_array_index_1085425_comb;
    p47_array_index_1085426 <= p47_array_index_1085426_comb;
    p47_array_index_1085427 <= p47_array_index_1085427_comb;
    p47_array_index_1085428 <= p47_array_index_1085428_comb;
    p47_array_index_1085429 <= p47_array_index_1085429_comb;
    p47_array_index_1085430 <= p47_array_index_1085430_comb;
    p47_res__35 <= p46_res__35;
    p48_arr <= p47_arr;
    p48_literal_1076345 <= p47_literal_1076345;
    p48_literal_1076347 <= p47_literal_1076347;
    p48_literal_1076349 <= p47_literal_1076349;
    p48_literal_1076351 <= p47_literal_1076351;
    p48_literal_1076353 <= p47_literal_1076353;
    p48_literal_1076355 <= p47_literal_1076355;
    p48_literal_1076358 <= p47_literal_1076358;
  end

  // ===== Pipe stage 48:
  wire [7:0] p48_res7__250_comb;
  wire [7:0] p48_array_index_1085565_comb;
  wire [7:0] p48_res7__251_comb;
  wire [7:0] p48_res7__252_comb;
  wire [7:0] p48_res7__253_comb;
  wire [7:0] p48_res7__254_comb;
  wire [7:0] p48_res7__255_comb;
  wire [127:0] p48_res__15_comb;
  wire [127:0] p48_k4_comb;
  wire [127:0] p48_addedKey__36_comb;
  wire [7:0] p48_bit_slice_1085607_comb;
  wire [7:0] p48_bit_slice_1085608_comb;
  wire [7:0] p48_bit_slice_1085609_comb;
  wire [7:0] p48_bit_slice_1085610_comb;
  wire [7:0] p48_bit_slice_1085611_comb;
  wire [7:0] p48_bit_slice_1085612_comb;
  wire [7:0] p48_bit_slice_1085613_comb;
  wire [7:0] p48_bit_slice_1085614_comb;
  wire [7:0] p48_bit_slice_1085615_comb;
  wire [7:0] p48_bit_slice_1085616_comb;
  wire [7:0] p48_bit_slice_1085617_comb;
  wire [7:0] p48_bit_slice_1085618_comb;
  wire [7:0] p48_bit_slice_1085619_comb;
  wire [7:0] p48_bit_slice_1085620_comb;
  wire [7:0] p48_bit_slice_1085621_comb;
  wire [7:0] p48_bit_slice_1085622_comb;
  assign p48_res7__250_comb = p47_array_index_1085422 ^ p47_array_index_1085423 ^ p47_array_index_1085424 ^ p47_array_index_1085425 ^ p47_array_index_1085426 ^ p47_array_index_1085427 ^ p47_res7__243 ^ p47_array_index_1085428 ^ p47_res7__241 ^ p47_array_index_1085381 ^ p47_array_index_1085250 ^ p47_array_index_1085221 ^ p47_array_index_1085189 ^ p47_array_index_1085429 ^ p47_array_index_1085430 ^ p47_array_index_1085176;
  assign p48_array_index_1085565_comb = p47_literal_1076355[p47_res7__245];
  assign p48_res7__251_comb = p47_literal_1076345[p48_res7__250_comb] ^ p47_literal_1076347[p47_res7__249] ^ p47_literal_1076349[p47_res7__248] ^ p47_literal_1076351[p47_res7__247] ^ p47_literal_1076353[p47_res7__246] ^ p48_array_index_1085565_comb ^ p47_res7__244 ^ p47_literal_1076358[p47_res7__243] ^ p47_res7__242 ^ p47_array_index_1085393 ^ p47_array_index_1085367 ^ p47_array_index_1085235 ^ p47_array_index_1085206 ^ p47_literal_1076347[p47_array_index_1085173] ^ p47_literal_1076345[p47_array_index_1085174] ^ p47_array_index_1085175;
  assign p48_res7__252_comb = p47_literal_1076345[p48_res7__251_comb] ^ p47_literal_1076347[p48_res7__250_comb] ^ p47_literal_1076349[p47_res7__249] ^ p47_literal_1076351[p47_res7__248] ^ p47_literal_1076353[p47_res7__247] ^ p47_literal_1076355[p47_res7__246] ^ p47_res7__245 ^ p47_literal_1076358[p47_res7__244] ^ p47_res7__243 ^ p47_array_index_1085405 ^ p47_array_index_1085380 ^ p47_array_index_1085249 ^ p47_array_index_1085220 ^ p47_array_index_1085188 ^ p47_literal_1076345[p47_array_index_1085173] ^ p47_array_index_1085174;
  assign p48_res7__253_comb = p47_literal_1076345[p48_res7__252_comb] ^ p47_literal_1076347[p48_res7__251_comb] ^ p47_literal_1076349[p48_res7__250_comb] ^ p47_literal_1076351[p47_res7__249] ^ p47_literal_1076353[p47_res7__248] ^ p47_literal_1076355[p47_res7__247] ^ p47_res7__246 ^ p47_literal_1076358[p47_res7__245] ^ p47_res7__244 ^ p47_array_index_1085416 ^ p47_array_index_1085392 ^ p47_array_index_1085366 ^ p47_array_index_1085234 ^ p47_array_index_1085205 ^ p47_literal_1076345[p47_array_index_1085172] ^ p47_array_index_1085173;
  assign p48_res7__254_comb = p47_literal_1076345[p48_res7__253_comb] ^ p47_literal_1076347[p48_res7__252_comb] ^ p47_literal_1076349[p48_res7__251_comb] ^ p47_literal_1076351[p48_res7__250_comb] ^ p47_literal_1076353[p47_res7__249] ^ p47_literal_1076355[p47_res7__248] ^ p47_res7__247 ^ p47_literal_1076358[p47_res7__246] ^ p47_res7__245 ^ p47_array_index_1085427 ^ p47_array_index_1085404 ^ p47_array_index_1085379 ^ p47_array_index_1085248 ^ p47_array_index_1085219 ^ p47_array_index_1085187 ^ p47_array_index_1085172;
  assign p48_res7__255_comb = p47_literal_1076345[p48_res7__254_comb] ^ p47_literal_1076347[p48_res7__253_comb] ^ p47_literal_1076349[p48_res7__252_comb] ^ p47_literal_1076351[p48_res7__251_comb] ^ p47_literal_1076353[p48_res7__250_comb] ^ p47_literal_1076355[p47_res7__249] ^ p47_res7__248 ^ p47_literal_1076358[p47_res7__247] ^ p47_res7__246 ^ p48_array_index_1085565_comb ^ p47_array_index_1085415 ^ p47_array_index_1085391 ^ p47_array_index_1085365 ^ p47_array_index_1085233 ^ p47_array_index_1085204 ^ p47_array_index_1085171;
  assign p48_res__15_comb = {p48_res7__255_comb, p48_res7__254_comb, p48_res7__253_comb, p48_res7__252_comb, p48_res7__251_comb, p48_res7__250_comb, p47_res7__249, p47_res7__248, p47_res7__247, p47_res7__246, p47_res7__245, p47_res7__244, p47_res7__243, p47_res7__242, p47_res7__241, p47_res7__240};
  assign p48_k4_comb = p48_res__15_comb ^ p47_xor_1084661;
  assign p48_addedKey__36_comb = p48_k4_comb ^ p47_res__35;
  assign p48_bit_slice_1085607_comb = p48_addedKey__36_comb[127:120];
  assign p48_bit_slice_1085608_comb = p48_addedKey__36_comb[119:112];
  assign p48_bit_slice_1085609_comb = p48_addedKey__36_comb[111:104];
  assign p48_bit_slice_1085610_comb = p48_addedKey__36_comb[103:96];
  assign p48_bit_slice_1085611_comb = p48_addedKey__36_comb[95:88];
  assign p48_bit_slice_1085612_comb = p48_addedKey__36_comb[87:80];
  assign p48_bit_slice_1085613_comb = p48_addedKey__36_comb[71:64];
  assign p48_bit_slice_1085614_comb = p48_addedKey__36_comb[55:48];
  assign p48_bit_slice_1085615_comb = p48_addedKey__36_comb[47:40];
  assign p48_bit_slice_1085616_comb = p48_addedKey__36_comb[39:32];
  assign p48_bit_slice_1085617_comb = p48_addedKey__36_comb[31:24];
  assign p48_bit_slice_1085618_comb = p48_addedKey__36_comb[23:16];
  assign p48_bit_slice_1085619_comb = p48_addedKey__36_comb[15:8];
  assign p48_bit_slice_1085620_comb = p48_addedKey__36_comb[79:72];
  assign p48_bit_slice_1085621_comb = p48_addedKey__36_comb[63:56];
  assign p48_bit_slice_1085622_comb = p48_addedKey__36_comb[7:0];

  // Registers for pipe stage 48:
  reg [127:0] p48_k5;
  reg [127:0] p48_k4;
  reg [7:0] p48_bit_slice_1085607;
  reg [7:0] p48_bit_slice_1085608;
  reg [7:0] p48_bit_slice_1085609;
  reg [7:0] p48_bit_slice_1085610;
  reg [7:0] p48_bit_slice_1085611;
  reg [7:0] p48_bit_slice_1085612;
  reg [7:0] p48_bit_slice_1085613;
  reg [7:0] p48_bit_slice_1085614;
  reg [7:0] p48_bit_slice_1085615;
  reg [7:0] p48_bit_slice_1085616;
  reg [7:0] p48_bit_slice_1085617;
  reg [7:0] p48_bit_slice_1085618;
  reg [7:0] p48_bit_slice_1085619;
  reg [7:0] p48_bit_slice_1085620;
  reg [7:0] p48_bit_slice_1085621;
  reg [7:0] p48_bit_slice_1085622;
  reg [7:0] p49_arr[256];
  reg [7:0] p49_literal_1076345[256];
  reg [7:0] p49_literal_1076347[256];
  reg [7:0] p49_literal_1076349[256];
  reg [7:0] p49_literal_1076351[256];
  reg [7:0] p49_literal_1076353[256];
  reg [7:0] p49_literal_1076355[256];
  reg [7:0] p49_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p48_k5 <= p47_k5;
    p48_k4 <= p48_k4_comb;
    p48_bit_slice_1085607 <= p48_bit_slice_1085607_comb;
    p48_bit_slice_1085608 <= p48_bit_slice_1085608_comb;
    p48_bit_slice_1085609 <= p48_bit_slice_1085609_comb;
    p48_bit_slice_1085610 <= p48_bit_slice_1085610_comb;
    p48_bit_slice_1085611 <= p48_bit_slice_1085611_comb;
    p48_bit_slice_1085612 <= p48_bit_slice_1085612_comb;
    p48_bit_slice_1085613 <= p48_bit_slice_1085613_comb;
    p48_bit_slice_1085614 <= p48_bit_slice_1085614_comb;
    p48_bit_slice_1085615 <= p48_bit_slice_1085615_comb;
    p48_bit_slice_1085616 <= p48_bit_slice_1085616_comb;
    p48_bit_slice_1085617 <= p48_bit_slice_1085617_comb;
    p48_bit_slice_1085618 <= p48_bit_slice_1085618_comb;
    p48_bit_slice_1085619 <= p48_bit_slice_1085619_comb;
    p48_bit_slice_1085620 <= p48_bit_slice_1085620_comb;
    p48_bit_slice_1085621 <= p48_bit_slice_1085621_comb;
    p48_bit_slice_1085622 <= p48_bit_slice_1085622_comb;
    p49_arr <= p48_arr;
    p49_literal_1076345 <= p48_literal_1076345;
    p49_literal_1076347 <= p48_literal_1076347;
    p49_literal_1076349 <= p48_literal_1076349;
    p49_literal_1076351 <= p48_literal_1076351;
    p49_literal_1076353 <= p48_literal_1076353;
    p49_literal_1076355 <= p48_literal_1076355;
    p49_literal_1076358 <= p48_literal_1076358;
  end

  // ===== Pipe stage 49:
  wire [127:0] p49_addedKey__57_comb;
  wire [7:0] p49_array_index_1085690_comb;
  wire [7:0] p49_array_index_1085691_comb;
  wire [7:0] p49_array_index_1085692_comb;
  wire [7:0] p49_array_index_1085693_comb;
  wire [7:0] p49_array_index_1085694_comb;
  wire [7:0] p49_array_index_1085695_comb;
  wire [7:0] p49_array_index_1085697_comb;
  wire [7:0] p49_array_index_1085699_comb;
  wire [7:0] p49_array_index_1085700_comb;
  wire [7:0] p49_array_index_1085701_comb;
  wire [7:0] p49_array_index_1085702_comb;
  wire [7:0] p49_array_index_1085703_comb;
  wire [7:0] p49_array_index_1085704_comb;
  wire [7:0] p49_array_index_1085778_comb;
  wire [7:0] p49_array_index_1085779_comb;
  wire [7:0] p49_array_index_1085780_comb;
  wire [7:0] p49_array_index_1085781_comb;
  wire [7:0] p49_array_index_1085782_comb;
  wire [7:0] p49_array_index_1085783_comb;
  wire [7:0] p49_array_index_1085784_comb;
  wire [7:0] p49_array_index_1085785_comb;
  wire [7:0] p49_array_index_1085786_comb;
  wire [7:0] p49_array_index_1085787_comb;
  wire [7:0] p49_array_index_1085788_comb;
  wire [7:0] p49_array_index_1085789_comb;
  wire [7:0] p49_array_index_1085790_comb;
  wire [7:0] p49_array_index_1085706_comb;
  wire [7:0] p49_array_index_1085707_comb;
  wire [7:0] p49_array_index_1085708_comb;
  wire [7:0] p49_array_index_1085709_comb;
  wire [7:0] p49_array_index_1085710_comb;
  wire [7:0] p49_array_index_1085711_comb;
  wire [7:0] p49_array_index_1085712_comb;
  wire [7:0] p49_array_index_1085714_comb;
  wire [7:0] p49_array_index_1085791_comb;
  wire [7:0] p49_array_index_1085792_comb;
  wire [7:0] p49_array_index_1085793_comb;
  wire [7:0] p49_array_index_1085794_comb;
  wire [7:0] p49_array_index_1085795_comb;
  wire [7:0] p49_array_index_1085796_comb;
  wire [7:0] p49_array_index_1085797_comb;
  wire [7:0] p49_array_index_1085799_comb;
  wire [7:0] p49_res7__256_comb;
  wire [7:0] p49_res7__576_comb;
  wire [7:0] p49_array_index_1085723_comb;
  wire [7:0] p49_array_index_1085724_comb;
  wire [7:0] p49_array_index_1085725_comb;
  wire [7:0] p49_array_index_1085726_comb;
  wire [7:0] p49_array_index_1085727_comb;
  wire [7:0] p49_array_index_1085728_comb;
  wire [7:0] p49_array_index_1085808_comb;
  wire [7:0] p49_array_index_1085809_comb;
  wire [7:0] p49_array_index_1085810_comb;
  wire [7:0] p49_array_index_1085811_comb;
  wire [7:0] p49_array_index_1085812_comb;
  wire [7:0] p49_array_index_1085813_comb;
  wire [7:0] p49_res7__257_comb;
  wire [7:0] p49_res7__577_comb;
  wire [7:0] p49_array_index_1085738_comb;
  wire [7:0] p49_array_index_1085739_comb;
  wire [7:0] p49_array_index_1085740_comb;
  wire [7:0] p49_array_index_1085741_comb;
  wire [7:0] p49_array_index_1085742_comb;
  wire [7:0] p49_array_index_1085823_comb;
  wire [7:0] p49_array_index_1085824_comb;
  wire [7:0] p49_array_index_1085825_comb;
  wire [7:0] p49_array_index_1085826_comb;
  wire [7:0] p49_array_index_1085827_comb;
  wire [7:0] p49_res7__258_comb;
  wire [7:0] p49_res7__578_comb;
  wire [7:0] p49_array_index_1085752_comb;
  wire [7:0] p49_array_index_1085753_comb;
  wire [7:0] p49_array_index_1085754_comb;
  wire [7:0] p49_array_index_1085755_comb;
  wire [7:0] p49_array_index_1085756_comb;
  wire [7:0] p49_array_index_1085837_comb;
  wire [7:0] p49_array_index_1085838_comb;
  wire [7:0] p49_array_index_1085839_comb;
  wire [7:0] p49_array_index_1085840_comb;
  wire [7:0] p49_array_index_1085841_comb;
  wire [7:0] p49_res7__259_comb;
  wire [7:0] p49_res7__579_comb;
  wire [7:0] p49_array_index_1085767_comb;
  wire [7:0] p49_array_index_1085768_comb;
  wire [7:0] p49_array_index_1085769_comb;
  wire [7:0] p49_array_index_1085770_comb;
  wire [7:0] p49_array_index_1085852_comb;
  wire [7:0] p49_array_index_1085853_comb;
  wire [7:0] p49_array_index_1085854_comb;
  wire [7:0] p49_array_index_1085855_comb;
  wire [7:0] p49_res7__260_comb;
  wire [7:0] p49_res7__580_comb;
  assign p49_addedKey__57_comb = p48_k4 ^ 128'h4110_1a5e_6342_d669_c412_3cd3_9313_c011;
  assign p49_array_index_1085690_comb = p48_arr[p49_addedKey__57_comb[127:120]];
  assign p49_array_index_1085691_comb = p48_arr[p49_addedKey__57_comb[119:112]];
  assign p49_array_index_1085692_comb = p48_arr[p49_addedKey__57_comb[111:104]];
  assign p49_array_index_1085693_comb = p48_arr[p49_addedKey__57_comb[103:96]];
  assign p49_array_index_1085694_comb = p48_arr[p49_addedKey__57_comb[95:88]];
  assign p49_array_index_1085695_comb = p48_arr[p49_addedKey__57_comb[87:80]];
  assign p49_array_index_1085697_comb = p48_arr[p49_addedKey__57_comb[71:64]];
  assign p49_array_index_1085699_comb = p48_arr[p49_addedKey__57_comb[55:48]];
  assign p49_array_index_1085700_comb = p48_arr[p49_addedKey__57_comb[47:40]];
  assign p49_array_index_1085701_comb = p48_arr[p49_addedKey__57_comb[39:32]];
  assign p49_array_index_1085702_comb = p48_arr[p49_addedKey__57_comb[31:24]];
  assign p49_array_index_1085703_comb = p48_arr[p49_addedKey__57_comb[23:16]];
  assign p49_array_index_1085704_comb = p48_arr[p49_addedKey__57_comb[15:8]];
  assign p49_array_index_1085778_comb = p48_arr[p48_bit_slice_1085607];
  assign p49_array_index_1085779_comb = p48_arr[p48_bit_slice_1085608];
  assign p49_array_index_1085780_comb = p48_arr[p48_bit_slice_1085609];
  assign p49_array_index_1085781_comb = p48_arr[p48_bit_slice_1085610];
  assign p49_array_index_1085782_comb = p48_arr[p48_bit_slice_1085611];
  assign p49_array_index_1085783_comb = p48_arr[p48_bit_slice_1085612];
  assign p49_array_index_1085784_comb = p48_arr[p48_bit_slice_1085613];
  assign p49_array_index_1085785_comb = p48_arr[p48_bit_slice_1085614];
  assign p49_array_index_1085786_comb = p48_arr[p48_bit_slice_1085615];
  assign p49_array_index_1085787_comb = p48_arr[p48_bit_slice_1085616];
  assign p49_array_index_1085788_comb = p48_arr[p48_bit_slice_1085617];
  assign p49_array_index_1085789_comb = p48_arr[p48_bit_slice_1085618];
  assign p49_array_index_1085790_comb = p48_arr[p48_bit_slice_1085619];
  assign p49_array_index_1085706_comb = p48_literal_1076345[p49_array_index_1085690_comb];
  assign p49_array_index_1085707_comb = p48_literal_1076347[p49_array_index_1085691_comb];
  assign p49_array_index_1085708_comb = p48_literal_1076349[p49_array_index_1085692_comb];
  assign p49_array_index_1085709_comb = p48_literal_1076351[p49_array_index_1085693_comb];
  assign p49_array_index_1085710_comb = p48_literal_1076353[p49_array_index_1085694_comb];
  assign p49_array_index_1085711_comb = p48_literal_1076355[p49_array_index_1085695_comb];
  assign p49_array_index_1085712_comb = p48_arr[p49_addedKey__57_comb[79:72]];
  assign p49_array_index_1085714_comb = p48_arr[p49_addedKey__57_comb[63:56]];
  assign p49_array_index_1085791_comb = p48_literal_1076345[p49_array_index_1085778_comb];
  assign p49_array_index_1085792_comb = p48_literal_1076347[p49_array_index_1085779_comb];
  assign p49_array_index_1085793_comb = p48_literal_1076349[p49_array_index_1085780_comb];
  assign p49_array_index_1085794_comb = p48_literal_1076351[p49_array_index_1085781_comb];
  assign p49_array_index_1085795_comb = p48_literal_1076353[p49_array_index_1085782_comb];
  assign p49_array_index_1085796_comb = p48_literal_1076355[p49_array_index_1085783_comb];
  assign p49_array_index_1085797_comb = p48_arr[p48_bit_slice_1085620];
  assign p49_array_index_1085799_comb = p48_arr[p48_bit_slice_1085621];
  assign p49_res7__256_comb = p49_array_index_1085706_comb ^ p49_array_index_1085707_comb ^ p49_array_index_1085708_comb ^ p49_array_index_1085709_comb ^ p49_array_index_1085710_comb ^ p49_array_index_1085711_comb ^ p49_array_index_1085712_comb ^ p48_literal_1076358[p49_array_index_1085697_comb] ^ p49_array_index_1085714_comb ^ p48_literal_1076355[p49_array_index_1085699_comb] ^ p48_literal_1076353[p49_array_index_1085700_comb] ^ p48_literal_1076351[p49_array_index_1085701_comb] ^ p48_literal_1076349[p49_array_index_1085702_comb] ^ p48_literal_1076347[p49_array_index_1085703_comb] ^ p48_literal_1076345[p49_array_index_1085704_comb] ^ p48_arr[p49_addedKey__57_comb[7:0]];
  assign p49_res7__576_comb = p49_array_index_1085791_comb ^ p49_array_index_1085792_comb ^ p49_array_index_1085793_comb ^ p49_array_index_1085794_comb ^ p49_array_index_1085795_comb ^ p49_array_index_1085796_comb ^ p49_array_index_1085797_comb ^ p48_literal_1076358[p49_array_index_1085784_comb] ^ p49_array_index_1085799_comb ^ p48_literal_1076355[p49_array_index_1085785_comb] ^ p48_literal_1076353[p49_array_index_1085786_comb] ^ p48_literal_1076351[p49_array_index_1085787_comb] ^ p48_literal_1076349[p49_array_index_1085788_comb] ^ p48_literal_1076347[p49_array_index_1085789_comb] ^ p48_literal_1076345[p49_array_index_1085790_comb] ^ p48_arr[p48_bit_slice_1085622];
  assign p49_array_index_1085723_comb = p48_literal_1076345[p49_res7__256_comb];
  assign p49_array_index_1085724_comb = p48_literal_1076347[p49_array_index_1085690_comb];
  assign p49_array_index_1085725_comb = p48_literal_1076349[p49_array_index_1085691_comb];
  assign p49_array_index_1085726_comb = p48_literal_1076351[p49_array_index_1085692_comb];
  assign p49_array_index_1085727_comb = p48_literal_1076353[p49_array_index_1085693_comb];
  assign p49_array_index_1085728_comb = p48_literal_1076355[p49_array_index_1085694_comb];
  assign p49_array_index_1085808_comb = p48_literal_1076345[p49_res7__576_comb];
  assign p49_array_index_1085809_comb = p48_literal_1076347[p49_array_index_1085778_comb];
  assign p49_array_index_1085810_comb = p48_literal_1076349[p49_array_index_1085779_comb];
  assign p49_array_index_1085811_comb = p48_literal_1076351[p49_array_index_1085780_comb];
  assign p49_array_index_1085812_comb = p48_literal_1076353[p49_array_index_1085781_comb];
  assign p49_array_index_1085813_comb = p48_literal_1076355[p49_array_index_1085782_comb];
  assign p49_res7__257_comb = p49_array_index_1085723_comb ^ p49_array_index_1085724_comb ^ p49_array_index_1085725_comb ^ p49_array_index_1085726_comb ^ p49_array_index_1085727_comb ^ p49_array_index_1085728_comb ^ p49_array_index_1085695_comb ^ p48_literal_1076358[p49_array_index_1085712_comb] ^ p49_array_index_1085697_comb ^ p48_literal_1076355[p49_array_index_1085714_comb] ^ p48_literal_1076353[p49_array_index_1085699_comb] ^ p48_literal_1076351[p49_array_index_1085700_comb] ^ p48_literal_1076349[p49_array_index_1085701_comb] ^ p48_literal_1076347[p49_array_index_1085702_comb] ^ p48_literal_1076345[p49_array_index_1085703_comb] ^ p49_array_index_1085704_comb;
  assign p49_res7__577_comb = p49_array_index_1085808_comb ^ p49_array_index_1085809_comb ^ p49_array_index_1085810_comb ^ p49_array_index_1085811_comb ^ p49_array_index_1085812_comb ^ p49_array_index_1085813_comb ^ p49_array_index_1085783_comb ^ p48_literal_1076358[p49_array_index_1085797_comb] ^ p49_array_index_1085784_comb ^ p48_literal_1076355[p49_array_index_1085799_comb] ^ p48_literal_1076353[p49_array_index_1085785_comb] ^ p48_literal_1076351[p49_array_index_1085786_comb] ^ p48_literal_1076349[p49_array_index_1085787_comb] ^ p48_literal_1076347[p49_array_index_1085788_comb] ^ p48_literal_1076345[p49_array_index_1085789_comb] ^ p49_array_index_1085790_comb;
  assign p49_array_index_1085738_comb = p48_literal_1076347[p49_res7__256_comb];
  assign p49_array_index_1085739_comb = p48_literal_1076349[p49_array_index_1085690_comb];
  assign p49_array_index_1085740_comb = p48_literal_1076351[p49_array_index_1085691_comb];
  assign p49_array_index_1085741_comb = p48_literal_1076353[p49_array_index_1085692_comb];
  assign p49_array_index_1085742_comb = p48_literal_1076355[p49_array_index_1085693_comb];
  assign p49_array_index_1085823_comb = p48_literal_1076347[p49_res7__576_comb];
  assign p49_array_index_1085824_comb = p48_literal_1076349[p49_array_index_1085778_comb];
  assign p49_array_index_1085825_comb = p48_literal_1076351[p49_array_index_1085779_comb];
  assign p49_array_index_1085826_comb = p48_literal_1076353[p49_array_index_1085780_comb];
  assign p49_array_index_1085827_comb = p48_literal_1076355[p49_array_index_1085781_comb];
  assign p49_res7__258_comb = p48_literal_1076345[p49_res7__257_comb] ^ p49_array_index_1085738_comb ^ p49_array_index_1085739_comb ^ p49_array_index_1085740_comb ^ p49_array_index_1085741_comb ^ p49_array_index_1085742_comb ^ p49_array_index_1085694_comb ^ p48_literal_1076358[p49_array_index_1085695_comb] ^ p49_array_index_1085712_comb ^ p48_literal_1076355[p49_array_index_1085697_comb] ^ p48_literal_1076353[p49_array_index_1085714_comb] ^ p48_literal_1076351[p49_array_index_1085699_comb] ^ p48_literal_1076349[p49_array_index_1085700_comb] ^ p48_literal_1076347[p49_array_index_1085701_comb] ^ p48_literal_1076345[p49_array_index_1085702_comb] ^ p49_array_index_1085703_comb;
  assign p49_res7__578_comb = p48_literal_1076345[p49_res7__577_comb] ^ p49_array_index_1085823_comb ^ p49_array_index_1085824_comb ^ p49_array_index_1085825_comb ^ p49_array_index_1085826_comb ^ p49_array_index_1085827_comb ^ p49_array_index_1085782_comb ^ p48_literal_1076358[p49_array_index_1085783_comb] ^ p49_array_index_1085797_comb ^ p48_literal_1076355[p49_array_index_1085784_comb] ^ p48_literal_1076353[p49_array_index_1085799_comb] ^ p48_literal_1076351[p49_array_index_1085785_comb] ^ p48_literal_1076349[p49_array_index_1085786_comb] ^ p48_literal_1076347[p49_array_index_1085787_comb] ^ p48_literal_1076345[p49_array_index_1085788_comb] ^ p49_array_index_1085789_comb;
  assign p49_array_index_1085752_comb = p48_literal_1076347[p49_res7__257_comb];
  assign p49_array_index_1085753_comb = p48_literal_1076349[p49_res7__256_comb];
  assign p49_array_index_1085754_comb = p48_literal_1076351[p49_array_index_1085690_comb];
  assign p49_array_index_1085755_comb = p48_literal_1076353[p49_array_index_1085691_comb];
  assign p49_array_index_1085756_comb = p48_literal_1076355[p49_array_index_1085692_comb];
  assign p49_array_index_1085837_comb = p48_literal_1076347[p49_res7__577_comb];
  assign p49_array_index_1085838_comb = p48_literal_1076349[p49_res7__576_comb];
  assign p49_array_index_1085839_comb = p48_literal_1076351[p49_array_index_1085778_comb];
  assign p49_array_index_1085840_comb = p48_literal_1076353[p49_array_index_1085779_comb];
  assign p49_array_index_1085841_comb = p48_literal_1076355[p49_array_index_1085780_comb];
  assign p49_res7__259_comb = p48_literal_1076345[p49_res7__258_comb] ^ p49_array_index_1085752_comb ^ p49_array_index_1085753_comb ^ p49_array_index_1085754_comb ^ p49_array_index_1085755_comb ^ p49_array_index_1085756_comb ^ p49_array_index_1085693_comb ^ p48_literal_1076358[p49_array_index_1085694_comb] ^ p49_array_index_1085695_comb ^ p48_literal_1076355[p49_array_index_1085712_comb] ^ p48_literal_1076353[p49_array_index_1085697_comb] ^ p48_literal_1076351[p49_array_index_1085714_comb] ^ p48_literal_1076349[p49_array_index_1085699_comb] ^ p48_literal_1076347[p49_array_index_1085700_comb] ^ p48_literal_1076345[p49_array_index_1085701_comb] ^ p49_array_index_1085702_comb;
  assign p49_res7__579_comb = p48_literal_1076345[p49_res7__578_comb] ^ p49_array_index_1085837_comb ^ p49_array_index_1085838_comb ^ p49_array_index_1085839_comb ^ p49_array_index_1085840_comb ^ p49_array_index_1085841_comb ^ p49_array_index_1085781_comb ^ p48_literal_1076358[p49_array_index_1085782_comb] ^ p49_array_index_1085783_comb ^ p48_literal_1076355[p49_array_index_1085797_comb] ^ p48_literal_1076353[p49_array_index_1085784_comb] ^ p48_literal_1076351[p49_array_index_1085799_comb] ^ p48_literal_1076349[p49_array_index_1085785_comb] ^ p48_literal_1076347[p49_array_index_1085786_comb] ^ p48_literal_1076345[p49_array_index_1085787_comb] ^ p49_array_index_1085788_comb;
  assign p49_array_index_1085767_comb = p48_literal_1076349[p49_res7__257_comb];
  assign p49_array_index_1085768_comb = p48_literal_1076351[p49_res7__256_comb];
  assign p49_array_index_1085769_comb = p48_literal_1076353[p49_array_index_1085690_comb];
  assign p49_array_index_1085770_comb = p48_literal_1076355[p49_array_index_1085691_comb];
  assign p49_array_index_1085852_comb = p48_literal_1076349[p49_res7__577_comb];
  assign p49_array_index_1085853_comb = p48_literal_1076351[p49_res7__576_comb];
  assign p49_array_index_1085854_comb = p48_literal_1076353[p49_array_index_1085778_comb];
  assign p49_array_index_1085855_comb = p48_literal_1076355[p49_array_index_1085779_comb];
  assign p49_res7__260_comb = p48_literal_1076345[p49_res7__259_comb] ^ p48_literal_1076347[p49_res7__258_comb] ^ p49_array_index_1085767_comb ^ p49_array_index_1085768_comb ^ p49_array_index_1085769_comb ^ p49_array_index_1085770_comb ^ p49_array_index_1085692_comb ^ p48_literal_1076358[p49_array_index_1085693_comb] ^ p49_array_index_1085694_comb ^ p49_array_index_1085711_comb ^ p48_literal_1076353[p49_array_index_1085712_comb] ^ p48_literal_1076351[p49_array_index_1085697_comb] ^ p48_literal_1076349[p49_array_index_1085714_comb] ^ p48_literal_1076347[p49_array_index_1085699_comb] ^ p48_literal_1076345[p49_array_index_1085700_comb] ^ p49_array_index_1085701_comb;
  assign p49_res7__580_comb = p48_literal_1076345[p49_res7__579_comb] ^ p48_literal_1076347[p49_res7__578_comb] ^ p49_array_index_1085852_comb ^ p49_array_index_1085853_comb ^ p49_array_index_1085854_comb ^ p49_array_index_1085855_comb ^ p49_array_index_1085780_comb ^ p48_literal_1076358[p49_array_index_1085781_comb] ^ p49_array_index_1085782_comb ^ p49_array_index_1085796_comb ^ p48_literal_1076353[p49_array_index_1085797_comb] ^ p48_literal_1076351[p49_array_index_1085784_comb] ^ p48_literal_1076349[p49_array_index_1085799_comb] ^ p48_literal_1076347[p49_array_index_1085785_comb] ^ p48_literal_1076345[p49_array_index_1085786_comb] ^ p49_array_index_1085787_comb;

  // Registers for pipe stage 49:
  reg [127:0] p49_k5;
  reg [127:0] p49_k4;
  reg [7:0] p49_array_index_1085690;
  reg [7:0] p49_array_index_1085691;
  reg [7:0] p49_array_index_1085692;
  reg [7:0] p49_array_index_1085693;
  reg [7:0] p49_array_index_1085694;
  reg [7:0] p49_array_index_1085695;
  reg [7:0] p49_array_index_1085697;
  reg [7:0] p49_array_index_1085699;
  reg [7:0] p49_array_index_1085700;
  reg [7:0] p49_array_index_1085706;
  reg [7:0] p49_array_index_1085707;
  reg [7:0] p49_array_index_1085708;
  reg [7:0] p49_array_index_1085709;
  reg [7:0] p49_array_index_1085710;
  reg [7:0] p49_array_index_1085712;
  reg [7:0] p49_array_index_1085714;
  reg [7:0] p49_res7__256;
  reg [7:0] p49_array_index_1085723;
  reg [7:0] p49_array_index_1085724;
  reg [7:0] p49_array_index_1085725;
  reg [7:0] p49_array_index_1085726;
  reg [7:0] p49_array_index_1085727;
  reg [7:0] p49_array_index_1085728;
  reg [7:0] p49_res7__257;
  reg [7:0] p49_array_index_1085738;
  reg [7:0] p49_array_index_1085739;
  reg [7:0] p49_array_index_1085740;
  reg [7:0] p49_array_index_1085741;
  reg [7:0] p49_array_index_1085742;
  reg [7:0] p49_res7__258;
  reg [7:0] p49_array_index_1085752;
  reg [7:0] p49_array_index_1085753;
  reg [7:0] p49_array_index_1085754;
  reg [7:0] p49_array_index_1085755;
  reg [7:0] p49_array_index_1085756;
  reg [7:0] p49_res7__259;
  reg [7:0] p49_array_index_1085767;
  reg [7:0] p49_array_index_1085768;
  reg [7:0] p49_array_index_1085769;
  reg [7:0] p49_array_index_1085770;
  reg [7:0] p49_res7__260;
  reg [7:0] p49_array_index_1085778;
  reg [7:0] p49_array_index_1085779;
  reg [7:0] p49_array_index_1085780;
  reg [7:0] p49_array_index_1085781;
  reg [7:0] p49_array_index_1085782;
  reg [7:0] p49_array_index_1085783;
  reg [7:0] p49_array_index_1085784;
  reg [7:0] p49_array_index_1085785;
  reg [7:0] p49_array_index_1085786;
  reg [7:0] p49_array_index_1085791;
  reg [7:0] p49_array_index_1085792;
  reg [7:0] p49_array_index_1085793;
  reg [7:0] p49_array_index_1085794;
  reg [7:0] p49_array_index_1085795;
  reg [7:0] p49_array_index_1085797;
  reg [7:0] p49_array_index_1085799;
  reg [7:0] p49_res7__576;
  reg [7:0] p49_array_index_1085808;
  reg [7:0] p49_array_index_1085809;
  reg [7:0] p49_array_index_1085810;
  reg [7:0] p49_array_index_1085811;
  reg [7:0] p49_array_index_1085812;
  reg [7:0] p49_array_index_1085813;
  reg [7:0] p49_res7__577;
  reg [7:0] p49_array_index_1085823;
  reg [7:0] p49_array_index_1085824;
  reg [7:0] p49_array_index_1085825;
  reg [7:0] p49_array_index_1085826;
  reg [7:0] p49_array_index_1085827;
  reg [7:0] p49_res7__578;
  reg [7:0] p49_array_index_1085837;
  reg [7:0] p49_array_index_1085838;
  reg [7:0] p49_array_index_1085839;
  reg [7:0] p49_array_index_1085840;
  reg [7:0] p49_array_index_1085841;
  reg [7:0] p49_res7__579;
  reg [7:0] p49_array_index_1085852;
  reg [7:0] p49_array_index_1085853;
  reg [7:0] p49_array_index_1085854;
  reg [7:0] p49_array_index_1085855;
  reg [7:0] p49_res7__580;
  reg [7:0] p50_arr[256];
  reg [7:0] p50_literal_1076345[256];
  reg [7:0] p50_literal_1076347[256];
  reg [7:0] p50_literal_1076349[256];
  reg [7:0] p50_literal_1076351[256];
  reg [7:0] p50_literal_1076353[256];
  reg [7:0] p50_literal_1076355[256];
  reg [7:0] p50_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p49_k5 <= p48_k5;
    p49_k4 <= p48_k4;
    p49_array_index_1085690 <= p49_array_index_1085690_comb;
    p49_array_index_1085691 <= p49_array_index_1085691_comb;
    p49_array_index_1085692 <= p49_array_index_1085692_comb;
    p49_array_index_1085693 <= p49_array_index_1085693_comb;
    p49_array_index_1085694 <= p49_array_index_1085694_comb;
    p49_array_index_1085695 <= p49_array_index_1085695_comb;
    p49_array_index_1085697 <= p49_array_index_1085697_comb;
    p49_array_index_1085699 <= p49_array_index_1085699_comb;
    p49_array_index_1085700 <= p49_array_index_1085700_comb;
    p49_array_index_1085706 <= p49_array_index_1085706_comb;
    p49_array_index_1085707 <= p49_array_index_1085707_comb;
    p49_array_index_1085708 <= p49_array_index_1085708_comb;
    p49_array_index_1085709 <= p49_array_index_1085709_comb;
    p49_array_index_1085710 <= p49_array_index_1085710_comb;
    p49_array_index_1085712 <= p49_array_index_1085712_comb;
    p49_array_index_1085714 <= p49_array_index_1085714_comb;
    p49_res7__256 <= p49_res7__256_comb;
    p49_array_index_1085723 <= p49_array_index_1085723_comb;
    p49_array_index_1085724 <= p49_array_index_1085724_comb;
    p49_array_index_1085725 <= p49_array_index_1085725_comb;
    p49_array_index_1085726 <= p49_array_index_1085726_comb;
    p49_array_index_1085727 <= p49_array_index_1085727_comb;
    p49_array_index_1085728 <= p49_array_index_1085728_comb;
    p49_res7__257 <= p49_res7__257_comb;
    p49_array_index_1085738 <= p49_array_index_1085738_comb;
    p49_array_index_1085739 <= p49_array_index_1085739_comb;
    p49_array_index_1085740 <= p49_array_index_1085740_comb;
    p49_array_index_1085741 <= p49_array_index_1085741_comb;
    p49_array_index_1085742 <= p49_array_index_1085742_comb;
    p49_res7__258 <= p49_res7__258_comb;
    p49_array_index_1085752 <= p49_array_index_1085752_comb;
    p49_array_index_1085753 <= p49_array_index_1085753_comb;
    p49_array_index_1085754 <= p49_array_index_1085754_comb;
    p49_array_index_1085755 <= p49_array_index_1085755_comb;
    p49_array_index_1085756 <= p49_array_index_1085756_comb;
    p49_res7__259 <= p49_res7__259_comb;
    p49_array_index_1085767 <= p49_array_index_1085767_comb;
    p49_array_index_1085768 <= p49_array_index_1085768_comb;
    p49_array_index_1085769 <= p49_array_index_1085769_comb;
    p49_array_index_1085770 <= p49_array_index_1085770_comb;
    p49_res7__260 <= p49_res7__260_comb;
    p49_array_index_1085778 <= p49_array_index_1085778_comb;
    p49_array_index_1085779 <= p49_array_index_1085779_comb;
    p49_array_index_1085780 <= p49_array_index_1085780_comb;
    p49_array_index_1085781 <= p49_array_index_1085781_comb;
    p49_array_index_1085782 <= p49_array_index_1085782_comb;
    p49_array_index_1085783 <= p49_array_index_1085783_comb;
    p49_array_index_1085784 <= p49_array_index_1085784_comb;
    p49_array_index_1085785 <= p49_array_index_1085785_comb;
    p49_array_index_1085786 <= p49_array_index_1085786_comb;
    p49_array_index_1085791 <= p49_array_index_1085791_comb;
    p49_array_index_1085792 <= p49_array_index_1085792_comb;
    p49_array_index_1085793 <= p49_array_index_1085793_comb;
    p49_array_index_1085794 <= p49_array_index_1085794_comb;
    p49_array_index_1085795 <= p49_array_index_1085795_comb;
    p49_array_index_1085797 <= p49_array_index_1085797_comb;
    p49_array_index_1085799 <= p49_array_index_1085799_comb;
    p49_res7__576 <= p49_res7__576_comb;
    p49_array_index_1085808 <= p49_array_index_1085808_comb;
    p49_array_index_1085809 <= p49_array_index_1085809_comb;
    p49_array_index_1085810 <= p49_array_index_1085810_comb;
    p49_array_index_1085811 <= p49_array_index_1085811_comb;
    p49_array_index_1085812 <= p49_array_index_1085812_comb;
    p49_array_index_1085813 <= p49_array_index_1085813_comb;
    p49_res7__577 <= p49_res7__577_comb;
    p49_array_index_1085823 <= p49_array_index_1085823_comb;
    p49_array_index_1085824 <= p49_array_index_1085824_comb;
    p49_array_index_1085825 <= p49_array_index_1085825_comb;
    p49_array_index_1085826 <= p49_array_index_1085826_comb;
    p49_array_index_1085827 <= p49_array_index_1085827_comb;
    p49_res7__578 <= p49_res7__578_comb;
    p49_array_index_1085837 <= p49_array_index_1085837_comb;
    p49_array_index_1085838 <= p49_array_index_1085838_comb;
    p49_array_index_1085839 <= p49_array_index_1085839_comb;
    p49_array_index_1085840 <= p49_array_index_1085840_comb;
    p49_array_index_1085841 <= p49_array_index_1085841_comb;
    p49_res7__579 <= p49_res7__579_comb;
    p49_array_index_1085852 <= p49_array_index_1085852_comb;
    p49_array_index_1085853 <= p49_array_index_1085853_comb;
    p49_array_index_1085854 <= p49_array_index_1085854_comb;
    p49_array_index_1085855 <= p49_array_index_1085855_comb;
    p49_res7__580 <= p49_res7__580_comb;
    p50_arr <= p49_arr;
    p50_literal_1076345 <= p49_literal_1076345;
    p50_literal_1076347 <= p49_literal_1076347;
    p50_literal_1076349 <= p49_literal_1076349;
    p50_literal_1076351 <= p49_literal_1076351;
    p50_literal_1076353 <= p49_literal_1076353;
    p50_literal_1076355 <= p49_literal_1076355;
    p50_literal_1076358 <= p49_literal_1076358;
  end

  // ===== Pipe stage 50:
  wire [7:0] p50_array_index_1086049_comb;
  wire [7:0] p50_array_index_1086050_comb;
  wire [7:0] p50_array_index_1086051_comb;
  wire [7:0] p50_array_index_1086052_comb;
  wire [7:0] p50_array_index_1086117_comb;
  wire [7:0] p50_array_index_1086118_comb;
  wire [7:0] p50_array_index_1086119_comb;
  wire [7:0] p50_array_index_1086120_comb;
  wire [7:0] p50_res7__261_comb;
  wire [7:0] p50_res7__581_comb;
  wire [7:0] p50_array_index_1086063_comb;
  wire [7:0] p50_array_index_1086064_comb;
  wire [7:0] p50_array_index_1086065_comb;
  wire [7:0] p50_array_index_1086131_comb;
  wire [7:0] p50_array_index_1086132_comb;
  wire [7:0] p50_array_index_1086133_comb;
  wire [7:0] p50_res7__262_comb;
  wire [7:0] p50_res7__582_comb;
  wire [7:0] p50_array_index_1086075_comb;
  wire [7:0] p50_array_index_1086076_comb;
  wire [7:0] p50_array_index_1086077_comb;
  wire [7:0] p50_array_index_1086143_comb;
  wire [7:0] p50_array_index_1086144_comb;
  wire [7:0] p50_array_index_1086145_comb;
  wire [7:0] p50_res7__263_comb;
  wire [7:0] p50_res7__583_comb;
  wire [7:0] p50_array_index_1086088_comb;
  wire [7:0] p50_array_index_1086089_comb;
  wire [7:0] p50_array_index_1086156_comb;
  wire [7:0] p50_array_index_1086157_comb;
  wire [7:0] p50_res7__264_comb;
  wire [7:0] p50_res7__584_comb;
  wire [7:0] p50_array_index_1086099_comb;
  wire [7:0] p50_array_index_1086100_comb;
  wire [7:0] p50_array_index_1086167_comb;
  wire [7:0] p50_array_index_1086168_comb;
  wire [7:0] p50_res7__265_comb;
  wire [7:0] p50_res7__585_comb;
  wire [7:0] p50_array_index_1086106_comb;
  wire [7:0] p50_array_index_1086107_comb;
  wire [7:0] p50_array_index_1086108_comb;
  wire [7:0] p50_array_index_1086109_comb;
  wire [7:0] p50_array_index_1086110_comb;
  wire [7:0] p50_array_index_1086111_comb;
  wire [7:0] p50_array_index_1086112_comb;
  wire [7:0] p50_array_index_1086113_comb;
  wire [7:0] p50_array_index_1086114_comb;
  wire [7:0] p50_array_index_1086174_comb;
  wire [7:0] p50_array_index_1086175_comb;
  wire [7:0] p50_array_index_1086176_comb;
  wire [7:0] p50_array_index_1086177_comb;
  wire [7:0] p50_array_index_1086178_comb;
  wire [7:0] p50_array_index_1086179_comb;
  wire [7:0] p50_array_index_1086180_comb;
  wire [7:0] p50_array_index_1086181_comb;
  wire [7:0] p50_array_index_1086182_comb;
  assign p50_array_index_1086049_comb = p49_literal_1076349[p49_res7__258];
  assign p50_array_index_1086050_comb = p49_literal_1076351[p49_res7__257];
  assign p50_array_index_1086051_comb = p49_literal_1076353[p49_res7__256];
  assign p50_array_index_1086052_comb = p49_literal_1076355[p49_array_index_1085690];
  assign p50_array_index_1086117_comb = p49_literal_1076349[p49_res7__578];
  assign p50_array_index_1086118_comb = p49_literal_1076351[p49_res7__577];
  assign p50_array_index_1086119_comb = p49_literal_1076353[p49_res7__576];
  assign p50_array_index_1086120_comb = p49_literal_1076355[p49_array_index_1085778];
  assign p50_res7__261_comb = p49_literal_1076345[p49_res7__260] ^ p49_literal_1076347[p49_res7__259] ^ p50_array_index_1086049_comb ^ p50_array_index_1086050_comb ^ p50_array_index_1086051_comb ^ p50_array_index_1086052_comb ^ p49_array_index_1085691 ^ p49_literal_1076358[p49_array_index_1085692] ^ p49_array_index_1085693 ^ p49_array_index_1085728 ^ p49_literal_1076353[p49_array_index_1085695] ^ p49_literal_1076351[p49_array_index_1085712] ^ p49_literal_1076349[p49_array_index_1085697] ^ p49_literal_1076347[p49_array_index_1085714] ^ p49_literal_1076345[p49_array_index_1085699] ^ p49_array_index_1085700;
  assign p50_res7__581_comb = p49_literal_1076345[p49_res7__580] ^ p49_literal_1076347[p49_res7__579] ^ p50_array_index_1086117_comb ^ p50_array_index_1086118_comb ^ p50_array_index_1086119_comb ^ p50_array_index_1086120_comb ^ p49_array_index_1085779 ^ p49_literal_1076358[p49_array_index_1085780] ^ p49_array_index_1085781 ^ p49_array_index_1085813 ^ p49_literal_1076353[p49_array_index_1085783] ^ p49_literal_1076351[p49_array_index_1085797] ^ p49_literal_1076349[p49_array_index_1085784] ^ p49_literal_1076347[p49_array_index_1085799] ^ p49_literal_1076345[p49_array_index_1085785] ^ p49_array_index_1085786;
  assign p50_array_index_1086063_comb = p49_literal_1076351[p49_res7__258];
  assign p50_array_index_1086064_comb = p49_literal_1076353[p49_res7__257];
  assign p50_array_index_1086065_comb = p49_literal_1076355[p49_res7__256];
  assign p50_array_index_1086131_comb = p49_literal_1076351[p49_res7__578];
  assign p50_array_index_1086132_comb = p49_literal_1076353[p49_res7__577];
  assign p50_array_index_1086133_comb = p49_literal_1076355[p49_res7__576];
  assign p50_res7__262_comb = p49_literal_1076345[p50_res7__261_comb] ^ p49_literal_1076347[p49_res7__260] ^ p49_literal_1076349[p49_res7__259] ^ p50_array_index_1086063_comb ^ p50_array_index_1086064_comb ^ p50_array_index_1086065_comb ^ p49_array_index_1085690 ^ p49_literal_1076358[p49_array_index_1085691] ^ p49_array_index_1085692 ^ p49_array_index_1085742 ^ p49_array_index_1085710 ^ p49_literal_1076351[p49_array_index_1085695] ^ p49_literal_1076349[p49_array_index_1085712] ^ p49_literal_1076347[p49_array_index_1085697] ^ p49_literal_1076345[p49_array_index_1085714] ^ p49_array_index_1085699;
  assign p50_res7__582_comb = p49_literal_1076345[p50_res7__581_comb] ^ p49_literal_1076347[p49_res7__580] ^ p49_literal_1076349[p49_res7__579] ^ p50_array_index_1086131_comb ^ p50_array_index_1086132_comb ^ p50_array_index_1086133_comb ^ p49_array_index_1085778 ^ p49_literal_1076358[p49_array_index_1085779] ^ p49_array_index_1085780 ^ p49_array_index_1085827 ^ p49_array_index_1085795 ^ p49_literal_1076351[p49_array_index_1085783] ^ p49_literal_1076349[p49_array_index_1085797] ^ p49_literal_1076347[p49_array_index_1085784] ^ p49_literal_1076345[p49_array_index_1085799] ^ p49_array_index_1085785;
  assign p50_array_index_1086075_comb = p49_literal_1076351[p49_res7__259];
  assign p50_array_index_1086076_comb = p49_literal_1076353[p49_res7__258];
  assign p50_array_index_1086077_comb = p49_literal_1076355[p49_res7__257];
  assign p50_array_index_1086143_comb = p49_literal_1076351[p49_res7__579];
  assign p50_array_index_1086144_comb = p49_literal_1076353[p49_res7__578];
  assign p50_array_index_1086145_comb = p49_literal_1076355[p49_res7__577];
  assign p50_res7__263_comb = p49_literal_1076345[p50_res7__262_comb] ^ p49_literal_1076347[p50_res7__261_comb] ^ p49_literal_1076349[p49_res7__260] ^ p50_array_index_1086075_comb ^ p50_array_index_1086076_comb ^ p50_array_index_1086077_comb ^ p49_res7__256 ^ p49_literal_1076358[p49_array_index_1085690] ^ p49_array_index_1085691 ^ p49_array_index_1085756 ^ p49_array_index_1085727 ^ p49_literal_1076351[p49_array_index_1085694] ^ p49_literal_1076349[p49_array_index_1085695] ^ p49_literal_1076347[p49_array_index_1085712] ^ p49_literal_1076345[p49_array_index_1085697] ^ p49_array_index_1085714;
  assign p50_res7__583_comb = p49_literal_1076345[p50_res7__582_comb] ^ p49_literal_1076347[p50_res7__581_comb] ^ p49_literal_1076349[p49_res7__580] ^ p50_array_index_1086143_comb ^ p50_array_index_1086144_comb ^ p50_array_index_1086145_comb ^ p49_res7__576 ^ p49_literal_1076358[p49_array_index_1085778] ^ p49_array_index_1085779 ^ p49_array_index_1085841 ^ p49_array_index_1085812 ^ p49_literal_1076351[p49_array_index_1085782] ^ p49_literal_1076349[p49_array_index_1085783] ^ p49_literal_1076347[p49_array_index_1085797] ^ p49_literal_1076345[p49_array_index_1085784] ^ p49_array_index_1085799;
  assign p50_array_index_1086088_comb = p49_literal_1076353[p49_res7__259];
  assign p50_array_index_1086089_comb = p49_literal_1076355[p49_res7__258];
  assign p50_array_index_1086156_comb = p49_literal_1076353[p49_res7__579];
  assign p50_array_index_1086157_comb = p49_literal_1076355[p49_res7__578];
  assign p50_res7__264_comb = p49_literal_1076345[p50_res7__263_comb] ^ p49_literal_1076347[p50_res7__262_comb] ^ p49_literal_1076349[p50_res7__261_comb] ^ p49_literal_1076351[p49_res7__260] ^ p50_array_index_1086088_comb ^ p50_array_index_1086089_comb ^ p49_res7__257 ^ p49_literal_1076358[p49_res7__256] ^ p49_array_index_1085690 ^ p49_array_index_1085770 ^ p49_array_index_1085741 ^ p49_array_index_1085709 ^ p49_literal_1076349[p49_array_index_1085694] ^ p49_literal_1076347[p49_array_index_1085695] ^ p49_literal_1076345[p49_array_index_1085712] ^ p49_array_index_1085697;
  assign p50_res7__584_comb = p49_literal_1076345[p50_res7__583_comb] ^ p49_literal_1076347[p50_res7__582_comb] ^ p49_literal_1076349[p50_res7__581_comb] ^ p49_literal_1076351[p49_res7__580] ^ p50_array_index_1086156_comb ^ p50_array_index_1086157_comb ^ p49_res7__577 ^ p49_literal_1076358[p49_res7__576] ^ p49_array_index_1085778 ^ p49_array_index_1085855 ^ p49_array_index_1085826 ^ p49_array_index_1085794 ^ p49_literal_1076349[p49_array_index_1085782] ^ p49_literal_1076347[p49_array_index_1085783] ^ p49_literal_1076345[p49_array_index_1085797] ^ p49_array_index_1085784;
  assign p50_array_index_1086099_comb = p49_literal_1076353[p49_res7__260];
  assign p50_array_index_1086100_comb = p49_literal_1076355[p49_res7__259];
  assign p50_array_index_1086167_comb = p49_literal_1076353[p49_res7__580];
  assign p50_array_index_1086168_comb = p49_literal_1076355[p49_res7__579];
  assign p50_res7__265_comb = p49_literal_1076345[p50_res7__264_comb] ^ p49_literal_1076347[p50_res7__263_comb] ^ p49_literal_1076349[p50_res7__262_comb] ^ p49_literal_1076351[p50_res7__261_comb] ^ p50_array_index_1086099_comb ^ p50_array_index_1086100_comb ^ p49_res7__258 ^ p49_literal_1076358[p49_res7__257] ^ p49_res7__256 ^ p50_array_index_1086052_comb ^ p49_array_index_1085755 ^ p49_array_index_1085726 ^ p49_literal_1076349[p49_array_index_1085693] ^ p49_literal_1076347[p49_array_index_1085694] ^ p49_literal_1076345[p49_array_index_1085695] ^ p49_array_index_1085712;
  assign p50_res7__585_comb = p49_literal_1076345[p50_res7__584_comb] ^ p49_literal_1076347[p50_res7__583_comb] ^ p49_literal_1076349[p50_res7__582_comb] ^ p49_literal_1076351[p50_res7__581_comb] ^ p50_array_index_1086167_comb ^ p50_array_index_1086168_comb ^ p49_res7__578 ^ p49_literal_1076358[p49_res7__577] ^ p49_res7__576 ^ p50_array_index_1086120_comb ^ p49_array_index_1085840 ^ p49_array_index_1085811 ^ p49_literal_1076349[p49_array_index_1085781] ^ p49_literal_1076347[p49_array_index_1085782] ^ p49_literal_1076345[p49_array_index_1085783] ^ p49_array_index_1085797;
  assign p50_array_index_1086106_comb = p49_literal_1076345[p50_res7__265_comb];
  assign p50_array_index_1086107_comb = p49_literal_1076347[p50_res7__264_comb];
  assign p50_array_index_1086108_comb = p49_literal_1076349[p50_res7__263_comb];
  assign p50_array_index_1086109_comb = p49_literal_1076351[p50_res7__262_comb];
  assign p50_array_index_1086110_comb = p49_literal_1076353[p50_res7__261_comb];
  assign p50_array_index_1086111_comb = p49_literal_1076355[p49_res7__260];
  assign p50_array_index_1086112_comb = p49_literal_1076358[p49_res7__258];
  assign p50_array_index_1086113_comb = p49_literal_1076347[p49_array_index_1085693];
  assign p50_array_index_1086114_comb = p49_literal_1076345[p49_array_index_1085694];
  assign p50_array_index_1086174_comb = p49_literal_1076345[p50_res7__585_comb];
  assign p50_array_index_1086175_comb = p49_literal_1076347[p50_res7__584_comb];
  assign p50_array_index_1086176_comb = p49_literal_1076349[p50_res7__583_comb];
  assign p50_array_index_1086177_comb = p49_literal_1076351[p50_res7__582_comb];
  assign p50_array_index_1086178_comb = p49_literal_1076353[p50_res7__581_comb];
  assign p50_array_index_1086179_comb = p49_literal_1076355[p49_res7__580];
  assign p50_array_index_1086180_comb = p49_literal_1076358[p49_res7__578];
  assign p50_array_index_1086181_comb = p49_literal_1076347[p49_array_index_1085781];
  assign p50_array_index_1086182_comb = p49_literal_1076345[p49_array_index_1085782];

  // Registers for pipe stage 50:
  reg [127:0] p50_k5;
  reg [127:0] p50_k4;
  reg [7:0] p50_array_index_1085690;
  reg [7:0] p50_array_index_1085691;
  reg [7:0] p50_array_index_1085692;
  reg [7:0] p50_array_index_1085693;
  reg [7:0] p50_array_index_1085694;
  reg [7:0] p50_array_index_1085695;
  reg [7:0] p50_array_index_1085706;
  reg [7:0] p50_array_index_1085707;
  reg [7:0] p50_array_index_1085708;
  reg [7:0] p50_res7__256;
  reg [7:0] p50_array_index_1085723;
  reg [7:0] p50_array_index_1085724;
  reg [7:0] p50_array_index_1085725;
  reg [7:0] p50_res7__257;
  reg [7:0] p50_array_index_1085738;
  reg [7:0] p50_array_index_1085739;
  reg [7:0] p50_array_index_1085740;
  reg [7:0] p50_res7__258;
  reg [7:0] p50_array_index_1085752;
  reg [7:0] p50_array_index_1085753;
  reg [7:0] p50_array_index_1085754;
  reg [7:0] p50_res7__259;
  reg [7:0] p50_array_index_1085767;
  reg [7:0] p50_array_index_1085768;
  reg [7:0] p50_array_index_1085769;
  reg [7:0] p50_res7__260;
  reg [7:0] p50_array_index_1086049;
  reg [7:0] p50_array_index_1086050;
  reg [7:0] p50_array_index_1086051;
  reg [7:0] p50_res7__261;
  reg [7:0] p50_array_index_1086063;
  reg [7:0] p50_array_index_1086064;
  reg [7:0] p50_array_index_1086065;
  reg [7:0] p50_res7__262;
  reg [7:0] p50_array_index_1086075;
  reg [7:0] p50_array_index_1086076;
  reg [7:0] p50_array_index_1086077;
  reg [7:0] p50_res7__263;
  reg [7:0] p50_array_index_1086088;
  reg [7:0] p50_array_index_1086089;
  reg [7:0] p50_res7__264;
  reg [7:0] p50_array_index_1086099;
  reg [7:0] p50_array_index_1086100;
  reg [7:0] p50_res7__265;
  reg [7:0] p50_array_index_1086106;
  reg [7:0] p50_array_index_1086107;
  reg [7:0] p50_array_index_1086108;
  reg [7:0] p50_array_index_1086109;
  reg [7:0] p50_array_index_1086110;
  reg [7:0] p50_array_index_1086111;
  reg [7:0] p50_array_index_1086112;
  reg [7:0] p50_array_index_1086113;
  reg [7:0] p50_array_index_1086114;
  reg [7:0] p50_array_index_1085778;
  reg [7:0] p50_array_index_1085779;
  reg [7:0] p50_array_index_1085780;
  reg [7:0] p50_array_index_1085781;
  reg [7:0] p50_array_index_1085782;
  reg [7:0] p50_array_index_1085783;
  reg [7:0] p50_array_index_1085791;
  reg [7:0] p50_array_index_1085792;
  reg [7:0] p50_array_index_1085793;
  reg [7:0] p50_res7__576;
  reg [7:0] p50_array_index_1085808;
  reg [7:0] p50_array_index_1085809;
  reg [7:0] p50_array_index_1085810;
  reg [7:0] p50_res7__577;
  reg [7:0] p50_array_index_1085823;
  reg [7:0] p50_array_index_1085824;
  reg [7:0] p50_array_index_1085825;
  reg [7:0] p50_res7__578;
  reg [7:0] p50_array_index_1085837;
  reg [7:0] p50_array_index_1085838;
  reg [7:0] p50_array_index_1085839;
  reg [7:0] p50_res7__579;
  reg [7:0] p50_array_index_1085852;
  reg [7:0] p50_array_index_1085853;
  reg [7:0] p50_array_index_1085854;
  reg [7:0] p50_res7__580;
  reg [7:0] p50_array_index_1086117;
  reg [7:0] p50_array_index_1086118;
  reg [7:0] p50_array_index_1086119;
  reg [7:0] p50_res7__581;
  reg [7:0] p50_array_index_1086131;
  reg [7:0] p50_array_index_1086132;
  reg [7:0] p50_array_index_1086133;
  reg [7:0] p50_res7__582;
  reg [7:0] p50_array_index_1086143;
  reg [7:0] p50_array_index_1086144;
  reg [7:0] p50_array_index_1086145;
  reg [7:0] p50_res7__583;
  reg [7:0] p50_array_index_1086156;
  reg [7:0] p50_array_index_1086157;
  reg [7:0] p50_res7__584;
  reg [7:0] p50_array_index_1086167;
  reg [7:0] p50_array_index_1086168;
  reg [7:0] p50_res7__585;
  reg [7:0] p50_array_index_1086174;
  reg [7:0] p50_array_index_1086175;
  reg [7:0] p50_array_index_1086176;
  reg [7:0] p50_array_index_1086177;
  reg [7:0] p50_array_index_1086178;
  reg [7:0] p50_array_index_1086179;
  reg [7:0] p50_array_index_1086180;
  reg [7:0] p50_array_index_1086181;
  reg [7:0] p50_array_index_1086182;
  reg [7:0] p51_arr[256];
  reg [7:0] p51_literal_1076345[256];
  reg [7:0] p51_literal_1076347[256];
  reg [7:0] p51_literal_1076349[256];
  reg [7:0] p51_literal_1076351[256];
  reg [7:0] p51_literal_1076353[256];
  reg [7:0] p51_literal_1076355[256];
  reg [7:0] p51_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p50_k5 <= p49_k5;
    p50_k4 <= p49_k4;
    p50_array_index_1085690 <= p49_array_index_1085690;
    p50_array_index_1085691 <= p49_array_index_1085691;
    p50_array_index_1085692 <= p49_array_index_1085692;
    p50_array_index_1085693 <= p49_array_index_1085693;
    p50_array_index_1085694 <= p49_array_index_1085694;
    p50_array_index_1085695 <= p49_array_index_1085695;
    p50_array_index_1085706 <= p49_array_index_1085706;
    p50_array_index_1085707 <= p49_array_index_1085707;
    p50_array_index_1085708 <= p49_array_index_1085708;
    p50_res7__256 <= p49_res7__256;
    p50_array_index_1085723 <= p49_array_index_1085723;
    p50_array_index_1085724 <= p49_array_index_1085724;
    p50_array_index_1085725 <= p49_array_index_1085725;
    p50_res7__257 <= p49_res7__257;
    p50_array_index_1085738 <= p49_array_index_1085738;
    p50_array_index_1085739 <= p49_array_index_1085739;
    p50_array_index_1085740 <= p49_array_index_1085740;
    p50_res7__258 <= p49_res7__258;
    p50_array_index_1085752 <= p49_array_index_1085752;
    p50_array_index_1085753 <= p49_array_index_1085753;
    p50_array_index_1085754 <= p49_array_index_1085754;
    p50_res7__259 <= p49_res7__259;
    p50_array_index_1085767 <= p49_array_index_1085767;
    p50_array_index_1085768 <= p49_array_index_1085768;
    p50_array_index_1085769 <= p49_array_index_1085769;
    p50_res7__260 <= p49_res7__260;
    p50_array_index_1086049 <= p50_array_index_1086049_comb;
    p50_array_index_1086050 <= p50_array_index_1086050_comb;
    p50_array_index_1086051 <= p50_array_index_1086051_comb;
    p50_res7__261 <= p50_res7__261_comb;
    p50_array_index_1086063 <= p50_array_index_1086063_comb;
    p50_array_index_1086064 <= p50_array_index_1086064_comb;
    p50_array_index_1086065 <= p50_array_index_1086065_comb;
    p50_res7__262 <= p50_res7__262_comb;
    p50_array_index_1086075 <= p50_array_index_1086075_comb;
    p50_array_index_1086076 <= p50_array_index_1086076_comb;
    p50_array_index_1086077 <= p50_array_index_1086077_comb;
    p50_res7__263 <= p50_res7__263_comb;
    p50_array_index_1086088 <= p50_array_index_1086088_comb;
    p50_array_index_1086089 <= p50_array_index_1086089_comb;
    p50_res7__264 <= p50_res7__264_comb;
    p50_array_index_1086099 <= p50_array_index_1086099_comb;
    p50_array_index_1086100 <= p50_array_index_1086100_comb;
    p50_res7__265 <= p50_res7__265_comb;
    p50_array_index_1086106 <= p50_array_index_1086106_comb;
    p50_array_index_1086107 <= p50_array_index_1086107_comb;
    p50_array_index_1086108 <= p50_array_index_1086108_comb;
    p50_array_index_1086109 <= p50_array_index_1086109_comb;
    p50_array_index_1086110 <= p50_array_index_1086110_comb;
    p50_array_index_1086111 <= p50_array_index_1086111_comb;
    p50_array_index_1086112 <= p50_array_index_1086112_comb;
    p50_array_index_1086113 <= p50_array_index_1086113_comb;
    p50_array_index_1086114 <= p50_array_index_1086114_comb;
    p50_array_index_1085778 <= p49_array_index_1085778;
    p50_array_index_1085779 <= p49_array_index_1085779;
    p50_array_index_1085780 <= p49_array_index_1085780;
    p50_array_index_1085781 <= p49_array_index_1085781;
    p50_array_index_1085782 <= p49_array_index_1085782;
    p50_array_index_1085783 <= p49_array_index_1085783;
    p50_array_index_1085791 <= p49_array_index_1085791;
    p50_array_index_1085792 <= p49_array_index_1085792;
    p50_array_index_1085793 <= p49_array_index_1085793;
    p50_res7__576 <= p49_res7__576;
    p50_array_index_1085808 <= p49_array_index_1085808;
    p50_array_index_1085809 <= p49_array_index_1085809;
    p50_array_index_1085810 <= p49_array_index_1085810;
    p50_res7__577 <= p49_res7__577;
    p50_array_index_1085823 <= p49_array_index_1085823;
    p50_array_index_1085824 <= p49_array_index_1085824;
    p50_array_index_1085825 <= p49_array_index_1085825;
    p50_res7__578 <= p49_res7__578;
    p50_array_index_1085837 <= p49_array_index_1085837;
    p50_array_index_1085838 <= p49_array_index_1085838;
    p50_array_index_1085839 <= p49_array_index_1085839;
    p50_res7__579 <= p49_res7__579;
    p50_array_index_1085852 <= p49_array_index_1085852;
    p50_array_index_1085853 <= p49_array_index_1085853;
    p50_array_index_1085854 <= p49_array_index_1085854;
    p50_res7__580 <= p49_res7__580;
    p50_array_index_1086117 <= p50_array_index_1086117_comb;
    p50_array_index_1086118 <= p50_array_index_1086118_comb;
    p50_array_index_1086119 <= p50_array_index_1086119_comb;
    p50_res7__581 <= p50_res7__581_comb;
    p50_array_index_1086131 <= p50_array_index_1086131_comb;
    p50_array_index_1086132 <= p50_array_index_1086132_comb;
    p50_array_index_1086133 <= p50_array_index_1086133_comb;
    p50_res7__582 <= p50_res7__582_comb;
    p50_array_index_1086143 <= p50_array_index_1086143_comb;
    p50_array_index_1086144 <= p50_array_index_1086144_comb;
    p50_array_index_1086145 <= p50_array_index_1086145_comb;
    p50_res7__583 <= p50_res7__583_comb;
    p50_array_index_1086156 <= p50_array_index_1086156_comb;
    p50_array_index_1086157 <= p50_array_index_1086157_comb;
    p50_res7__584 <= p50_res7__584_comb;
    p50_array_index_1086167 <= p50_array_index_1086167_comb;
    p50_array_index_1086168 <= p50_array_index_1086168_comb;
    p50_res7__585 <= p50_res7__585_comb;
    p50_array_index_1086174 <= p50_array_index_1086174_comb;
    p50_array_index_1086175 <= p50_array_index_1086175_comb;
    p50_array_index_1086176 <= p50_array_index_1086176_comb;
    p50_array_index_1086177 <= p50_array_index_1086177_comb;
    p50_array_index_1086178 <= p50_array_index_1086178_comb;
    p50_array_index_1086179 <= p50_array_index_1086179_comb;
    p50_array_index_1086180 <= p50_array_index_1086180_comb;
    p50_array_index_1086181 <= p50_array_index_1086181_comb;
    p50_array_index_1086182 <= p50_array_index_1086182_comb;
    p51_arr <= p50_arr;
    p51_literal_1076345 <= p50_literal_1076345;
    p51_literal_1076347 <= p50_literal_1076347;
    p51_literal_1076349 <= p50_literal_1076349;
    p51_literal_1076351 <= p50_literal_1076351;
    p51_literal_1076353 <= p50_literal_1076353;
    p51_literal_1076355 <= p50_literal_1076355;
    p51_literal_1076358 <= p50_literal_1076358;
  end

  // ===== Pipe stage 51:
  wire [7:0] p51_res7__586_comb;
  wire [7:0] p51_res7__266_comb;
  wire [7:0] p51_array_index_1086468_comb;
  wire [7:0] p51_array_index_1086421_comb;
  wire [7:0] p51_res7__587_comb;
  wire [7:0] p51_res7__267_comb;
  wire [7:0] p51_res7__588_comb;
  wire [7:0] p51_res7__268_comb;
  wire [7:0] p51_res7__589_comb;
  wire [7:0] p51_res7__269_comb;
  wire [7:0] p51_res7__590_comb;
  wire [7:0] p51_res7__270_comb;
  wire [7:0] p51_res7__591_comb;
  wire [7:0] p51_res7__271_comb;
  wire [127:0] p51_res__36_comb;
  wire [127:0] p51_res__16_comb;
  wire [127:0] p51_addedKey__37_comb;
  wire [127:0] p51_xor_1086461_comb;
  wire [7:0] p51_bit_slice_1086509_comb;
  wire [7:0] p51_bit_slice_1086510_comb;
  wire [7:0] p51_bit_slice_1086511_comb;
  wire [7:0] p51_bit_slice_1086512_comb;
  wire [7:0] p51_bit_slice_1086513_comb;
  wire [7:0] p51_bit_slice_1086514_comb;
  wire [7:0] p51_bit_slice_1086515_comb;
  wire [7:0] p51_bit_slice_1086516_comb;
  wire [7:0] p51_bit_slice_1086517_comb;
  wire [7:0] p51_bit_slice_1086518_comb;
  wire [7:0] p51_bit_slice_1086519_comb;
  wire [7:0] p51_bit_slice_1086520_comb;
  wire [7:0] p51_bit_slice_1086521_comb;
  wire [7:0] p51_bit_slice_1086522_comb;
  wire [7:0] p51_bit_slice_1086523_comb;
  wire [7:0] p51_bit_slice_1086524_comb;
  assign p51_res7__586_comb = p50_array_index_1086174 ^ p50_array_index_1086175 ^ p50_array_index_1086176 ^ p50_array_index_1086177 ^ p50_array_index_1086178 ^ p50_array_index_1086179 ^ p50_res7__579 ^ p50_array_index_1086180 ^ p50_res7__577 ^ p50_array_index_1086133 ^ p50_array_index_1085854 ^ p50_array_index_1085825 ^ p50_array_index_1085793 ^ p50_array_index_1086181 ^ p50_array_index_1086182 ^ p50_array_index_1085783;
  assign p51_res7__266_comb = p50_array_index_1086106 ^ p50_array_index_1086107 ^ p50_array_index_1086108 ^ p50_array_index_1086109 ^ p50_array_index_1086110 ^ p50_array_index_1086111 ^ p50_res7__259 ^ p50_array_index_1086112 ^ p50_res7__257 ^ p50_array_index_1086065 ^ p50_array_index_1085769 ^ p50_array_index_1085740 ^ p50_array_index_1085708 ^ p50_array_index_1086113 ^ p50_array_index_1086114 ^ p50_array_index_1085695;
  assign p51_array_index_1086468_comb = p50_literal_1076355[p50_res7__581];
  assign p51_array_index_1086421_comb = p50_literal_1076355[p50_res7__261];
  assign p51_res7__587_comb = p50_literal_1076345[p51_res7__586_comb] ^ p50_literal_1076347[p50_res7__585] ^ p50_literal_1076349[p50_res7__584] ^ p50_literal_1076351[p50_res7__583] ^ p50_literal_1076353[p50_res7__582] ^ p51_array_index_1086468_comb ^ p50_res7__580 ^ p50_literal_1076358[p50_res7__579] ^ p50_res7__578 ^ p50_array_index_1086145 ^ p50_array_index_1086119 ^ p50_array_index_1085839 ^ p50_array_index_1085810 ^ p50_literal_1076347[p50_array_index_1085780] ^ p50_literal_1076345[p50_array_index_1085781] ^ p50_array_index_1085782;
  assign p51_res7__267_comb = p50_literal_1076345[p51_res7__266_comb] ^ p50_literal_1076347[p50_res7__265] ^ p50_literal_1076349[p50_res7__264] ^ p50_literal_1076351[p50_res7__263] ^ p50_literal_1076353[p50_res7__262] ^ p51_array_index_1086421_comb ^ p50_res7__260 ^ p50_literal_1076358[p50_res7__259] ^ p50_res7__258 ^ p50_array_index_1086077 ^ p50_array_index_1086051 ^ p50_array_index_1085754 ^ p50_array_index_1085725 ^ p50_literal_1076347[p50_array_index_1085692] ^ p50_literal_1076345[p50_array_index_1085693] ^ p50_array_index_1085694;
  assign p51_res7__588_comb = p50_literal_1076345[p51_res7__587_comb] ^ p50_literal_1076347[p51_res7__586_comb] ^ p50_literal_1076349[p50_res7__585] ^ p50_literal_1076351[p50_res7__584] ^ p50_literal_1076353[p50_res7__583] ^ p50_literal_1076355[p50_res7__582] ^ p50_res7__581 ^ p50_literal_1076358[p50_res7__580] ^ p50_res7__579 ^ p50_array_index_1086157 ^ p50_array_index_1086132 ^ p50_array_index_1085853 ^ p50_array_index_1085824 ^ p50_array_index_1085792 ^ p50_literal_1076345[p50_array_index_1085780] ^ p50_array_index_1085781;
  assign p51_res7__268_comb = p50_literal_1076345[p51_res7__267_comb] ^ p50_literal_1076347[p51_res7__266_comb] ^ p50_literal_1076349[p50_res7__265] ^ p50_literal_1076351[p50_res7__264] ^ p50_literal_1076353[p50_res7__263] ^ p50_literal_1076355[p50_res7__262] ^ p50_res7__261 ^ p50_literal_1076358[p50_res7__260] ^ p50_res7__259 ^ p50_array_index_1086089 ^ p50_array_index_1086064 ^ p50_array_index_1085768 ^ p50_array_index_1085739 ^ p50_array_index_1085707 ^ p50_literal_1076345[p50_array_index_1085692] ^ p50_array_index_1085693;
  assign p51_res7__589_comb = p50_literal_1076345[p51_res7__588_comb] ^ p50_literal_1076347[p51_res7__587_comb] ^ p50_literal_1076349[p51_res7__586_comb] ^ p50_literal_1076351[p50_res7__585] ^ p50_literal_1076353[p50_res7__584] ^ p50_literal_1076355[p50_res7__583] ^ p50_res7__582 ^ p50_literal_1076358[p50_res7__581] ^ p50_res7__580 ^ p50_array_index_1086168 ^ p50_array_index_1086144 ^ p50_array_index_1086118 ^ p50_array_index_1085838 ^ p50_array_index_1085809 ^ p50_literal_1076345[p50_array_index_1085779] ^ p50_array_index_1085780;
  assign p51_res7__269_comb = p50_literal_1076345[p51_res7__268_comb] ^ p50_literal_1076347[p51_res7__267_comb] ^ p50_literal_1076349[p51_res7__266_comb] ^ p50_literal_1076351[p50_res7__265] ^ p50_literal_1076353[p50_res7__264] ^ p50_literal_1076355[p50_res7__263] ^ p50_res7__262 ^ p50_literal_1076358[p50_res7__261] ^ p50_res7__260 ^ p50_array_index_1086100 ^ p50_array_index_1086076 ^ p50_array_index_1086050 ^ p50_array_index_1085753 ^ p50_array_index_1085724 ^ p50_literal_1076345[p50_array_index_1085691] ^ p50_array_index_1085692;
  assign p51_res7__590_comb = p50_literal_1076345[p51_res7__589_comb] ^ p50_literal_1076347[p51_res7__588_comb] ^ p50_literal_1076349[p51_res7__587_comb] ^ p50_literal_1076351[p51_res7__586_comb] ^ p50_literal_1076353[p50_res7__585] ^ p50_literal_1076355[p50_res7__584] ^ p50_res7__583 ^ p50_literal_1076358[p50_res7__582] ^ p50_res7__581 ^ p50_array_index_1086179 ^ p50_array_index_1086156 ^ p50_array_index_1086131 ^ p50_array_index_1085852 ^ p50_array_index_1085823 ^ p50_array_index_1085791 ^ p50_array_index_1085779;
  assign p51_res7__270_comb = p50_literal_1076345[p51_res7__269_comb] ^ p50_literal_1076347[p51_res7__268_comb] ^ p50_literal_1076349[p51_res7__267_comb] ^ p50_literal_1076351[p51_res7__266_comb] ^ p50_literal_1076353[p50_res7__265] ^ p50_literal_1076355[p50_res7__264] ^ p50_res7__263 ^ p50_literal_1076358[p50_res7__262] ^ p50_res7__261 ^ p50_array_index_1086111 ^ p50_array_index_1086088 ^ p50_array_index_1086063 ^ p50_array_index_1085767 ^ p50_array_index_1085738 ^ p50_array_index_1085706 ^ p50_array_index_1085691;
  assign p51_res7__591_comb = p50_literal_1076345[p51_res7__590_comb] ^ p50_literal_1076347[p51_res7__589_comb] ^ p50_literal_1076349[p51_res7__588_comb] ^ p50_literal_1076351[p51_res7__587_comb] ^ p50_literal_1076353[p51_res7__586_comb] ^ p50_literal_1076355[p50_res7__585] ^ p50_res7__584 ^ p50_literal_1076358[p50_res7__583] ^ p50_res7__582 ^ p51_array_index_1086468_comb ^ p50_array_index_1086167 ^ p50_array_index_1086143 ^ p50_array_index_1086117 ^ p50_array_index_1085837 ^ p50_array_index_1085808 ^ p50_array_index_1085778;
  assign p51_res7__271_comb = p50_literal_1076345[p51_res7__270_comb] ^ p50_literal_1076347[p51_res7__269_comb] ^ p50_literal_1076349[p51_res7__268_comb] ^ p50_literal_1076351[p51_res7__267_comb] ^ p50_literal_1076353[p51_res7__266_comb] ^ p50_literal_1076355[p50_res7__265] ^ p50_res7__264 ^ p50_literal_1076358[p50_res7__263] ^ p50_res7__262 ^ p51_array_index_1086421_comb ^ p50_array_index_1086099 ^ p50_array_index_1086075 ^ p50_array_index_1086049 ^ p50_array_index_1085752 ^ p50_array_index_1085723 ^ p50_array_index_1085690;
  assign p51_res__36_comb = {p51_res7__591_comb, p51_res7__590_comb, p51_res7__589_comb, p51_res7__588_comb, p51_res7__587_comb, p51_res7__586_comb, p50_res7__585, p50_res7__584, p50_res7__583, p50_res7__582, p50_res7__581, p50_res7__580, p50_res7__579, p50_res7__578, p50_res7__577, p50_res7__576};
  assign p51_res__16_comb = {p51_res7__271_comb, p51_res7__270_comb, p51_res7__269_comb, p51_res7__268_comb, p51_res7__267_comb, p51_res7__266_comb, p50_res7__265, p50_res7__264, p50_res7__263, p50_res7__262, p50_res7__261, p50_res7__260, p50_res7__259, p50_res7__258, p50_res7__257, p50_res7__256};
  assign p51_addedKey__37_comb = p50_k5 ^ p51_res__36_comb;
  assign p51_xor_1086461_comb = p51_res__16_comb ^ p50_k5;
  assign p51_bit_slice_1086509_comb = p51_addedKey__37_comb[127:120];
  assign p51_bit_slice_1086510_comb = p51_addedKey__37_comb[119:112];
  assign p51_bit_slice_1086511_comb = p51_addedKey__37_comb[111:104];
  assign p51_bit_slice_1086512_comb = p51_addedKey__37_comb[103:96];
  assign p51_bit_slice_1086513_comb = p51_addedKey__37_comb[95:88];
  assign p51_bit_slice_1086514_comb = p51_addedKey__37_comb[87:80];
  assign p51_bit_slice_1086515_comb = p51_addedKey__37_comb[71:64];
  assign p51_bit_slice_1086516_comb = p51_addedKey__37_comb[55:48];
  assign p51_bit_slice_1086517_comb = p51_addedKey__37_comb[47:40];
  assign p51_bit_slice_1086518_comb = p51_addedKey__37_comb[39:32];
  assign p51_bit_slice_1086519_comb = p51_addedKey__37_comb[31:24];
  assign p51_bit_slice_1086520_comb = p51_addedKey__37_comb[23:16];
  assign p51_bit_slice_1086521_comb = p51_addedKey__37_comb[15:8];
  assign p51_bit_slice_1086522_comb = p51_addedKey__37_comb[79:72];
  assign p51_bit_slice_1086523_comb = p51_addedKey__37_comb[63:56];
  assign p51_bit_slice_1086524_comb = p51_addedKey__37_comb[7:0];

  // Registers for pipe stage 51:
  reg [127:0] p51_k4;
  reg [127:0] p51_xor_1086461;
  reg [7:0] p51_bit_slice_1086509;
  reg [7:0] p51_bit_slice_1086510;
  reg [7:0] p51_bit_slice_1086511;
  reg [7:0] p51_bit_slice_1086512;
  reg [7:0] p51_bit_slice_1086513;
  reg [7:0] p51_bit_slice_1086514;
  reg [7:0] p51_bit_slice_1086515;
  reg [7:0] p51_bit_slice_1086516;
  reg [7:0] p51_bit_slice_1086517;
  reg [7:0] p51_bit_slice_1086518;
  reg [7:0] p51_bit_slice_1086519;
  reg [7:0] p51_bit_slice_1086520;
  reg [7:0] p51_bit_slice_1086521;
  reg [7:0] p51_bit_slice_1086522;
  reg [7:0] p51_bit_slice_1086523;
  reg [7:0] p51_bit_slice_1086524;
  reg [7:0] p52_arr[256];
  reg [7:0] p52_literal_1076345[256];
  reg [7:0] p52_literal_1076347[256];
  reg [7:0] p52_literal_1076349[256];
  reg [7:0] p52_literal_1076351[256];
  reg [7:0] p52_literal_1076353[256];
  reg [7:0] p52_literal_1076355[256];
  reg [7:0] p52_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p51_k4 <= p50_k4;
    p51_xor_1086461 <= p51_xor_1086461_comb;
    p51_bit_slice_1086509 <= p51_bit_slice_1086509_comb;
    p51_bit_slice_1086510 <= p51_bit_slice_1086510_comb;
    p51_bit_slice_1086511 <= p51_bit_slice_1086511_comb;
    p51_bit_slice_1086512 <= p51_bit_slice_1086512_comb;
    p51_bit_slice_1086513 <= p51_bit_slice_1086513_comb;
    p51_bit_slice_1086514 <= p51_bit_slice_1086514_comb;
    p51_bit_slice_1086515 <= p51_bit_slice_1086515_comb;
    p51_bit_slice_1086516 <= p51_bit_slice_1086516_comb;
    p51_bit_slice_1086517 <= p51_bit_slice_1086517_comb;
    p51_bit_slice_1086518 <= p51_bit_slice_1086518_comb;
    p51_bit_slice_1086519 <= p51_bit_slice_1086519_comb;
    p51_bit_slice_1086520 <= p51_bit_slice_1086520_comb;
    p51_bit_slice_1086521 <= p51_bit_slice_1086521_comb;
    p51_bit_slice_1086522 <= p51_bit_slice_1086522_comb;
    p51_bit_slice_1086523 <= p51_bit_slice_1086523_comb;
    p51_bit_slice_1086524 <= p51_bit_slice_1086524_comb;
    p52_arr <= p51_arr;
    p52_literal_1076345 <= p51_literal_1076345;
    p52_literal_1076347 <= p51_literal_1076347;
    p52_literal_1076349 <= p51_literal_1076349;
    p52_literal_1076351 <= p51_literal_1076351;
    p52_literal_1076353 <= p51_literal_1076353;
    p52_literal_1076355 <= p51_literal_1076355;
    p52_literal_1076358 <= p51_literal_1076358;
  end

  // ===== Pipe stage 52:
  wire [127:0] p52_addedKey__58_comb;
  wire [7:0] p52_array_index_1086592_comb;
  wire [7:0] p52_array_index_1086593_comb;
  wire [7:0] p52_array_index_1086594_comb;
  wire [7:0] p52_array_index_1086595_comb;
  wire [7:0] p52_array_index_1086596_comb;
  wire [7:0] p52_array_index_1086597_comb;
  wire [7:0] p52_array_index_1086599_comb;
  wire [7:0] p52_array_index_1086601_comb;
  wire [7:0] p52_array_index_1086602_comb;
  wire [7:0] p52_array_index_1086603_comb;
  wire [7:0] p52_array_index_1086604_comb;
  wire [7:0] p52_array_index_1086605_comb;
  wire [7:0] p52_array_index_1086606_comb;
  wire [7:0] p52_array_index_1086680_comb;
  wire [7:0] p52_array_index_1086681_comb;
  wire [7:0] p52_array_index_1086682_comb;
  wire [7:0] p52_array_index_1086683_comb;
  wire [7:0] p52_array_index_1086684_comb;
  wire [7:0] p52_array_index_1086685_comb;
  wire [7:0] p52_array_index_1086686_comb;
  wire [7:0] p52_array_index_1086687_comb;
  wire [7:0] p52_array_index_1086688_comb;
  wire [7:0] p52_array_index_1086689_comb;
  wire [7:0] p52_array_index_1086690_comb;
  wire [7:0] p52_array_index_1086691_comb;
  wire [7:0] p52_array_index_1086692_comb;
  wire [7:0] p52_array_index_1086608_comb;
  wire [7:0] p52_array_index_1086609_comb;
  wire [7:0] p52_array_index_1086610_comb;
  wire [7:0] p52_array_index_1086611_comb;
  wire [7:0] p52_array_index_1086612_comb;
  wire [7:0] p52_array_index_1086613_comb;
  wire [7:0] p52_array_index_1086614_comb;
  wire [7:0] p52_array_index_1086616_comb;
  wire [7:0] p52_array_index_1086693_comb;
  wire [7:0] p52_array_index_1086694_comb;
  wire [7:0] p52_array_index_1086695_comb;
  wire [7:0] p52_array_index_1086696_comb;
  wire [7:0] p52_array_index_1086697_comb;
  wire [7:0] p52_array_index_1086698_comb;
  wire [7:0] p52_array_index_1086699_comb;
  wire [7:0] p52_array_index_1086701_comb;
  wire [7:0] p52_res7__272_comb;
  wire [7:0] p52_res7__592_comb;
  wire [7:0] p52_array_index_1086625_comb;
  wire [7:0] p52_array_index_1086626_comb;
  wire [7:0] p52_array_index_1086627_comb;
  wire [7:0] p52_array_index_1086628_comb;
  wire [7:0] p52_array_index_1086629_comb;
  wire [7:0] p52_array_index_1086630_comb;
  wire [7:0] p52_array_index_1086710_comb;
  wire [7:0] p52_array_index_1086711_comb;
  wire [7:0] p52_array_index_1086712_comb;
  wire [7:0] p52_array_index_1086713_comb;
  wire [7:0] p52_array_index_1086714_comb;
  wire [7:0] p52_array_index_1086715_comb;
  wire [7:0] p52_res7__273_comb;
  wire [7:0] p52_res7__593_comb;
  wire [7:0] p52_array_index_1086640_comb;
  wire [7:0] p52_array_index_1086641_comb;
  wire [7:0] p52_array_index_1086642_comb;
  wire [7:0] p52_array_index_1086643_comb;
  wire [7:0] p52_array_index_1086644_comb;
  wire [7:0] p52_array_index_1086725_comb;
  wire [7:0] p52_array_index_1086726_comb;
  wire [7:0] p52_array_index_1086727_comb;
  wire [7:0] p52_array_index_1086728_comb;
  wire [7:0] p52_array_index_1086729_comb;
  wire [7:0] p52_res7__274_comb;
  wire [7:0] p52_res7__594_comb;
  wire [7:0] p52_array_index_1086654_comb;
  wire [7:0] p52_array_index_1086655_comb;
  wire [7:0] p52_array_index_1086656_comb;
  wire [7:0] p52_array_index_1086657_comb;
  wire [7:0] p52_array_index_1086658_comb;
  wire [7:0] p52_array_index_1086739_comb;
  wire [7:0] p52_array_index_1086740_comb;
  wire [7:0] p52_array_index_1086741_comb;
  wire [7:0] p52_array_index_1086742_comb;
  wire [7:0] p52_array_index_1086743_comb;
  wire [7:0] p52_res7__275_comb;
  wire [7:0] p52_res7__595_comb;
  wire [7:0] p52_array_index_1086669_comb;
  wire [7:0] p52_array_index_1086670_comb;
  wire [7:0] p52_array_index_1086671_comb;
  wire [7:0] p52_array_index_1086672_comb;
  wire [7:0] p52_array_index_1086754_comb;
  wire [7:0] p52_array_index_1086755_comb;
  wire [7:0] p52_array_index_1086756_comb;
  wire [7:0] p52_array_index_1086757_comb;
  wire [7:0] p52_res7__276_comb;
  wire [7:0] p52_res7__596_comb;
  assign p52_addedKey__58_comb = p51_xor_1086461 ^ 128'hf335_80c8_d79a_5862_237b_38e3_375c_bf12;
  assign p52_array_index_1086592_comb = p51_arr[p52_addedKey__58_comb[127:120]];
  assign p52_array_index_1086593_comb = p51_arr[p52_addedKey__58_comb[119:112]];
  assign p52_array_index_1086594_comb = p51_arr[p52_addedKey__58_comb[111:104]];
  assign p52_array_index_1086595_comb = p51_arr[p52_addedKey__58_comb[103:96]];
  assign p52_array_index_1086596_comb = p51_arr[p52_addedKey__58_comb[95:88]];
  assign p52_array_index_1086597_comb = p51_arr[p52_addedKey__58_comb[87:80]];
  assign p52_array_index_1086599_comb = p51_arr[p52_addedKey__58_comb[71:64]];
  assign p52_array_index_1086601_comb = p51_arr[p52_addedKey__58_comb[55:48]];
  assign p52_array_index_1086602_comb = p51_arr[p52_addedKey__58_comb[47:40]];
  assign p52_array_index_1086603_comb = p51_arr[p52_addedKey__58_comb[39:32]];
  assign p52_array_index_1086604_comb = p51_arr[p52_addedKey__58_comb[31:24]];
  assign p52_array_index_1086605_comb = p51_arr[p52_addedKey__58_comb[23:16]];
  assign p52_array_index_1086606_comb = p51_arr[p52_addedKey__58_comb[15:8]];
  assign p52_array_index_1086680_comb = p51_arr[p51_bit_slice_1086509];
  assign p52_array_index_1086681_comb = p51_arr[p51_bit_slice_1086510];
  assign p52_array_index_1086682_comb = p51_arr[p51_bit_slice_1086511];
  assign p52_array_index_1086683_comb = p51_arr[p51_bit_slice_1086512];
  assign p52_array_index_1086684_comb = p51_arr[p51_bit_slice_1086513];
  assign p52_array_index_1086685_comb = p51_arr[p51_bit_slice_1086514];
  assign p52_array_index_1086686_comb = p51_arr[p51_bit_slice_1086515];
  assign p52_array_index_1086687_comb = p51_arr[p51_bit_slice_1086516];
  assign p52_array_index_1086688_comb = p51_arr[p51_bit_slice_1086517];
  assign p52_array_index_1086689_comb = p51_arr[p51_bit_slice_1086518];
  assign p52_array_index_1086690_comb = p51_arr[p51_bit_slice_1086519];
  assign p52_array_index_1086691_comb = p51_arr[p51_bit_slice_1086520];
  assign p52_array_index_1086692_comb = p51_arr[p51_bit_slice_1086521];
  assign p52_array_index_1086608_comb = p51_literal_1076345[p52_array_index_1086592_comb];
  assign p52_array_index_1086609_comb = p51_literal_1076347[p52_array_index_1086593_comb];
  assign p52_array_index_1086610_comb = p51_literal_1076349[p52_array_index_1086594_comb];
  assign p52_array_index_1086611_comb = p51_literal_1076351[p52_array_index_1086595_comb];
  assign p52_array_index_1086612_comb = p51_literal_1076353[p52_array_index_1086596_comb];
  assign p52_array_index_1086613_comb = p51_literal_1076355[p52_array_index_1086597_comb];
  assign p52_array_index_1086614_comb = p51_arr[p52_addedKey__58_comb[79:72]];
  assign p52_array_index_1086616_comb = p51_arr[p52_addedKey__58_comb[63:56]];
  assign p52_array_index_1086693_comb = p51_literal_1076345[p52_array_index_1086680_comb];
  assign p52_array_index_1086694_comb = p51_literal_1076347[p52_array_index_1086681_comb];
  assign p52_array_index_1086695_comb = p51_literal_1076349[p52_array_index_1086682_comb];
  assign p52_array_index_1086696_comb = p51_literal_1076351[p52_array_index_1086683_comb];
  assign p52_array_index_1086697_comb = p51_literal_1076353[p52_array_index_1086684_comb];
  assign p52_array_index_1086698_comb = p51_literal_1076355[p52_array_index_1086685_comb];
  assign p52_array_index_1086699_comb = p51_arr[p51_bit_slice_1086522];
  assign p52_array_index_1086701_comb = p51_arr[p51_bit_slice_1086523];
  assign p52_res7__272_comb = p52_array_index_1086608_comb ^ p52_array_index_1086609_comb ^ p52_array_index_1086610_comb ^ p52_array_index_1086611_comb ^ p52_array_index_1086612_comb ^ p52_array_index_1086613_comb ^ p52_array_index_1086614_comb ^ p51_literal_1076358[p52_array_index_1086599_comb] ^ p52_array_index_1086616_comb ^ p51_literal_1076355[p52_array_index_1086601_comb] ^ p51_literal_1076353[p52_array_index_1086602_comb] ^ p51_literal_1076351[p52_array_index_1086603_comb] ^ p51_literal_1076349[p52_array_index_1086604_comb] ^ p51_literal_1076347[p52_array_index_1086605_comb] ^ p51_literal_1076345[p52_array_index_1086606_comb] ^ p51_arr[p52_addedKey__58_comb[7:0]];
  assign p52_res7__592_comb = p52_array_index_1086693_comb ^ p52_array_index_1086694_comb ^ p52_array_index_1086695_comb ^ p52_array_index_1086696_comb ^ p52_array_index_1086697_comb ^ p52_array_index_1086698_comb ^ p52_array_index_1086699_comb ^ p51_literal_1076358[p52_array_index_1086686_comb] ^ p52_array_index_1086701_comb ^ p51_literal_1076355[p52_array_index_1086687_comb] ^ p51_literal_1076353[p52_array_index_1086688_comb] ^ p51_literal_1076351[p52_array_index_1086689_comb] ^ p51_literal_1076349[p52_array_index_1086690_comb] ^ p51_literal_1076347[p52_array_index_1086691_comb] ^ p51_literal_1076345[p52_array_index_1086692_comb] ^ p51_arr[p51_bit_slice_1086524];
  assign p52_array_index_1086625_comb = p51_literal_1076345[p52_res7__272_comb];
  assign p52_array_index_1086626_comb = p51_literal_1076347[p52_array_index_1086592_comb];
  assign p52_array_index_1086627_comb = p51_literal_1076349[p52_array_index_1086593_comb];
  assign p52_array_index_1086628_comb = p51_literal_1076351[p52_array_index_1086594_comb];
  assign p52_array_index_1086629_comb = p51_literal_1076353[p52_array_index_1086595_comb];
  assign p52_array_index_1086630_comb = p51_literal_1076355[p52_array_index_1086596_comb];
  assign p52_array_index_1086710_comb = p51_literal_1076345[p52_res7__592_comb];
  assign p52_array_index_1086711_comb = p51_literal_1076347[p52_array_index_1086680_comb];
  assign p52_array_index_1086712_comb = p51_literal_1076349[p52_array_index_1086681_comb];
  assign p52_array_index_1086713_comb = p51_literal_1076351[p52_array_index_1086682_comb];
  assign p52_array_index_1086714_comb = p51_literal_1076353[p52_array_index_1086683_comb];
  assign p52_array_index_1086715_comb = p51_literal_1076355[p52_array_index_1086684_comb];
  assign p52_res7__273_comb = p52_array_index_1086625_comb ^ p52_array_index_1086626_comb ^ p52_array_index_1086627_comb ^ p52_array_index_1086628_comb ^ p52_array_index_1086629_comb ^ p52_array_index_1086630_comb ^ p52_array_index_1086597_comb ^ p51_literal_1076358[p52_array_index_1086614_comb] ^ p52_array_index_1086599_comb ^ p51_literal_1076355[p52_array_index_1086616_comb] ^ p51_literal_1076353[p52_array_index_1086601_comb] ^ p51_literal_1076351[p52_array_index_1086602_comb] ^ p51_literal_1076349[p52_array_index_1086603_comb] ^ p51_literal_1076347[p52_array_index_1086604_comb] ^ p51_literal_1076345[p52_array_index_1086605_comb] ^ p52_array_index_1086606_comb;
  assign p52_res7__593_comb = p52_array_index_1086710_comb ^ p52_array_index_1086711_comb ^ p52_array_index_1086712_comb ^ p52_array_index_1086713_comb ^ p52_array_index_1086714_comb ^ p52_array_index_1086715_comb ^ p52_array_index_1086685_comb ^ p51_literal_1076358[p52_array_index_1086699_comb] ^ p52_array_index_1086686_comb ^ p51_literal_1076355[p52_array_index_1086701_comb] ^ p51_literal_1076353[p52_array_index_1086687_comb] ^ p51_literal_1076351[p52_array_index_1086688_comb] ^ p51_literal_1076349[p52_array_index_1086689_comb] ^ p51_literal_1076347[p52_array_index_1086690_comb] ^ p51_literal_1076345[p52_array_index_1086691_comb] ^ p52_array_index_1086692_comb;
  assign p52_array_index_1086640_comb = p51_literal_1076347[p52_res7__272_comb];
  assign p52_array_index_1086641_comb = p51_literal_1076349[p52_array_index_1086592_comb];
  assign p52_array_index_1086642_comb = p51_literal_1076351[p52_array_index_1086593_comb];
  assign p52_array_index_1086643_comb = p51_literal_1076353[p52_array_index_1086594_comb];
  assign p52_array_index_1086644_comb = p51_literal_1076355[p52_array_index_1086595_comb];
  assign p52_array_index_1086725_comb = p51_literal_1076347[p52_res7__592_comb];
  assign p52_array_index_1086726_comb = p51_literal_1076349[p52_array_index_1086680_comb];
  assign p52_array_index_1086727_comb = p51_literal_1076351[p52_array_index_1086681_comb];
  assign p52_array_index_1086728_comb = p51_literal_1076353[p52_array_index_1086682_comb];
  assign p52_array_index_1086729_comb = p51_literal_1076355[p52_array_index_1086683_comb];
  assign p52_res7__274_comb = p51_literal_1076345[p52_res7__273_comb] ^ p52_array_index_1086640_comb ^ p52_array_index_1086641_comb ^ p52_array_index_1086642_comb ^ p52_array_index_1086643_comb ^ p52_array_index_1086644_comb ^ p52_array_index_1086596_comb ^ p51_literal_1076358[p52_array_index_1086597_comb] ^ p52_array_index_1086614_comb ^ p51_literal_1076355[p52_array_index_1086599_comb] ^ p51_literal_1076353[p52_array_index_1086616_comb] ^ p51_literal_1076351[p52_array_index_1086601_comb] ^ p51_literal_1076349[p52_array_index_1086602_comb] ^ p51_literal_1076347[p52_array_index_1086603_comb] ^ p51_literal_1076345[p52_array_index_1086604_comb] ^ p52_array_index_1086605_comb;
  assign p52_res7__594_comb = p51_literal_1076345[p52_res7__593_comb] ^ p52_array_index_1086725_comb ^ p52_array_index_1086726_comb ^ p52_array_index_1086727_comb ^ p52_array_index_1086728_comb ^ p52_array_index_1086729_comb ^ p52_array_index_1086684_comb ^ p51_literal_1076358[p52_array_index_1086685_comb] ^ p52_array_index_1086699_comb ^ p51_literal_1076355[p52_array_index_1086686_comb] ^ p51_literal_1076353[p52_array_index_1086701_comb] ^ p51_literal_1076351[p52_array_index_1086687_comb] ^ p51_literal_1076349[p52_array_index_1086688_comb] ^ p51_literal_1076347[p52_array_index_1086689_comb] ^ p51_literal_1076345[p52_array_index_1086690_comb] ^ p52_array_index_1086691_comb;
  assign p52_array_index_1086654_comb = p51_literal_1076347[p52_res7__273_comb];
  assign p52_array_index_1086655_comb = p51_literal_1076349[p52_res7__272_comb];
  assign p52_array_index_1086656_comb = p51_literal_1076351[p52_array_index_1086592_comb];
  assign p52_array_index_1086657_comb = p51_literal_1076353[p52_array_index_1086593_comb];
  assign p52_array_index_1086658_comb = p51_literal_1076355[p52_array_index_1086594_comb];
  assign p52_array_index_1086739_comb = p51_literal_1076347[p52_res7__593_comb];
  assign p52_array_index_1086740_comb = p51_literal_1076349[p52_res7__592_comb];
  assign p52_array_index_1086741_comb = p51_literal_1076351[p52_array_index_1086680_comb];
  assign p52_array_index_1086742_comb = p51_literal_1076353[p52_array_index_1086681_comb];
  assign p52_array_index_1086743_comb = p51_literal_1076355[p52_array_index_1086682_comb];
  assign p52_res7__275_comb = p51_literal_1076345[p52_res7__274_comb] ^ p52_array_index_1086654_comb ^ p52_array_index_1086655_comb ^ p52_array_index_1086656_comb ^ p52_array_index_1086657_comb ^ p52_array_index_1086658_comb ^ p52_array_index_1086595_comb ^ p51_literal_1076358[p52_array_index_1086596_comb] ^ p52_array_index_1086597_comb ^ p51_literal_1076355[p52_array_index_1086614_comb] ^ p51_literal_1076353[p52_array_index_1086599_comb] ^ p51_literal_1076351[p52_array_index_1086616_comb] ^ p51_literal_1076349[p52_array_index_1086601_comb] ^ p51_literal_1076347[p52_array_index_1086602_comb] ^ p51_literal_1076345[p52_array_index_1086603_comb] ^ p52_array_index_1086604_comb;
  assign p52_res7__595_comb = p51_literal_1076345[p52_res7__594_comb] ^ p52_array_index_1086739_comb ^ p52_array_index_1086740_comb ^ p52_array_index_1086741_comb ^ p52_array_index_1086742_comb ^ p52_array_index_1086743_comb ^ p52_array_index_1086683_comb ^ p51_literal_1076358[p52_array_index_1086684_comb] ^ p52_array_index_1086685_comb ^ p51_literal_1076355[p52_array_index_1086699_comb] ^ p51_literal_1076353[p52_array_index_1086686_comb] ^ p51_literal_1076351[p52_array_index_1086701_comb] ^ p51_literal_1076349[p52_array_index_1086687_comb] ^ p51_literal_1076347[p52_array_index_1086688_comb] ^ p51_literal_1076345[p52_array_index_1086689_comb] ^ p52_array_index_1086690_comb;
  assign p52_array_index_1086669_comb = p51_literal_1076349[p52_res7__273_comb];
  assign p52_array_index_1086670_comb = p51_literal_1076351[p52_res7__272_comb];
  assign p52_array_index_1086671_comb = p51_literal_1076353[p52_array_index_1086592_comb];
  assign p52_array_index_1086672_comb = p51_literal_1076355[p52_array_index_1086593_comb];
  assign p52_array_index_1086754_comb = p51_literal_1076349[p52_res7__593_comb];
  assign p52_array_index_1086755_comb = p51_literal_1076351[p52_res7__592_comb];
  assign p52_array_index_1086756_comb = p51_literal_1076353[p52_array_index_1086680_comb];
  assign p52_array_index_1086757_comb = p51_literal_1076355[p52_array_index_1086681_comb];
  assign p52_res7__276_comb = p51_literal_1076345[p52_res7__275_comb] ^ p51_literal_1076347[p52_res7__274_comb] ^ p52_array_index_1086669_comb ^ p52_array_index_1086670_comb ^ p52_array_index_1086671_comb ^ p52_array_index_1086672_comb ^ p52_array_index_1086594_comb ^ p51_literal_1076358[p52_array_index_1086595_comb] ^ p52_array_index_1086596_comb ^ p52_array_index_1086613_comb ^ p51_literal_1076353[p52_array_index_1086614_comb] ^ p51_literal_1076351[p52_array_index_1086599_comb] ^ p51_literal_1076349[p52_array_index_1086616_comb] ^ p51_literal_1076347[p52_array_index_1086601_comb] ^ p51_literal_1076345[p52_array_index_1086602_comb] ^ p52_array_index_1086603_comb;
  assign p52_res7__596_comb = p51_literal_1076345[p52_res7__595_comb] ^ p51_literal_1076347[p52_res7__594_comb] ^ p52_array_index_1086754_comb ^ p52_array_index_1086755_comb ^ p52_array_index_1086756_comb ^ p52_array_index_1086757_comb ^ p52_array_index_1086682_comb ^ p51_literal_1076358[p52_array_index_1086683_comb] ^ p52_array_index_1086684_comb ^ p52_array_index_1086698_comb ^ p51_literal_1076353[p52_array_index_1086699_comb] ^ p51_literal_1076351[p52_array_index_1086686_comb] ^ p51_literal_1076349[p52_array_index_1086701_comb] ^ p51_literal_1076347[p52_array_index_1086687_comb] ^ p51_literal_1076345[p52_array_index_1086688_comb] ^ p52_array_index_1086689_comb;

  // Registers for pipe stage 52:
  reg [127:0] p52_k4;
  reg [127:0] p52_xor_1086461;
  reg [7:0] p52_array_index_1086592;
  reg [7:0] p52_array_index_1086593;
  reg [7:0] p52_array_index_1086594;
  reg [7:0] p52_array_index_1086595;
  reg [7:0] p52_array_index_1086596;
  reg [7:0] p52_array_index_1086597;
  reg [7:0] p52_array_index_1086599;
  reg [7:0] p52_array_index_1086601;
  reg [7:0] p52_array_index_1086602;
  reg [7:0] p52_array_index_1086608;
  reg [7:0] p52_array_index_1086609;
  reg [7:0] p52_array_index_1086610;
  reg [7:0] p52_array_index_1086611;
  reg [7:0] p52_array_index_1086612;
  reg [7:0] p52_array_index_1086614;
  reg [7:0] p52_array_index_1086616;
  reg [7:0] p52_res7__272;
  reg [7:0] p52_array_index_1086625;
  reg [7:0] p52_array_index_1086626;
  reg [7:0] p52_array_index_1086627;
  reg [7:0] p52_array_index_1086628;
  reg [7:0] p52_array_index_1086629;
  reg [7:0] p52_array_index_1086630;
  reg [7:0] p52_res7__273;
  reg [7:0] p52_array_index_1086640;
  reg [7:0] p52_array_index_1086641;
  reg [7:0] p52_array_index_1086642;
  reg [7:0] p52_array_index_1086643;
  reg [7:0] p52_array_index_1086644;
  reg [7:0] p52_res7__274;
  reg [7:0] p52_array_index_1086654;
  reg [7:0] p52_array_index_1086655;
  reg [7:0] p52_array_index_1086656;
  reg [7:0] p52_array_index_1086657;
  reg [7:0] p52_array_index_1086658;
  reg [7:0] p52_res7__275;
  reg [7:0] p52_array_index_1086669;
  reg [7:0] p52_array_index_1086670;
  reg [7:0] p52_array_index_1086671;
  reg [7:0] p52_array_index_1086672;
  reg [7:0] p52_res7__276;
  reg [7:0] p52_array_index_1086680;
  reg [7:0] p52_array_index_1086681;
  reg [7:0] p52_array_index_1086682;
  reg [7:0] p52_array_index_1086683;
  reg [7:0] p52_array_index_1086684;
  reg [7:0] p52_array_index_1086685;
  reg [7:0] p52_array_index_1086686;
  reg [7:0] p52_array_index_1086687;
  reg [7:0] p52_array_index_1086688;
  reg [7:0] p52_array_index_1086693;
  reg [7:0] p52_array_index_1086694;
  reg [7:0] p52_array_index_1086695;
  reg [7:0] p52_array_index_1086696;
  reg [7:0] p52_array_index_1086697;
  reg [7:0] p52_array_index_1086699;
  reg [7:0] p52_array_index_1086701;
  reg [7:0] p52_res7__592;
  reg [7:0] p52_array_index_1086710;
  reg [7:0] p52_array_index_1086711;
  reg [7:0] p52_array_index_1086712;
  reg [7:0] p52_array_index_1086713;
  reg [7:0] p52_array_index_1086714;
  reg [7:0] p52_array_index_1086715;
  reg [7:0] p52_res7__593;
  reg [7:0] p52_array_index_1086725;
  reg [7:0] p52_array_index_1086726;
  reg [7:0] p52_array_index_1086727;
  reg [7:0] p52_array_index_1086728;
  reg [7:0] p52_array_index_1086729;
  reg [7:0] p52_res7__594;
  reg [7:0] p52_array_index_1086739;
  reg [7:0] p52_array_index_1086740;
  reg [7:0] p52_array_index_1086741;
  reg [7:0] p52_array_index_1086742;
  reg [7:0] p52_array_index_1086743;
  reg [7:0] p52_res7__595;
  reg [7:0] p52_array_index_1086754;
  reg [7:0] p52_array_index_1086755;
  reg [7:0] p52_array_index_1086756;
  reg [7:0] p52_array_index_1086757;
  reg [7:0] p52_res7__596;
  reg [7:0] p53_arr[256];
  reg [7:0] p53_literal_1076345[256];
  reg [7:0] p53_literal_1076347[256];
  reg [7:0] p53_literal_1076349[256];
  reg [7:0] p53_literal_1076351[256];
  reg [7:0] p53_literal_1076353[256];
  reg [7:0] p53_literal_1076355[256];
  reg [7:0] p53_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p52_k4 <= p51_k4;
    p52_xor_1086461 <= p51_xor_1086461;
    p52_array_index_1086592 <= p52_array_index_1086592_comb;
    p52_array_index_1086593 <= p52_array_index_1086593_comb;
    p52_array_index_1086594 <= p52_array_index_1086594_comb;
    p52_array_index_1086595 <= p52_array_index_1086595_comb;
    p52_array_index_1086596 <= p52_array_index_1086596_comb;
    p52_array_index_1086597 <= p52_array_index_1086597_comb;
    p52_array_index_1086599 <= p52_array_index_1086599_comb;
    p52_array_index_1086601 <= p52_array_index_1086601_comb;
    p52_array_index_1086602 <= p52_array_index_1086602_comb;
    p52_array_index_1086608 <= p52_array_index_1086608_comb;
    p52_array_index_1086609 <= p52_array_index_1086609_comb;
    p52_array_index_1086610 <= p52_array_index_1086610_comb;
    p52_array_index_1086611 <= p52_array_index_1086611_comb;
    p52_array_index_1086612 <= p52_array_index_1086612_comb;
    p52_array_index_1086614 <= p52_array_index_1086614_comb;
    p52_array_index_1086616 <= p52_array_index_1086616_comb;
    p52_res7__272 <= p52_res7__272_comb;
    p52_array_index_1086625 <= p52_array_index_1086625_comb;
    p52_array_index_1086626 <= p52_array_index_1086626_comb;
    p52_array_index_1086627 <= p52_array_index_1086627_comb;
    p52_array_index_1086628 <= p52_array_index_1086628_comb;
    p52_array_index_1086629 <= p52_array_index_1086629_comb;
    p52_array_index_1086630 <= p52_array_index_1086630_comb;
    p52_res7__273 <= p52_res7__273_comb;
    p52_array_index_1086640 <= p52_array_index_1086640_comb;
    p52_array_index_1086641 <= p52_array_index_1086641_comb;
    p52_array_index_1086642 <= p52_array_index_1086642_comb;
    p52_array_index_1086643 <= p52_array_index_1086643_comb;
    p52_array_index_1086644 <= p52_array_index_1086644_comb;
    p52_res7__274 <= p52_res7__274_comb;
    p52_array_index_1086654 <= p52_array_index_1086654_comb;
    p52_array_index_1086655 <= p52_array_index_1086655_comb;
    p52_array_index_1086656 <= p52_array_index_1086656_comb;
    p52_array_index_1086657 <= p52_array_index_1086657_comb;
    p52_array_index_1086658 <= p52_array_index_1086658_comb;
    p52_res7__275 <= p52_res7__275_comb;
    p52_array_index_1086669 <= p52_array_index_1086669_comb;
    p52_array_index_1086670 <= p52_array_index_1086670_comb;
    p52_array_index_1086671 <= p52_array_index_1086671_comb;
    p52_array_index_1086672 <= p52_array_index_1086672_comb;
    p52_res7__276 <= p52_res7__276_comb;
    p52_array_index_1086680 <= p52_array_index_1086680_comb;
    p52_array_index_1086681 <= p52_array_index_1086681_comb;
    p52_array_index_1086682 <= p52_array_index_1086682_comb;
    p52_array_index_1086683 <= p52_array_index_1086683_comb;
    p52_array_index_1086684 <= p52_array_index_1086684_comb;
    p52_array_index_1086685 <= p52_array_index_1086685_comb;
    p52_array_index_1086686 <= p52_array_index_1086686_comb;
    p52_array_index_1086687 <= p52_array_index_1086687_comb;
    p52_array_index_1086688 <= p52_array_index_1086688_comb;
    p52_array_index_1086693 <= p52_array_index_1086693_comb;
    p52_array_index_1086694 <= p52_array_index_1086694_comb;
    p52_array_index_1086695 <= p52_array_index_1086695_comb;
    p52_array_index_1086696 <= p52_array_index_1086696_comb;
    p52_array_index_1086697 <= p52_array_index_1086697_comb;
    p52_array_index_1086699 <= p52_array_index_1086699_comb;
    p52_array_index_1086701 <= p52_array_index_1086701_comb;
    p52_res7__592 <= p52_res7__592_comb;
    p52_array_index_1086710 <= p52_array_index_1086710_comb;
    p52_array_index_1086711 <= p52_array_index_1086711_comb;
    p52_array_index_1086712 <= p52_array_index_1086712_comb;
    p52_array_index_1086713 <= p52_array_index_1086713_comb;
    p52_array_index_1086714 <= p52_array_index_1086714_comb;
    p52_array_index_1086715 <= p52_array_index_1086715_comb;
    p52_res7__593 <= p52_res7__593_comb;
    p52_array_index_1086725 <= p52_array_index_1086725_comb;
    p52_array_index_1086726 <= p52_array_index_1086726_comb;
    p52_array_index_1086727 <= p52_array_index_1086727_comb;
    p52_array_index_1086728 <= p52_array_index_1086728_comb;
    p52_array_index_1086729 <= p52_array_index_1086729_comb;
    p52_res7__594 <= p52_res7__594_comb;
    p52_array_index_1086739 <= p52_array_index_1086739_comb;
    p52_array_index_1086740 <= p52_array_index_1086740_comb;
    p52_array_index_1086741 <= p52_array_index_1086741_comb;
    p52_array_index_1086742 <= p52_array_index_1086742_comb;
    p52_array_index_1086743 <= p52_array_index_1086743_comb;
    p52_res7__595 <= p52_res7__595_comb;
    p52_array_index_1086754 <= p52_array_index_1086754_comb;
    p52_array_index_1086755 <= p52_array_index_1086755_comb;
    p52_array_index_1086756 <= p52_array_index_1086756_comb;
    p52_array_index_1086757 <= p52_array_index_1086757_comb;
    p52_res7__596 <= p52_res7__596_comb;
    p53_arr <= p52_arr;
    p53_literal_1076345 <= p52_literal_1076345;
    p53_literal_1076347 <= p52_literal_1076347;
    p53_literal_1076349 <= p52_literal_1076349;
    p53_literal_1076351 <= p52_literal_1076351;
    p53_literal_1076353 <= p52_literal_1076353;
    p53_literal_1076355 <= p52_literal_1076355;
    p53_literal_1076358 <= p52_literal_1076358;
  end

  // ===== Pipe stage 53:
  wire [7:0] p53_array_index_1086951_comb;
  wire [7:0] p53_array_index_1086952_comb;
  wire [7:0] p53_array_index_1086953_comb;
  wire [7:0] p53_array_index_1086954_comb;
  wire [7:0] p53_res7__277_comb;
  wire [7:0] p53_array_index_1087019_comb;
  wire [7:0] p53_array_index_1087020_comb;
  wire [7:0] p53_array_index_1087021_comb;
  wire [7:0] p53_array_index_1087022_comb;
  wire [7:0] p53_array_index_1086965_comb;
  wire [7:0] p53_array_index_1086966_comb;
  wire [7:0] p53_array_index_1086967_comb;
  wire [7:0] p53_res7__597_comb;
  wire [7:0] p53_res7__278_comb;
  wire [7:0] p53_array_index_1087033_comb;
  wire [7:0] p53_array_index_1087034_comb;
  wire [7:0] p53_array_index_1087035_comb;
  wire [7:0] p53_array_index_1086977_comb;
  wire [7:0] p53_array_index_1086978_comb;
  wire [7:0] p53_array_index_1086979_comb;
  wire [7:0] p53_res7__598_comb;
  wire [7:0] p53_res7__279_comb;
  wire [7:0] p53_array_index_1087045_comb;
  wire [7:0] p53_array_index_1087046_comb;
  wire [7:0] p53_array_index_1087047_comb;
  wire [7:0] p53_array_index_1086990_comb;
  wire [7:0] p53_array_index_1086991_comb;
  wire [7:0] p53_res7__599_comb;
  wire [7:0] p53_res7__280_comb;
  wire [7:0] p53_array_index_1087058_comb;
  wire [7:0] p53_array_index_1087059_comb;
  wire [7:0] p53_array_index_1087001_comb;
  wire [7:0] p53_array_index_1087002_comb;
  wire [7:0] p53_res7__600_comb;
  wire [7:0] p53_res7__281_comb;
  wire [7:0] p53_array_index_1087069_comb;
  wire [7:0] p53_array_index_1087070_comb;
  wire [7:0] p53_array_index_1087008_comb;
  wire [7:0] p53_array_index_1087009_comb;
  wire [7:0] p53_array_index_1087010_comb;
  wire [7:0] p53_array_index_1087011_comb;
  wire [7:0] p53_array_index_1087012_comb;
  wire [7:0] p53_array_index_1087013_comb;
  wire [7:0] p53_array_index_1087014_comb;
  wire [7:0] p53_array_index_1087015_comb;
  wire [7:0] p53_array_index_1087016_comb;
  wire [7:0] p53_res7__601_comb;
  assign p53_array_index_1086951_comb = p52_literal_1076349[p52_res7__274];
  assign p53_array_index_1086952_comb = p52_literal_1076351[p52_res7__273];
  assign p53_array_index_1086953_comb = p52_literal_1076353[p52_res7__272];
  assign p53_array_index_1086954_comb = p52_literal_1076355[p52_array_index_1086592];
  assign p53_res7__277_comb = p52_literal_1076345[p52_res7__276] ^ p52_literal_1076347[p52_res7__275] ^ p53_array_index_1086951_comb ^ p53_array_index_1086952_comb ^ p53_array_index_1086953_comb ^ p53_array_index_1086954_comb ^ p52_array_index_1086593 ^ p52_literal_1076358[p52_array_index_1086594] ^ p52_array_index_1086595 ^ p52_array_index_1086630 ^ p52_literal_1076353[p52_array_index_1086597] ^ p52_literal_1076351[p52_array_index_1086614] ^ p52_literal_1076349[p52_array_index_1086599] ^ p52_literal_1076347[p52_array_index_1086616] ^ p52_literal_1076345[p52_array_index_1086601] ^ p52_array_index_1086602;
  assign p53_array_index_1087019_comb = p52_literal_1076349[p52_res7__594];
  assign p53_array_index_1087020_comb = p52_literal_1076351[p52_res7__593];
  assign p53_array_index_1087021_comb = p52_literal_1076353[p52_res7__592];
  assign p53_array_index_1087022_comb = p52_literal_1076355[p52_array_index_1086680];
  assign p53_array_index_1086965_comb = p52_literal_1076351[p52_res7__274];
  assign p53_array_index_1086966_comb = p52_literal_1076353[p52_res7__273];
  assign p53_array_index_1086967_comb = p52_literal_1076355[p52_res7__272];
  assign p53_res7__597_comb = p52_literal_1076345[p52_res7__596] ^ p52_literal_1076347[p52_res7__595] ^ p53_array_index_1087019_comb ^ p53_array_index_1087020_comb ^ p53_array_index_1087021_comb ^ p53_array_index_1087022_comb ^ p52_array_index_1086681 ^ p52_literal_1076358[p52_array_index_1086682] ^ p52_array_index_1086683 ^ p52_array_index_1086715 ^ p52_literal_1076353[p52_array_index_1086685] ^ p52_literal_1076351[p52_array_index_1086699] ^ p52_literal_1076349[p52_array_index_1086686] ^ p52_literal_1076347[p52_array_index_1086701] ^ p52_literal_1076345[p52_array_index_1086687] ^ p52_array_index_1086688;
  assign p53_res7__278_comb = p52_literal_1076345[p53_res7__277_comb] ^ p52_literal_1076347[p52_res7__276] ^ p52_literal_1076349[p52_res7__275] ^ p53_array_index_1086965_comb ^ p53_array_index_1086966_comb ^ p53_array_index_1086967_comb ^ p52_array_index_1086592 ^ p52_literal_1076358[p52_array_index_1086593] ^ p52_array_index_1086594 ^ p52_array_index_1086644 ^ p52_array_index_1086612 ^ p52_literal_1076351[p52_array_index_1086597] ^ p52_literal_1076349[p52_array_index_1086614] ^ p52_literal_1076347[p52_array_index_1086599] ^ p52_literal_1076345[p52_array_index_1086616] ^ p52_array_index_1086601;
  assign p53_array_index_1087033_comb = p52_literal_1076351[p52_res7__594];
  assign p53_array_index_1087034_comb = p52_literal_1076353[p52_res7__593];
  assign p53_array_index_1087035_comb = p52_literal_1076355[p52_res7__592];
  assign p53_array_index_1086977_comb = p52_literal_1076351[p52_res7__275];
  assign p53_array_index_1086978_comb = p52_literal_1076353[p52_res7__274];
  assign p53_array_index_1086979_comb = p52_literal_1076355[p52_res7__273];
  assign p53_res7__598_comb = p52_literal_1076345[p53_res7__597_comb] ^ p52_literal_1076347[p52_res7__596] ^ p52_literal_1076349[p52_res7__595] ^ p53_array_index_1087033_comb ^ p53_array_index_1087034_comb ^ p53_array_index_1087035_comb ^ p52_array_index_1086680 ^ p52_literal_1076358[p52_array_index_1086681] ^ p52_array_index_1086682 ^ p52_array_index_1086729 ^ p52_array_index_1086697 ^ p52_literal_1076351[p52_array_index_1086685] ^ p52_literal_1076349[p52_array_index_1086699] ^ p52_literal_1076347[p52_array_index_1086686] ^ p52_literal_1076345[p52_array_index_1086701] ^ p52_array_index_1086687;
  assign p53_res7__279_comb = p52_literal_1076345[p53_res7__278_comb] ^ p52_literal_1076347[p53_res7__277_comb] ^ p52_literal_1076349[p52_res7__276] ^ p53_array_index_1086977_comb ^ p53_array_index_1086978_comb ^ p53_array_index_1086979_comb ^ p52_res7__272 ^ p52_literal_1076358[p52_array_index_1086592] ^ p52_array_index_1086593 ^ p52_array_index_1086658 ^ p52_array_index_1086629 ^ p52_literal_1076351[p52_array_index_1086596] ^ p52_literal_1076349[p52_array_index_1086597] ^ p52_literal_1076347[p52_array_index_1086614] ^ p52_literal_1076345[p52_array_index_1086599] ^ p52_array_index_1086616;
  assign p53_array_index_1087045_comb = p52_literal_1076351[p52_res7__595];
  assign p53_array_index_1087046_comb = p52_literal_1076353[p52_res7__594];
  assign p53_array_index_1087047_comb = p52_literal_1076355[p52_res7__593];
  assign p53_array_index_1086990_comb = p52_literal_1076353[p52_res7__275];
  assign p53_array_index_1086991_comb = p52_literal_1076355[p52_res7__274];
  assign p53_res7__599_comb = p52_literal_1076345[p53_res7__598_comb] ^ p52_literal_1076347[p53_res7__597_comb] ^ p52_literal_1076349[p52_res7__596] ^ p53_array_index_1087045_comb ^ p53_array_index_1087046_comb ^ p53_array_index_1087047_comb ^ p52_res7__592 ^ p52_literal_1076358[p52_array_index_1086680] ^ p52_array_index_1086681 ^ p52_array_index_1086743 ^ p52_array_index_1086714 ^ p52_literal_1076351[p52_array_index_1086684] ^ p52_literal_1076349[p52_array_index_1086685] ^ p52_literal_1076347[p52_array_index_1086699] ^ p52_literal_1076345[p52_array_index_1086686] ^ p52_array_index_1086701;
  assign p53_res7__280_comb = p52_literal_1076345[p53_res7__279_comb] ^ p52_literal_1076347[p53_res7__278_comb] ^ p52_literal_1076349[p53_res7__277_comb] ^ p52_literal_1076351[p52_res7__276] ^ p53_array_index_1086990_comb ^ p53_array_index_1086991_comb ^ p52_res7__273 ^ p52_literal_1076358[p52_res7__272] ^ p52_array_index_1086592 ^ p52_array_index_1086672 ^ p52_array_index_1086643 ^ p52_array_index_1086611 ^ p52_literal_1076349[p52_array_index_1086596] ^ p52_literal_1076347[p52_array_index_1086597] ^ p52_literal_1076345[p52_array_index_1086614] ^ p52_array_index_1086599;
  assign p53_array_index_1087058_comb = p52_literal_1076353[p52_res7__595];
  assign p53_array_index_1087059_comb = p52_literal_1076355[p52_res7__594];
  assign p53_array_index_1087001_comb = p52_literal_1076353[p52_res7__276];
  assign p53_array_index_1087002_comb = p52_literal_1076355[p52_res7__275];
  assign p53_res7__600_comb = p52_literal_1076345[p53_res7__599_comb] ^ p52_literal_1076347[p53_res7__598_comb] ^ p52_literal_1076349[p53_res7__597_comb] ^ p52_literal_1076351[p52_res7__596] ^ p53_array_index_1087058_comb ^ p53_array_index_1087059_comb ^ p52_res7__593 ^ p52_literal_1076358[p52_res7__592] ^ p52_array_index_1086680 ^ p52_array_index_1086757 ^ p52_array_index_1086728 ^ p52_array_index_1086696 ^ p52_literal_1076349[p52_array_index_1086684] ^ p52_literal_1076347[p52_array_index_1086685] ^ p52_literal_1076345[p52_array_index_1086699] ^ p52_array_index_1086686;
  assign p53_res7__281_comb = p52_literal_1076345[p53_res7__280_comb] ^ p52_literal_1076347[p53_res7__279_comb] ^ p52_literal_1076349[p53_res7__278_comb] ^ p52_literal_1076351[p53_res7__277_comb] ^ p53_array_index_1087001_comb ^ p53_array_index_1087002_comb ^ p52_res7__274 ^ p52_literal_1076358[p52_res7__273] ^ p52_res7__272 ^ p53_array_index_1086954_comb ^ p52_array_index_1086657 ^ p52_array_index_1086628 ^ p52_literal_1076349[p52_array_index_1086595] ^ p52_literal_1076347[p52_array_index_1086596] ^ p52_literal_1076345[p52_array_index_1086597] ^ p52_array_index_1086614;
  assign p53_array_index_1087069_comb = p52_literal_1076353[p52_res7__596];
  assign p53_array_index_1087070_comb = p52_literal_1076355[p52_res7__595];
  assign p53_array_index_1087008_comb = p52_literal_1076345[p53_res7__281_comb];
  assign p53_array_index_1087009_comb = p52_literal_1076347[p53_res7__280_comb];
  assign p53_array_index_1087010_comb = p52_literal_1076349[p53_res7__279_comb];
  assign p53_array_index_1087011_comb = p52_literal_1076351[p53_res7__278_comb];
  assign p53_array_index_1087012_comb = p52_literal_1076353[p53_res7__277_comb];
  assign p53_array_index_1087013_comb = p52_literal_1076355[p52_res7__276];
  assign p53_array_index_1087014_comb = p52_literal_1076358[p52_res7__274];
  assign p53_array_index_1087015_comb = p52_literal_1076347[p52_array_index_1086595];
  assign p53_array_index_1087016_comb = p52_literal_1076345[p52_array_index_1086596];
  assign p53_res7__601_comb = p52_literal_1076345[p53_res7__600_comb] ^ p52_literal_1076347[p53_res7__599_comb] ^ p52_literal_1076349[p53_res7__598_comb] ^ p52_literal_1076351[p53_res7__597_comb] ^ p53_array_index_1087069_comb ^ p53_array_index_1087070_comb ^ p52_res7__594 ^ p52_literal_1076358[p52_res7__593] ^ p52_res7__592 ^ p53_array_index_1087022_comb ^ p52_array_index_1086742 ^ p52_array_index_1086713 ^ p52_literal_1076349[p52_array_index_1086683] ^ p52_literal_1076347[p52_array_index_1086684] ^ p52_literal_1076345[p52_array_index_1086685] ^ p52_array_index_1086699;

  // Registers for pipe stage 53:
  reg [127:0] p53_k4;
  reg [127:0] p53_xor_1086461;
  reg [7:0] p53_array_index_1086592;
  reg [7:0] p53_array_index_1086593;
  reg [7:0] p53_array_index_1086594;
  reg [7:0] p53_array_index_1086595;
  reg [7:0] p53_array_index_1086596;
  reg [7:0] p53_array_index_1086597;
  reg [7:0] p53_array_index_1086608;
  reg [7:0] p53_array_index_1086609;
  reg [7:0] p53_array_index_1086610;
  reg [7:0] p53_res7__272;
  reg [7:0] p53_array_index_1086625;
  reg [7:0] p53_array_index_1086626;
  reg [7:0] p53_array_index_1086627;
  reg [7:0] p53_res7__273;
  reg [7:0] p53_array_index_1086640;
  reg [7:0] p53_array_index_1086641;
  reg [7:0] p53_array_index_1086642;
  reg [7:0] p53_res7__274;
  reg [7:0] p53_array_index_1086654;
  reg [7:0] p53_array_index_1086655;
  reg [7:0] p53_array_index_1086656;
  reg [7:0] p53_res7__275;
  reg [7:0] p53_array_index_1086669;
  reg [7:0] p53_array_index_1086670;
  reg [7:0] p53_array_index_1086671;
  reg [7:0] p53_res7__276;
  reg [7:0] p53_array_index_1086951;
  reg [7:0] p53_array_index_1086952;
  reg [7:0] p53_array_index_1086953;
  reg [7:0] p53_res7__277;
  reg [7:0] p53_array_index_1086965;
  reg [7:0] p53_array_index_1086966;
  reg [7:0] p53_array_index_1086967;
  reg [7:0] p53_res7__278;
  reg [7:0] p53_array_index_1086977;
  reg [7:0] p53_array_index_1086978;
  reg [7:0] p53_array_index_1086979;
  reg [7:0] p53_res7__279;
  reg [7:0] p53_array_index_1086990;
  reg [7:0] p53_array_index_1086991;
  reg [7:0] p53_res7__280;
  reg [7:0] p53_array_index_1087001;
  reg [7:0] p53_array_index_1087002;
  reg [7:0] p53_res7__281;
  reg [7:0] p53_array_index_1087008;
  reg [7:0] p53_array_index_1087009;
  reg [7:0] p53_array_index_1087010;
  reg [7:0] p53_array_index_1087011;
  reg [7:0] p53_array_index_1087012;
  reg [7:0] p53_array_index_1087013;
  reg [7:0] p53_array_index_1087014;
  reg [7:0] p53_array_index_1087015;
  reg [7:0] p53_array_index_1087016;
  reg [7:0] p53_array_index_1086680;
  reg [7:0] p53_array_index_1086681;
  reg [7:0] p53_array_index_1086682;
  reg [7:0] p53_array_index_1086683;
  reg [7:0] p53_array_index_1086684;
  reg [7:0] p53_array_index_1086685;
  reg [7:0] p53_array_index_1086693;
  reg [7:0] p53_array_index_1086694;
  reg [7:0] p53_array_index_1086695;
  reg [7:0] p53_res7__592;
  reg [7:0] p53_array_index_1086710;
  reg [7:0] p53_array_index_1086711;
  reg [7:0] p53_array_index_1086712;
  reg [7:0] p53_res7__593;
  reg [7:0] p53_array_index_1086725;
  reg [7:0] p53_array_index_1086726;
  reg [7:0] p53_array_index_1086727;
  reg [7:0] p53_res7__594;
  reg [7:0] p53_array_index_1086739;
  reg [7:0] p53_array_index_1086740;
  reg [7:0] p53_array_index_1086741;
  reg [7:0] p53_res7__595;
  reg [7:0] p53_array_index_1086754;
  reg [7:0] p53_array_index_1086755;
  reg [7:0] p53_array_index_1086756;
  reg [7:0] p53_res7__596;
  reg [7:0] p53_array_index_1087019;
  reg [7:0] p53_array_index_1087020;
  reg [7:0] p53_array_index_1087021;
  reg [7:0] p53_res7__597;
  reg [7:0] p53_array_index_1087033;
  reg [7:0] p53_array_index_1087034;
  reg [7:0] p53_array_index_1087035;
  reg [7:0] p53_res7__598;
  reg [7:0] p53_array_index_1087045;
  reg [7:0] p53_array_index_1087046;
  reg [7:0] p53_array_index_1087047;
  reg [7:0] p53_res7__599;
  reg [7:0] p53_array_index_1087058;
  reg [7:0] p53_array_index_1087059;
  reg [7:0] p53_res7__600;
  reg [7:0] p53_array_index_1087069;
  reg [7:0] p53_array_index_1087070;
  reg [7:0] p53_res7__601;
  reg [7:0] p54_arr[256];
  reg [7:0] p54_literal_1076345[256];
  reg [7:0] p54_literal_1076347[256];
  reg [7:0] p54_literal_1076349[256];
  reg [7:0] p54_literal_1076351[256];
  reg [7:0] p54_literal_1076353[256];
  reg [7:0] p54_literal_1076355[256];
  reg [7:0] p54_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p53_k4 <= p52_k4;
    p53_xor_1086461 <= p52_xor_1086461;
    p53_array_index_1086592 <= p52_array_index_1086592;
    p53_array_index_1086593 <= p52_array_index_1086593;
    p53_array_index_1086594 <= p52_array_index_1086594;
    p53_array_index_1086595 <= p52_array_index_1086595;
    p53_array_index_1086596 <= p52_array_index_1086596;
    p53_array_index_1086597 <= p52_array_index_1086597;
    p53_array_index_1086608 <= p52_array_index_1086608;
    p53_array_index_1086609 <= p52_array_index_1086609;
    p53_array_index_1086610 <= p52_array_index_1086610;
    p53_res7__272 <= p52_res7__272;
    p53_array_index_1086625 <= p52_array_index_1086625;
    p53_array_index_1086626 <= p52_array_index_1086626;
    p53_array_index_1086627 <= p52_array_index_1086627;
    p53_res7__273 <= p52_res7__273;
    p53_array_index_1086640 <= p52_array_index_1086640;
    p53_array_index_1086641 <= p52_array_index_1086641;
    p53_array_index_1086642 <= p52_array_index_1086642;
    p53_res7__274 <= p52_res7__274;
    p53_array_index_1086654 <= p52_array_index_1086654;
    p53_array_index_1086655 <= p52_array_index_1086655;
    p53_array_index_1086656 <= p52_array_index_1086656;
    p53_res7__275 <= p52_res7__275;
    p53_array_index_1086669 <= p52_array_index_1086669;
    p53_array_index_1086670 <= p52_array_index_1086670;
    p53_array_index_1086671 <= p52_array_index_1086671;
    p53_res7__276 <= p52_res7__276;
    p53_array_index_1086951 <= p53_array_index_1086951_comb;
    p53_array_index_1086952 <= p53_array_index_1086952_comb;
    p53_array_index_1086953 <= p53_array_index_1086953_comb;
    p53_res7__277 <= p53_res7__277_comb;
    p53_array_index_1086965 <= p53_array_index_1086965_comb;
    p53_array_index_1086966 <= p53_array_index_1086966_comb;
    p53_array_index_1086967 <= p53_array_index_1086967_comb;
    p53_res7__278 <= p53_res7__278_comb;
    p53_array_index_1086977 <= p53_array_index_1086977_comb;
    p53_array_index_1086978 <= p53_array_index_1086978_comb;
    p53_array_index_1086979 <= p53_array_index_1086979_comb;
    p53_res7__279 <= p53_res7__279_comb;
    p53_array_index_1086990 <= p53_array_index_1086990_comb;
    p53_array_index_1086991 <= p53_array_index_1086991_comb;
    p53_res7__280 <= p53_res7__280_comb;
    p53_array_index_1087001 <= p53_array_index_1087001_comb;
    p53_array_index_1087002 <= p53_array_index_1087002_comb;
    p53_res7__281 <= p53_res7__281_comb;
    p53_array_index_1087008 <= p53_array_index_1087008_comb;
    p53_array_index_1087009 <= p53_array_index_1087009_comb;
    p53_array_index_1087010 <= p53_array_index_1087010_comb;
    p53_array_index_1087011 <= p53_array_index_1087011_comb;
    p53_array_index_1087012 <= p53_array_index_1087012_comb;
    p53_array_index_1087013 <= p53_array_index_1087013_comb;
    p53_array_index_1087014 <= p53_array_index_1087014_comb;
    p53_array_index_1087015 <= p53_array_index_1087015_comb;
    p53_array_index_1087016 <= p53_array_index_1087016_comb;
    p53_array_index_1086680 <= p52_array_index_1086680;
    p53_array_index_1086681 <= p52_array_index_1086681;
    p53_array_index_1086682 <= p52_array_index_1086682;
    p53_array_index_1086683 <= p52_array_index_1086683;
    p53_array_index_1086684 <= p52_array_index_1086684;
    p53_array_index_1086685 <= p52_array_index_1086685;
    p53_array_index_1086693 <= p52_array_index_1086693;
    p53_array_index_1086694 <= p52_array_index_1086694;
    p53_array_index_1086695 <= p52_array_index_1086695;
    p53_res7__592 <= p52_res7__592;
    p53_array_index_1086710 <= p52_array_index_1086710;
    p53_array_index_1086711 <= p52_array_index_1086711;
    p53_array_index_1086712 <= p52_array_index_1086712;
    p53_res7__593 <= p52_res7__593;
    p53_array_index_1086725 <= p52_array_index_1086725;
    p53_array_index_1086726 <= p52_array_index_1086726;
    p53_array_index_1086727 <= p52_array_index_1086727;
    p53_res7__594 <= p52_res7__594;
    p53_array_index_1086739 <= p52_array_index_1086739;
    p53_array_index_1086740 <= p52_array_index_1086740;
    p53_array_index_1086741 <= p52_array_index_1086741;
    p53_res7__595 <= p52_res7__595;
    p53_array_index_1086754 <= p52_array_index_1086754;
    p53_array_index_1086755 <= p52_array_index_1086755;
    p53_array_index_1086756 <= p52_array_index_1086756;
    p53_res7__596 <= p52_res7__596;
    p53_array_index_1087019 <= p53_array_index_1087019_comb;
    p53_array_index_1087020 <= p53_array_index_1087020_comb;
    p53_array_index_1087021 <= p53_array_index_1087021_comb;
    p53_res7__597 <= p53_res7__597_comb;
    p53_array_index_1087033 <= p53_array_index_1087033_comb;
    p53_array_index_1087034 <= p53_array_index_1087034_comb;
    p53_array_index_1087035 <= p53_array_index_1087035_comb;
    p53_res7__598 <= p53_res7__598_comb;
    p53_array_index_1087045 <= p53_array_index_1087045_comb;
    p53_array_index_1087046 <= p53_array_index_1087046_comb;
    p53_array_index_1087047 <= p53_array_index_1087047_comb;
    p53_res7__599 <= p53_res7__599_comb;
    p53_array_index_1087058 <= p53_array_index_1087058_comb;
    p53_array_index_1087059 <= p53_array_index_1087059_comb;
    p53_res7__600 <= p53_res7__600_comb;
    p53_array_index_1087069 <= p53_array_index_1087069_comb;
    p53_array_index_1087070 <= p53_array_index_1087070_comb;
    p53_res7__601 <= p53_res7__601_comb;
    p54_arr <= p53_arr;
    p54_literal_1076345 <= p53_literal_1076345;
    p54_literal_1076347 <= p53_literal_1076347;
    p54_literal_1076349 <= p53_literal_1076349;
    p54_literal_1076351 <= p53_literal_1076351;
    p54_literal_1076353 <= p53_literal_1076353;
    p54_literal_1076355 <= p53_literal_1076355;
    p54_literal_1076358 <= p53_literal_1076358;
  end

  // ===== Pipe stage 54:
  wire [7:0] p54_res7__282_comb;
  wire [7:0] p54_array_index_1087296_comb;
  wire [7:0] p54_res7__283_comb;
  wire [7:0] p54_array_index_1087342_comb;
  wire [7:0] p54_res7__284_comb;
  wire [7:0] p54_res7__602_comb;
  wire [7:0] p54_array_index_1087352_comb;
  wire [7:0] p54_res7__285_comb;
  wire [7:0] p54_res7__603_comb;
  wire [7:0] p54_res7__286_comb;
  wire [7:0] p54_res7__604_comb;
  wire [7:0] p54_res7__287_comb;
  wire [7:0] p54_res7__605_comb;
  wire [127:0] p54_res__17_comb;
  wire [127:0] p54_xor_1087336_comb;
  wire [7:0] p54_res7__606_comb;
  assign p54_res7__282_comb = p53_array_index_1087008 ^ p53_array_index_1087009 ^ p53_array_index_1087010 ^ p53_array_index_1087011 ^ p53_array_index_1087012 ^ p53_array_index_1087013 ^ p53_res7__275 ^ p53_array_index_1087014 ^ p53_res7__273 ^ p53_array_index_1086967 ^ p53_array_index_1086671 ^ p53_array_index_1086642 ^ p53_array_index_1086610 ^ p53_array_index_1087015 ^ p53_array_index_1087016 ^ p53_array_index_1086597;
  assign p54_array_index_1087296_comb = p53_literal_1076355[p53_res7__277];
  assign p54_res7__283_comb = p53_literal_1076345[p54_res7__282_comb] ^ p53_literal_1076347[p53_res7__281] ^ p53_literal_1076349[p53_res7__280] ^ p53_literal_1076351[p53_res7__279] ^ p53_literal_1076353[p53_res7__278] ^ p54_array_index_1087296_comb ^ p53_res7__276 ^ p53_literal_1076358[p53_res7__275] ^ p53_res7__274 ^ p53_array_index_1086979 ^ p53_array_index_1086953 ^ p53_array_index_1086656 ^ p53_array_index_1086627 ^ p53_literal_1076347[p53_array_index_1086594] ^ p53_literal_1076345[p53_array_index_1086595] ^ p53_array_index_1086596;
  assign p54_array_index_1087342_comb = p53_literal_1076355[p53_res7__596];
  assign p54_res7__284_comb = p53_literal_1076345[p54_res7__283_comb] ^ p53_literal_1076347[p54_res7__282_comb] ^ p53_literal_1076349[p53_res7__281] ^ p53_literal_1076351[p53_res7__280] ^ p53_literal_1076353[p53_res7__279] ^ p53_literal_1076355[p53_res7__278] ^ p53_res7__277 ^ p53_literal_1076358[p53_res7__276] ^ p53_res7__275 ^ p53_array_index_1086991 ^ p53_array_index_1086966 ^ p53_array_index_1086670 ^ p53_array_index_1086641 ^ p53_array_index_1086609 ^ p53_literal_1076345[p53_array_index_1086594] ^ p53_array_index_1086595;
  assign p54_res7__602_comb = p53_literal_1076345[p53_res7__601] ^ p53_literal_1076347[p53_res7__600] ^ p53_literal_1076349[p53_res7__599] ^ p53_literal_1076351[p53_res7__598] ^ p53_literal_1076353[p53_res7__597] ^ p54_array_index_1087342_comb ^ p53_res7__595 ^ p53_literal_1076358[p53_res7__594] ^ p53_res7__593 ^ p53_array_index_1087035 ^ p53_array_index_1086756 ^ p53_array_index_1086727 ^ p53_array_index_1086695 ^ p53_literal_1076347[p53_array_index_1086683] ^ p53_literal_1076345[p53_array_index_1086684] ^ p53_array_index_1086685;
  assign p54_array_index_1087352_comb = p53_literal_1076355[p53_res7__597];
  assign p54_res7__285_comb = p53_literal_1076345[p54_res7__284_comb] ^ p53_literal_1076347[p54_res7__283_comb] ^ p53_literal_1076349[p54_res7__282_comb] ^ p53_literal_1076351[p53_res7__281] ^ p53_literal_1076353[p53_res7__280] ^ p53_literal_1076355[p53_res7__279] ^ p53_res7__278 ^ p53_literal_1076358[p53_res7__277] ^ p53_res7__276 ^ p53_array_index_1087002 ^ p53_array_index_1086978 ^ p53_array_index_1086952 ^ p53_array_index_1086655 ^ p53_array_index_1086626 ^ p53_literal_1076345[p53_array_index_1086593] ^ p53_array_index_1086594;
  assign p54_res7__603_comb = p53_literal_1076345[p54_res7__602_comb] ^ p53_literal_1076347[p53_res7__601] ^ p53_literal_1076349[p53_res7__600] ^ p53_literal_1076351[p53_res7__599] ^ p53_literal_1076353[p53_res7__598] ^ p54_array_index_1087352_comb ^ p53_res7__596 ^ p53_literal_1076358[p53_res7__595] ^ p53_res7__594 ^ p53_array_index_1087047 ^ p53_array_index_1087021 ^ p53_array_index_1086741 ^ p53_array_index_1086712 ^ p53_literal_1076347[p53_array_index_1086682] ^ p53_literal_1076345[p53_array_index_1086683] ^ p53_array_index_1086684;
  assign p54_res7__286_comb = p53_literal_1076345[p54_res7__285_comb] ^ p53_literal_1076347[p54_res7__284_comb] ^ p53_literal_1076349[p54_res7__283_comb] ^ p53_literal_1076351[p54_res7__282_comb] ^ p53_literal_1076353[p53_res7__281] ^ p53_literal_1076355[p53_res7__280] ^ p53_res7__279 ^ p53_literal_1076358[p53_res7__278] ^ p53_res7__277 ^ p53_array_index_1087013 ^ p53_array_index_1086990 ^ p53_array_index_1086965 ^ p53_array_index_1086669 ^ p53_array_index_1086640 ^ p53_array_index_1086608 ^ p53_array_index_1086593;
  assign p54_res7__604_comb = p53_literal_1076345[p54_res7__603_comb] ^ p53_literal_1076347[p54_res7__602_comb] ^ p53_literal_1076349[p53_res7__601] ^ p53_literal_1076351[p53_res7__600] ^ p53_literal_1076353[p53_res7__599] ^ p53_literal_1076355[p53_res7__598] ^ p53_res7__597 ^ p53_literal_1076358[p53_res7__596] ^ p53_res7__595 ^ p53_array_index_1087059 ^ p53_array_index_1087034 ^ p53_array_index_1086755 ^ p53_array_index_1086726 ^ p53_array_index_1086694 ^ p53_literal_1076345[p53_array_index_1086682] ^ p53_array_index_1086683;
  assign p54_res7__287_comb = p53_literal_1076345[p54_res7__286_comb] ^ p53_literal_1076347[p54_res7__285_comb] ^ p53_literal_1076349[p54_res7__284_comb] ^ p53_literal_1076351[p54_res7__283_comb] ^ p53_literal_1076353[p54_res7__282_comb] ^ p53_literal_1076355[p53_res7__281] ^ p53_res7__280 ^ p53_literal_1076358[p53_res7__279] ^ p53_res7__278 ^ p54_array_index_1087296_comb ^ p53_array_index_1087001 ^ p53_array_index_1086977 ^ p53_array_index_1086951 ^ p53_array_index_1086654 ^ p53_array_index_1086625 ^ p53_array_index_1086592;
  assign p54_res7__605_comb = p53_literal_1076345[p54_res7__604_comb] ^ p53_literal_1076347[p54_res7__603_comb] ^ p53_literal_1076349[p54_res7__602_comb] ^ p53_literal_1076351[p53_res7__601] ^ p53_literal_1076353[p53_res7__600] ^ p53_literal_1076355[p53_res7__599] ^ p53_res7__598 ^ p53_literal_1076358[p53_res7__597] ^ p53_res7__596 ^ p53_array_index_1087070 ^ p53_array_index_1087046 ^ p53_array_index_1087020 ^ p53_array_index_1086740 ^ p53_array_index_1086711 ^ p53_literal_1076345[p53_array_index_1086681] ^ p53_array_index_1086682;
  assign p54_res__17_comb = {p54_res7__287_comb, p54_res7__286_comb, p54_res7__285_comb, p54_res7__284_comb, p54_res7__283_comb, p54_res7__282_comb, p53_res7__281, p53_res7__280, p53_res7__279, p53_res7__278, p53_res7__277, p53_res7__276, p53_res7__275, p53_res7__274, p53_res7__273, p53_res7__272};
  assign p54_xor_1087336_comb = p54_res__17_comb ^ p53_k4;
  assign p54_res7__606_comb = p53_literal_1076345[p54_res7__605_comb] ^ p53_literal_1076347[p54_res7__604_comb] ^ p53_literal_1076349[p54_res7__603_comb] ^ p53_literal_1076351[p54_res7__602_comb] ^ p53_literal_1076353[p53_res7__601] ^ p53_literal_1076355[p53_res7__600] ^ p53_res7__599 ^ p53_literal_1076358[p53_res7__598] ^ p53_res7__597 ^ p54_array_index_1087342_comb ^ p53_array_index_1087058 ^ p53_array_index_1087033 ^ p53_array_index_1086754 ^ p53_array_index_1086725 ^ p53_array_index_1086693 ^ p53_array_index_1086681;

  // Registers for pipe stage 54:
  reg [127:0] p54_xor_1086461;
  reg [127:0] p54_xor_1087336;
  reg [7:0] p54_array_index_1086680;
  reg [7:0] p54_res7__592;
  reg [7:0] p54_array_index_1086710;
  reg [7:0] p54_res7__593;
  reg [7:0] p54_res7__594;
  reg [7:0] p54_array_index_1086739;
  reg [7:0] p54_res7__595;
  reg [7:0] p54_res7__596;
  reg [7:0] p54_array_index_1087019;
  reg [7:0] p54_res7__597;
  reg [7:0] p54_res7__598;
  reg [7:0] p54_array_index_1087045;
  reg [7:0] p54_res7__599;
  reg [7:0] p54_res7__600;
  reg [7:0] p54_array_index_1087069;
  reg [7:0] p54_res7__601;
  reg [7:0] p54_res7__602;
  reg [7:0] p54_array_index_1087352;
  reg [7:0] p54_res7__603;
  reg [7:0] p54_res7__604;
  reg [7:0] p54_res7__605;
  reg [7:0] p54_res7__606;
  reg [7:0] p55_arr[256];
  reg [7:0] p55_literal_1076345[256];
  reg [7:0] p55_literal_1076347[256];
  reg [7:0] p55_literal_1076349[256];
  reg [7:0] p55_literal_1076351[256];
  reg [7:0] p55_literal_1076353[256];
  reg [7:0] p55_literal_1076355[256];
  reg [7:0] p55_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p54_xor_1086461 <= p53_xor_1086461;
    p54_xor_1087336 <= p54_xor_1087336_comb;
    p54_array_index_1086680 <= p53_array_index_1086680;
    p54_res7__592 <= p53_res7__592;
    p54_array_index_1086710 <= p53_array_index_1086710;
    p54_res7__593 <= p53_res7__593;
    p54_res7__594 <= p53_res7__594;
    p54_array_index_1086739 <= p53_array_index_1086739;
    p54_res7__595 <= p53_res7__595;
    p54_res7__596 <= p53_res7__596;
    p54_array_index_1087019 <= p53_array_index_1087019;
    p54_res7__597 <= p53_res7__597;
    p54_res7__598 <= p53_res7__598;
    p54_array_index_1087045 <= p53_array_index_1087045;
    p54_res7__599 <= p53_res7__599;
    p54_res7__600 <= p53_res7__600;
    p54_array_index_1087069 <= p53_array_index_1087069;
    p54_res7__601 <= p53_res7__601;
    p54_res7__602 <= p54_res7__602_comb;
    p54_array_index_1087352 <= p54_array_index_1087352_comb;
    p54_res7__603 <= p54_res7__603_comb;
    p54_res7__604 <= p54_res7__604_comb;
    p54_res7__605 <= p54_res7__605_comb;
    p54_res7__606 <= p54_res7__606_comb;
    p55_arr <= p54_arr;
    p55_literal_1076345 <= p54_literal_1076345;
    p55_literal_1076347 <= p54_literal_1076347;
    p55_literal_1076349 <= p54_literal_1076349;
    p55_literal_1076351 <= p54_literal_1076351;
    p55_literal_1076353 <= p54_literal_1076353;
    p55_literal_1076355 <= p54_literal_1076355;
    p55_literal_1076358 <= p54_literal_1076358;
  end

  // ===== Pipe stage 55:
  wire [127:0] p55_addedKey__59_comb;
  wire [7:0] p55_array_index_1087462_comb;
  wire [7:0] p55_array_index_1087463_comb;
  wire [7:0] p55_array_index_1087464_comb;
  wire [7:0] p55_array_index_1087465_comb;
  wire [7:0] p55_array_index_1087466_comb;
  wire [7:0] p55_array_index_1087467_comb;
  wire [7:0] p55_array_index_1087469_comb;
  wire [7:0] p55_array_index_1087471_comb;
  wire [7:0] p55_array_index_1087472_comb;
  wire [7:0] p55_array_index_1087473_comb;
  wire [7:0] p55_array_index_1087474_comb;
  wire [7:0] p55_array_index_1087475_comb;
  wire [7:0] p55_array_index_1087476_comb;
  wire [7:0] p55_array_index_1087478_comb;
  wire [7:0] p55_array_index_1087479_comb;
  wire [7:0] p55_array_index_1087480_comb;
  wire [7:0] p55_array_index_1087481_comb;
  wire [7:0] p55_array_index_1087482_comb;
  wire [7:0] p55_array_index_1087483_comb;
  wire [7:0] p55_array_index_1087484_comb;
  wire [7:0] p55_array_index_1087486_comb;
  wire [7:0] p55_res7__288_comb;
  wire [7:0] p55_array_index_1087495_comb;
  wire [7:0] p55_array_index_1087496_comb;
  wire [7:0] p55_array_index_1087497_comb;
  wire [7:0] p55_array_index_1087498_comb;
  wire [7:0] p55_array_index_1087499_comb;
  wire [7:0] p55_array_index_1087500_comb;
  wire [7:0] p55_res7__289_comb;
  wire [7:0] p55_array_index_1087510_comb;
  wire [7:0] p55_array_index_1087511_comb;
  wire [7:0] p55_array_index_1087512_comb;
  wire [7:0] p55_array_index_1087513_comb;
  wire [7:0] p55_array_index_1087514_comb;
  wire [7:0] p55_res7__290_comb;
  wire [7:0] p55_array_index_1087524_comb;
  wire [7:0] p55_array_index_1087525_comb;
  wire [7:0] p55_array_index_1087526_comb;
  wire [7:0] p55_array_index_1087527_comb;
  wire [7:0] p55_array_index_1087528_comb;
  wire [7:0] p55_res7__291_comb;
  wire [7:0] p55_array_index_1087539_comb;
  wire [7:0] p55_array_index_1087540_comb;
  wire [7:0] p55_array_index_1087541_comb;
  wire [7:0] p55_array_index_1087542_comb;
  wire [7:0] p55_res7__607_comb;
  wire [7:0] p55_res7__292_comb;
  wire [127:0] p55_res__37_comb;
  assign p55_addedKey__59_comb = p54_xor_1087336 ^ 128'h9d97_f6ba_bbd2_22da_7e5c_85f3_ead8_2b13;
  assign p55_array_index_1087462_comb = p54_arr[p55_addedKey__59_comb[127:120]];
  assign p55_array_index_1087463_comb = p54_arr[p55_addedKey__59_comb[119:112]];
  assign p55_array_index_1087464_comb = p54_arr[p55_addedKey__59_comb[111:104]];
  assign p55_array_index_1087465_comb = p54_arr[p55_addedKey__59_comb[103:96]];
  assign p55_array_index_1087466_comb = p54_arr[p55_addedKey__59_comb[95:88]];
  assign p55_array_index_1087467_comb = p54_arr[p55_addedKey__59_comb[87:80]];
  assign p55_array_index_1087469_comb = p54_arr[p55_addedKey__59_comb[71:64]];
  assign p55_array_index_1087471_comb = p54_arr[p55_addedKey__59_comb[55:48]];
  assign p55_array_index_1087472_comb = p54_arr[p55_addedKey__59_comb[47:40]];
  assign p55_array_index_1087473_comb = p54_arr[p55_addedKey__59_comb[39:32]];
  assign p55_array_index_1087474_comb = p54_arr[p55_addedKey__59_comb[31:24]];
  assign p55_array_index_1087475_comb = p54_arr[p55_addedKey__59_comb[23:16]];
  assign p55_array_index_1087476_comb = p54_arr[p55_addedKey__59_comb[15:8]];
  assign p55_array_index_1087478_comb = p54_literal_1076345[p55_array_index_1087462_comb];
  assign p55_array_index_1087479_comb = p54_literal_1076347[p55_array_index_1087463_comb];
  assign p55_array_index_1087480_comb = p54_literal_1076349[p55_array_index_1087464_comb];
  assign p55_array_index_1087481_comb = p54_literal_1076351[p55_array_index_1087465_comb];
  assign p55_array_index_1087482_comb = p54_literal_1076353[p55_array_index_1087466_comb];
  assign p55_array_index_1087483_comb = p54_literal_1076355[p55_array_index_1087467_comb];
  assign p55_array_index_1087484_comb = p54_arr[p55_addedKey__59_comb[79:72]];
  assign p55_array_index_1087486_comb = p54_arr[p55_addedKey__59_comb[63:56]];
  assign p55_res7__288_comb = p55_array_index_1087478_comb ^ p55_array_index_1087479_comb ^ p55_array_index_1087480_comb ^ p55_array_index_1087481_comb ^ p55_array_index_1087482_comb ^ p55_array_index_1087483_comb ^ p55_array_index_1087484_comb ^ p54_literal_1076358[p55_array_index_1087469_comb] ^ p55_array_index_1087486_comb ^ p54_literal_1076355[p55_array_index_1087471_comb] ^ p54_literal_1076353[p55_array_index_1087472_comb] ^ p54_literal_1076351[p55_array_index_1087473_comb] ^ p54_literal_1076349[p55_array_index_1087474_comb] ^ p54_literal_1076347[p55_array_index_1087475_comb] ^ p54_literal_1076345[p55_array_index_1087476_comb] ^ p54_arr[p55_addedKey__59_comb[7:0]];
  assign p55_array_index_1087495_comb = p54_literal_1076345[p55_res7__288_comb];
  assign p55_array_index_1087496_comb = p54_literal_1076347[p55_array_index_1087462_comb];
  assign p55_array_index_1087497_comb = p54_literal_1076349[p55_array_index_1087463_comb];
  assign p55_array_index_1087498_comb = p54_literal_1076351[p55_array_index_1087464_comb];
  assign p55_array_index_1087499_comb = p54_literal_1076353[p55_array_index_1087465_comb];
  assign p55_array_index_1087500_comb = p54_literal_1076355[p55_array_index_1087466_comb];
  assign p55_res7__289_comb = p55_array_index_1087495_comb ^ p55_array_index_1087496_comb ^ p55_array_index_1087497_comb ^ p55_array_index_1087498_comb ^ p55_array_index_1087499_comb ^ p55_array_index_1087500_comb ^ p55_array_index_1087467_comb ^ p54_literal_1076358[p55_array_index_1087484_comb] ^ p55_array_index_1087469_comb ^ p54_literal_1076355[p55_array_index_1087486_comb] ^ p54_literal_1076353[p55_array_index_1087471_comb] ^ p54_literal_1076351[p55_array_index_1087472_comb] ^ p54_literal_1076349[p55_array_index_1087473_comb] ^ p54_literal_1076347[p55_array_index_1087474_comb] ^ p54_literal_1076345[p55_array_index_1087475_comb] ^ p55_array_index_1087476_comb;
  assign p55_array_index_1087510_comb = p54_literal_1076347[p55_res7__288_comb];
  assign p55_array_index_1087511_comb = p54_literal_1076349[p55_array_index_1087462_comb];
  assign p55_array_index_1087512_comb = p54_literal_1076351[p55_array_index_1087463_comb];
  assign p55_array_index_1087513_comb = p54_literal_1076353[p55_array_index_1087464_comb];
  assign p55_array_index_1087514_comb = p54_literal_1076355[p55_array_index_1087465_comb];
  assign p55_res7__290_comb = p54_literal_1076345[p55_res7__289_comb] ^ p55_array_index_1087510_comb ^ p55_array_index_1087511_comb ^ p55_array_index_1087512_comb ^ p55_array_index_1087513_comb ^ p55_array_index_1087514_comb ^ p55_array_index_1087466_comb ^ p54_literal_1076358[p55_array_index_1087467_comb] ^ p55_array_index_1087484_comb ^ p54_literal_1076355[p55_array_index_1087469_comb] ^ p54_literal_1076353[p55_array_index_1087486_comb] ^ p54_literal_1076351[p55_array_index_1087471_comb] ^ p54_literal_1076349[p55_array_index_1087472_comb] ^ p54_literal_1076347[p55_array_index_1087473_comb] ^ p54_literal_1076345[p55_array_index_1087474_comb] ^ p55_array_index_1087475_comb;
  assign p55_array_index_1087524_comb = p54_literal_1076347[p55_res7__289_comb];
  assign p55_array_index_1087525_comb = p54_literal_1076349[p55_res7__288_comb];
  assign p55_array_index_1087526_comb = p54_literal_1076351[p55_array_index_1087462_comb];
  assign p55_array_index_1087527_comb = p54_literal_1076353[p55_array_index_1087463_comb];
  assign p55_array_index_1087528_comb = p54_literal_1076355[p55_array_index_1087464_comb];
  assign p55_res7__291_comb = p54_literal_1076345[p55_res7__290_comb] ^ p55_array_index_1087524_comb ^ p55_array_index_1087525_comb ^ p55_array_index_1087526_comb ^ p55_array_index_1087527_comb ^ p55_array_index_1087528_comb ^ p55_array_index_1087465_comb ^ p54_literal_1076358[p55_array_index_1087466_comb] ^ p55_array_index_1087467_comb ^ p54_literal_1076355[p55_array_index_1087484_comb] ^ p54_literal_1076353[p55_array_index_1087469_comb] ^ p54_literal_1076351[p55_array_index_1087486_comb] ^ p54_literal_1076349[p55_array_index_1087471_comb] ^ p54_literal_1076347[p55_array_index_1087472_comb] ^ p54_literal_1076345[p55_array_index_1087473_comb] ^ p55_array_index_1087474_comb;
  assign p55_array_index_1087539_comb = p54_literal_1076349[p55_res7__289_comb];
  assign p55_array_index_1087540_comb = p54_literal_1076351[p55_res7__288_comb];
  assign p55_array_index_1087541_comb = p54_literal_1076353[p55_array_index_1087462_comb];
  assign p55_array_index_1087542_comb = p54_literal_1076355[p55_array_index_1087463_comb];
  assign p55_res7__607_comb = p54_literal_1076345[p54_res7__606] ^ p54_literal_1076347[p54_res7__605] ^ p54_literal_1076349[p54_res7__604] ^ p54_literal_1076351[p54_res7__603] ^ p54_literal_1076353[p54_res7__602] ^ p54_literal_1076355[p54_res7__601] ^ p54_res7__600 ^ p54_literal_1076358[p54_res7__599] ^ p54_res7__598 ^ p54_array_index_1087352 ^ p54_array_index_1087069 ^ p54_array_index_1087045 ^ p54_array_index_1087019 ^ p54_array_index_1086739 ^ p54_array_index_1086710 ^ p54_array_index_1086680;
  assign p55_res7__292_comb = p54_literal_1076345[p55_res7__291_comb] ^ p54_literal_1076347[p55_res7__290_comb] ^ p55_array_index_1087539_comb ^ p55_array_index_1087540_comb ^ p55_array_index_1087541_comb ^ p55_array_index_1087542_comb ^ p55_array_index_1087464_comb ^ p54_literal_1076358[p55_array_index_1087465_comb] ^ p55_array_index_1087466_comb ^ p55_array_index_1087483_comb ^ p54_literal_1076353[p55_array_index_1087484_comb] ^ p54_literal_1076351[p55_array_index_1087469_comb] ^ p54_literal_1076349[p55_array_index_1087486_comb] ^ p54_literal_1076347[p55_array_index_1087471_comb] ^ p54_literal_1076345[p55_array_index_1087472_comb] ^ p55_array_index_1087473_comb;
  assign p55_res__37_comb = {p55_res7__607_comb, p54_res7__606, p54_res7__605, p54_res7__604, p54_res7__603, p54_res7__602, p54_res7__601, p54_res7__600, p54_res7__599, p54_res7__598, p54_res7__597, p54_res7__596, p54_res7__595, p54_res7__594, p54_res7__593, p54_res7__592};

  // Registers for pipe stage 55:
  reg [127:0] p55_xor_1086461;
  reg [127:0] p55_xor_1087336;
  reg [7:0] p55_array_index_1087462;
  reg [7:0] p55_array_index_1087463;
  reg [7:0] p55_array_index_1087464;
  reg [7:0] p55_array_index_1087465;
  reg [7:0] p55_array_index_1087466;
  reg [7:0] p55_array_index_1087467;
  reg [7:0] p55_array_index_1087469;
  reg [7:0] p55_array_index_1087471;
  reg [7:0] p55_array_index_1087472;
  reg [7:0] p55_array_index_1087478;
  reg [7:0] p55_array_index_1087479;
  reg [7:0] p55_array_index_1087480;
  reg [7:0] p55_array_index_1087481;
  reg [7:0] p55_array_index_1087482;
  reg [7:0] p55_array_index_1087484;
  reg [7:0] p55_array_index_1087486;
  reg [7:0] p55_res7__288;
  reg [7:0] p55_array_index_1087495;
  reg [7:0] p55_array_index_1087496;
  reg [7:0] p55_array_index_1087497;
  reg [7:0] p55_array_index_1087498;
  reg [7:0] p55_array_index_1087499;
  reg [7:0] p55_array_index_1087500;
  reg [7:0] p55_res7__289;
  reg [7:0] p55_array_index_1087510;
  reg [7:0] p55_array_index_1087511;
  reg [7:0] p55_array_index_1087512;
  reg [7:0] p55_array_index_1087513;
  reg [7:0] p55_array_index_1087514;
  reg [7:0] p55_res7__290;
  reg [7:0] p55_array_index_1087524;
  reg [7:0] p55_array_index_1087525;
  reg [7:0] p55_array_index_1087526;
  reg [7:0] p55_array_index_1087527;
  reg [7:0] p55_array_index_1087528;
  reg [7:0] p55_res7__291;
  reg [7:0] p55_array_index_1087539;
  reg [7:0] p55_array_index_1087540;
  reg [7:0] p55_array_index_1087541;
  reg [7:0] p55_array_index_1087542;
  reg [7:0] p55_res7__292;
  reg [127:0] p55_res__37;
  reg [7:0] p56_arr[256];
  reg [7:0] p56_literal_1076345[256];
  reg [7:0] p56_literal_1076347[256];
  reg [7:0] p56_literal_1076349[256];
  reg [7:0] p56_literal_1076351[256];
  reg [7:0] p56_literal_1076353[256];
  reg [7:0] p56_literal_1076355[256];
  reg [7:0] p56_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p55_xor_1086461 <= p54_xor_1086461;
    p55_xor_1087336 <= p54_xor_1087336;
    p55_array_index_1087462 <= p55_array_index_1087462_comb;
    p55_array_index_1087463 <= p55_array_index_1087463_comb;
    p55_array_index_1087464 <= p55_array_index_1087464_comb;
    p55_array_index_1087465 <= p55_array_index_1087465_comb;
    p55_array_index_1087466 <= p55_array_index_1087466_comb;
    p55_array_index_1087467 <= p55_array_index_1087467_comb;
    p55_array_index_1087469 <= p55_array_index_1087469_comb;
    p55_array_index_1087471 <= p55_array_index_1087471_comb;
    p55_array_index_1087472 <= p55_array_index_1087472_comb;
    p55_array_index_1087478 <= p55_array_index_1087478_comb;
    p55_array_index_1087479 <= p55_array_index_1087479_comb;
    p55_array_index_1087480 <= p55_array_index_1087480_comb;
    p55_array_index_1087481 <= p55_array_index_1087481_comb;
    p55_array_index_1087482 <= p55_array_index_1087482_comb;
    p55_array_index_1087484 <= p55_array_index_1087484_comb;
    p55_array_index_1087486 <= p55_array_index_1087486_comb;
    p55_res7__288 <= p55_res7__288_comb;
    p55_array_index_1087495 <= p55_array_index_1087495_comb;
    p55_array_index_1087496 <= p55_array_index_1087496_comb;
    p55_array_index_1087497 <= p55_array_index_1087497_comb;
    p55_array_index_1087498 <= p55_array_index_1087498_comb;
    p55_array_index_1087499 <= p55_array_index_1087499_comb;
    p55_array_index_1087500 <= p55_array_index_1087500_comb;
    p55_res7__289 <= p55_res7__289_comb;
    p55_array_index_1087510 <= p55_array_index_1087510_comb;
    p55_array_index_1087511 <= p55_array_index_1087511_comb;
    p55_array_index_1087512 <= p55_array_index_1087512_comb;
    p55_array_index_1087513 <= p55_array_index_1087513_comb;
    p55_array_index_1087514 <= p55_array_index_1087514_comb;
    p55_res7__290 <= p55_res7__290_comb;
    p55_array_index_1087524 <= p55_array_index_1087524_comb;
    p55_array_index_1087525 <= p55_array_index_1087525_comb;
    p55_array_index_1087526 <= p55_array_index_1087526_comb;
    p55_array_index_1087527 <= p55_array_index_1087527_comb;
    p55_array_index_1087528 <= p55_array_index_1087528_comb;
    p55_res7__291 <= p55_res7__291_comb;
    p55_array_index_1087539 <= p55_array_index_1087539_comb;
    p55_array_index_1087540 <= p55_array_index_1087540_comb;
    p55_array_index_1087541 <= p55_array_index_1087541_comb;
    p55_array_index_1087542 <= p55_array_index_1087542_comb;
    p55_res7__292 <= p55_res7__292_comb;
    p55_res__37 <= p55_res__37_comb;
    p56_arr <= p55_arr;
    p56_literal_1076345 <= p55_literal_1076345;
    p56_literal_1076347 <= p55_literal_1076347;
    p56_literal_1076349 <= p55_literal_1076349;
    p56_literal_1076351 <= p55_literal_1076351;
    p56_literal_1076353 <= p55_literal_1076353;
    p56_literal_1076355 <= p55_literal_1076355;
    p56_literal_1076358 <= p55_literal_1076358;
  end

  // ===== Pipe stage 56:
  wire [7:0] p56_array_index_1087665_comb;
  wire [7:0] p56_array_index_1087666_comb;
  wire [7:0] p56_array_index_1087667_comb;
  wire [7:0] p56_array_index_1087668_comb;
  wire [7:0] p56_res7__293_comb;
  wire [7:0] p56_array_index_1087679_comb;
  wire [7:0] p56_array_index_1087680_comb;
  wire [7:0] p56_array_index_1087681_comb;
  wire [7:0] p56_res7__294_comb;
  wire [7:0] p56_array_index_1087691_comb;
  wire [7:0] p56_array_index_1087692_comb;
  wire [7:0] p56_array_index_1087693_comb;
  wire [7:0] p56_res7__295_comb;
  wire [7:0] p56_array_index_1087704_comb;
  wire [7:0] p56_array_index_1087705_comb;
  wire [7:0] p56_res7__296_comb;
  wire [7:0] p56_array_index_1087715_comb;
  wire [7:0] p56_array_index_1087716_comb;
  wire [7:0] p56_res7__297_comb;
  wire [7:0] p56_array_index_1087722_comb;
  wire [7:0] p56_array_index_1087723_comb;
  wire [7:0] p56_array_index_1087724_comb;
  wire [7:0] p56_array_index_1087725_comb;
  wire [7:0] p56_array_index_1087726_comb;
  wire [7:0] p56_array_index_1087727_comb;
  wire [7:0] p56_array_index_1087728_comb;
  wire [7:0] p56_array_index_1087729_comb;
  wire [7:0] p56_array_index_1087730_comb;
  assign p56_array_index_1087665_comb = p55_literal_1076349[p55_res7__290];
  assign p56_array_index_1087666_comb = p55_literal_1076351[p55_res7__289];
  assign p56_array_index_1087667_comb = p55_literal_1076353[p55_res7__288];
  assign p56_array_index_1087668_comb = p55_literal_1076355[p55_array_index_1087462];
  assign p56_res7__293_comb = p55_literal_1076345[p55_res7__292] ^ p55_literal_1076347[p55_res7__291] ^ p56_array_index_1087665_comb ^ p56_array_index_1087666_comb ^ p56_array_index_1087667_comb ^ p56_array_index_1087668_comb ^ p55_array_index_1087463 ^ p55_literal_1076358[p55_array_index_1087464] ^ p55_array_index_1087465 ^ p55_array_index_1087500 ^ p55_literal_1076353[p55_array_index_1087467] ^ p55_literal_1076351[p55_array_index_1087484] ^ p55_literal_1076349[p55_array_index_1087469] ^ p55_literal_1076347[p55_array_index_1087486] ^ p55_literal_1076345[p55_array_index_1087471] ^ p55_array_index_1087472;
  assign p56_array_index_1087679_comb = p55_literal_1076351[p55_res7__290];
  assign p56_array_index_1087680_comb = p55_literal_1076353[p55_res7__289];
  assign p56_array_index_1087681_comb = p55_literal_1076355[p55_res7__288];
  assign p56_res7__294_comb = p55_literal_1076345[p56_res7__293_comb] ^ p55_literal_1076347[p55_res7__292] ^ p55_literal_1076349[p55_res7__291] ^ p56_array_index_1087679_comb ^ p56_array_index_1087680_comb ^ p56_array_index_1087681_comb ^ p55_array_index_1087462 ^ p55_literal_1076358[p55_array_index_1087463] ^ p55_array_index_1087464 ^ p55_array_index_1087514 ^ p55_array_index_1087482 ^ p55_literal_1076351[p55_array_index_1087467] ^ p55_literal_1076349[p55_array_index_1087484] ^ p55_literal_1076347[p55_array_index_1087469] ^ p55_literal_1076345[p55_array_index_1087486] ^ p55_array_index_1087471;
  assign p56_array_index_1087691_comb = p55_literal_1076351[p55_res7__291];
  assign p56_array_index_1087692_comb = p55_literal_1076353[p55_res7__290];
  assign p56_array_index_1087693_comb = p55_literal_1076355[p55_res7__289];
  assign p56_res7__295_comb = p55_literal_1076345[p56_res7__294_comb] ^ p55_literal_1076347[p56_res7__293_comb] ^ p55_literal_1076349[p55_res7__292] ^ p56_array_index_1087691_comb ^ p56_array_index_1087692_comb ^ p56_array_index_1087693_comb ^ p55_res7__288 ^ p55_literal_1076358[p55_array_index_1087462] ^ p55_array_index_1087463 ^ p55_array_index_1087528 ^ p55_array_index_1087499 ^ p55_literal_1076351[p55_array_index_1087466] ^ p55_literal_1076349[p55_array_index_1087467] ^ p55_literal_1076347[p55_array_index_1087484] ^ p55_literal_1076345[p55_array_index_1087469] ^ p55_array_index_1087486;
  assign p56_array_index_1087704_comb = p55_literal_1076353[p55_res7__291];
  assign p56_array_index_1087705_comb = p55_literal_1076355[p55_res7__290];
  assign p56_res7__296_comb = p55_literal_1076345[p56_res7__295_comb] ^ p55_literal_1076347[p56_res7__294_comb] ^ p55_literal_1076349[p56_res7__293_comb] ^ p55_literal_1076351[p55_res7__292] ^ p56_array_index_1087704_comb ^ p56_array_index_1087705_comb ^ p55_res7__289 ^ p55_literal_1076358[p55_res7__288] ^ p55_array_index_1087462 ^ p55_array_index_1087542 ^ p55_array_index_1087513 ^ p55_array_index_1087481 ^ p55_literal_1076349[p55_array_index_1087466] ^ p55_literal_1076347[p55_array_index_1087467] ^ p55_literal_1076345[p55_array_index_1087484] ^ p55_array_index_1087469;
  assign p56_array_index_1087715_comb = p55_literal_1076353[p55_res7__292];
  assign p56_array_index_1087716_comb = p55_literal_1076355[p55_res7__291];
  assign p56_res7__297_comb = p55_literal_1076345[p56_res7__296_comb] ^ p55_literal_1076347[p56_res7__295_comb] ^ p55_literal_1076349[p56_res7__294_comb] ^ p55_literal_1076351[p56_res7__293_comb] ^ p56_array_index_1087715_comb ^ p56_array_index_1087716_comb ^ p55_res7__290 ^ p55_literal_1076358[p55_res7__289] ^ p55_res7__288 ^ p56_array_index_1087668_comb ^ p55_array_index_1087527 ^ p55_array_index_1087498 ^ p55_literal_1076349[p55_array_index_1087465] ^ p55_literal_1076347[p55_array_index_1087466] ^ p55_literal_1076345[p55_array_index_1087467] ^ p55_array_index_1087484;
  assign p56_array_index_1087722_comb = p55_literal_1076345[p56_res7__297_comb];
  assign p56_array_index_1087723_comb = p55_literal_1076347[p56_res7__296_comb];
  assign p56_array_index_1087724_comb = p55_literal_1076349[p56_res7__295_comb];
  assign p56_array_index_1087725_comb = p55_literal_1076351[p56_res7__294_comb];
  assign p56_array_index_1087726_comb = p55_literal_1076353[p56_res7__293_comb];
  assign p56_array_index_1087727_comb = p55_literal_1076355[p55_res7__292];
  assign p56_array_index_1087728_comb = p55_literal_1076358[p55_res7__290];
  assign p56_array_index_1087729_comb = p55_literal_1076347[p55_array_index_1087465];
  assign p56_array_index_1087730_comb = p55_literal_1076345[p55_array_index_1087466];

  // Registers for pipe stage 56:
  reg [127:0] p56_xor_1086461;
  reg [127:0] p56_xor_1087336;
  reg [7:0] p56_array_index_1087462;
  reg [7:0] p56_array_index_1087463;
  reg [7:0] p56_array_index_1087464;
  reg [7:0] p56_array_index_1087465;
  reg [7:0] p56_array_index_1087466;
  reg [7:0] p56_array_index_1087467;
  reg [7:0] p56_array_index_1087478;
  reg [7:0] p56_array_index_1087479;
  reg [7:0] p56_array_index_1087480;
  reg [7:0] p56_res7__288;
  reg [7:0] p56_array_index_1087495;
  reg [7:0] p56_array_index_1087496;
  reg [7:0] p56_array_index_1087497;
  reg [7:0] p56_res7__289;
  reg [7:0] p56_array_index_1087510;
  reg [7:0] p56_array_index_1087511;
  reg [7:0] p56_array_index_1087512;
  reg [7:0] p56_res7__290;
  reg [7:0] p56_array_index_1087524;
  reg [7:0] p56_array_index_1087525;
  reg [7:0] p56_array_index_1087526;
  reg [7:0] p56_res7__291;
  reg [7:0] p56_array_index_1087539;
  reg [7:0] p56_array_index_1087540;
  reg [7:0] p56_array_index_1087541;
  reg [7:0] p56_res7__292;
  reg [7:0] p56_array_index_1087665;
  reg [7:0] p56_array_index_1087666;
  reg [7:0] p56_array_index_1087667;
  reg [7:0] p56_res7__293;
  reg [7:0] p56_array_index_1087679;
  reg [7:0] p56_array_index_1087680;
  reg [7:0] p56_array_index_1087681;
  reg [7:0] p56_res7__294;
  reg [7:0] p56_array_index_1087691;
  reg [7:0] p56_array_index_1087692;
  reg [7:0] p56_array_index_1087693;
  reg [7:0] p56_res7__295;
  reg [7:0] p56_array_index_1087704;
  reg [7:0] p56_array_index_1087705;
  reg [7:0] p56_res7__296;
  reg [7:0] p56_array_index_1087715;
  reg [7:0] p56_array_index_1087716;
  reg [7:0] p56_res7__297;
  reg [7:0] p56_array_index_1087722;
  reg [7:0] p56_array_index_1087723;
  reg [7:0] p56_array_index_1087724;
  reg [7:0] p56_array_index_1087725;
  reg [7:0] p56_array_index_1087726;
  reg [7:0] p56_array_index_1087727;
  reg [7:0] p56_array_index_1087728;
  reg [7:0] p56_array_index_1087729;
  reg [7:0] p56_array_index_1087730;
  reg [127:0] p56_res__37;
  reg [7:0] p57_arr[256];
  reg [7:0] p57_literal_1076345[256];
  reg [7:0] p57_literal_1076347[256];
  reg [7:0] p57_literal_1076349[256];
  reg [7:0] p57_literal_1076351[256];
  reg [7:0] p57_literal_1076353[256];
  reg [7:0] p57_literal_1076355[256];
  reg [7:0] p57_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p56_xor_1086461 <= p55_xor_1086461;
    p56_xor_1087336 <= p55_xor_1087336;
    p56_array_index_1087462 <= p55_array_index_1087462;
    p56_array_index_1087463 <= p55_array_index_1087463;
    p56_array_index_1087464 <= p55_array_index_1087464;
    p56_array_index_1087465 <= p55_array_index_1087465;
    p56_array_index_1087466 <= p55_array_index_1087466;
    p56_array_index_1087467 <= p55_array_index_1087467;
    p56_array_index_1087478 <= p55_array_index_1087478;
    p56_array_index_1087479 <= p55_array_index_1087479;
    p56_array_index_1087480 <= p55_array_index_1087480;
    p56_res7__288 <= p55_res7__288;
    p56_array_index_1087495 <= p55_array_index_1087495;
    p56_array_index_1087496 <= p55_array_index_1087496;
    p56_array_index_1087497 <= p55_array_index_1087497;
    p56_res7__289 <= p55_res7__289;
    p56_array_index_1087510 <= p55_array_index_1087510;
    p56_array_index_1087511 <= p55_array_index_1087511;
    p56_array_index_1087512 <= p55_array_index_1087512;
    p56_res7__290 <= p55_res7__290;
    p56_array_index_1087524 <= p55_array_index_1087524;
    p56_array_index_1087525 <= p55_array_index_1087525;
    p56_array_index_1087526 <= p55_array_index_1087526;
    p56_res7__291 <= p55_res7__291;
    p56_array_index_1087539 <= p55_array_index_1087539;
    p56_array_index_1087540 <= p55_array_index_1087540;
    p56_array_index_1087541 <= p55_array_index_1087541;
    p56_res7__292 <= p55_res7__292;
    p56_array_index_1087665 <= p56_array_index_1087665_comb;
    p56_array_index_1087666 <= p56_array_index_1087666_comb;
    p56_array_index_1087667 <= p56_array_index_1087667_comb;
    p56_res7__293 <= p56_res7__293_comb;
    p56_array_index_1087679 <= p56_array_index_1087679_comb;
    p56_array_index_1087680 <= p56_array_index_1087680_comb;
    p56_array_index_1087681 <= p56_array_index_1087681_comb;
    p56_res7__294 <= p56_res7__294_comb;
    p56_array_index_1087691 <= p56_array_index_1087691_comb;
    p56_array_index_1087692 <= p56_array_index_1087692_comb;
    p56_array_index_1087693 <= p56_array_index_1087693_comb;
    p56_res7__295 <= p56_res7__295_comb;
    p56_array_index_1087704 <= p56_array_index_1087704_comb;
    p56_array_index_1087705 <= p56_array_index_1087705_comb;
    p56_res7__296 <= p56_res7__296_comb;
    p56_array_index_1087715 <= p56_array_index_1087715_comb;
    p56_array_index_1087716 <= p56_array_index_1087716_comb;
    p56_res7__297 <= p56_res7__297_comb;
    p56_array_index_1087722 <= p56_array_index_1087722_comb;
    p56_array_index_1087723 <= p56_array_index_1087723_comb;
    p56_array_index_1087724 <= p56_array_index_1087724_comb;
    p56_array_index_1087725 <= p56_array_index_1087725_comb;
    p56_array_index_1087726 <= p56_array_index_1087726_comb;
    p56_array_index_1087727 <= p56_array_index_1087727_comb;
    p56_array_index_1087728 <= p56_array_index_1087728_comb;
    p56_array_index_1087729 <= p56_array_index_1087729_comb;
    p56_array_index_1087730 <= p56_array_index_1087730_comb;
    p56_res__37 <= p55_res__37;
    p57_arr <= p56_arr;
    p57_literal_1076345 <= p56_literal_1076345;
    p57_literal_1076347 <= p56_literal_1076347;
    p57_literal_1076349 <= p56_literal_1076349;
    p57_literal_1076351 <= p56_literal_1076351;
    p57_literal_1076353 <= p56_literal_1076353;
    p57_literal_1076355 <= p56_literal_1076355;
    p57_literal_1076358 <= p56_literal_1076358;
  end

  // ===== Pipe stage 57:
  wire [7:0] p57_res7__298_comb;
  wire [7:0] p57_array_index_1087865_comb;
  wire [7:0] p57_res7__299_comb;
  wire [7:0] p57_res7__300_comb;
  wire [7:0] p57_res7__301_comb;
  wire [7:0] p57_res7__302_comb;
  wire [7:0] p57_res7__303_comb;
  wire [127:0] p57_res__18_comb;
  wire [127:0] p57_xor_1087905_comb;
  assign p57_res7__298_comb = p56_array_index_1087722 ^ p56_array_index_1087723 ^ p56_array_index_1087724 ^ p56_array_index_1087725 ^ p56_array_index_1087726 ^ p56_array_index_1087727 ^ p56_res7__291 ^ p56_array_index_1087728 ^ p56_res7__289 ^ p56_array_index_1087681 ^ p56_array_index_1087541 ^ p56_array_index_1087512 ^ p56_array_index_1087480 ^ p56_array_index_1087729 ^ p56_array_index_1087730 ^ p56_array_index_1087467;
  assign p57_array_index_1087865_comb = p56_literal_1076355[p56_res7__293];
  assign p57_res7__299_comb = p56_literal_1076345[p57_res7__298_comb] ^ p56_literal_1076347[p56_res7__297] ^ p56_literal_1076349[p56_res7__296] ^ p56_literal_1076351[p56_res7__295] ^ p56_literal_1076353[p56_res7__294] ^ p57_array_index_1087865_comb ^ p56_res7__292 ^ p56_literal_1076358[p56_res7__291] ^ p56_res7__290 ^ p56_array_index_1087693 ^ p56_array_index_1087667 ^ p56_array_index_1087526 ^ p56_array_index_1087497 ^ p56_literal_1076347[p56_array_index_1087464] ^ p56_literal_1076345[p56_array_index_1087465] ^ p56_array_index_1087466;
  assign p57_res7__300_comb = p56_literal_1076345[p57_res7__299_comb] ^ p56_literal_1076347[p57_res7__298_comb] ^ p56_literal_1076349[p56_res7__297] ^ p56_literal_1076351[p56_res7__296] ^ p56_literal_1076353[p56_res7__295] ^ p56_literal_1076355[p56_res7__294] ^ p56_res7__293 ^ p56_literal_1076358[p56_res7__292] ^ p56_res7__291 ^ p56_array_index_1087705 ^ p56_array_index_1087680 ^ p56_array_index_1087540 ^ p56_array_index_1087511 ^ p56_array_index_1087479 ^ p56_literal_1076345[p56_array_index_1087464] ^ p56_array_index_1087465;
  assign p57_res7__301_comb = p56_literal_1076345[p57_res7__300_comb] ^ p56_literal_1076347[p57_res7__299_comb] ^ p56_literal_1076349[p57_res7__298_comb] ^ p56_literal_1076351[p56_res7__297] ^ p56_literal_1076353[p56_res7__296] ^ p56_literal_1076355[p56_res7__295] ^ p56_res7__294 ^ p56_literal_1076358[p56_res7__293] ^ p56_res7__292 ^ p56_array_index_1087716 ^ p56_array_index_1087692 ^ p56_array_index_1087666 ^ p56_array_index_1087525 ^ p56_array_index_1087496 ^ p56_literal_1076345[p56_array_index_1087463] ^ p56_array_index_1087464;
  assign p57_res7__302_comb = p56_literal_1076345[p57_res7__301_comb] ^ p56_literal_1076347[p57_res7__300_comb] ^ p56_literal_1076349[p57_res7__299_comb] ^ p56_literal_1076351[p57_res7__298_comb] ^ p56_literal_1076353[p56_res7__297] ^ p56_literal_1076355[p56_res7__296] ^ p56_res7__295 ^ p56_literal_1076358[p56_res7__294] ^ p56_res7__293 ^ p56_array_index_1087727 ^ p56_array_index_1087704 ^ p56_array_index_1087679 ^ p56_array_index_1087539 ^ p56_array_index_1087510 ^ p56_array_index_1087478 ^ p56_array_index_1087463;
  assign p57_res7__303_comb = p56_literal_1076345[p57_res7__302_comb] ^ p56_literal_1076347[p57_res7__301_comb] ^ p56_literal_1076349[p57_res7__300_comb] ^ p56_literal_1076351[p57_res7__299_comb] ^ p56_literal_1076353[p57_res7__298_comb] ^ p56_literal_1076355[p56_res7__297] ^ p56_res7__296 ^ p56_literal_1076358[p56_res7__295] ^ p56_res7__294 ^ p57_array_index_1087865_comb ^ p56_array_index_1087715 ^ p56_array_index_1087691 ^ p56_array_index_1087665 ^ p56_array_index_1087524 ^ p56_array_index_1087495 ^ p56_array_index_1087462;
  assign p57_res__18_comb = {p57_res7__303_comb, p57_res7__302_comb, p57_res7__301_comb, p57_res7__300_comb, p57_res7__299_comb, p57_res7__298_comb, p56_res7__297, p56_res7__296, p56_res7__295, p56_res7__294, p56_res7__293, p56_res7__292, p56_res7__291, p56_res7__290, p56_res7__289, p56_res7__288};
  assign p57_xor_1087905_comb = p57_res__18_comb ^ p56_xor_1086461;

  // Registers for pipe stage 57:
  reg [127:0] p57_xor_1087336;
  reg [127:0] p57_xor_1087905;
  reg [127:0] p57_res__37;
  reg [7:0] p58_arr[256];
  reg [7:0] p58_literal_1076345[256];
  reg [7:0] p58_literal_1076347[256];
  reg [7:0] p58_literal_1076349[256];
  reg [7:0] p58_literal_1076351[256];
  reg [7:0] p58_literal_1076353[256];
  reg [7:0] p58_literal_1076355[256];
  reg [7:0] p58_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p57_xor_1087336 <= p56_xor_1087336;
    p57_xor_1087905 <= p57_xor_1087905_comb;
    p57_res__37 <= p56_res__37;
    p58_arr <= p57_arr;
    p58_literal_1076345 <= p57_literal_1076345;
    p58_literal_1076347 <= p57_literal_1076347;
    p58_literal_1076349 <= p57_literal_1076349;
    p58_literal_1076351 <= p57_literal_1076351;
    p58_literal_1076353 <= p57_literal_1076353;
    p58_literal_1076355 <= p57_literal_1076355;
    p58_literal_1076358 <= p57_literal_1076358;
  end

  // ===== Pipe stage 58:
  wire [127:0] p58_addedKey__60_comb;
  wire [7:0] p58_array_index_1087943_comb;
  wire [7:0] p58_array_index_1087944_comb;
  wire [7:0] p58_array_index_1087945_comb;
  wire [7:0] p58_array_index_1087946_comb;
  wire [7:0] p58_array_index_1087947_comb;
  wire [7:0] p58_array_index_1087948_comb;
  wire [7:0] p58_array_index_1087950_comb;
  wire [7:0] p58_array_index_1087952_comb;
  wire [7:0] p58_array_index_1087953_comb;
  wire [7:0] p58_array_index_1087954_comb;
  wire [7:0] p58_array_index_1087955_comb;
  wire [7:0] p58_array_index_1087956_comb;
  wire [7:0] p58_array_index_1087957_comb;
  wire [7:0] p58_array_index_1087959_comb;
  wire [7:0] p58_array_index_1087960_comb;
  wire [7:0] p58_array_index_1087961_comb;
  wire [7:0] p58_array_index_1087962_comb;
  wire [7:0] p58_array_index_1087963_comb;
  wire [7:0] p58_array_index_1087964_comb;
  wire [7:0] p58_array_index_1087965_comb;
  wire [7:0] p58_array_index_1087967_comb;
  wire [7:0] p58_res7__304_comb;
  wire [7:0] p58_array_index_1087976_comb;
  wire [7:0] p58_array_index_1087977_comb;
  wire [7:0] p58_array_index_1087978_comb;
  wire [7:0] p58_array_index_1087979_comb;
  wire [7:0] p58_array_index_1087980_comb;
  wire [7:0] p58_array_index_1087981_comb;
  wire [7:0] p58_res7__305_comb;
  wire [7:0] p58_array_index_1087991_comb;
  wire [7:0] p58_array_index_1087992_comb;
  wire [7:0] p58_array_index_1087993_comb;
  wire [7:0] p58_array_index_1087994_comb;
  wire [7:0] p58_array_index_1087995_comb;
  wire [7:0] p58_res7__306_comb;
  wire [7:0] p58_array_index_1088005_comb;
  wire [7:0] p58_array_index_1088006_comb;
  wire [7:0] p58_array_index_1088007_comb;
  wire [7:0] p58_array_index_1088008_comb;
  wire [7:0] p58_array_index_1088009_comb;
  wire [7:0] p58_res7__307_comb;
  wire [7:0] p58_array_index_1088020_comb;
  wire [7:0] p58_array_index_1088021_comb;
  wire [7:0] p58_array_index_1088022_comb;
  wire [7:0] p58_array_index_1088023_comb;
  wire [7:0] p58_res7__308_comb;
  assign p58_addedKey__60_comb = p57_xor_1087905 ^ 128'h547f_7727_7ce9_8774_2ea9_3083_bcc2_4114;
  assign p58_array_index_1087943_comb = p57_arr[p58_addedKey__60_comb[127:120]];
  assign p58_array_index_1087944_comb = p57_arr[p58_addedKey__60_comb[119:112]];
  assign p58_array_index_1087945_comb = p57_arr[p58_addedKey__60_comb[111:104]];
  assign p58_array_index_1087946_comb = p57_arr[p58_addedKey__60_comb[103:96]];
  assign p58_array_index_1087947_comb = p57_arr[p58_addedKey__60_comb[95:88]];
  assign p58_array_index_1087948_comb = p57_arr[p58_addedKey__60_comb[87:80]];
  assign p58_array_index_1087950_comb = p57_arr[p58_addedKey__60_comb[71:64]];
  assign p58_array_index_1087952_comb = p57_arr[p58_addedKey__60_comb[55:48]];
  assign p58_array_index_1087953_comb = p57_arr[p58_addedKey__60_comb[47:40]];
  assign p58_array_index_1087954_comb = p57_arr[p58_addedKey__60_comb[39:32]];
  assign p58_array_index_1087955_comb = p57_arr[p58_addedKey__60_comb[31:24]];
  assign p58_array_index_1087956_comb = p57_arr[p58_addedKey__60_comb[23:16]];
  assign p58_array_index_1087957_comb = p57_arr[p58_addedKey__60_comb[15:8]];
  assign p58_array_index_1087959_comb = p57_literal_1076345[p58_array_index_1087943_comb];
  assign p58_array_index_1087960_comb = p57_literal_1076347[p58_array_index_1087944_comb];
  assign p58_array_index_1087961_comb = p57_literal_1076349[p58_array_index_1087945_comb];
  assign p58_array_index_1087962_comb = p57_literal_1076351[p58_array_index_1087946_comb];
  assign p58_array_index_1087963_comb = p57_literal_1076353[p58_array_index_1087947_comb];
  assign p58_array_index_1087964_comb = p57_literal_1076355[p58_array_index_1087948_comb];
  assign p58_array_index_1087965_comb = p57_arr[p58_addedKey__60_comb[79:72]];
  assign p58_array_index_1087967_comb = p57_arr[p58_addedKey__60_comb[63:56]];
  assign p58_res7__304_comb = p58_array_index_1087959_comb ^ p58_array_index_1087960_comb ^ p58_array_index_1087961_comb ^ p58_array_index_1087962_comb ^ p58_array_index_1087963_comb ^ p58_array_index_1087964_comb ^ p58_array_index_1087965_comb ^ p57_literal_1076358[p58_array_index_1087950_comb] ^ p58_array_index_1087967_comb ^ p57_literal_1076355[p58_array_index_1087952_comb] ^ p57_literal_1076353[p58_array_index_1087953_comb] ^ p57_literal_1076351[p58_array_index_1087954_comb] ^ p57_literal_1076349[p58_array_index_1087955_comb] ^ p57_literal_1076347[p58_array_index_1087956_comb] ^ p57_literal_1076345[p58_array_index_1087957_comb] ^ p57_arr[p58_addedKey__60_comb[7:0]];
  assign p58_array_index_1087976_comb = p57_literal_1076345[p58_res7__304_comb];
  assign p58_array_index_1087977_comb = p57_literal_1076347[p58_array_index_1087943_comb];
  assign p58_array_index_1087978_comb = p57_literal_1076349[p58_array_index_1087944_comb];
  assign p58_array_index_1087979_comb = p57_literal_1076351[p58_array_index_1087945_comb];
  assign p58_array_index_1087980_comb = p57_literal_1076353[p58_array_index_1087946_comb];
  assign p58_array_index_1087981_comb = p57_literal_1076355[p58_array_index_1087947_comb];
  assign p58_res7__305_comb = p58_array_index_1087976_comb ^ p58_array_index_1087977_comb ^ p58_array_index_1087978_comb ^ p58_array_index_1087979_comb ^ p58_array_index_1087980_comb ^ p58_array_index_1087981_comb ^ p58_array_index_1087948_comb ^ p57_literal_1076358[p58_array_index_1087965_comb] ^ p58_array_index_1087950_comb ^ p57_literal_1076355[p58_array_index_1087967_comb] ^ p57_literal_1076353[p58_array_index_1087952_comb] ^ p57_literal_1076351[p58_array_index_1087953_comb] ^ p57_literal_1076349[p58_array_index_1087954_comb] ^ p57_literal_1076347[p58_array_index_1087955_comb] ^ p57_literal_1076345[p58_array_index_1087956_comb] ^ p58_array_index_1087957_comb;
  assign p58_array_index_1087991_comb = p57_literal_1076347[p58_res7__304_comb];
  assign p58_array_index_1087992_comb = p57_literal_1076349[p58_array_index_1087943_comb];
  assign p58_array_index_1087993_comb = p57_literal_1076351[p58_array_index_1087944_comb];
  assign p58_array_index_1087994_comb = p57_literal_1076353[p58_array_index_1087945_comb];
  assign p58_array_index_1087995_comb = p57_literal_1076355[p58_array_index_1087946_comb];
  assign p58_res7__306_comb = p57_literal_1076345[p58_res7__305_comb] ^ p58_array_index_1087991_comb ^ p58_array_index_1087992_comb ^ p58_array_index_1087993_comb ^ p58_array_index_1087994_comb ^ p58_array_index_1087995_comb ^ p58_array_index_1087947_comb ^ p57_literal_1076358[p58_array_index_1087948_comb] ^ p58_array_index_1087965_comb ^ p57_literal_1076355[p58_array_index_1087950_comb] ^ p57_literal_1076353[p58_array_index_1087967_comb] ^ p57_literal_1076351[p58_array_index_1087952_comb] ^ p57_literal_1076349[p58_array_index_1087953_comb] ^ p57_literal_1076347[p58_array_index_1087954_comb] ^ p57_literal_1076345[p58_array_index_1087955_comb] ^ p58_array_index_1087956_comb;
  assign p58_array_index_1088005_comb = p57_literal_1076347[p58_res7__305_comb];
  assign p58_array_index_1088006_comb = p57_literal_1076349[p58_res7__304_comb];
  assign p58_array_index_1088007_comb = p57_literal_1076351[p58_array_index_1087943_comb];
  assign p58_array_index_1088008_comb = p57_literal_1076353[p58_array_index_1087944_comb];
  assign p58_array_index_1088009_comb = p57_literal_1076355[p58_array_index_1087945_comb];
  assign p58_res7__307_comb = p57_literal_1076345[p58_res7__306_comb] ^ p58_array_index_1088005_comb ^ p58_array_index_1088006_comb ^ p58_array_index_1088007_comb ^ p58_array_index_1088008_comb ^ p58_array_index_1088009_comb ^ p58_array_index_1087946_comb ^ p57_literal_1076358[p58_array_index_1087947_comb] ^ p58_array_index_1087948_comb ^ p57_literal_1076355[p58_array_index_1087965_comb] ^ p57_literal_1076353[p58_array_index_1087950_comb] ^ p57_literal_1076351[p58_array_index_1087967_comb] ^ p57_literal_1076349[p58_array_index_1087952_comb] ^ p57_literal_1076347[p58_array_index_1087953_comb] ^ p57_literal_1076345[p58_array_index_1087954_comb] ^ p58_array_index_1087955_comb;
  assign p58_array_index_1088020_comb = p57_literal_1076349[p58_res7__305_comb];
  assign p58_array_index_1088021_comb = p57_literal_1076351[p58_res7__304_comb];
  assign p58_array_index_1088022_comb = p57_literal_1076353[p58_array_index_1087943_comb];
  assign p58_array_index_1088023_comb = p57_literal_1076355[p58_array_index_1087944_comb];
  assign p58_res7__308_comb = p57_literal_1076345[p58_res7__307_comb] ^ p57_literal_1076347[p58_res7__306_comb] ^ p58_array_index_1088020_comb ^ p58_array_index_1088021_comb ^ p58_array_index_1088022_comb ^ p58_array_index_1088023_comb ^ p58_array_index_1087945_comb ^ p57_literal_1076358[p58_array_index_1087946_comb] ^ p58_array_index_1087947_comb ^ p58_array_index_1087964_comb ^ p57_literal_1076353[p58_array_index_1087965_comb] ^ p57_literal_1076351[p58_array_index_1087950_comb] ^ p57_literal_1076349[p58_array_index_1087967_comb] ^ p57_literal_1076347[p58_array_index_1087952_comb] ^ p57_literal_1076345[p58_array_index_1087953_comb] ^ p58_array_index_1087954_comb;

  // Registers for pipe stage 58:
  reg [127:0] p58_xor_1087336;
  reg [127:0] p58_xor_1087905;
  reg [7:0] p58_array_index_1087943;
  reg [7:0] p58_array_index_1087944;
  reg [7:0] p58_array_index_1087945;
  reg [7:0] p58_array_index_1087946;
  reg [7:0] p58_array_index_1087947;
  reg [7:0] p58_array_index_1087948;
  reg [7:0] p58_array_index_1087950;
  reg [7:0] p58_array_index_1087952;
  reg [7:0] p58_array_index_1087953;
  reg [7:0] p58_array_index_1087959;
  reg [7:0] p58_array_index_1087960;
  reg [7:0] p58_array_index_1087961;
  reg [7:0] p58_array_index_1087962;
  reg [7:0] p58_array_index_1087963;
  reg [7:0] p58_array_index_1087965;
  reg [7:0] p58_array_index_1087967;
  reg [7:0] p58_res7__304;
  reg [7:0] p58_array_index_1087976;
  reg [7:0] p58_array_index_1087977;
  reg [7:0] p58_array_index_1087978;
  reg [7:0] p58_array_index_1087979;
  reg [7:0] p58_array_index_1087980;
  reg [7:0] p58_array_index_1087981;
  reg [7:0] p58_res7__305;
  reg [7:0] p58_array_index_1087991;
  reg [7:0] p58_array_index_1087992;
  reg [7:0] p58_array_index_1087993;
  reg [7:0] p58_array_index_1087994;
  reg [7:0] p58_array_index_1087995;
  reg [7:0] p58_res7__306;
  reg [7:0] p58_array_index_1088005;
  reg [7:0] p58_array_index_1088006;
  reg [7:0] p58_array_index_1088007;
  reg [7:0] p58_array_index_1088008;
  reg [7:0] p58_array_index_1088009;
  reg [7:0] p58_res7__307;
  reg [7:0] p58_array_index_1088020;
  reg [7:0] p58_array_index_1088021;
  reg [7:0] p58_array_index_1088022;
  reg [7:0] p58_array_index_1088023;
  reg [7:0] p58_res7__308;
  reg [127:0] p58_res__37;
  reg [7:0] p59_arr[256];
  reg [7:0] p59_literal_1076345[256];
  reg [7:0] p59_literal_1076347[256];
  reg [7:0] p59_literal_1076349[256];
  reg [7:0] p59_literal_1076351[256];
  reg [7:0] p59_literal_1076353[256];
  reg [7:0] p59_literal_1076355[256];
  reg [7:0] p59_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p58_xor_1087336 <= p57_xor_1087336;
    p58_xor_1087905 <= p57_xor_1087905;
    p58_array_index_1087943 <= p58_array_index_1087943_comb;
    p58_array_index_1087944 <= p58_array_index_1087944_comb;
    p58_array_index_1087945 <= p58_array_index_1087945_comb;
    p58_array_index_1087946 <= p58_array_index_1087946_comb;
    p58_array_index_1087947 <= p58_array_index_1087947_comb;
    p58_array_index_1087948 <= p58_array_index_1087948_comb;
    p58_array_index_1087950 <= p58_array_index_1087950_comb;
    p58_array_index_1087952 <= p58_array_index_1087952_comb;
    p58_array_index_1087953 <= p58_array_index_1087953_comb;
    p58_array_index_1087959 <= p58_array_index_1087959_comb;
    p58_array_index_1087960 <= p58_array_index_1087960_comb;
    p58_array_index_1087961 <= p58_array_index_1087961_comb;
    p58_array_index_1087962 <= p58_array_index_1087962_comb;
    p58_array_index_1087963 <= p58_array_index_1087963_comb;
    p58_array_index_1087965 <= p58_array_index_1087965_comb;
    p58_array_index_1087967 <= p58_array_index_1087967_comb;
    p58_res7__304 <= p58_res7__304_comb;
    p58_array_index_1087976 <= p58_array_index_1087976_comb;
    p58_array_index_1087977 <= p58_array_index_1087977_comb;
    p58_array_index_1087978 <= p58_array_index_1087978_comb;
    p58_array_index_1087979 <= p58_array_index_1087979_comb;
    p58_array_index_1087980 <= p58_array_index_1087980_comb;
    p58_array_index_1087981 <= p58_array_index_1087981_comb;
    p58_res7__305 <= p58_res7__305_comb;
    p58_array_index_1087991 <= p58_array_index_1087991_comb;
    p58_array_index_1087992 <= p58_array_index_1087992_comb;
    p58_array_index_1087993 <= p58_array_index_1087993_comb;
    p58_array_index_1087994 <= p58_array_index_1087994_comb;
    p58_array_index_1087995 <= p58_array_index_1087995_comb;
    p58_res7__306 <= p58_res7__306_comb;
    p58_array_index_1088005 <= p58_array_index_1088005_comb;
    p58_array_index_1088006 <= p58_array_index_1088006_comb;
    p58_array_index_1088007 <= p58_array_index_1088007_comb;
    p58_array_index_1088008 <= p58_array_index_1088008_comb;
    p58_array_index_1088009 <= p58_array_index_1088009_comb;
    p58_res7__307 <= p58_res7__307_comb;
    p58_array_index_1088020 <= p58_array_index_1088020_comb;
    p58_array_index_1088021 <= p58_array_index_1088021_comb;
    p58_array_index_1088022 <= p58_array_index_1088022_comb;
    p58_array_index_1088023 <= p58_array_index_1088023_comb;
    p58_res7__308 <= p58_res7__308_comb;
    p58_res__37 <= p57_res__37;
    p59_arr <= p58_arr;
    p59_literal_1076345 <= p58_literal_1076345;
    p59_literal_1076347 <= p58_literal_1076347;
    p59_literal_1076349 <= p58_literal_1076349;
    p59_literal_1076351 <= p58_literal_1076351;
    p59_literal_1076353 <= p58_literal_1076353;
    p59_literal_1076355 <= p58_literal_1076355;
    p59_literal_1076358 <= p58_literal_1076358;
  end

  // ===== Pipe stage 59:
  wire [7:0] p59_array_index_1088137_comb;
  wire [7:0] p59_array_index_1088138_comb;
  wire [7:0] p59_array_index_1088139_comb;
  wire [7:0] p59_array_index_1088140_comb;
  wire [7:0] p59_res7__309_comb;
  wire [7:0] p59_array_index_1088151_comb;
  wire [7:0] p59_array_index_1088152_comb;
  wire [7:0] p59_array_index_1088153_comb;
  wire [7:0] p59_res7__310_comb;
  wire [7:0] p59_array_index_1088163_comb;
  wire [7:0] p59_array_index_1088164_comb;
  wire [7:0] p59_array_index_1088165_comb;
  wire [7:0] p59_res7__311_comb;
  wire [7:0] p59_array_index_1088176_comb;
  wire [7:0] p59_array_index_1088177_comb;
  wire [7:0] p59_res7__312_comb;
  wire [7:0] p59_array_index_1088187_comb;
  wire [7:0] p59_array_index_1088188_comb;
  wire [7:0] p59_res7__313_comb;
  wire [7:0] p59_array_index_1088194_comb;
  wire [7:0] p59_array_index_1088195_comb;
  wire [7:0] p59_array_index_1088196_comb;
  wire [7:0] p59_array_index_1088197_comb;
  wire [7:0] p59_array_index_1088198_comb;
  wire [7:0] p59_array_index_1088199_comb;
  wire [7:0] p59_array_index_1088200_comb;
  wire [7:0] p59_array_index_1088201_comb;
  wire [7:0] p59_array_index_1088202_comb;
  assign p59_array_index_1088137_comb = p58_literal_1076349[p58_res7__306];
  assign p59_array_index_1088138_comb = p58_literal_1076351[p58_res7__305];
  assign p59_array_index_1088139_comb = p58_literal_1076353[p58_res7__304];
  assign p59_array_index_1088140_comb = p58_literal_1076355[p58_array_index_1087943];
  assign p59_res7__309_comb = p58_literal_1076345[p58_res7__308] ^ p58_literal_1076347[p58_res7__307] ^ p59_array_index_1088137_comb ^ p59_array_index_1088138_comb ^ p59_array_index_1088139_comb ^ p59_array_index_1088140_comb ^ p58_array_index_1087944 ^ p58_literal_1076358[p58_array_index_1087945] ^ p58_array_index_1087946 ^ p58_array_index_1087981 ^ p58_literal_1076353[p58_array_index_1087948] ^ p58_literal_1076351[p58_array_index_1087965] ^ p58_literal_1076349[p58_array_index_1087950] ^ p58_literal_1076347[p58_array_index_1087967] ^ p58_literal_1076345[p58_array_index_1087952] ^ p58_array_index_1087953;
  assign p59_array_index_1088151_comb = p58_literal_1076351[p58_res7__306];
  assign p59_array_index_1088152_comb = p58_literal_1076353[p58_res7__305];
  assign p59_array_index_1088153_comb = p58_literal_1076355[p58_res7__304];
  assign p59_res7__310_comb = p58_literal_1076345[p59_res7__309_comb] ^ p58_literal_1076347[p58_res7__308] ^ p58_literal_1076349[p58_res7__307] ^ p59_array_index_1088151_comb ^ p59_array_index_1088152_comb ^ p59_array_index_1088153_comb ^ p58_array_index_1087943 ^ p58_literal_1076358[p58_array_index_1087944] ^ p58_array_index_1087945 ^ p58_array_index_1087995 ^ p58_array_index_1087963 ^ p58_literal_1076351[p58_array_index_1087948] ^ p58_literal_1076349[p58_array_index_1087965] ^ p58_literal_1076347[p58_array_index_1087950] ^ p58_literal_1076345[p58_array_index_1087967] ^ p58_array_index_1087952;
  assign p59_array_index_1088163_comb = p58_literal_1076351[p58_res7__307];
  assign p59_array_index_1088164_comb = p58_literal_1076353[p58_res7__306];
  assign p59_array_index_1088165_comb = p58_literal_1076355[p58_res7__305];
  assign p59_res7__311_comb = p58_literal_1076345[p59_res7__310_comb] ^ p58_literal_1076347[p59_res7__309_comb] ^ p58_literal_1076349[p58_res7__308] ^ p59_array_index_1088163_comb ^ p59_array_index_1088164_comb ^ p59_array_index_1088165_comb ^ p58_res7__304 ^ p58_literal_1076358[p58_array_index_1087943] ^ p58_array_index_1087944 ^ p58_array_index_1088009 ^ p58_array_index_1087980 ^ p58_literal_1076351[p58_array_index_1087947] ^ p58_literal_1076349[p58_array_index_1087948] ^ p58_literal_1076347[p58_array_index_1087965] ^ p58_literal_1076345[p58_array_index_1087950] ^ p58_array_index_1087967;
  assign p59_array_index_1088176_comb = p58_literal_1076353[p58_res7__307];
  assign p59_array_index_1088177_comb = p58_literal_1076355[p58_res7__306];
  assign p59_res7__312_comb = p58_literal_1076345[p59_res7__311_comb] ^ p58_literal_1076347[p59_res7__310_comb] ^ p58_literal_1076349[p59_res7__309_comb] ^ p58_literal_1076351[p58_res7__308] ^ p59_array_index_1088176_comb ^ p59_array_index_1088177_comb ^ p58_res7__305 ^ p58_literal_1076358[p58_res7__304] ^ p58_array_index_1087943 ^ p58_array_index_1088023 ^ p58_array_index_1087994 ^ p58_array_index_1087962 ^ p58_literal_1076349[p58_array_index_1087947] ^ p58_literal_1076347[p58_array_index_1087948] ^ p58_literal_1076345[p58_array_index_1087965] ^ p58_array_index_1087950;
  assign p59_array_index_1088187_comb = p58_literal_1076353[p58_res7__308];
  assign p59_array_index_1088188_comb = p58_literal_1076355[p58_res7__307];
  assign p59_res7__313_comb = p58_literal_1076345[p59_res7__312_comb] ^ p58_literal_1076347[p59_res7__311_comb] ^ p58_literal_1076349[p59_res7__310_comb] ^ p58_literal_1076351[p59_res7__309_comb] ^ p59_array_index_1088187_comb ^ p59_array_index_1088188_comb ^ p58_res7__306 ^ p58_literal_1076358[p58_res7__305] ^ p58_res7__304 ^ p59_array_index_1088140_comb ^ p58_array_index_1088008 ^ p58_array_index_1087979 ^ p58_literal_1076349[p58_array_index_1087946] ^ p58_literal_1076347[p58_array_index_1087947] ^ p58_literal_1076345[p58_array_index_1087948] ^ p58_array_index_1087965;
  assign p59_array_index_1088194_comb = p58_literal_1076345[p59_res7__313_comb];
  assign p59_array_index_1088195_comb = p58_literal_1076347[p59_res7__312_comb];
  assign p59_array_index_1088196_comb = p58_literal_1076349[p59_res7__311_comb];
  assign p59_array_index_1088197_comb = p58_literal_1076351[p59_res7__310_comb];
  assign p59_array_index_1088198_comb = p58_literal_1076353[p59_res7__309_comb];
  assign p59_array_index_1088199_comb = p58_literal_1076355[p58_res7__308];
  assign p59_array_index_1088200_comb = p58_literal_1076358[p58_res7__306];
  assign p59_array_index_1088201_comb = p58_literal_1076347[p58_array_index_1087946];
  assign p59_array_index_1088202_comb = p58_literal_1076345[p58_array_index_1087947];

  // Registers for pipe stage 59:
  reg [127:0] p59_xor_1087336;
  reg [127:0] p59_xor_1087905;
  reg [7:0] p59_array_index_1087943;
  reg [7:0] p59_array_index_1087944;
  reg [7:0] p59_array_index_1087945;
  reg [7:0] p59_array_index_1087946;
  reg [7:0] p59_array_index_1087947;
  reg [7:0] p59_array_index_1087948;
  reg [7:0] p59_array_index_1087959;
  reg [7:0] p59_array_index_1087960;
  reg [7:0] p59_array_index_1087961;
  reg [7:0] p59_res7__304;
  reg [7:0] p59_array_index_1087976;
  reg [7:0] p59_array_index_1087977;
  reg [7:0] p59_array_index_1087978;
  reg [7:0] p59_res7__305;
  reg [7:0] p59_array_index_1087991;
  reg [7:0] p59_array_index_1087992;
  reg [7:0] p59_array_index_1087993;
  reg [7:0] p59_res7__306;
  reg [7:0] p59_array_index_1088005;
  reg [7:0] p59_array_index_1088006;
  reg [7:0] p59_array_index_1088007;
  reg [7:0] p59_res7__307;
  reg [7:0] p59_array_index_1088020;
  reg [7:0] p59_array_index_1088021;
  reg [7:0] p59_array_index_1088022;
  reg [7:0] p59_res7__308;
  reg [7:0] p59_array_index_1088137;
  reg [7:0] p59_array_index_1088138;
  reg [7:0] p59_array_index_1088139;
  reg [7:0] p59_res7__309;
  reg [7:0] p59_array_index_1088151;
  reg [7:0] p59_array_index_1088152;
  reg [7:0] p59_array_index_1088153;
  reg [7:0] p59_res7__310;
  reg [7:0] p59_array_index_1088163;
  reg [7:0] p59_array_index_1088164;
  reg [7:0] p59_array_index_1088165;
  reg [7:0] p59_res7__311;
  reg [7:0] p59_array_index_1088176;
  reg [7:0] p59_array_index_1088177;
  reg [7:0] p59_res7__312;
  reg [7:0] p59_array_index_1088187;
  reg [7:0] p59_array_index_1088188;
  reg [7:0] p59_res7__313;
  reg [7:0] p59_array_index_1088194;
  reg [7:0] p59_array_index_1088195;
  reg [7:0] p59_array_index_1088196;
  reg [7:0] p59_array_index_1088197;
  reg [7:0] p59_array_index_1088198;
  reg [7:0] p59_array_index_1088199;
  reg [7:0] p59_array_index_1088200;
  reg [7:0] p59_array_index_1088201;
  reg [7:0] p59_array_index_1088202;
  reg [127:0] p59_res__37;
  reg [7:0] p60_arr[256];
  reg [7:0] p60_literal_1076345[256];
  reg [7:0] p60_literal_1076347[256];
  reg [7:0] p60_literal_1076349[256];
  reg [7:0] p60_literal_1076351[256];
  reg [7:0] p60_literal_1076353[256];
  reg [7:0] p60_literal_1076355[256];
  reg [7:0] p60_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p59_xor_1087336 <= p58_xor_1087336;
    p59_xor_1087905 <= p58_xor_1087905;
    p59_array_index_1087943 <= p58_array_index_1087943;
    p59_array_index_1087944 <= p58_array_index_1087944;
    p59_array_index_1087945 <= p58_array_index_1087945;
    p59_array_index_1087946 <= p58_array_index_1087946;
    p59_array_index_1087947 <= p58_array_index_1087947;
    p59_array_index_1087948 <= p58_array_index_1087948;
    p59_array_index_1087959 <= p58_array_index_1087959;
    p59_array_index_1087960 <= p58_array_index_1087960;
    p59_array_index_1087961 <= p58_array_index_1087961;
    p59_res7__304 <= p58_res7__304;
    p59_array_index_1087976 <= p58_array_index_1087976;
    p59_array_index_1087977 <= p58_array_index_1087977;
    p59_array_index_1087978 <= p58_array_index_1087978;
    p59_res7__305 <= p58_res7__305;
    p59_array_index_1087991 <= p58_array_index_1087991;
    p59_array_index_1087992 <= p58_array_index_1087992;
    p59_array_index_1087993 <= p58_array_index_1087993;
    p59_res7__306 <= p58_res7__306;
    p59_array_index_1088005 <= p58_array_index_1088005;
    p59_array_index_1088006 <= p58_array_index_1088006;
    p59_array_index_1088007 <= p58_array_index_1088007;
    p59_res7__307 <= p58_res7__307;
    p59_array_index_1088020 <= p58_array_index_1088020;
    p59_array_index_1088021 <= p58_array_index_1088021;
    p59_array_index_1088022 <= p58_array_index_1088022;
    p59_res7__308 <= p58_res7__308;
    p59_array_index_1088137 <= p59_array_index_1088137_comb;
    p59_array_index_1088138 <= p59_array_index_1088138_comb;
    p59_array_index_1088139 <= p59_array_index_1088139_comb;
    p59_res7__309 <= p59_res7__309_comb;
    p59_array_index_1088151 <= p59_array_index_1088151_comb;
    p59_array_index_1088152 <= p59_array_index_1088152_comb;
    p59_array_index_1088153 <= p59_array_index_1088153_comb;
    p59_res7__310 <= p59_res7__310_comb;
    p59_array_index_1088163 <= p59_array_index_1088163_comb;
    p59_array_index_1088164 <= p59_array_index_1088164_comb;
    p59_array_index_1088165 <= p59_array_index_1088165_comb;
    p59_res7__311 <= p59_res7__311_comb;
    p59_array_index_1088176 <= p59_array_index_1088176_comb;
    p59_array_index_1088177 <= p59_array_index_1088177_comb;
    p59_res7__312 <= p59_res7__312_comb;
    p59_array_index_1088187 <= p59_array_index_1088187_comb;
    p59_array_index_1088188 <= p59_array_index_1088188_comb;
    p59_res7__313 <= p59_res7__313_comb;
    p59_array_index_1088194 <= p59_array_index_1088194_comb;
    p59_array_index_1088195 <= p59_array_index_1088195_comb;
    p59_array_index_1088196 <= p59_array_index_1088196_comb;
    p59_array_index_1088197 <= p59_array_index_1088197_comb;
    p59_array_index_1088198 <= p59_array_index_1088198_comb;
    p59_array_index_1088199 <= p59_array_index_1088199_comb;
    p59_array_index_1088200 <= p59_array_index_1088200_comb;
    p59_array_index_1088201 <= p59_array_index_1088201_comb;
    p59_array_index_1088202 <= p59_array_index_1088202_comb;
    p59_res__37 <= p58_res__37;
    p60_arr <= p59_arr;
    p60_literal_1076345 <= p59_literal_1076345;
    p60_literal_1076347 <= p59_literal_1076347;
    p60_literal_1076349 <= p59_literal_1076349;
    p60_literal_1076351 <= p59_literal_1076351;
    p60_literal_1076353 <= p59_literal_1076353;
    p60_literal_1076355 <= p59_literal_1076355;
    p60_literal_1076358 <= p59_literal_1076358;
  end

  // ===== Pipe stage 60:
  wire [7:0] p60_res7__314_comb;
  wire [7:0] p60_array_index_1088337_comb;
  wire [7:0] p60_res7__315_comb;
  wire [7:0] p60_res7__316_comb;
  wire [7:0] p60_res7__317_comb;
  wire [7:0] p60_res7__318_comb;
  wire [7:0] p60_res7__319_comb;
  wire [127:0] p60_res__19_comb;
  wire [127:0] p60_xor_1088377_comb;
  assign p60_res7__314_comb = p59_array_index_1088194 ^ p59_array_index_1088195 ^ p59_array_index_1088196 ^ p59_array_index_1088197 ^ p59_array_index_1088198 ^ p59_array_index_1088199 ^ p59_res7__307 ^ p59_array_index_1088200 ^ p59_res7__305 ^ p59_array_index_1088153 ^ p59_array_index_1088022 ^ p59_array_index_1087993 ^ p59_array_index_1087961 ^ p59_array_index_1088201 ^ p59_array_index_1088202 ^ p59_array_index_1087948;
  assign p60_array_index_1088337_comb = p59_literal_1076355[p59_res7__309];
  assign p60_res7__315_comb = p59_literal_1076345[p60_res7__314_comb] ^ p59_literal_1076347[p59_res7__313] ^ p59_literal_1076349[p59_res7__312] ^ p59_literal_1076351[p59_res7__311] ^ p59_literal_1076353[p59_res7__310] ^ p60_array_index_1088337_comb ^ p59_res7__308 ^ p59_literal_1076358[p59_res7__307] ^ p59_res7__306 ^ p59_array_index_1088165 ^ p59_array_index_1088139 ^ p59_array_index_1088007 ^ p59_array_index_1087978 ^ p59_literal_1076347[p59_array_index_1087945] ^ p59_literal_1076345[p59_array_index_1087946] ^ p59_array_index_1087947;
  assign p60_res7__316_comb = p59_literal_1076345[p60_res7__315_comb] ^ p59_literal_1076347[p60_res7__314_comb] ^ p59_literal_1076349[p59_res7__313] ^ p59_literal_1076351[p59_res7__312] ^ p59_literal_1076353[p59_res7__311] ^ p59_literal_1076355[p59_res7__310] ^ p59_res7__309 ^ p59_literal_1076358[p59_res7__308] ^ p59_res7__307 ^ p59_array_index_1088177 ^ p59_array_index_1088152 ^ p59_array_index_1088021 ^ p59_array_index_1087992 ^ p59_array_index_1087960 ^ p59_literal_1076345[p59_array_index_1087945] ^ p59_array_index_1087946;
  assign p60_res7__317_comb = p59_literal_1076345[p60_res7__316_comb] ^ p59_literal_1076347[p60_res7__315_comb] ^ p59_literal_1076349[p60_res7__314_comb] ^ p59_literal_1076351[p59_res7__313] ^ p59_literal_1076353[p59_res7__312] ^ p59_literal_1076355[p59_res7__311] ^ p59_res7__310 ^ p59_literal_1076358[p59_res7__309] ^ p59_res7__308 ^ p59_array_index_1088188 ^ p59_array_index_1088164 ^ p59_array_index_1088138 ^ p59_array_index_1088006 ^ p59_array_index_1087977 ^ p59_literal_1076345[p59_array_index_1087944] ^ p59_array_index_1087945;
  assign p60_res7__318_comb = p59_literal_1076345[p60_res7__317_comb] ^ p59_literal_1076347[p60_res7__316_comb] ^ p59_literal_1076349[p60_res7__315_comb] ^ p59_literal_1076351[p60_res7__314_comb] ^ p59_literal_1076353[p59_res7__313] ^ p59_literal_1076355[p59_res7__312] ^ p59_res7__311 ^ p59_literal_1076358[p59_res7__310] ^ p59_res7__309 ^ p59_array_index_1088199 ^ p59_array_index_1088176 ^ p59_array_index_1088151 ^ p59_array_index_1088020 ^ p59_array_index_1087991 ^ p59_array_index_1087959 ^ p59_array_index_1087944;
  assign p60_res7__319_comb = p59_literal_1076345[p60_res7__318_comb] ^ p59_literal_1076347[p60_res7__317_comb] ^ p59_literal_1076349[p60_res7__316_comb] ^ p59_literal_1076351[p60_res7__315_comb] ^ p59_literal_1076353[p60_res7__314_comb] ^ p59_literal_1076355[p59_res7__313] ^ p59_res7__312 ^ p59_literal_1076358[p59_res7__311] ^ p59_res7__310 ^ p60_array_index_1088337_comb ^ p59_array_index_1088187 ^ p59_array_index_1088163 ^ p59_array_index_1088137 ^ p59_array_index_1088005 ^ p59_array_index_1087976 ^ p59_array_index_1087943;
  assign p60_res__19_comb = {p60_res7__319_comb, p60_res7__318_comb, p60_res7__317_comb, p60_res7__316_comb, p60_res7__315_comb, p60_res7__314_comb, p59_res7__313, p59_res7__312, p59_res7__311, p59_res7__310, p59_res7__309, p59_res7__308, p59_res7__307, p59_res7__306, p59_res7__305, p59_res7__304};
  assign p60_xor_1088377_comb = p60_res__19_comb ^ p59_xor_1087336;

  // Registers for pipe stage 60:
  reg [127:0] p60_xor_1087905;
  reg [127:0] p60_xor_1088377;
  reg [127:0] p60_res__37;
  reg [7:0] p61_arr[256];
  reg [7:0] p61_literal_1076345[256];
  reg [7:0] p61_literal_1076347[256];
  reg [7:0] p61_literal_1076349[256];
  reg [7:0] p61_literal_1076351[256];
  reg [7:0] p61_literal_1076353[256];
  reg [7:0] p61_literal_1076355[256];
  reg [7:0] p61_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p60_xor_1087905 <= p59_xor_1087905;
    p60_xor_1088377 <= p60_xor_1088377_comb;
    p60_res__37 <= p59_res__37;
    p61_arr <= p60_arr;
    p61_literal_1076345 <= p60_literal_1076345;
    p61_literal_1076347 <= p60_literal_1076347;
    p61_literal_1076349 <= p60_literal_1076349;
    p61_literal_1076351 <= p60_literal_1076351;
    p61_literal_1076353 <= p60_literal_1076353;
    p61_literal_1076355 <= p60_literal_1076355;
    p61_literal_1076358 <= p60_literal_1076358;
  end

  // ===== Pipe stage 61:
  wire [127:0] p61_addedKey__61_comb;
  wire [7:0] p61_array_index_1088415_comb;
  wire [7:0] p61_array_index_1088416_comb;
  wire [7:0] p61_array_index_1088417_comb;
  wire [7:0] p61_array_index_1088418_comb;
  wire [7:0] p61_array_index_1088419_comb;
  wire [7:0] p61_array_index_1088420_comb;
  wire [7:0] p61_array_index_1088422_comb;
  wire [7:0] p61_array_index_1088424_comb;
  wire [7:0] p61_array_index_1088425_comb;
  wire [7:0] p61_array_index_1088426_comb;
  wire [7:0] p61_array_index_1088427_comb;
  wire [7:0] p61_array_index_1088428_comb;
  wire [7:0] p61_array_index_1088429_comb;
  wire [7:0] p61_array_index_1088431_comb;
  wire [7:0] p61_array_index_1088432_comb;
  wire [7:0] p61_array_index_1088433_comb;
  wire [7:0] p61_array_index_1088434_comb;
  wire [7:0] p61_array_index_1088435_comb;
  wire [7:0] p61_array_index_1088436_comb;
  wire [7:0] p61_array_index_1088437_comb;
  wire [7:0] p61_array_index_1088439_comb;
  wire [7:0] p61_res7__320_comb;
  wire [7:0] p61_array_index_1088448_comb;
  wire [7:0] p61_array_index_1088449_comb;
  wire [7:0] p61_array_index_1088450_comb;
  wire [7:0] p61_array_index_1088451_comb;
  wire [7:0] p61_array_index_1088452_comb;
  wire [7:0] p61_array_index_1088453_comb;
  wire [7:0] p61_res7__321_comb;
  wire [7:0] p61_array_index_1088463_comb;
  wire [7:0] p61_array_index_1088464_comb;
  wire [7:0] p61_array_index_1088465_comb;
  wire [7:0] p61_array_index_1088466_comb;
  wire [7:0] p61_array_index_1088467_comb;
  wire [7:0] p61_res7__322_comb;
  wire [7:0] p61_array_index_1088477_comb;
  wire [7:0] p61_array_index_1088478_comb;
  wire [7:0] p61_array_index_1088479_comb;
  wire [7:0] p61_array_index_1088480_comb;
  wire [7:0] p61_array_index_1088481_comb;
  wire [7:0] p61_res7__323_comb;
  wire [7:0] p61_array_index_1088492_comb;
  wire [7:0] p61_array_index_1088493_comb;
  wire [7:0] p61_array_index_1088494_comb;
  wire [7:0] p61_array_index_1088495_comb;
  wire [7:0] p61_res7__324_comb;
  assign p61_addedKey__61_comb = p60_xor_1088377 ^ 128'h3add_0155_10a1_fdcc_738e_8d93_6146_d515;
  assign p61_array_index_1088415_comb = p60_arr[p61_addedKey__61_comb[127:120]];
  assign p61_array_index_1088416_comb = p60_arr[p61_addedKey__61_comb[119:112]];
  assign p61_array_index_1088417_comb = p60_arr[p61_addedKey__61_comb[111:104]];
  assign p61_array_index_1088418_comb = p60_arr[p61_addedKey__61_comb[103:96]];
  assign p61_array_index_1088419_comb = p60_arr[p61_addedKey__61_comb[95:88]];
  assign p61_array_index_1088420_comb = p60_arr[p61_addedKey__61_comb[87:80]];
  assign p61_array_index_1088422_comb = p60_arr[p61_addedKey__61_comb[71:64]];
  assign p61_array_index_1088424_comb = p60_arr[p61_addedKey__61_comb[55:48]];
  assign p61_array_index_1088425_comb = p60_arr[p61_addedKey__61_comb[47:40]];
  assign p61_array_index_1088426_comb = p60_arr[p61_addedKey__61_comb[39:32]];
  assign p61_array_index_1088427_comb = p60_arr[p61_addedKey__61_comb[31:24]];
  assign p61_array_index_1088428_comb = p60_arr[p61_addedKey__61_comb[23:16]];
  assign p61_array_index_1088429_comb = p60_arr[p61_addedKey__61_comb[15:8]];
  assign p61_array_index_1088431_comb = p60_literal_1076345[p61_array_index_1088415_comb];
  assign p61_array_index_1088432_comb = p60_literal_1076347[p61_array_index_1088416_comb];
  assign p61_array_index_1088433_comb = p60_literal_1076349[p61_array_index_1088417_comb];
  assign p61_array_index_1088434_comb = p60_literal_1076351[p61_array_index_1088418_comb];
  assign p61_array_index_1088435_comb = p60_literal_1076353[p61_array_index_1088419_comb];
  assign p61_array_index_1088436_comb = p60_literal_1076355[p61_array_index_1088420_comb];
  assign p61_array_index_1088437_comb = p60_arr[p61_addedKey__61_comb[79:72]];
  assign p61_array_index_1088439_comb = p60_arr[p61_addedKey__61_comb[63:56]];
  assign p61_res7__320_comb = p61_array_index_1088431_comb ^ p61_array_index_1088432_comb ^ p61_array_index_1088433_comb ^ p61_array_index_1088434_comb ^ p61_array_index_1088435_comb ^ p61_array_index_1088436_comb ^ p61_array_index_1088437_comb ^ p60_literal_1076358[p61_array_index_1088422_comb] ^ p61_array_index_1088439_comb ^ p60_literal_1076355[p61_array_index_1088424_comb] ^ p60_literal_1076353[p61_array_index_1088425_comb] ^ p60_literal_1076351[p61_array_index_1088426_comb] ^ p60_literal_1076349[p61_array_index_1088427_comb] ^ p60_literal_1076347[p61_array_index_1088428_comb] ^ p60_literal_1076345[p61_array_index_1088429_comb] ^ p60_arr[p61_addedKey__61_comb[7:0]];
  assign p61_array_index_1088448_comb = p60_literal_1076345[p61_res7__320_comb];
  assign p61_array_index_1088449_comb = p60_literal_1076347[p61_array_index_1088415_comb];
  assign p61_array_index_1088450_comb = p60_literal_1076349[p61_array_index_1088416_comb];
  assign p61_array_index_1088451_comb = p60_literal_1076351[p61_array_index_1088417_comb];
  assign p61_array_index_1088452_comb = p60_literal_1076353[p61_array_index_1088418_comb];
  assign p61_array_index_1088453_comb = p60_literal_1076355[p61_array_index_1088419_comb];
  assign p61_res7__321_comb = p61_array_index_1088448_comb ^ p61_array_index_1088449_comb ^ p61_array_index_1088450_comb ^ p61_array_index_1088451_comb ^ p61_array_index_1088452_comb ^ p61_array_index_1088453_comb ^ p61_array_index_1088420_comb ^ p60_literal_1076358[p61_array_index_1088437_comb] ^ p61_array_index_1088422_comb ^ p60_literal_1076355[p61_array_index_1088439_comb] ^ p60_literal_1076353[p61_array_index_1088424_comb] ^ p60_literal_1076351[p61_array_index_1088425_comb] ^ p60_literal_1076349[p61_array_index_1088426_comb] ^ p60_literal_1076347[p61_array_index_1088427_comb] ^ p60_literal_1076345[p61_array_index_1088428_comb] ^ p61_array_index_1088429_comb;
  assign p61_array_index_1088463_comb = p60_literal_1076347[p61_res7__320_comb];
  assign p61_array_index_1088464_comb = p60_literal_1076349[p61_array_index_1088415_comb];
  assign p61_array_index_1088465_comb = p60_literal_1076351[p61_array_index_1088416_comb];
  assign p61_array_index_1088466_comb = p60_literal_1076353[p61_array_index_1088417_comb];
  assign p61_array_index_1088467_comb = p60_literal_1076355[p61_array_index_1088418_comb];
  assign p61_res7__322_comb = p60_literal_1076345[p61_res7__321_comb] ^ p61_array_index_1088463_comb ^ p61_array_index_1088464_comb ^ p61_array_index_1088465_comb ^ p61_array_index_1088466_comb ^ p61_array_index_1088467_comb ^ p61_array_index_1088419_comb ^ p60_literal_1076358[p61_array_index_1088420_comb] ^ p61_array_index_1088437_comb ^ p60_literal_1076355[p61_array_index_1088422_comb] ^ p60_literal_1076353[p61_array_index_1088439_comb] ^ p60_literal_1076351[p61_array_index_1088424_comb] ^ p60_literal_1076349[p61_array_index_1088425_comb] ^ p60_literal_1076347[p61_array_index_1088426_comb] ^ p60_literal_1076345[p61_array_index_1088427_comb] ^ p61_array_index_1088428_comb;
  assign p61_array_index_1088477_comb = p60_literal_1076347[p61_res7__321_comb];
  assign p61_array_index_1088478_comb = p60_literal_1076349[p61_res7__320_comb];
  assign p61_array_index_1088479_comb = p60_literal_1076351[p61_array_index_1088415_comb];
  assign p61_array_index_1088480_comb = p60_literal_1076353[p61_array_index_1088416_comb];
  assign p61_array_index_1088481_comb = p60_literal_1076355[p61_array_index_1088417_comb];
  assign p61_res7__323_comb = p60_literal_1076345[p61_res7__322_comb] ^ p61_array_index_1088477_comb ^ p61_array_index_1088478_comb ^ p61_array_index_1088479_comb ^ p61_array_index_1088480_comb ^ p61_array_index_1088481_comb ^ p61_array_index_1088418_comb ^ p60_literal_1076358[p61_array_index_1088419_comb] ^ p61_array_index_1088420_comb ^ p60_literal_1076355[p61_array_index_1088437_comb] ^ p60_literal_1076353[p61_array_index_1088422_comb] ^ p60_literal_1076351[p61_array_index_1088439_comb] ^ p60_literal_1076349[p61_array_index_1088424_comb] ^ p60_literal_1076347[p61_array_index_1088425_comb] ^ p60_literal_1076345[p61_array_index_1088426_comb] ^ p61_array_index_1088427_comb;
  assign p61_array_index_1088492_comb = p60_literal_1076349[p61_res7__321_comb];
  assign p61_array_index_1088493_comb = p60_literal_1076351[p61_res7__320_comb];
  assign p61_array_index_1088494_comb = p60_literal_1076353[p61_array_index_1088415_comb];
  assign p61_array_index_1088495_comb = p60_literal_1076355[p61_array_index_1088416_comb];
  assign p61_res7__324_comb = p60_literal_1076345[p61_res7__323_comb] ^ p60_literal_1076347[p61_res7__322_comb] ^ p61_array_index_1088492_comb ^ p61_array_index_1088493_comb ^ p61_array_index_1088494_comb ^ p61_array_index_1088495_comb ^ p61_array_index_1088417_comb ^ p60_literal_1076358[p61_array_index_1088418_comb] ^ p61_array_index_1088419_comb ^ p61_array_index_1088436_comb ^ p60_literal_1076353[p61_array_index_1088437_comb] ^ p60_literal_1076351[p61_array_index_1088422_comb] ^ p60_literal_1076349[p61_array_index_1088439_comb] ^ p60_literal_1076347[p61_array_index_1088424_comb] ^ p60_literal_1076345[p61_array_index_1088425_comb] ^ p61_array_index_1088426_comb;

  // Registers for pipe stage 61:
  reg [127:0] p61_xor_1087905;
  reg [127:0] p61_xor_1088377;
  reg [7:0] p61_array_index_1088415;
  reg [7:0] p61_array_index_1088416;
  reg [7:0] p61_array_index_1088417;
  reg [7:0] p61_array_index_1088418;
  reg [7:0] p61_array_index_1088419;
  reg [7:0] p61_array_index_1088420;
  reg [7:0] p61_array_index_1088422;
  reg [7:0] p61_array_index_1088424;
  reg [7:0] p61_array_index_1088425;
  reg [7:0] p61_array_index_1088431;
  reg [7:0] p61_array_index_1088432;
  reg [7:0] p61_array_index_1088433;
  reg [7:0] p61_array_index_1088434;
  reg [7:0] p61_array_index_1088435;
  reg [7:0] p61_array_index_1088437;
  reg [7:0] p61_array_index_1088439;
  reg [7:0] p61_res7__320;
  reg [7:0] p61_array_index_1088448;
  reg [7:0] p61_array_index_1088449;
  reg [7:0] p61_array_index_1088450;
  reg [7:0] p61_array_index_1088451;
  reg [7:0] p61_array_index_1088452;
  reg [7:0] p61_array_index_1088453;
  reg [7:0] p61_res7__321;
  reg [7:0] p61_array_index_1088463;
  reg [7:0] p61_array_index_1088464;
  reg [7:0] p61_array_index_1088465;
  reg [7:0] p61_array_index_1088466;
  reg [7:0] p61_array_index_1088467;
  reg [7:0] p61_res7__322;
  reg [7:0] p61_array_index_1088477;
  reg [7:0] p61_array_index_1088478;
  reg [7:0] p61_array_index_1088479;
  reg [7:0] p61_array_index_1088480;
  reg [7:0] p61_array_index_1088481;
  reg [7:0] p61_res7__323;
  reg [7:0] p61_array_index_1088492;
  reg [7:0] p61_array_index_1088493;
  reg [7:0] p61_array_index_1088494;
  reg [7:0] p61_array_index_1088495;
  reg [7:0] p61_res7__324;
  reg [127:0] p61_res__37;
  reg [7:0] p62_arr[256];
  reg [7:0] p62_literal_1076345[256];
  reg [7:0] p62_literal_1076347[256];
  reg [7:0] p62_literal_1076349[256];
  reg [7:0] p62_literal_1076351[256];
  reg [7:0] p62_literal_1076353[256];
  reg [7:0] p62_literal_1076355[256];
  reg [7:0] p62_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p61_xor_1087905 <= p60_xor_1087905;
    p61_xor_1088377 <= p60_xor_1088377;
    p61_array_index_1088415 <= p61_array_index_1088415_comb;
    p61_array_index_1088416 <= p61_array_index_1088416_comb;
    p61_array_index_1088417 <= p61_array_index_1088417_comb;
    p61_array_index_1088418 <= p61_array_index_1088418_comb;
    p61_array_index_1088419 <= p61_array_index_1088419_comb;
    p61_array_index_1088420 <= p61_array_index_1088420_comb;
    p61_array_index_1088422 <= p61_array_index_1088422_comb;
    p61_array_index_1088424 <= p61_array_index_1088424_comb;
    p61_array_index_1088425 <= p61_array_index_1088425_comb;
    p61_array_index_1088431 <= p61_array_index_1088431_comb;
    p61_array_index_1088432 <= p61_array_index_1088432_comb;
    p61_array_index_1088433 <= p61_array_index_1088433_comb;
    p61_array_index_1088434 <= p61_array_index_1088434_comb;
    p61_array_index_1088435 <= p61_array_index_1088435_comb;
    p61_array_index_1088437 <= p61_array_index_1088437_comb;
    p61_array_index_1088439 <= p61_array_index_1088439_comb;
    p61_res7__320 <= p61_res7__320_comb;
    p61_array_index_1088448 <= p61_array_index_1088448_comb;
    p61_array_index_1088449 <= p61_array_index_1088449_comb;
    p61_array_index_1088450 <= p61_array_index_1088450_comb;
    p61_array_index_1088451 <= p61_array_index_1088451_comb;
    p61_array_index_1088452 <= p61_array_index_1088452_comb;
    p61_array_index_1088453 <= p61_array_index_1088453_comb;
    p61_res7__321 <= p61_res7__321_comb;
    p61_array_index_1088463 <= p61_array_index_1088463_comb;
    p61_array_index_1088464 <= p61_array_index_1088464_comb;
    p61_array_index_1088465 <= p61_array_index_1088465_comb;
    p61_array_index_1088466 <= p61_array_index_1088466_comb;
    p61_array_index_1088467 <= p61_array_index_1088467_comb;
    p61_res7__322 <= p61_res7__322_comb;
    p61_array_index_1088477 <= p61_array_index_1088477_comb;
    p61_array_index_1088478 <= p61_array_index_1088478_comb;
    p61_array_index_1088479 <= p61_array_index_1088479_comb;
    p61_array_index_1088480 <= p61_array_index_1088480_comb;
    p61_array_index_1088481 <= p61_array_index_1088481_comb;
    p61_res7__323 <= p61_res7__323_comb;
    p61_array_index_1088492 <= p61_array_index_1088492_comb;
    p61_array_index_1088493 <= p61_array_index_1088493_comb;
    p61_array_index_1088494 <= p61_array_index_1088494_comb;
    p61_array_index_1088495 <= p61_array_index_1088495_comb;
    p61_res7__324 <= p61_res7__324_comb;
    p61_res__37 <= p60_res__37;
    p62_arr <= p61_arr;
    p62_literal_1076345 <= p61_literal_1076345;
    p62_literal_1076347 <= p61_literal_1076347;
    p62_literal_1076349 <= p61_literal_1076349;
    p62_literal_1076351 <= p61_literal_1076351;
    p62_literal_1076353 <= p61_literal_1076353;
    p62_literal_1076355 <= p61_literal_1076355;
    p62_literal_1076358 <= p61_literal_1076358;
  end

  // ===== Pipe stage 62:
  wire [7:0] p62_array_index_1088609_comb;
  wire [7:0] p62_array_index_1088610_comb;
  wire [7:0] p62_array_index_1088611_comb;
  wire [7:0] p62_array_index_1088612_comb;
  wire [7:0] p62_res7__325_comb;
  wire [7:0] p62_array_index_1088623_comb;
  wire [7:0] p62_array_index_1088624_comb;
  wire [7:0] p62_array_index_1088625_comb;
  wire [7:0] p62_res7__326_comb;
  wire [7:0] p62_array_index_1088635_comb;
  wire [7:0] p62_array_index_1088636_comb;
  wire [7:0] p62_array_index_1088637_comb;
  wire [7:0] p62_res7__327_comb;
  wire [7:0] p62_array_index_1088648_comb;
  wire [7:0] p62_array_index_1088649_comb;
  wire [7:0] p62_res7__328_comb;
  wire [7:0] p62_array_index_1088659_comb;
  wire [7:0] p62_array_index_1088660_comb;
  wire [7:0] p62_res7__329_comb;
  wire [7:0] p62_array_index_1088666_comb;
  wire [7:0] p62_array_index_1088667_comb;
  wire [7:0] p62_array_index_1088668_comb;
  wire [7:0] p62_array_index_1088669_comb;
  wire [7:0] p62_array_index_1088670_comb;
  wire [7:0] p62_array_index_1088671_comb;
  wire [7:0] p62_array_index_1088672_comb;
  wire [7:0] p62_array_index_1088673_comb;
  wire [7:0] p62_array_index_1088674_comb;
  assign p62_array_index_1088609_comb = p61_literal_1076349[p61_res7__322];
  assign p62_array_index_1088610_comb = p61_literal_1076351[p61_res7__321];
  assign p62_array_index_1088611_comb = p61_literal_1076353[p61_res7__320];
  assign p62_array_index_1088612_comb = p61_literal_1076355[p61_array_index_1088415];
  assign p62_res7__325_comb = p61_literal_1076345[p61_res7__324] ^ p61_literal_1076347[p61_res7__323] ^ p62_array_index_1088609_comb ^ p62_array_index_1088610_comb ^ p62_array_index_1088611_comb ^ p62_array_index_1088612_comb ^ p61_array_index_1088416 ^ p61_literal_1076358[p61_array_index_1088417] ^ p61_array_index_1088418 ^ p61_array_index_1088453 ^ p61_literal_1076353[p61_array_index_1088420] ^ p61_literal_1076351[p61_array_index_1088437] ^ p61_literal_1076349[p61_array_index_1088422] ^ p61_literal_1076347[p61_array_index_1088439] ^ p61_literal_1076345[p61_array_index_1088424] ^ p61_array_index_1088425;
  assign p62_array_index_1088623_comb = p61_literal_1076351[p61_res7__322];
  assign p62_array_index_1088624_comb = p61_literal_1076353[p61_res7__321];
  assign p62_array_index_1088625_comb = p61_literal_1076355[p61_res7__320];
  assign p62_res7__326_comb = p61_literal_1076345[p62_res7__325_comb] ^ p61_literal_1076347[p61_res7__324] ^ p61_literal_1076349[p61_res7__323] ^ p62_array_index_1088623_comb ^ p62_array_index_1088624_comb ^ p62_array_index_1088625_comb ^ p61_array_index_1088415 ^ p61_literal_1076358[p61_array_index_1088416] ^ p61_array_index_1088417 ^ p61_array_index_1088467 ^ p61_array_index_1088435 ^ p61_literal_1076351[p61_array_index_1088420] ^ p61_literal_1076349[p61_array_index_1088437] ^ p61_literal_1076347[p61_array_index_1088422] ^ p61_literal_1076345[p61_array_index_1088439] ^ p61_array_index_1088424;
  assign p62_array_index_1088635_comb = p61_literal_1076351[p61_res7__323];
  assign p62_array_index_1088636_comb = p61_literal_1076353[p61_res7__322];
  assign p62_array_index_1088637_comb = p61_literal_1076355[p61_res7__321];
  assign p62_res7__327_comb = p61_literal_1076345[p62_res7__326_comb] ^ p61_literal_1076347[p62_res7__325_comb] ^ p61_literal_1076349[p61_res7__324] ^ p62_array_index_1088635_comb ^ p62_array_index_1088636_comb ^ p62_array_index_1088637_comb ^ p61_res7__320 ^ p61_literal_1076358[p61_array_index_1088415] ^ p61_array_index_1088416 ^ p61_array_index_1088481 ^ p61_array_index_1088452 ^ p61_literal_1076351[p61_array_index_1088419] ^ p61_literal_1076349[p61_array_index_1088420] ^ p61_literal_1076347[p61_array_index_1088437] ^ p61_literal_1076345[p61_array_index_1088422] ^ p61_array_index_1088439;
  assign p62_array_index_1088648_comb = p61_literal_1076353[p61_res7__323];
  assign p62_array_index_1088649_comb = p61_literal_1076355[p61_res7__322];
  assign p62_res7__328_comb = p61_literal_1076345[p62_res7__327_comb] ^ p61_literal_1076347[p62_res7__326_comb] ^ p61_literal_1076349[p62_res7__325_comb] ^ p61_literal_1076351[p61_res7__324] ^ p62_array_index_1088648_comb ^ p62_array_index_1088649_comb ^ p61_res7__321 ^ p61_literal_1076358[p61_res7__320] ^ p61_array_index_1088415 ^ p61_array_index_1088495 ^ p61_array_index_1088466 ^ p61_array_index_1088434 ^ p61_literal_1076349[p61_array_index_1088419] ^ p61_literal_1076347[p61_array_index_1088420] ^ p61_literal_1076345[p61_array_index_1088437] ^ p61_array_index_1088422;
  assign p62_array_index_1088659_comb = p61_literal_1076353[p61_res7__324];
  assign p62_array_index_1088660_comb = p61_literal_1076355[p61_res7__323];
  assign p62_res7__329_comb = p61_literal_1076345[p62_res7__328_comb] ^ p61_literal_1076347[p62_res7__327_comb] ^ p61_literal_1076349[p62_res7__326_comb] ^ p61_literal_1076351[p62_res7__325_comb] ^ p62_array_index_1088659_comb ^ p62_array_index_1088660_comb ^ p61_res7__322 ^ p61_literal_1076358[p61_res7__321] ^ p61_res7__320 ^ p62_array_index_1088612_comb ^ p61_array_index_1088480 ^ p61_array_index_1088451 ^ p61_literal_1076349[p61_array_index_1088418] ^ p61_literal_1076347[p61_array_index_1088419] ^ p61_literal_1076345[p61_array_index_1088420] ^ p61_array_index_1088437;
  assign p62_array_index_1088666_comb = p61_literal_1076345[p62_res7__329_comb];
  assign p62_array_index_1088667_comb = p61_literal_1076347[p62_res7__328_comb];
  assign p62_array_index_1088668_comb = p61_literal_1076349[p62_res7__327_comb];
  assign p62_array_index_1088669_comb = p61_literal_1076351[p62_res7__326_comb];
  assign p62_array_index_1088670_comb = p61_literal_1076353[p62_res7__325_comb];
  assign p62_array_index_1088671_comb = p61_literal_1076355[p61_res7__324];
  assign p62_array_index_1088672_comb = p61_literal_1076358[p61_res7__322];
  assign p62_array_index_1088673_comb = p61_literal_1076347[p61_array_index_1088418];
  assign p62_array_index_1088674_comb = p61_literal_1076345[p61_array_index_1088419];

  // Registers for pipe stage 62:
  reg [127:0] p62_xor_1087905;
  reg [127:0] p62_xor_1088377;
  reg [7:0] p62_array_index_1088415;
  reg [7:0] p62_array_index_1088416;
  reg [7:0] p62_array_index_1088417;
  reg [7:0] p62_array_index_1088418;
  reg [7:0] p62_array_index_1088419;
  reg [7:0] p62_array_index_1088420;
  reg [7:0] p62_array_index_1088431;
  reg [7:0] p62_array_index_1088432;
  reg [7:0] p62_array_index_1088433;
  reg [7:0] p62_res7__320;
  reg [7:0] p62_array_index_1088448;
  reg [7:0] p62_array_index_1088449;
  reg [7:0] p62_array_index_1088450;
  reg [7:0] p62_res7__321;
  reg [7:0] p62_array_index_1088463;
  reg [7:0] p62_array_index_1088464;
  reg [7:0] p62_array_index_1088465;
  reg [7:0] p62_res7__322;
  reg [7:0] p62_array_index_1088477;
  reg [7:0] p62_array_index_1088478;
  reg [7:0] p62_array_index_1088479;
  reg [7:0] p62_res7__323;
  reg [7:0] p62_array_index_1088492;
  reg [7:0] p62_array_index_1088493;
  reg [7:0] p62_array_index_1088494;
  reg [7:0] p62_res7__324;
  reg [7:0] p62_array_index_1088609;
  reg [7:0] p62_array_index_1088610;
  reg [7:0] p62_array_index_1088611;
  reg [7:0] p62_res7__325;
  reg [7:0] p62_array_index_1088623;
  reg [7:0] p62_array_index_1088624;
  reg [7:0] p62_array_index_1088625;
  reg [7:0] p62_res7__326;
  reg [7:0] p62_array_index_1088635;
  reg [7:0] p62_array_index_1088636;
  reg [7:0] p62_array_index_1088637;
  reg [7:0] p62_res7__327;
  reg [7:0] p62_array_index_1088648;
  reg [7:0] p62_array_index_1088649;
  reg [7:0] p62_res7__328;
  reg [7:0] p62_array_index_1088659;
  reg [7:0] p62_array_index_1088660;
  reg [7:0] p62_res7__329;
  reg [7:0] p62_array_index_1088666;
  reg [7:0] p62_array_index_1088667;
  reg [7:0] p62_array_index_1088668;
  reg [7:0] p62_array_index_1088669;
  reg [7:0] p62_array_index_1088670;
  reg [7:0] p62_array_index_1088671;
  reg [7:0] p62_array_index_1088672;
  reg [7:0] p62_array_index_1088673;
  reg [7:0] p62_array_index_1088674;
  reg [127:0] p62_res__37;
  reg [7:0] p63_arr[256];
  reg [7:0] p63_literal_1076345[256];
  reg [7:0] p63_literal_1076347[256];
  reg [7:0] p63_literal_1076349[256];
  reg [7:0] p63_literal_1076351[256];
  reg [7:0] p63_literal_1076353[256];
  reg [7:0] p63_literal_1076355[256];
  reg [7:0] p63_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p62_xor_1087905 <= p61_xor_1087905;
    p62_xor_1088377 <= p61_xor_1088377;
    p62_array_index_1088415 <= p61_array_index_1088415;
    p62_array_index_1088416 <= p61_array_index_1088416;
    p62_array_index_1088417 <= p61_array_index_1088417;
    p62_array_index_1088418 <= p61_array_index_1088418;
    p62_array_index_1088419 <= p61_array_index_1088419;
    p62_array_index_1088420 <= p61_array_index_1088420;
    p62_array_index_1088431 <= p61_array_index_1088431;
    p62_array_index_1088432 <= p61_array_index_1088432;
    p62_array_index_1088433 <= p61_array_index_1088433;
    p62_res7__320 <= p61_res7__320;
    p62_array_index_1088448 <= p61_array_index_1088448;
    p62_array_index_1088449 <= p61_array_index_1088449;
    p62_array_index_1088450 <= p61_array_index_1088450;
    p62_res7__321 <= p61_res7__321;
    p62_array_index_1088463 <= p61_array_index_1088463;
    p62_array_index_1088464 <= p61_array_index_1088464;
    p62_array_index_1088465 <= p61_array_index_1088465;
    p62_res7__322 <= p61_res7__322;
    p62_array_index_1088477 <= p61_array_index_1088477;
    p62_array_index_1088478 <= p61_array_index_1088478;
    p62_array_index_1088479 <= p61_array_index_1088479;
    p62_res7__323 <= p61_res7__323;
    p62_array_index_1088492 <= p61_array_index_1088492;
    p62_array_index_1088493 <= p61_array_index_1088493;
    p62_array_index_1088494 <= p61_array_index_1088494;
    p62_res7__324 <= p61_res7__324;
    p62_array_index_1088609 <= p62_array_index_1088609_comb;
    p62_array_index_1088610 <= p62_array_index_1088610_comb;
    p62_array_index_1088611 <= p62_array_index_1088611_comb;
    p62_res7__325 <= p62_res7__325_comb;
    p62_array_index_1088623 <= p62_array_index_1088623_comb;
    p62_array_index_1088624 <= p62_array_index_1088624_comb;
    p62_array_index_1088625 <= p62_array_index_1088625_comb;
    p62_res7__326 <= p62_res7__326_comb;
    p62_array_index_1088635 <= p62_array_index_1088635_comb;
    p62_array_index_1088636 <= p62_array_index_1088636_comb;
    p62_array_index_1088637 <= p62_array_index_1088637_comb;
    p62_res7__327 <= p62_res7__327_comb;
    p62_array_index_1088648 <= p62_array_index_1088648_comb;
    p62_array_index_1088649 <= p62_array_index_1088649_comb;
    p62_res7__328 <= p62_res7__328_comb;
    p62_array_index_1088659 <= p62_array_index_1088659_comb;
    p62_array_index_1088660 <= p62_array_index_1088660_comb;
    p62_res7__329 <= p62_res7__329_comb;
    p62_array_index_1088666 <= p62_array_index_1088666_comb;
    p62_array_index_1088667 <= p62_array_index_1088667_comb;
    p62_array_index_1088668 <= p62_array_index_1088668_comb;
    p62_array_index_1088669 <= p62_array_index_1088669_comb;
    p62_array_index_1088670 <= p62_array_index_1088670_comb;
    p62_array_index_1088671 <= p62_array_index_1088671_comb;
    p62_array_index_1088672 <= p62_array_index_1088672_comb;
    p62_array_index_1088673 <= p62_array_index_1088673_comb;
    p62_array_index_1088674 <= p62_array_index_1088674_comb;
    p62_res__37 <= p61_res__37;
    p63_arr <= p62_arr;
    p63_literal_1076345 <= p62_literal_1076345;
    p63_literal_1076347 <= p62_literal_1076347;
    p63_literal_1076349 <= p62_literal_1076349;
    p63_literal_1076351 <= p62_literal_1076351;
    p63_literal_1076353 <= p62_literal_1076353;
    p63_literal_1076355 <= p62_literal_1076355;
    p63_literal_1076358 <= p62_literal_1076358;
  end

  // ===== Pipe stage 63:
  wire [7:0] p63_res7__330_comb;
  wire [7:0] p63_array_index_1088809_comb;
  wire [7:0] p63_res7__331_comb;
  wire [7:0] p63_res7__332_comb;
  wire [7:0] p63_res7__333_comb;
  wire [7:0] p63_res7__334_comb;
  wire [7:0] p63_res7__335_comb;
  wire [127:0] p63_res__20_comb;
  wire [127:0] p63_xor_1088849_comb;
  assign p63_res7__330_comb = p62_array_index_1088666 ^ p62_array_index_1088667 ^ p62_array_index_1088668 ^ p62_array_index_1088669 ^ p62_array_index_1088670 ^ p62_array_index_1088671 ^ p62_res7__323 ^ p62_array_index_1088672 ^ p62_res7__321 ^ p62_array_index_1088625 ^ p62_array_index_1088494 ^ p62_array_index_1088465 ^ p62_array_index_1088433 ^ p62_array_index_1088673 ^ p62_array_index_1088674 ^ p62_array_index_1088420;
  assign p63_array_index_1088809_comb = p62_literal_1076355[p62_res7__325];
  assign p63_res7__331_comb = p62_literal_1076345[p63_res7__330_comb] ^ p62_literal_1076347[p62_res7__329] ^ p62_literal_1076349[p62_res7__328] ^ p62_literal_1076351[p62_res7__327] ^ p62_literal_1076353[p62_res7__326] ^ p63_array_index_1088809_comb ^ p62_res7__324 ^ p62_literal_1076358[p62_res7__323] ^ p62_res7__322 ^ p62_array_index_1088637 ^ p62_array_index_1088611 ^ p62_array_index_1088479 ^ p62_array_index_1088450 ^ p62_literal_1076347[p62_array_index_1088417] ^ p62_literal_1076345[p62_array_index_1088418] ^ p62_array_index_1088419;
  assign p63_res7__332_comb = p62_literal_1076345[p63_res7__331_comb] ^ p62_literal_1076347[p63_res7__330_comb] ^ p62_literal_1076349[p62_res7__329] ^ p62_literal_1076351[p62_res7__328] ^ p62_literal_1076353[p62_res7__327] ^ p62_literal_1076355[p62_res7__326] ^ p62_res7__325 ^ p62_literal_1076358[p62_res7__324] ^ p62_res7__323 ^ p62_array_index_1088649 ^ p62_array_index_1088624 ^ p62_array_index_1088493 ^ p62_array_index_1088464 ^ p62_array_index_1088432 ^ p62_literal_1076345[p62_array_index_1088417] ^ p62_array_index_1088418;
  assign p63_res7__333_comb = p62_literal_1076345[p63_res7__332_comb] ^ p62_literal_1076347[p63_res7__331_comb] ^ p62_literal_1076349[p63_res7__330_comb] ^ p62_literal_1076351[p62_res7__329] ^ p62_literal_1076353[p62_res7__328] ^ p62_literal_1076355[p62_res7__327] ^ p62_res7__326 ^ p62_literal_1076358[p62_res7__325] ^ p62_res7__324 ^ p62_array_index_1088660 ^ p62_array_index_1088636 ^ p62_array_index_1088610 ^ p62_array_index_1088478 ^ p62_array_index_1088449 ^ p62_literal_1076345[p62_array_index_1088416] ^ p62_array_index_1088417;
  assign p63_res7__334_comb = p62_literal_1076345[p63_res7__333_comb] ^ p62_literal_1076347[p63_res7__332_comb] ^ p62_literal_1076349[p63_res7__331_comb] ^ p62_literal_1076351[p63_res7__330_comb] ^ p62_literal_1076353[p62_res7__329] ^ p62_literal_1076355[p62_res7__328] ^ p62_res7__327 ^ p62_literal_1076358[p62_res7__326] ^ p62_res7__325 ^ p62_array_index_1088671 ^ p62_array_index_1088648 ^ p62_array_index_1088623 ^ p62_array_index_1088492 ^ p62_array_index_1088463 ^ p62_array_index_1088431 ^ p62_array_index_1088416;
  assign p63_res7__335_comb = p62_literal_1076345[p63_res7__334_comb] ^ p62_literal_1076347[p63_res7__333_comb] ^ p62_literal_1076349[p63_res7__332_comb] ^ p62_literal_1076351[p63_res7__331_comb] ^ p62_literal_1076353[p63_res7__330_comb] ^ p62_literal_1076355[p62_res7__329] ^ p62_res7__328 ^ p62_literal_1076358[p62_res7__327] ^ p62_res7__326 ^ p63_array_index_1088809_comb ^ p62_array_index_1088659 ^ p62_array_index_1088635 ^ p62_array_index_1088609 ^ p62_array_index_1088477 ^ p62_array_index_1088448 ^ p62_array_index_1088415;
  assign p63_res__20_comb = {p63_res7__335_comb, p63_res7__334_comb, p63_res7__333_comb, p63_res7__332_comb, p63_res7__331_comb, p63_res7__330_comb, p62_res7__329, p62_res7__328, p62_res7__327, p62_res7__326, p62_res7__325, p62_res7__324, p62_res7__323, p62_res7__322, p62_res7__321, p62_res7__320};
  assign p63_xor_1088849_comb = p63_res__20_comb ^ p62_xor_1087905;

  // Registers for pipe stage 63:
  reg [127:0] p63_xor_1088377;
  reg [127:0] p63_xor_1088849;
  reg [127:0] p63_res__37;
  reg [7:0] p64_arr[256];
  reg [7:0] p64_literal_1076345[256];
  reg [7:0] p64_literal_1076347[256];
  reg [7:0] p64_literal_1076349[256];
  reg [7:0] p64_literal_1076351[256];
  reg [7:0] p64_literal_1076353[256];
  reg [7:0] p64_literal_1076355[256];
  reg [7:0] p64_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p63_xor_1088377 <= p62_xor_1088377;
    p63_xor_1088849 <= p63_xor_1088849_comb;
    p63_res__37 <= p62_res__37;
    p64_arr <= p63_arr;
    p64_literal_1076345 <= p63_literal_1076345;
    p64_literal_1076347 <= p63_literal_1076347;
    p64_literal_1076349 <= p63_literal_1076349;
    p64_literal_1076351 <= p63_literal_1076351;
    p64_literal_1076353 <= p63_literal_1076353;
    p64_literal_1076355 <= p63_literal_1076355;
    p64_literal_1076358 <= p63_literal_1076358;
  end

  // ===== Pipe stage 64:
  wire [127:0] p64_addedKey__62_comb;
  wire [7:0] p64_array_index_1088887_comb;
  wire [7:0] p64_array_index_1088888_comb;
  wire [7:0] p64_array_index_1088889_comb;
  wire [7:0] p64_array_index_1088890_comb;
  wire [7:0] p64_array_index_1088891_comb;
  wire [7:0] p64_array_index_1088892_comb;
  wire [7:0] p64_array_index_1088894_comb;
  wire [7:0] p64_array_index_1088896_comb;
  wire [7:0] p64_array_index_1088897_comb;
  wire [7:0] p64_array_index_1088898_comb;
  wire [7:0] p64_array_index_1088899_comb;
  wire [7:0] p64_array_index_1088900_comb;
  wire [7:0] p64_array_index_1088901_comb;
  wire [7:0] p64_array_index_1088903_comb;
  wire [7:0] p64_array_index_1088904_comb;
  wire [7:0] p64_array_index_1088905_comb;
  wire [7:0] p64_array_index_1088906_comb;
  wire [7:0] p64_array_index_1088907_comb;
  wire [7:0] p64_array_index_1088908_comb;
  wire [7:0] p64_array_index_1088909_comb;
  wire [7:0] p64_array_index_1088911_comb;
  wire [7:0] p64_res7__336_comb;
  wire [7:0] p64_array_index_1088920_comb;
  wire [7:0] p64_array_index_1088921_comb;
  wire [7:0] p64_array_index_1088922_comb;
  wire [7:0] p64_array_index_1088923_comb;
  wire [7:0] p64_array_index_1088924_comb;
  wire [7:0] p64_array_index_1088925_comb;
  wire [7:0] p64_res7__337_comb;
  wire [7:0] p64_array_index_1088935_comb;
  wire [7:0] p64_array_index_1088936_comb;
  wire [7:0] p64_array_index_1088937_comb;
  wire [7:0] p64_array_index_1088938_comb;
  wire [7:0] p64_array_index_1088939_comb;
  wire [7:0] p64_res7__338_comb;
  wire [7:0] p64_array_index_1088949_comb;
  wire [7:0] p64_array_index_1088950_comb;
  wire [7:0] p64_array_index_1088951_comb;
  wire [7:0] p64_array_index_1088952_comb;
  wire [7:0] p64_array_index_1088953_comb;
  wire [7:0] p64_res7__339_comb;
  wire [7:0] p64_array_index_1088964_comb;
  wire [7:0] p64_array_index_1088965_comb;
  wire [7:0] p64_array_index_1088966_comb;
  wire [7:0] p64_array_index_1088967_comb;
  wire [7:0] p64_res7__340_comb;
  assign p64_addedKey__62_comb = p63_xor_1088849 ^ 128'h88f8_9bc3_a479_73c7_94e7_89a3_c509_aa16;
  assign p64_array_index_1088887_comb = p63_arr[p64_addedKey__62_comb[127:120]];
  assign p64_array_index_1088888_comb = p63_arr[p64_addedKey__62_comb[119:112]];
  assign p64_array_index_1088889_comb = p63_arr[p64_addedKey__62_comb[111:104]];
  assign p64_array_index_1088890_comb = p63_arr[p64_addedKey__62_comb[103:96]];
  assign p64_array_index_1088891_comb = p63_arr[p64_addedKey__62_comb[95:88]];
  assign p64_array_index_1088892_comb = p63_arr[p64_addedKey__62_comb[87:80]];
  assign p64_array_index_1088894_comb = p63_arr[p64_addedKey__62_comb[71:64]];
  assign p64_array_index_1088896_comb = p63_arr[p64_addedKey__62_comb[55:48]];
  assign p64_array_index_1088897_comb = p63_arr[p64_addedKey__62_comb[47:40]];
  assign p64_array_index_1088898_comb = p63_arr[p64_addedKey__62_comb[39:32]];
  assign p64_array_index_1088899_comb = p63_arr[p64_addedKey__62_comb[31:24]];
  assign p64_array_index_1088900_comb = p63_arr[p64_addedKey__62_comb[23:16]];
  assign p64_array_index_1088901_comb = p63_arr[p64_addedKey__62_comb[15:8]];
  assign p64_array_index_1088903_comb = p63_literal_1076345[p64_array_index_1088887_comb];
  assign p64_array_index_1088904_comb = p63_literal_1076347[p64_array_index_1088888_comb];
  assign p64_array_index_1088905_comb = p63_literal_1076349[p64_array_index_1088889_comb];
  assign p64_array_index_1088906_comb = p63_literal_1076351[p64_array_index_1088890_comb];
  assign p64_array_index_1088907_comb = p63_literal_1076353[p64_array_index_1088891_comb];
  assign p64_array_index_1088908_comb = p63_literal_1076355[p64_array_index_1088892_comb];
  assign p64_array_index_1088909_comb = p63_arr[p64_addedKey__62_comb[79:72]];
  assign p64_array_index_1088911_comb = p63_arr[p64_addedKey__62_comb[63:56]];
  assign p64_res7__336_comb = p64_array_index_1088903_comb ^ p64_array_index_1088904_comb ^ p64_array_index_1088905_comb ^ p64_array_index_1088906_comb ^ p64_array_index_1088907_comb ^ p64_array_index_1088908_comb ^ p64_array_index_1088909_comb ^ p63_literal_1076358[p64_array_index_1088894_comb] ^ p64_array_index_1088911_comb ^ p63_literal_1076355[p64_array_index_1088896_comb] ^ p63_literal_1076353[p64_array_index_1088897_comb] ^ p63_literal_1076351[p64_array_index_1088898_comb] ^ p63_literal_1076349[p64_array_index_1088899_comb] ^ p63_literal_1076347[p64_array_index_1088900_comb] ^ p63_literal_1076345[p64_array_index_1088901_comb] ^ p63_arr[p64_addedKey__62_comb[7:0]];
  assign p64_array_index_1088920_comb = p63_literal_1076345[p64_res7__336_comb];
  assign p64_array_index_1088921_comb = p63_literal_1076347[p64_array_index_1088887_comb];
  assign p64_array_index_1088922_comb = p63_literal_1076349[p64_array_index_1088888_comb];
  assign p64_array_index_1088923_comb = p63_literal_1076351[p64_array_index_1088889_comb];
  assign p64_array_index_1088924_comb = p63_literal_1076353[p64_array_index_1088890_comb];
  assign p64_array_index_1088925_comb = p63_literal_1076355[p64_array_index_1088891_comb];
  assign p64_res7__337_comb = p64_array_index_1088920_comb ^ p64_array_index_1088921_comb ^ p64_array_index_1088922_comb ^ p64_array_index_1088923_comb ^ p64_array_index_1088924_comb ^ p64_array_index_1088925_comb ^ p64_array_index_1088892_comb ^ p63_literal_1076358[p64_array_index_1088909_comb] ^ p64_array_index_1088894_comb ^ p63_literal_1076355[p64_array_index_1088911_comb] ^ p63_literal_1076353[p64_array_index_1088896_comb] ^ p63_literal_1076351[p64_array_index_1088897_comb] ^ p63_literal_1076349[p64_array_index_1088898_comb] ^ p63_literal_1076347[p64_array_index_1088899_comb] ^ p63_literal_1076345[p64_array_index_1088900_comb] ^ p64_array_index_1088901_comb;
  assign p64_array_index_1088935_comb = p63_literal_1076347[p64_res7__336_comb];
  assign p64_array_index_1088936_comb = p63_literal_1076349[p64_array_index_1088887_comb];
  assign p64_array_index_1088937_comb = p63_literal_1076351[p64_array_index_1088888_comb];
  assign p64_array_index_1088938_comb = p63_literal_1076353[p64_array_index_1088889_comb];
  assign p64_array_index_1088939_comb = p63_literal_1076355[p64_array_index_1088890_comb];
  assign p64_res7__338_comb = p63_literal_1076345[p64_res7__337_comb] ^ p64_array_index_1088935_comb ^ p64_array_index_1088936_comb ^ p64_array_index_1088937_comb ^ p64_array_index_1088938_comb ^ p64_array_index_1088939_comb ^ p64_array_index_1088891_comb ^ p63_literal_1076358[p64_array_index_1088892_comb] ^ p64_array_index_1088909_comb ^ p63_literal_1076355[p64_array_index_1088894_comb] ^ p63_literal_1076353[p64_array_index_1088911_comb] ^ p63_literal_1076351[p64_array_index_1088896_comb] ^ p63_literal_1076349[p64_array_index_1088897_comb] ^ p63_literal_1076347[p64_array_index_1088898_comb] ^ p63_literal_1076345[p64_array_index_1088899_comb] ^ p64_array_index_1088900_comb;
  assign p64_array_index_1088949_comb = p63_literal_1076347[p64_res7__337_comb];
  assign p64_array_index_1088950_comb = p63_literal_1076349[p64_res7__336_comb];
  assign p64_array_index_1088951_comb = p63_literal_1076351[p64_array_index_1088887_comb];
  assign p64_array_index_1088952_comb = p63_literal_1076353[p64_array_index_1088888_comb];
  assign p64_array_index_1088953_comb = p63_literal_1076355[p64_array_index_1088889_comb];
  assign p64_res7__339_comb = p63_literal_1076345[p64_res7__338_comb] ^ p64_array_index_1088949_comb ^ p64_array_index_1088950_comb ^ p64_array_index_1088951_comb ^ p64_array_index_1088952_comb ^ p64_array_index_1088953_comb ^ p64_array_index_1088890_comb ^ p63_literal_1076358[p64_array_index_1088891_comb] ^ p64_array_index_1088892_comb ^ p63_literal_1076355[p64_array_index_1088909_comb] ^ p63_literal_1076353[p64_array_index_1088894_comb] ^ p63_literal_1076351[p64_array_index_1088911_comb] ^ p63_literal_1076349[p64_array_index_1088896_comb] ^ p63_literal_1076347[p64_array_index_1088897_comb] ^ p63_literal_1076345[p64_array_index_1088898_comb] ^ p64_array_index_1088899_comb;
  assign p64_array_index_1088964_comb = p63_literal_1076349[p64_res7__337_comb];
  assign p64_array_index_1088965_comb = p63_literal_1076351[p64_res7__336_comb];
  assign p64_array_index_1088966_comb = p63_literal_1076353[p64_array_index_1088887_comb];
  assign p64_array_index_1088967_comb = p63_literal_1076355[p64_array_index_1088888_comb];
  assign p64_res7__340_comb = p63_literal_1076345[p64_res7__339_comb] ^ p63_literal_1076347[p64_res7__338_comb] ^ p64_array_index_1088964_comb ^ p64_array_index_1088965_comb ^ p64_array_index_1088966_comb ^ p64_array_index_1088967_comb ^ p64_array_index_1088889_comb ^ p63_literal_1076358[p64_array_index_1088890_comb] ^ p64_array_index_1088891_comb ^ p64_array_index_1088908_comb ^ p63_literal_1076353[p64_array_index_1088909_comb] ^ p63_literal_1076351[p64_array_index_1088894_comb] ^ p63_literal_1076349[p64_array_index_1088911_comb] ^ p63_literal_1076347[p64_array_index_1088896_comb] ^ p63_literal_1076345[p64_array_index_1088897_comb] ^ p64_array_index_1088898_comb;

  // Registers for pipe stage 64:
  reg [127:0] p64_xor_1088377;
  reg [127:0] p64_xor_1088849;
  reg [7:0] p64_array_index_1088887;
  reg [7:0] p64_array_index_1088888;
  reg [7:0] p64_array_index_1088889;
  reg [7:0] p64_array_index_1088890;
  reg [7:0] p64_array_index_1088891;
  reg [7:0] p64_array_index_1088892;
  reg [7:0] p64_array_index_1088894;
  reg [7:0] p64_array_index_1088896;
  reg [7:0] p64_array_index_1088897;
  reg [7:0] p64_array_index_1088903;
  reg [7:0] p64_array_index_1088904;
  reg [7:0] p64_array_index_1088905;
  reg [7:0] p64_array_index_1088906;
  reg [7:0] p64_array_index_1088907;
  reg [7:0] p64_array_index_1088909;
  reg [7:0] p64_array_index_1088911;
  reg [7:0] p64_res7__336;
  reg [7:0] p64_array_index_1088920;
  reg [7:0] p64_array_index_1088921;
  reg [7:0] p64_array_index_1088922;
  reg [7:0] p64_array_index_1088923;
  reg [7:0] p64_array_index_1088924;
  reg [7:0] p64_array_index_1088925;
  reg [7:0] p64_res7__337;
  reg [7:0] p64_array_index_1088935;
  reg [7:0] p64_array_index_1088936;
  reg [7:0] p64_array_index_1088937;
  reg [7:0] p64_array_index_1088938;
  reg [7:0] p64_array_index_1088939;
  reg [7:0] p64_res7__338;
  reg [7:0] p64_array_index_1088949;
  reg [7:0] p64_array_index_1088950;
  reg [7:0] p64_array_index_1088951;
  reg [7:0] p64_array_index_1088952;
  reg [7:0] p64_array_index_1088953;
  reg [7:0] p64_res7__339;
  reg [7:0] p64_array_index_1088964;
  reg [7:0] p64_array_index_1088965;
  reg [7:0] p64_array_index_1088966;
  reg [7:0] p64_array_index_1088967;
  reg [7:0] p64_res7__340;
  reg [127:0] p64_res__37;
  reg [7:0] p65_arr[256];
  reg [7:0] p65_literal_1076345[256];
  reg [7:0] p65_literal_1076347[256];
  reg [7:0] p65_literal_1076349[256];
  reg [7:0] p65_literal_1076351[256];
  reg [7:0] p65_literal_1076353[256];
  reg [7:0] p65_literal_1076355[256];
  reg [7:0] p65_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p64_xor_1088377 <= p63_xor_1088377;
    p64_xor_1088849 <= p63_xor_1088849;
    p64_array_index_1088887 <= p64_array_index_1088887_comb;
    p64_array_index_1088888 <= p64_array_index_1088888_comb;
    p64_array_index_1088889 <= p64_array_index_1088889_comb;
    p64_array_index_1088890 <= p64_array_index_1088890_comb;
    p64_array_index_1088891 <= p64_array_index_1088891_comb;
    p64_array_index_1088892 <= p64_array_index_1088892_comb;
    p64_array_index_1088894 <= p64_array_index_1088894_comb;
    p64_array_index_1088896 <= p64_array_index_1088896_comb;
    p64_array_index_1088897 <= p64_array_index_1088897_comb;
    p64_array_index_1088903 <= p64_array_index_1088903_comb;
    p64_array_index_1088904 <= p64_array_index_1088904_comb;
    p64_array_index_1088905 <= p64_array_index_1088905_comb;
    p64_array_index_1088906 <= p64_array_index_1088906_comb;
    p64_array_index_1088907 <= p64_array_index_1088907_comb;
    p64_array_index_1088909 <= p64_array_index_1088909_comb;
    p64_array_index_1088911 <= p64_array_index_1088911_comb;
    p64_res7__336 <= p64_res7__336_comb;
    p64_array_index_1088920 <= p64_array_index_1088920_comb;
    p64_array_index_1088921 <= p64_array_index_1088921_comb;
    p64_array_index_1088922 <= p64_array_index_1088922_comb;
    p64_array_index_1088923 <= p64_array_index_1088923_comb;
    p64_array_index_1088924 <= p64_array_index_1088924_comb;
    p64_array_index_1088925 <= p64_array_index_1088925_comb;
    p64_res7__337 <= p64_res7__337_comb;
    p64_array_index_1088935 <= p64_array_index_1088935_comb;
    p64_array_index_1088936 <= p64_array_index_1088936_comb;
    p64_array_index_1088937 <= p64_array_index_1088937_comb;
    p64_array_index_1088938 <= p64_array_index_1088938_comb;
    p64_array_index_1088939 <= p64_array_index_1088939_comb;
    p64_res7__338 <= p64_res7__338_comb;
    p64_array_index_1088949 <= p64_array_index_1088949_comb;
    p64_array_index_1088950 <= p64_array_index_1088950_comb;
    p64_array_index_1088951 <= p64_array_index_1088951_comb;
    p64_array_index_1088952 <= p64_array_index_1088952_comb;
    p64_array_index_1088953 <= p64_array_index_1088953_comb;
    p64_res7__339 <= p64_res7__339_comb;
    p64_array_index_1088964 <= p64_array_index_1088964_comb;
    p64_array_index_1088965 <= p64_array_index_1088965_comb;
    p64_array_index_1088966 <= p64_array_index_1088966_comb;
    p64_array_index_1088967 <= p64_array_index_1088967_comb;
    p64_res7__340 <= p64_res7__340_comb;
    p64_res__37 <= p63_res__37;
    p65_arr <= p64_arr;
    p65_literal_1076345 <= p64_literal_1076345;
    p65_literal_1076347 <= p64_literal_1076347;
    p65_literal_1076349 <= p64_literal_1076349;
    p65_literal_1076351 <= p64_literal_1076351;
    p65_literal_1076353 <= p64_literal_1076353;
    p65_literal_1076355 <= p64_literal_1076355;
    p65_literal_1076358 <= p64_literal_1076358;
  end

  // ===== Pipe stage 65:
  wire [7:0] p65_array_index_1089081_comb;
  wire [7:0] p65_array_index_1089082_comb;
  wire [7:0] p65_array_index_1089083_comb;
  wire [7:0] p65_array_index_1089084_comb;
  wire [7:0] p65_res7__341_comb;
  wire [7:0] p65_array_index_1089095_comb;
  wire [7:0] p65_array_index_1089096_comb;
  wire [7:0] p65_array_index_1089097_comb;
  wire [7:0] p65_res7__342_comb;
  wire [7:0] p65_array_index_1089107_comb;
  wire [7:0] p65_array_index_1089108_comb;
  wire [7:0] p65_array_index_1089109_comb;
  wire [7:0] p65_res7__343_comb;
  wire [7:0] p65_array_index_1089120_comb;
  wire [7:0] p65_array_index_1089121_comb;
  wire [7:0] p65_res7__344_comb;
  wire [7:0] p65_array_index_1089131_comb;
  wire [7:0] p65_array_index_1089132_comb;
  wire [7:0] p65_res7__345_comb;
  wire [7:0] p65_array_index_1089138_comb;
  wire [7:0] p65_array_index_1089139_comb;
  wire [7:0] p65_array_index_1089140_comb;
  wire [7:0] p65_array_index_1089141_comb;
  wire [7:0] p65_array_index_1089142_comb;
  wire [7:0] p65_array_index_1089143_comb;
  wire [7:0] p65_array_index_1089144_comb;
  wire [7:0] p65_array_index_1089145_comb;
  wire [7:0] p65_array_index_1089146_comb;
  assign p65_array_index_1089081_comb = p64_literal_1076349[p64_res7__338];
  assign p65_array_index_1089082_comb = p64_literal_1076351[p64_res7__337];
  assign p65_array_index_1089083_comb = p64_literal_1076353[p64_res7__336];
  assign p65_array_index_1089084_comb = p64_literal_1076355[p64_array_index_1088887];
  assign p65_res7__341_comb = p64_literal_1076345[p64_res7__340] ^ p64_literal_1076347[p64_res7__339] ^ p65_array_index_1089081_comb ^ p65_array_index_1089082_comb ^ p65_array_index_1089083_comb ^ p65_array_index_1089084_comb ^ p64_array_index_1088888 ^ p64_literal_1076358[p64_array_index_1088889] ^ p64_array_index_1088890 ^ p64_array_index_1088925 ^ p64_literal_1076353[p64_array_index_1088892] ^ p64_literal_1076351[p64_array_index_1088909] ^ p64_literal_1076349[p64_array_index_1088894] ^ p64_literal_1076347[p64_array_index_1088911] ^ p64_literal_1076345[p64_array_index_1088896] ^ p64_array_index_1088897;
  assign p65_array_index_1089095_comb = p64_literal_1076351[p64_res7__338];
  assign p65_array_index_1089096_comb = p64_literal_1076353[p64_res7__337];
  assign p65_array_index_1089097_comb = p64_literal_1076355[p64_res7__336];
  assign p65_res7__342_comb = p64_literal_1076345[p65_res7__341_comb] ^ p64_literal_1076347[p64_res7__340] ^ p64_literal_1076349[p64_res7__339] ^ p65_array_index_1089095_comb ^ p65_array_index_1089096_comb ^ p65_array_index_1089097_comb ^ p64_array_index_1088887 ^ p64_literal_1076358[p64_array_index_1088888] ^ p64_array_index_1088889 ^ p64_array_index_1088939 ^ p64_array_index_1088907 ^ p64_literal_1076351[p64_array_index_1088892] ^ p64_literal_1076349[p64_array_index_1088909] ^ p64_literal_1076347[p64_array_index_1088894] ^ p64_literal_1076345[p64_array_index_1088911] ^ p64_array_index_1088896;
  assign p65_array_index_1089107_comb = p64_literal_1076351[p64_res7__339];
  assign p65_array_index_1089108_comb = p64_literal_1076353[p64_res7__338];
  assign p65_array_index_1089109_comb = p64_literal_1076355[p64_res7__337];
  assign p65_res7__343_comb = p64_literal_1076345[p65_res7__342_comb] ^ p64_literal_1076347[p65_res7__341_comb] ^ p64_literal_1076349[p64_res7__340] ^ p65_array_index_1089107_comb ^ p65_array_index_1089108_comb ^ p65_array_index_1089109_comb ^ p64_res7__336 ^ p64_literal_1076358[p64_array_index_1088887] ^ p64_array_index_1088888 ^ p64_array_index_1088953 ^ p64_array_index_1088924 ^ p64_literal_1076351[p64_array_index_1088891] ^ p64_literal_1076349[p64_array_index_1088892] ^ p64_literal_1076347[p64_array_index_1088909] ^ p64_literal_1076345[p64_array_index_1088894] ^ p64_array_index_1088911;
  assign p65_array_index_1089120_comb = p64_literal_1076353[p64_res7__339];
  assign p65_array_index_1089121_comb = p64_literal_1076355[p64_res7__338];
  assign p65_res7__344_comb = p64_literal_1076345[p65_res7__343_comb] ^ p64_literal_1076347[p65_res7__342_comb] ^ p64_literal_1076349[p65_res7__341_comb] ^ p64_literal_1076351[p64_res7__340] ^ p65_array_index_1089120_comb ^ p65_array_index_1089121_comb ^ p64_res7__337 ^ p64_literal_1076358[p64_res7__336] ^ p64_array_index_1088887 ^ p64_array_index_1088967 ^ p64_array_index_1088938 ^ p64_array_index_1088906 ^ p64_literal_1076349[p64_array_index_1088891] ^ p64_literal_1076347[p64_array_index_1088892] ^ p64_literal_1076345[p64_array_index_1088909] ^ p64_array_index_1088894;
  assign p65_array_index_1089131_comb = p64_literal_1076353[p64_res7__340];
  assign p65_array_index_1089132_comb = p64_literal_1076355[p64_res7__339];
  assign p65_res7__345_comb = p64_literal_1076345[p65_res7__344_comb] ^ p64_literal_1076347[p65_res7__343_comb] ^ p64_literal_1076349[p65_res7__342_comb] ^ p64_literal_1076351[p65_res7__341_comb] ^ p65_array_index_1089131_comb ^ p65_array_index_1089132_comb ^ p64_res7__338 ^ p64_literal_1076358[p64_res7__337] ^ p64_res7__336 ^ p65_array_index_1089084_comb ^ p64_array_index_1088952 ^ p64_array_index_1088923 ^ p64_literal_1076349[p64_array_index_1088890] ^ p64_literal_1076347[p64_array_index_1088891] ^ p64_literal_1076345[p64_array_index_1088892] ^ p64_array_index_1088909;
  assign p65_array_index_1089138_comb = p64_literal_1076345[p65_res7__345_comb];
  assign p65_array_index_1089139_comb = p64_literal_1076347[p65_res7__344_comb];
  assign p65_array_index_1089140_comb = p64_literal_1076349[p65_res7__343_comb];
  assign p65_array_index_1089141_comb = p64_literal_1076351[p65_res7__342_comb];
  assign p65_array_index_1089142_comb = p64_literal_1076353[p65_res7__341_comb];
  assign p65_array_index_1089143_comb = p64_literal_1076355[p64_res7__340];
  assign p65_array_index_1089144_comb = p64_literal_1076358[p64_res7__338];
  assign p65_array_index_1089145_comb = p64_literal_1076347[p64_array_index_1088890];
  assign p65_array_index_1089146_comb = p64_literal_1076345[p64_array_index_1088891];

  // Registers for pipe stage 65:
  reg [127:0] p65_xor_1088377;
  reg [127:0] p65_xor_1088849;
  reg [7:0] p65_array_index_1088887;
  reg [7:0] p65_array_index_1088888;
  reg [7:0] p65_array_index_1088889;
  reg [7:0] p65_array_index_1088890;
  reg [7:0] p65_array_index_1088891;
  reg [7:0] p65_array_index_1088892;
  reg [7:0] p65_array_index_1088903;
  reg [7:0] p65_array_index_1088904;
  reg [7:0] p65_array_index_1088905;
  reg [7:0] p65_res7__336;
  reg [7:0] p65_array_index_1088920;
  reg [7:0] p65_array_index_1088921;
  reg [7:0] p65_array_index_1088922;
  reg [7:0] p65_res7__337;
  reg [7:0] p65_array_index_1088935;
  reg [7:0] p65_array_index_1088936;
  reg [7:0] p65_array_index_1088937;
  reg [7:0] p65_res7__338;
  reg [7:0] p65_array_index_1088949;
  reg [7:0] p65_array_index_1088950;
  reg [7:0] p65_array_index_1088951;
  reg [7:0] p65_res7__339;
  reg [7:0] p65_array_index_1088964;
  reg [7:0] p65_array_index_1088965;
  reg [7:0] p65_array_index_1088966;
  reg [7:0] p65_res7__340;
  reg [7:0] p65_array_index_1089081;
  reg [7:0] p65_array_index_1089082;
  reg [7:0] p65_array_index_1089083;
  reg [7:0] p65_res7__341;
  reg [7:0] p65_array_index_1089095;
  reg [7:0] p65_array_index_1089096;
  reg [7:0] p65_array_index_1089097;
  reg [7:0] p65_res7__342;
  reg [7:0] p65_array_index_1089107;
  reg [7:0] p65_array_index_1089108;
  reg [7:0] p65_array_index_1089109;
  reg [7:0] p65_res7__343;
  reg [7:0] p65_array_index_1089120;
  reg [7:0] p65_array_index_1089121;
  reg [7:0] p65_res7__344;
  reg [7:0] p65_array_index_1089131;
  reg [7:0] p65_array_index_1089132;
  reg [7:0] p65_res7__345;
  reg [7:0] p65_array_index_1089138;
  reg [7:0] p65_array_index_1089139;
  reg [7:0] p65_array_index_1089140;
  reg [7:0] p65_array_index_1089141;
  reg [7:0] p65_array_index_1089142;
  reg [7:0] p65_array_index_1089143;
  reg [7:0] p65_array_index_1089144;
  reg [7:0] p65_array_index_1089145;
  reg [7:0] p65_array_index_1089146;
  reg [127:0] p65_res__37;
  reg [7:0] p66_arr[256];
  reg [7:0] p66_literal_1076345[256];
  reg [7:0] p66_literal_1076347[256];
  reg [7:0] p66_literal_1076349[256];
  reg [7:0] p66_literal_1076351[256];
  reg [7:0] p66_literal_1076353[256];
  reg [7:0] p66_literal_1076355[256];
  reg [7:0] p66_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p65_xor_1088377 <= p64_xor_1088377;
    p65_xor_1088849 <= p64_xor_1088849;
    p65_array_index_1088887 <= p64_array_index_1088887;
    p65_array_index_1088888 <= p64_array_index_1088888;
    p65_array_index_1088889 <= p64_array_index_1088889;
    p65_array_index_1088890 <= p64_array_index_1088890;
    p65_array_index_1088891 <= p64_array_index_1088891;
    p65_array_index_1088892 <= p64_array_index_1088892;
    p65_array_index_1088903 <= p64_array_index_1088903;
    p65_array_index_1088904 <= p64_array_index_1088904;
    p65_array_index_1088905 <= p64_array_index_1088905;
    p65_res7__336 <= p64_res7__336;
    p65_array_index_1088920 <= p64_array_index_1088920;
    p65_array_index_1088921 <= p64_array_index_1088921;
    p65_array_index_1088922 <= p64_array_index_1088922;
    p65_res7__337 <= p64_res7__337;
    p65_array_index_1088935 <= p64_array_index_1088935;
    p65_array_index_1088936 <= p64_array_index_1088936;
    p65_array_index_1088937 <= p64_array_index_1088937;
    p65_res7__338 <= p64_res7__338;
    p65_array_index_1088949 <= p64_array_index_1088949;
    p65_array_index_1088950 <= p64_array_index_1088950;
    p65_array_index_1088951 <= p64_array_index_1088951;
    p65_res7__339 <= p64_res7__339;
    p65_array_index_1088964 <= p64_array_index_1088964;
    p65_array_index_1088965 <= p64_array_index_1088965;
    p65_array_index_1088966 <= p64_array_index_1088966;
    p65_res7__340 <= p64_res7__340;
    p65_array_index_1089081 <= p65_array_index_1089081_comb;
    p65_array_index_1089082 <= p65_array_index_1089082_comb;
    p65_array_index_1089083 <= p65_array_index_1089083_comb;
    p65_res7__341 <= p65_res7__341_comb;
    p65_array_index_1089095 <= p65_array_index_1089095_comb;
    p65_array_index_1089096 <= p65_array_index_1089096_comb;
    p65_array_index_1089097 <= p65_array_index_1089097_comb;
    p65_res7__342 <= p65_res7__342_comb;
    p65_array_index_1089107 <= p65_array_index_1089107_comb;
    p65_array_index_1089108 <= p65_array_index_1089108_comb;
    p65_array_index_1089109 <= p65_array_index_1089109_comb;
    p65_res7__343 <= p65_res7__343_comb;
    p65_array_index_1089120 <= p65_array_index_1089120_comb;
    p65_array_index_1089121 <= p65_array_index_1089121_comb;
    p65_res7__344 <= p65_res7__344_comb;
    p65_array_index_1089131 <= p65_array_index_1089131_comb;
    p65_array_index_1089132 <= p65_array_index_1089132_comb;
    p65_res7__345 <= p65_res7__345_comb;
    p65_array_index_1089138 <= p65_array_index_1089138_comb;
    p65_array_index_1089139 <= p65_array_index_1089139_comb;
    p65_array_index_1089140 <= p65_array_index_1089140_comb;
    p65_array_index_1089141 <= p65_array_index_1089141_comb;
    p65_array_index_1089142 <= p65_array_index_1089142_comb;
    p65_array_index_1089143 <= p65_array_index_1089143_comb;
    p65_array_index_1089144 <= p65_array_index_1089144_comb;
    p65_array_index_1089145 <= p65_array_index_1089145_comb;
    p65_array_index_1089146 <= p65_array_index_1089146_comb;
    p65_res__37 <= p64_res__37;
    p66_arr <= p65_arr;
    p66_literal_1076345 <= p65_literal_1076345;
    p66_literal_1076347 <= p65_literal_1076347;
    p66_literal_1076349 <= p65_literal_1076349;
    p66_literal_1076351 <= p65_literal_1076351;
    p66_literal_1076353 <= p65_literal_1076353;
    p66_literal_1076355 <= p65_literal_1076355;
    p66_literal_1076358 <= p65_literal_1076358;
  end

  // ===== Pipe stage 66:
  wire [7:0] p66_res7__346_comb;
  wire [7:0] p66_array_index_1089281_comb;
  wire [7:0] p66_res7__347_comb;
  wire [7:0] p66_res7__348_comb;
  wire [7:0] p66_res7__349_comb;
  wire [7:0] p66_res7__350_comb;
  wire [7:0] p66_res7__351_comb;
  wire [127:0] p66_res__21_comb;
  wire [127:0] p66_xor_1089321_comb;
  assign p66_res7__346_comb = p65_array_index_1089138 ^ p65_array_index_1089139 ^ p65_array_index_1089140 ^ p65_array_index_1089141 ^ p65_array_index_1089142 ^ p65_array_index_1089143 ^ p65_res7__339 ^ p65_array_index_1089144 ^ p65_res7__337 ^ p65_array_index_1089097 ^ p65_array_index_1088966 ^ p65_array_index_1088937 ^ p65_array_index_1088905 ^ p65_array_index_1089145 ^ p65_array_index_1089146 ^ p65_array_index_1088892;
  assign p66_array_index_1089281_comb = p65_literal_1076355[p65_res7__341];
  assign p66_res7__347_comb = p65_literal_1076345[p66_res7__346_comb] ^ p65_literal_1076347[p65_res7__345] ^ p65_literal_1076349[p65_res7__344] ^ p65_literal_1076351[p65_res7__343] ^ p65_literal_1076353[p65_res7__342] ^ p66_array_index_1089281_comb ^ p65_res7__340 ^ p65_literal_1076358[p65_res7__339] ^ p65_res7__338 ^ p65_array_index_1089109 ^ p65_array_index_1089083 ^ p65_array_index_1088951 ^ p65_array_index_1088922 ^ p65_literal_1076347[p65_array_index_1088889] ^ p65_literal_1076345[p65_array_index_1088890] ^ p65_array_index_1088891;
  assign p66_res7__348_comb = p65_literal_1076345[p66_res7__347_comb] ^ p65_literal_1076347[p66_res7__346_comb] ^ p65_literal_1076349[p65_res7__345] ^ p65_literal_1076351[p65_res7__344] ^ p65_literal_1076353[p65_res7__343] ^ p65_literal_1076355[p65_res7__342] ^ p65_res7__341 ^ p65_literal_1076358[p65_res7__340] ^ p65_res7__339 ^ p65_array_index_1089121 ^ p65_array_index_1089096 ^ p65_array_index_1088965 ^ p65_array_index_1088936 ^ p65_array_index_1088904 ^ p65_literal_1076345[p65_array_index_1088889] ^ p65_array_index_1088890;
  assign p66_res7__349_comb = p65_literal_1076345[p66_res7__348_comb] ^ p65_literal_1076347[p66_res7__347_comb] ^ p65_literal_1076349[p66_res7__346_comb] ^ p65_literal_1076351[p65_res7__345] ^ p65_literal_1076353[p65_res7__344] ^ p65_literal_1076355[p65_res7__343] ^ p65_res7__342 ^ p65_literal_1076358[p65_res7__341] ^ p65_res7__340 ^ p65_array_index_1089132 ^ p65_array_index_1089108 ^ p65_array_index_1089082 ^ p65_array_index_1088950 ^ p65_array_index_1088921 ^ p65_literal_1076345[p65_array_index_1088888] ^ p65_array_index_1088889;
  assign p66_res7__350_comb = p65_literal_1076345[p66_res7__349_comb] ^ p65_literal_1076347[p66_res7__348_comb] ^ p65_literal_1076349[p66_res7__347_comb] ^ p65_literal_1076351[p66_res7__346_comb] ^ p65_literal_1076353[p65_res7__345] ^ p65_literal_1076355[p65_res7__344] ^ p65_res7__343 ^ p65_literal_1076358[p65_res7__342] ^ p65_res7__341 ^ p65_array_index_1089143 ^ p65_array_index_1089120 ^ p65_array_index_1089095 ^ p65_array_index_1088964 ^ p65_array_index_1088935 ^ p65_array_index_1088903 ^ p65_array_index_1088888;
  assign p66_res7__351_comb = p65_literal_1076345[p66_res7__350_comb] ^ p65_literal_1076347[p66_res7__349_comb] ^ p65_literal_1076349[p66_res7__348_comb] ^ p65_literal_1076351[p66_res7__347_comb] ^ p65_literal_1076353[p66_res7__346_comb] ^ p65_literal_1076355[p65_res7__345] ^ p65_res7__344 ^ p65_literal_1076358[p65_res7__343] ^ p65_res7__342 ^ p66_array_index_1089281_comb ^ p65_array_index_1089131 ^ p65_array_index_1089107 ^ p65_array_index_1089081 ^ p65_array_index_1088949 ^ p65_array_index_1088920 ^ p65_array_index_1088887;
  assign p66_res__21_comb = {p66_res7__351_comb, p66_res7__350_comb, p66_res7__349_comb, p66_res7__348_comb, p66_res7__347_comb, p66_res7__346_comb, p65_res7__345, p65_res7__344, p65_res7__343, p65_res7__342, p65_res7__341, p65_res7__340, p65_res7__339, p65_res7__338, p65_res7__337, p65_res7__336};
  assign p66_xor_1089321_comb = p66_res__21_comb ^ p65_xor_1088377;

  // Registers for pipe stage 66:
  reg [127:0] p66_xor_1088849;
  reg [127:0] p66_xor_1089321;
  reg [127:0] p66_res__37;
  reg [7:0] p67_arr[256];
  reg [7:0] p67_literal_1076345[256];
  reg [7:0] p67_literal_1076347[256];
  reg [7:0] p67_literal_1076349[256];
  reg [7:0] p67_literal_1076351[256];
  reg [7:0] p67_literal_1076353[256];
  reg [7:0] p67_literal_1076355[256];
  reg [7:0] p67_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p66_xor_1088849 <= p65_xor_1088849;
    p66_xor_1089321 <= p66_xor_1089321_comb;
    p66_res__37 <= p65_res__37;
    p67_arr <= p66_arr;
    p67_literal_1076345 <= p66_literal_1076345;
    p67_literal_1076347 <= p66_literal_1076347;
    p67_literal_1076349 <= p66_literal_1076349;
    p67_literal_1076351 <= p66_literal_1076351;
    p67_literal_1076353 <= p66_literal_1076353;
    p67_literal_1076355 <= p66_literal_1076355;
    p67_literal_1076358 <= p66_literal_1076358;
  end

  // ===== Pipe stage 67:
  wire [127:0] p67_addedKey__63_comb;
  wire [7:0] p67_array_index_1089359_comb;
  wire [7:0] p67_array_index_1089360_comb;
  wire [7:0] p67_array_index_1089361_comb;
  wire [7:0] p67_array_index_1089362_comb;
  wire [7:0] p67_array_index_1089363_comb;
  wire [7:0] p67_array_index_1089364_comb;
  wire [7:0] p67_array_index_1089366_comb;
  wire [7:0] p67_array_index_1089368_comb;
  wire [7:0] p67_array_index_1089369_comb;
  wire [7:0] p67_array_index_1089370_comb;
  wire [7:0] p67_array_index_1089371_comb;
  wire [7:0] p67_array_index_1089372_comb;
  wire [7:0] p67_array_index_1089373_comb;
  wire [7:0] p67_array_index_1089375_comb;
  wire [7:0] p67_array_index_1089376_comb;
  wire [7:0] p67_array_index_1089377_comb;
  wire [7:0] p67_array_index_1089378_comb;
  wire [7:0] p67_array_index_1089379_comb;
  wire [7:0] p67_array_index_1089380_comb;
  wire [7:0] p67_array_index_1089381_comb;
  wire [7:0] p67_array_index_1089383_comb;
  wire [7:0] p67_res7__352_comb;
  wire [7:0] p67_array_index_1089392_comb;
  wire [7:0] p67_array_index_1089393_comb;
  wire [7:0] p67_array_index_1089394_comb;
  wire [7:0] p67_array_index_1089395_comb;
  wire [7:0] p67_array_index_1089396_comb;
  wire [7:0] p67_array_index_1089397_comb;
  wire [7:0] p67_res7__353_comb;
  wire [7:0] p67_array_index_1089407_comb;
  wire [7:0] p67_array_index_1089408_comb;
  wire [7:0] p67_array_index_1089409_comb;
  wire [7:0] p67_array_index_1089410_comb;
  wire [7:0] p67_array_index_1089411_comb;
  wire [7:0] p67_res7__354_comb;
  wire [7:0] p67_array_index_1089421_comb;
  wire [7:0] p67_array_index_1089422_comb;
  wire [7:0] p67_array_index_1089423_comb;
  wire [7:0] p67_array_index_1089424_comb;
  wire [7:0] p67_array_index_1089425_comb;
  wire [7:0] p67_res7__355_comb;
  wire [7:0] p67_array_index_1089436_comb;
  wire [7:0] p67_array_index_1089437_comb;
  wire [7:0] p67_array_index_1089438_comb;
  wire [7:0] p67_array_index_1089439_comb;
  wire [7:0] p67_res7__356_comb;
  assign p67_addedKey__63_comb = p66_xor_1089321 ^ 128'he65a_edb1_c831_097f_c9c0_34b3_188d_3e17;
  assign p67_array_index_1089359_comb = p66_arr[p67_addedKey__63_comb[127:120]];
  assign p67_array_index_1089360_comb = p66_arr[p67_addedKey__63_comb[119:112]];
  assign p67_array_index_1089361_comb = p66_arr[p67_addedKey__63_comb[111:104]];
  assign p67_array_index_1089362_comb = p66_arr[p67_addedKey__63_comb[103:96]];
  assign p67_array_index_1089363_comb = p66_arr[p67_addedKey__63_comb[95:88]];
  assign p67_array_index_1089364_comb = p66_arr[p67_addedKey__63_comb[87:80]];
  assign p67_array_index_1089366_comb = p66_arr[p67_addedKey__63_comb[71:64]];
  assign p67_array_index_1089368_comb = p66_arr[p67_addedKey__63_comb[55:48]];
  assign p67_array_index_1089369_comb = p66_arr[p67_addedKey__63_comb[47:40]];
  assign p67_array_index_1089370_comb = p66_arr[p67_addedKey__63_comb[39:32]];
  assign p67_array_index_1089371_comb = p66_arr[p67_addedKey__63_comb[31:24]];
  assign p67_array_index_1089372_comb = p66_arr[p67_addedKey__63_comb[23:16]];
  assign p67_array_index_1089373_comb = p66_arr[p67_addedKey__63_comb[15:8]];
  assign p67_array_index_1089375_comb = p66_literal_1076345[p67_array_index_1089359_comb];
  assign p67_array_index_1089376_comb = p66_literal_1076347[p67_array_index_1089360_comb];
  assign p67_array_index_1089377_comb = p66_literal_1076349[p67_array_index_1089361_comb];
  assign p67_array_index_1089378_comb = p66_literal_1076351[p67_array_index_1089362_comb];
  assign p67_array_index_1089379_comb = p66_literal_1076353[p67_array_index_1089363_comb];
  assign p67_array_index_1089380_comb = p66_literal_1076355[p67_array_index_1089364_comb];
  assign p67_array_index_1089381_comb = p66_arr[p67_addedKey__63_comb[79:72]];
  assign p67_array_index_1089383_comb = p66_arr[p67_addedKey__63_comb[63:56]];
  assign p67_res7__352_comb = p67_array_index_1089375_comb ^ p67_array_index_1089376_comb ^ p67_array_index_1089377_comb ^ p67_array_index_1089378_comb ^ p67_array_index_1089379_comb ^ p67_array_index_1089380_comb ^ p67_array_index_1089381_comb ^ p66_literal_1076358[p67_array_index_1089366_comb] ^ p67_array_index_1089383_comb ^ p66_literal_1076355[p67_array_index_1089368_comb] ^ p66_literal_1076353[p67_array_index_1089369_comb] ^ p66_literal_1076351[p67_array_index_1089370_comb] ^ p66_literal_1076349[p67_array_index_1089371_comb] ^ p66_literal_1076347[p67_array_index_1089372_comb] ^ p66_literal_1076345[p67_array_index_1089373_comb] ^ p66_arr[p67_addedKey__63_comb[7:0]];
  assign p67_array_index_1089392_comb = p66_literal_1076345[p67_res7__352_comb];
  assign p67_array_index_1089393_comb = p66_literal_1076347[p67_array_index_1089359_comb];
  assign p67_array_index_1089394_comb = p66_literal_1076349[p67_array_index_1089360_comb];
  assign p67_array_index_1089395_comb = p66_literal_1076351[p67_array_index_1089361_comb];
  assign p67_array_index_1089396_comb = p66_literal_1076353[p67_array_index_1089362_comb];
  assign p67_array_index_1089397_comb = p66_literal_1076355[p67_array_index_1089363_comb];
  assign p67_res7__353_comb = p67_array_index_1089392_comb ^ p67_array_index_1089393_comb ^ p67_array_index_1089394_comb ^ p67_array_index_1089395_comb ^ p67_array_index_1089396_comb ^ p67_array_index_1089397_comb ^ p67_array_index_1089364_comb ^ p66_literal_1076358[p67_array_index_1089381_comb] ^ p67_array_index_1089366_comb ^ p66_literal_1076355[p67_array_index_1089383_comb] ^ p66_literal_1076353[p67_array_index_1089368_comb] ^ p66_literal_1076351[p67_array_index_1089369_comb] ^ p66_literal_1076349[p67_array_index_1089370_comb] ^ p66_literal_1076347[p67_array_index_1089371_comb] ^ p66_literal_1076345[p67_array_index_1089372_comb] ^ p67_array_index_1089373_comb;
  assign p67_array_index_1089407_comb = p66_literal_1076347[p67_res7__352_comb];
  assign p67_array_index_1089408_comb = p66_literal_1076349[p67_array_index_1089359_comb];
  assign p67_array_index_1089409_comb = p66_literal_1076351[p67_array_index_1089360_comb];
  assign p67_array_index_1089410_comb = p66_literal_1076353[p67_array_index_1089361_comb];
  assign p67_array_index_1089411_comb = p66_literal_1076355[p67_array_index_1089362_comb];
  assign p67_res7__354_comb = p66_literal_1076345[p67_res7__353_comb] ^ p67_array_index_1089407_comb ^ p67_array_index_1089408_comb ^ p67_array_index_1089409_comb ^ p67_array_index_1089410_comb ^ p67_array_index_1089411_comb ^ p67_array_index_1089363_comb ^ p66_literal_1076358[p67_array_index_1089364_comb] ^ p67_array_index_1089381_comb ^ p66_literal_1076355[p67_array_index_1089366_comb] ^ p66_literal_1076353[p67_array_index_1089383_comb] ^ p66_literal_1076351[p67_array_index_1089368_comb] ^ p66_literal_1076349[p67_array_index_1089369_comb] ^ p66_literal_1076347[p67_array_index_1089370_comb] ^ p66_literal_1076345[p67_array_index_1089371_comb] ^ p67_array_index_1089372_comb;
  assign p67_array_index_1089421_comb = p66_literal_1076347[p67_res7__353_comb];
  assign p67_array_index_1089422_comb = p66_literal_1076349[p67_res7__352_comb];
  assign p67_array_index_1089423_comb = p66_literal_1076351[p67_array_index_1089359_comb];
  assign p67_array_index_1089424_comb = p66_literal_1076353[p67_array_index_1089360_comb];
  assign p67_array_index_1089425_comb = p66_literal_1076355[p67_array_index_1089361_comb];
  assign p67_res7__355_comb = p66_literal_1076345[p67_res7__354_comb] ^ p67_array_index_1089421_comb ^ p67_array_index_1089422_comb ^ p67_array_index_1089423_comb ^ p67_array_index_1089424_comb ^ p67_array_index_1089425_comb ^ p67_array_index_1089362_comb ^ p66_literal_1076358[p67_array_index_1089363_comb] ^ p67_array_index_1089364_comb ^ p66_literal_1076355[p67_array_index_1089381_comb] ^ p66_literal_1076353[p67_array_index_1089366_comb] ^ p66_literal_1076351[p67_array_index_1089383_comb] ^ p66_literal_1076349[p67_array_index_1089368_comb] ^ p66_literal_1076347[p67_array_index_1089369_comb] ^ p66_literal_1076345[p67_array_index_1089370_comb] ^ p67_array_index_1089371_comb;
  assign p67_array_index_1089436_comb = p66_literal_1076349[p67_res7__353_comb];
  assign p67_array_index_1089437_comb = p66_literal_1076351[p67_res7__352_comb];
  assign p67_array_index_1089438_comb = p66_literal_1076353[p67_array_index_1089359_comb];
  assign p67_array_index_1089439_comb = p66_literal_1076355[p67_array_index_1089360_comb];
  assign p67_res7__356_comb = p66_literal_1076345[p67_res7__355_comb] ^ p66_literal_1076347[p67_res7__354_comb] ^ p67_array_index_1089436_comb ^ p67_array_index_1089437_comb ^ p67_array_index_1089438_comb ^ p67_array_index_1089439_comb ^ p67_array_index_1089361_comb ^ p66_literal_1076358[p67_array_index_1089362_comb] ^ p67_array_index_1089363_comb ^ p67_array_index_1089380_comb ^ p66_literal_1076353[p67_array_index_1089381_comb] ^ p66_literal_1076351[p67_array_index_1089366_comb] ^ p66_literal_1076349[p67_array_index_1089383_comb] ^ p66_literal_1076347[p67_array_index_1089368_comb] ^ p66_literal_1076345[p67_array_index_1089369_comb] ^ p67_array_index_1089370_comb;

  // Registers for pipe stage 67:
  reg [127:0] p67_xor_1088849;
  reg [127:0] p67_xor_1089321;
  reg [7:0] p67_array_index_1089359;
  reg [7:0] p67_array_index_1089360;
  reg [7:0] p67_array_index_1089361;
  reg [7:0] p67_array_index_1089362;
  reg [7:0] p67_array_index_1089363;
  reg [7:0] p67_array_index_1089364;
  reg [7:0] p67_array_index_1089366;
  reg [7:0] p67_array_index_1089368;
  reg [7:0] p67_array_index_1089369;
  reg [7:0] p67_array_index_1089375;
  reg [7:0] p67_array_index_1089376;
  reg [7:0] p67_array_index_1089377;
  reg [7:0] p67_array_index_1089378;
  reg [7:0] p67_array_index_1089379;
  reg [7:0] p67_array_index_1089381;
  reg [7:0] p67_array_index_1089383;
  reg [7:0] p67_res7__352;
  reg [7:0] p67_array_index_1089392;
  reg [7:0] p67_array_index_1089393;
  reg [7:0] p67_array_index_1089394;
  reg [7:0] p67_array_index_1089395;
  reg [7:0] p67_array_index_1089396;
  reg [7:0] p67_array_index_1089397;
  reg [7:0] p67_res7__353;
  reg [7:0] p67_array_index_1089407;
  reg [7:0] p67_array_index_1089408;
  reg [7:0] p67_array_index_1089409;
  reg [7:0] p67_array_index_1089410;
  reg [7:0] p67_array_index_1089411;
  reg [7:0] p67_res7__354;
  reg [7:0] p67_array_index_1089421;
  reg [7:0] p67_array_index_1089422;
  reg [7:0] p67_array_index_1089423;
  reg [7:0] p67_array_index_1089424;
  reg [7:0] p67_array_index_1089425;
  reg [7:0] p67_res7__355;
  reg [7:0] p67_array_index_1089436;
  reg [7:0] p67_array_index_1089437;
  reg [7:0] p67_array_index_1089438;
  reg [7:0] p67_array_index_1089439;
  reg [7:0] p67_res7__356;
  reg [127:0] p67_res__37;
  reg [7:0] p68_arr[256];
  reg [7:0] p68_literal_1076345[256];
  reg [7:0] p68_literal_1076347[256];
  reg [7:0] p68_literal_1076349[256];
  reg [7:0] p68_literal_1076351[256];
  reg [7:0] p68_literal_1076353[256];
  reg [7:0] p68_literal_1076355[256];
  reg [7:0] p68_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p67_xor_1088849 <= p66_xor_1088849;
    p67_xor_1089321 <= p66_xor_1089321;
    p67_array_index_1089359 <= p67_array_index_1089359_comb;
    p67_array_index_1089360 <= p67_array_index_1089360_comb;
    p67_array_index_1089361 <= p67_array_index_1089361_comb;
    p67_array_index_1089362 <= p67_array_index_1089362_comb;
    p67_array_index_1089363 <= p67_array_index_1089363_comb;
    p67_array_index_1089364 <= p67_array_index_1089364_comb;
    p67_array_index_1089366 <= p67_array_index_1089366_comb;
    p67_array_index_1089368 <= p67_array_index_1089368_comb;
    p67_array_index_1089369 <= p67_array_index_1089369_comb;
    p67_array_index_1089375 <= p67_array_index_1089375_comb;
    p67_array_index_1089376 <= p67_array_index_1089376_comb;
    p67_array_index_1089377 <= p67_array_index_1089377_comb;
    p67_array_index_1089378 <= p67_array_index_1089378_comb;
    p67_array_index_1089379 <= p67_array_index_1089379_comb;
    p67_array_index_1089381 <= p67_array_index_1089381_comb;
    p67_array_index_1089383 <= p67_array_index_1089383_comb;
    p67_res7__352 <= p67_res7__352_comb;
    p67_array_index_1089392 <= p67_array_index_1089392_comb;
    p67_array_index_1089393 <= p67_array_index_1089393_comb;
    p67_array_index_1089394 <= p67_array_index_1089394_comb;
    p67_array_index_1089395 <= p67_array_index_1089395_comb;
    p67_array_index_1089396 <= p67_array_index_1089396_comb;
    p67_array_index_1089397 <= p67_array_index_1089397_comb;
    p67_res7__353 <= p67_res7__353_comb;
    p67_array_index_1089407 <= p67_array_index_1089407_comb;
    p67_array_index_1089408 <= p67_array_index_1089408_comb;
    p67_array_index_1089409 <= p67_array_index_1089409_comb;
    p67_array_index_1089410 <= p67_array_index_1089410_comb;
    p67_array_index_1089411 <= p67_array_index_1089411_comb;
    p67_res7__354 <= p67_res7__354_comb;
    p67_array_index_1089421 <= p67_array_index_1089421_comb;
    p67_array_index_1089422 <= p67_array_index_1089422_comb;
    p67_array_index_1089423 <= p67_array_index_1089423_comb;
    p67_array_index_1089424 <= p67_array_index_1089424_comb;
    p67_array_index_1089425 <= p67_array_index_1089425_comb;
    p67_res7__355 <= p67_res7__355_comb;
    p67_array_index_1089436 <= p67_array_index_1089436_comb;
    p67_array_index_1089437 <= p67_array_index_1089437_comb;
    p67_array_index_1089438 <= p67_array_index_1089438_comb;
    p67_array_index_1089439 <= p67_array_index_1089439_comb;
    p67_res7__356 <= p67_res7__356_comb;
    p67_res__37 <= p66_res__37;
    p68_arr <= p67_arr;
    p68_literal_1076345 <= p67_literal_1076345;
    p68_literal_1076347 <= p67_literal_1076347;
    p68_literal_1076349 <= p67_literal_1076349;
    p68_literal_1076351 <= p67_literal_1076351;
    p68_literal_1076353 <= p67_literal_1076353;
    p68_literal_1076355 <= p67_literal_1076355;
    p68_literal_1076358 <= p67_literal_1076358;
  end

  // ===== Pipe stage 68:
  wire [7:0] p68_array_index_1089553_comb;
  wire [7:0] p68_array_index_1089554_comb;
  wire [7:0] p68_array_index_1089555_comb;
  wire [7:0] p68_array_index_1089556_comb;
  wire [7:0] p68_res7__357_comb;
  wire [7:0] p68_array_index_1089567_comb;
  wire [7:0] p68_array_index_1089568_comb;
  wire [7:0] p68_array_index_1089569_comb;
  wire [7:0] p68_res7__358_comb;
  wire [7:0] p68_array_index_1089579_comb;
  wire [7:0] p68_array_index_1089580_comb;
  wire [7:0] p68_array_index_1089581_comb;
  wire [7:0] p68_res7__359_comb;
  wire [7:0] p68_array_index_1089592_comb;
  wire [7:0] p68_array_index_1089593_comb;
  wire [7:0] p68_res7__360_comb;
  wire [7:0] p68_array_index_1089603_comb;
  wire [7:0] p68_array_index_1089604_comb;
  wire [7:0] p68_res7__361_comb;
  wire [7:0] p68_array_index_1089610_comb;
  wire [7:0] p68_array_index_1089611_comb;
  wire [7:0] p68_array_index_1089612_comb;
  wire [7:0] p68_array_index_1089613_comb;
  wire [7:0] p68_array_index_1089614_comb;
  wire [7:0] p68_array_index_1089615_comb;
  wire [7:0] p68_array_index_1089616_comb;
  wire [7:0] p68_array_index_1089617_comb;
  wire [7:0] p68_array_index_1089618_comb;
  assign p68_array_index_1089553_comb = p67_literal_1076349[p67_res7__354];
  assign p68_array_index_1089554_comb = p67_literal_1076351[p67_res7__353];
  assign p68_array_index_1089555_comb = p67_literal_1076353[p67_res7__352];
  assign p68_array_index_1089556_comb = p67_literal_1076355[p67_array_index_1089359];
  assign p68_res7__357_comb = p67_literal_1076345[p67_res7__356] ^ p67_literal_1076347[p67_res7__355] ^ p68_array_index_1089553_comb ^ p68_array_index_1089554_comb ^ p68_array_index_1089555_comb ^ p68_array_index_1089556_comb ^ p67_array_index_1089360 ^ p67_literal_1076358[p67_array_index_1089361] ^ p67_array_index_1089362 ^ p67_array_index_1089397 ^ p67_literal_1076353[p67_array_index_1089364] ^ p67_literal_1076351[p67_array_index_1089381] ^ p67_literal_1076349[p67_array_index_1089366] ^ p67_literal_1076347[p67_array_index_1089383] ^ p67_literal_1076345[p67_array_index_1089368] ^ p67_array_index_1089369;
  assign p68_array_index_1089567_comb = p67_literal_1076351[p67_res7__354];
  assign p68_array_index_1089568_comb = p67_literal_1076353[p67_res7__353];
  assign p68_array_index_1089569_comb = p67_literal_1076355[p67_res7__352];
  assign p68_res7__358_comb = p67_literal_1076345[p68_res7__357_comb] ^ p67_literal_1076347[p67_res7__356] ^ p67_literal_1076349[p67_res7__355] ^ p68_array_index_1089567_comb ^ p68_array_index_1089568_comb ^ p68_array_index_1089569_comb ^ p67_array_index_1089359 ^ p67_literal_1076358[p67_array_index_1089360] ^ p67_array_index_1089361 ^ p67_array_index_1089411 ^ p67_array_index_1089379 ^ p67_literal_1076351[p67_array_index_1089364] ^ p67_literal_1076349[p67_array_index_1089381] ^ p67_literal_1076347[p67_array_index_1089366] ^ p67_literal_1076345[p67_array_index_1089383] ^ p67_array_index_1089368;
  assign p68_array_index_1089579_comb = p67_literal_1076351[p67_res7__355];
  assign p68_array_index_1089580_comb = p67_literal_1076353[p67_res7__354];
  assign p68_array_index_1089581_comb = p67_literal_1076355[p67_res7__353];
  assign p68_res7__359_comb = p67_literal_1076345[p68_res7__358_comb] ^ p67_literal_1076347[p68_res7__357_comb] ^ p67_literal_1076349[p67_res7__356] ^ p68_array_index_1089579_comb ^ p68_array_index_1089580_comb ^ p68_array_index_1089581_comb ^ p67_res7__352 ^ p67_literal_1076358[p67_array_index_1089359] ^ p67_array_index_1089360 ^ p67_array_index_1089425 ^ p67_array_index_1089396 ^ p67_literal_1076351[p67_array_index_1089363] ^ p67_literal_1076349[p67_array_index_1089364] ^ p67_literal_1076347[p67_array_index_1089381] ^ p67_literal_1076345[p67_array_index_1089366] ^ p67_array_index_1089383;
  assign p68_array_index_1089592_comb = p67_literal_1076353[p67_res7__355];
  assign p68_array_index_1089593_comb = p67_literal_1076355[p67_res7__354];
  assign p68_res7__360_comb = p67_literal_1076345[p68_res7__359_comb] ^ p67_literal_1076347[p68_res7__358_comb] ^ p67_literal_1076349[p68_res7__357_comb] ^ p67_literal_1076351[p67_res7__356] ^ p68_array_index_1089592_comb ^ p68_array_index_1089593_comb ^ p67_res7__353 ^ p67_literal_1076358[p67_res7__352] ^ p67_array_index_1089359 ^ p67_array_index_1089439 ^ p67_array_index_1089410 ^ p67_array_index_1089378 ^ p67_literal_1076349[p67_array_index_1089363] ^ p67_literal_1076347[p67_array_index_1089364] ^ p67_literal_1076345[p67_array_index_1089381] ^ p67_array_index_1089366;
  assign p68_array_index_1089603_comb = p67_literal_1076353[p67_res7__356];
  assign p68_array_index_1089604_comb = p67_literal_1076355[p67_res7__355];
  assign p68_res7__361_comb = p67_literal_1076345[p68_res7__360_comb] ^ p67_literal_1076347[p68_res7__359_comb] ^ p67_literal_1076349[p68_res7__358_comb] ^ p67_literal_1076351[p68_res7__357_comb] ^ p68_array_index_1089603_comb ^ p68_array_index_1089604_comb ^ p67_res7__354 ^ p67_literal_1076358[p67_res7__353] ^ p67_res7__352 ^ p68_array_index_1089556_comb ^ p67_array_index_1089424 ^ p67_array_index_1089395 ^ p67_literal_1076349[p67_array_index_1089362] ^ p67_literal_1076347[p67_array_index_1089363] ^ p67_literal_1076345[p67_array_index_1089364] ^ p67_array_index_1089381;
  assign p68_array_index_1089610_comb = p67_literal_1076345[p68_res7__361_comb];
  assign p68_array_index_1089611_comb = p67_literal_1076347[p68_res7__360_comb];
  assign p68_array_index_1089612_comb = p67_literal_1076349[p68_res7__359_comb];
  assign p68_array_index_1089613_comb = p67_literal_1076351[p68_res7__358_comb];
  assign p68_array_index_1089614_comb = p67_literal_1076353[p68_res7__357_comb];
  assign p68_array_index_1089615_comb = p67_literal_1076355[p67_res7__356];
  assign p68_array_index_1089616_comb = p67_literal_1076358[p67_res7__354];
  assign p68_array_index_1089617_comb = p67_literal_1076347[p67_array_index_1089362];
  assign p68_array_index_1089618_comb = p67_literal_1076345[p67_array_index_1089363];

  // Registers for pipe stage 68:
  reg [127:0] p68_xor_1088849;
  reg [127:0] p68_xor_1089321;
  reg [7:0] p68_array_index_1089359;
  reg [7:0] p68_array_index_1089360;
  reg [7:0] p68_array_index_1089361;
  reg [7:0] p68_array_index_1089362;
  reg [7:0] p68_array_index_1089363;
  reg [7:0] p68_array_index_1089364;
  reg [7:0] p68_array_index_1089375;
  reg [7:0] p68_array_index_1089376;
  reg [7:0] p68_array_index_1089377;
  reg [7:0] p68_res7__352;
  reg [7:0] p68_array_index_1089392;
  reg [7:0] p68_array_index_1089393;
  reg [7:0] p68_array_index_1089394;
  reg [7:0] p68_res7__353;
  reg [7:0] p68_array_index_1089407;
  reg [7:0] p68_array_index_1089408;
  reg [7:0] p68_array_index_1089409;
  reg [7:0] p68_res7__354;
  reg [7:0] p68_array_index_1089421;
  reg [7:0] p68_array_index_1089422;
  reg [7:0] p68_array_index_1089423;
  reg [7:0] p68_res7__355;
  reg [7:0] p68_array_index_1089436;
  reg [7:0] p68_array_index_1089437;
  reg [7:0] p68_array_index_1089438;
  reg [7:0] p68_res7__356;
  reg [7:0] p68_array_index_1089553;
  reg [7:0] p68_array_index_1089554;
  reg [7:0] p68_array_index_1089555;
  reg [7:0] p68_res7__357;
  reg [7:0] p68_array_index_1089567;
  reg [7:0] p68_array_index_1089568;
  reg [7:0] p68_array_index_1089569;
  reg [7:0] p68_res7__358;
  reg [7:0] p68_array_index_1089579;
  reg [7:0] p68_array_index_1089580;
  reg [7:0] p68_array_index_1089581;
  reg [7:0] p68_res7__359;
  reg [7:0] p68_array_index_1089592;
  reg [7:0] p68_array_index_1089593;
  reg [7:0] p68_res7__360;
  reg [7:0] p68_array_index_1089603;
  reg [7:0] p68_array_index_1089604;
  reg [7:0] p68_res7__361;
  reg [7:0] p68_array_index_1089610;
  reg [7:0] p68_array_index_1089611;
  reg [7:0] p68_array_index_1089612;
  reg [7:0] p68_array_index_1089613;
  reg [7:0] p68_array_index_1089614;
  reg [7:0] p68_array_index_1089615;
  reg [7:0] p68_array_index_1089616;
  reg [7:0] p68_array_index_1089617;
  reg [7:0] p68_array_index_1089618;
  reg [127:0] p68_res__37;
  reg [7:0] p69_arr[256];
  reg [7:0] p69_literal_1076345[256];
  reg [7:0] p69_literal_1076347[256];
  reg [7:0] p69_literal_1076349[256];
  reg [7:0] p69_literal_1076351[256];
  reg [7:0] p69_literal_1076353[256];
  reg [7:0] p69_literal_1076355[256];
  reg [7:0] p69_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p68_xor_1088849 <= p67_xor_1088849;
    p68_xor_1089321 <= p67_xor_1089321;
    p68_array_index_1089359 <= p67_array_index_1089359;
    p68_array_index_1089360 <= p67_array_index_1089360;
    p68_array_index_1089361 <= p67_array_index_1089361;
    p68_array_index_1089362 <= p67_array_index_1089362;
    p68_array_index_1089363 <= p67_array_index_1089363;
    p68_array_index_1089364 <= p67_array_index_1089364;
    p68_array_index_1089375 <= p67_array_index_1089375;
    p68_array_index_1089376 <= p67_array_index_1089376;
    p68_array_index_1089377 <= p67_array_index_1089377;
    p68_res7__352 <= p67_res7__352;
    p68_array_index_1089392 <= p67_array_index_1089392;
    p68_array_index_1089393 <= p67_array_index_1089393;
    p68_array_index_1089394 <= p67_array_index_1089394;
    p68_res7__353 <= p67_res7__353;
    p68_array_index_1089407 <= p67_array_index_1089407;
    p68_array_index_1089408 <= p67_array_index_1089408;
    p68_array_index_1089409 <= p67_array_index_1089409;
    p68_res7__354 <= p67_res7__354;
    p68_array_index_1089421 <= p67_array_index_1089421;
    p68_array_index_1089422 <= p67_array_index_1089422;
    p68_array_index_1089423 <= p67_array_index_1089423;
    p68_res7__355 <= p67_res7__355;
    p68_array_index_1089436 <= p67_array_index_1089436;
    p68_array_index_1089437 <= p67_array_index_1089437;
    p68_array_index_1089438 <= p67_array_index_1089438;
    p68_res7__356 <= p67_res7__356;
    p68_array_index_1089553 <= p68_array_index_1089553_comb;
    p68_array_index_1089554 <= p68_array_index_1089554_comb;
    p68_array_index_1089555 <= p68_array_index_1089555_comb;
    p68_res7__357 <= p68_res7__357_comb;
    p68_array_index_1089567 <= p68_array_index_1089567_comb;
    p68_array_index_1089568 <= p68_array_index_1089568_comb;
    p68_array_index_1089569 <= p68_array_index_1089569_comb;
    p68_res7__358 <= p68_res7__358_comb;
    p68_array_index_1089579 <= p68_array_index_1089579_comb;
    p68_array_index_1089580 <= p68_array_index_1089580_comb;
    p68_array_index_1089581 <= p68_array_index_1089581_comb;
    p68_res7__359 <= p68_res7__359_comb;
    p68_array_index_1089592 <= p68_array_index_1089592_comb;
    p68_array_index_1089593 <= p68_array_index_1089593_comb;
    p68_res7__360 <= p68_res7__360_comb;
    p68_array_index_1089603 <= p68_array_index_1089603_comb;
    p68_array_index_1089604 <= p68_array_index_1089604_comb;
    p68_res7__361 <= p68_res7__361_comb;
    p68_array_index_1089610 <= p68_array_index_1089610_comb;
    p68_array_index_1089611 <= p68_array_index_1089611_comb;
    p68_array_index_1089612 <= p68_array_index_1089612_comb;
    p68_array_index_1089613 <= p68_array_index_1089613_comb;
    p68_array_index_1089614 <= p68_array_index_1089614_comb;
    p68_array_index_1089615 <= p68_array_index_1089615_comb;
    p68_array_index_1089616 <= p68_array_index_1089616_comb;
    p68_array_index_1089617 <= p68_array_index_1089617_comb;
    p68_array_index_1089618 <= p68_array_index_1089618_comb;
    p68_res__37 <= p67_res__37;
    p69_arr <= p68_arr;
    p69_literal_1076345 <= p68_literal_1076345;
    p69_literal_1076347 <= p68_literal_1076347;
    p69_literal_1076349 <= p68_literal_1076349;
    p69_literal_1076351 <= p68_literal_1076351;
    p69_literal_1076353 <= p68_literal_1076353;
    p69_literal_1076355 <= p68_literal_1076355;
    p69_literal_1076358 <= p68_literal_1076358;
  end

  // ===== Pipe stage 69:
  wire [7:0] p69_res7__362_comb;
  wire [7:0] p69_array_index_1089753_comb;
  wire [7:0] p69_res7__363_comb;
  wire [7:0] p69_res7__364_comb;
  wire [7:0] p69_res7__365_comb;
  wire [7:0] p69_res7__366_comb;
  wire [7:0] p69_res7__367_comb;
  wire [127:0] p69_res__22_comb;
  wire [127:0] p69_k7_comb;
  assign p69_res7__362_comb = p68_array_index_1089610 ^ p68_array_index_1089611 ^ p68_array_index_1089612 ^ p68_array_index_1089613 ^ p68_array_index_1089614 ^ p68_array_index_1089615 ^ p68_res7__355 ^ p68_array_index_1089616 ^ p68_res7__353 ^ p68_array_index_1089569 ^ p68_array_index_1089438 ^ p68_array_index_1089409 ^ p68_array_index_1089377 ^ p68_array_index_1089617 ^ p68_array_index_1089618 ^ p68_array_index_1089364;
  assign p69_array_index_1089753_comb = p68_literal_1076355[p68_res7__357];
  assign p69_res7__363_comb = p68_literal_1076345[p69_res7__362_comb] ^ p68_literal_1076347[p68_res7__361] ^ p68_literal_1076349[p68_res7__360] ^ p68_literal_1076351[p68_res7__359] ^ p68_literal_1076353[p68_res7__358] ^ p69_array_index_1089753_comb ^ p68_res7__356 ^ p68_literal_1076358[p68_res7__355] ^ p68_res7__354 ^ p68_array_index_1089581 ^ p68_array_index_1089555 ^ p68_array_index_1089423 ^ p68_array_index_1089394 ^ p68_literal_1076347[p68_array_index_1089361] ^ p68_literal_1076345[p68_array_index_1089362] ^ p68_array_index_1089363;
  assign p69_res7__364_comb = p68_literal_1076345[p69_res7__363_comb] ^ p68_literal_1076347[p69_res7__362_comb] ^ p68_literal_1076349[p68_res7__361] ^ p68_literal_1076351[p68_res7__360] ^ p68_literal_1076353[p68_res7__359] ^ p68_literal_1076355[p68_res7__358] ^ p68_res7__357 ^ p68_literal_1076358[p68_res7__356] ^ p68_res7__355 ^ p68_array_index_1089593 ^ p68_array_index_1089568 ^ p68_array_index_1089437 ^ p68_array_index_1089408 ^ p68_array_index_1089376 ^ p68_literal_1076345[p68_array_index_1089361] ^ p68_array_index_1089362;
  assign p69_res7__365_comb = p68_literal_1076345[p69_res7__364_comb] ^ p68_literal_1076347[p69_res7__363_comb] ^ p68_literal_1076349[p69_res7__362_comb] ^ p68_literal_1076351[p68_res7__361] ^ p68_literal_1076353[p68_res7__360] ^ p68_literal_1076355[p68_res7__359] ^ p68_res7__358 ^ p68_literal_1076358[p68_res7__357] ^ p68_res7__356 ^ p68_array_index_1089604 ^ p68_array_index_1089580 ^ p68_array_index_1089554 ^ p68_array_index_1089422 ^ p68_array_index_1089393 ^ p68_literal_1076345[p68_array_index_1089360] ^ p68_array_index_1089361;
  assign p69_res7__366_comb = p68_literal_1076345[p69_res7__365_comb] ^ p68_literal_1076347[p69_res7__364_comb] ^ p68_literal_1076349[p69_res7__363_comb] ^ p68_literal_1076351[p69_res7__362_comb] ^ p68_literal_1076353[p68_res7__361] ^ p68_literal_1076355[p68_res7__360] ^ p68_res7__359 ^ p68_literal_1076358[p68_res7__358] ^ p68_res7__357 ^ p68_array_index_1089615 ^ p68_array_index_1089592 ^ p68_array_index_1089567 ^ p68_array_index_1089436 ^ p68_array_index_1089407 ^ p68_array_index_1089375 ^ p68_array_index_1089360;
  assign p69_res7__367_comb = p68_literal_1076345[p69_res7__366_comb] ^ p68_literal_1076347[p69_res7__365_comb] ^ p68_literal_1076349[p69_res7__364_comb] ^ p68_literal_1076351[p69_res7__363_comb] ^ p68_literal_1076353[p69_res7__362_comb] ^ p68_literal_1076355[p68_res7__361] ^ p68_res7__360 ^ p68_literal_1076358[p68_res7__359] ^ p68_res7__358 ^ p69_array_index_1089753_comb ^ p68_array_index_1089603 ^ p68_array_index_1089579 ^ p68_array_index_1089553 ^ p68_array_index_1089421 ^ p68_array_index_1089392 ^ p68_array_index_1089359;
  assign p69_res__22_comb = {p69_res7__367_comb, p69_res7__366_comb, p69_res7__365_comb, p69_res7__364_comb, p69_res7__363_comb, p69_res7__362_comb, p68_res7__361, p68_res7__360, p68_res7__359, p68_res7__358, p68_res7__357, p68_res7__356, p68_res7__355, p68_res7__354, p68_res7__353, p68_res7__352};
  assign p69_k7_comb = p69_res__22_comb ^ p68_xor_1088849;

  // Registers for pipe stage 69:
  reg [127:0] p69_xor_1089321;
  reg [127:0] p69_k7;
  reg [127:0] p69_res__37;
  reg [7:0] p70_arr[256];
  reg [7:0] p70_literal_1076345[256];
  reg [7:0] p70_literal_1076347[256];
  reg [7:0] p70_literal_1076349[256];
  reg [7:0] p70_literal_1076351[256];
  reg [7:0] p70_literal_1076353[256];
  reg [7:0] p70_literal_1076355[256];
  reg [7:0] p70_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p69_xor_1089321 <= p68_xor_1089321;
    p69_k7 <= p69_k7_comb;
    p69_res__37 <= p68_res__37;
    p70_arr <= p69_arr;
    p70_literal_1076345 <= p69_literal_1076345;
    p70_literal_1076347 <= p69_literal_1076347;
    p70_literal_1076349 <= p69_literal_1076349;
    p70_literal_1076351 <= p69_literal_1076351;
    p70_literal_1076353 <= p69_literal_1076353;
    p70_literal_1076355 <= p69_literal_1076355;
    p70_literal_1076358 <= p69_literal_1076358;
  end

  // ===== Pipe stage 70:
  wire [127:0] p70_addedKey__64_comb;
  wire [7:0] p70_array_index_1089831_comb;
  wire [7:0] p70_array_index_1089832_comb;
  wire [7:0] p70_array_index_1089833_comb;
  wire [7:0] p70_array_index_1089834_comb;
  wire [7:0] p70_array_index_1089835_comb;
  wire [7:0] p70_array_index_1089836_comb;
  wire [7:0] p70_array_index_1089838_comb;
  wire [7:0] p70_array_index_1089840_comb;
  wire [7:0] p70_array_index_1089841_comb;
  wire [7:0] p70_array_index_1089842_comb;
  wire [7:0] p70_array_index_1089843_comb;
  wire [7:0] p70_array_index_1089844_comb;
  wire [7:0] p70_array_index_1089845_comb;
  wire [7:0] p70_array_index_1089847_comb;
  wire [7:0] p70_array_index_1089848_comb;
  wire [7:0] p70_array_index_1089849_comb;
  wire [7:0] p70_array_index_1089850_comb;
  wire [7:0] p70_array_index_1089851_comb;
  wire [7:0] p70_array_index_1089852_comb;
  wire [7:0] p70_array_index_1089853_comb;
  wire [7:0] p70_array_index_1089855_comb;
  wire [7:0] p70_res7__368_comb;
  wire [7:0] p70_array_index_1089864_comb;
  wire [7:0] p70_array_index_1089865_comb;
  wire [7:0] p70_array_index_1089866_comb;
  wire [7:0] p70_array_index_1089867_comb;
  wire [7:0] p70_array_index_1089868_comb;
  wire [7:0] p70_array_index_1089869_comb;
  wire [7:0] p70_res7__369_comb;
  wire [7:0] p70_array_index_1089879_comb;
  wire [7:0] p70_array_index_1089880_comb;
  wire [7:0] p70_array_index_1089881_comb;
  wire [7:0] p70_array_index_1089882_comb;
  wire [7:0] p70_array_index_1089883_comb;
  wire [7:0] p70_res7__370_comb;
  wire [7:0] p70_array_index_1089893_comb;
  wire [7:0] p70_array_index_1089894_comb;
  wire [7:0] p70_array_index_1089895_comb;
  wire [7:0] p70_array_index_1089896_comb;
  wire [7:0] p70_array_index_1089897_comb;
  wire [7:0] p70_res7__371_comb;
  wire [7:0] p70_array_index_1089908_comb;
  wire [7:0] p70_array_index_1089909_comb;
  wire [7:0] p70_array_index_1089910_comb;
  wire [7:0] p70_array_index_1089911_comb;
  wire [7:0] p70_res7__372_comb;
  assign p70_addedKey__64_comb = p69_k7 ^ 128'hd9eb_5a3a_e90f_fa58_34ce_2043_693d_7e18;
  assign p70_array_index_1089831_comb = p69_arr[p70_addedKey__64_comb[127:120]];
  assign p70_array_index_1089832_comb = p69_arr[p70_addedKey__64_comb[119:112]];
  assign p70_array_index_1089833_comb = p69_arr[p70_addedKey__64_comb[111:104]];
  assign p70_array_index_1089834_comb = p69_arr[p70_addedKey__64_comb[103:96]];
  assign p70_array_index_1089835_comb = p69_arr[p70_addedKey__64_comb[95:88]];
  assign p70_array_index_1089836_comb = p69_arr[p70_addedKey__64_comb[87:80]];
  assign p70_array_index_1089838_comb = p69_arr[p70_addedKey__64_comb[71:64]];
  assign p70_array_index_1089840_comb = p69_arr[p70_addedKey__64_comb[55:48]];
  assign p70_array_index_1089841_comb = p69_arr[p70_addedKey__64_comb[47:40]];
  assign p70_array_index_1089842_comb = p69_arr[p70_addedKey__64_comb[39:32]];
  assign p70_array_index_1089843_comb = p69_arr[p70_addedKey__64_comb[31:24]];
  assign p70_array_index_1089844_comb = p69_arr[p70_addedKey__64_comb[23:16]];
  assign p70_array_index_1089845_comb = p69_arr[p70_addedKey__64_comb[15:8]];
  assign p70_array_index_1089847_comb = p69_literal_1076345[p70_array_index_1089831_comb];
  assign p70_array_index_1089848_comb = p69_literal_1076347[p70_array_index_1089832_comb];
  assign p70_array_index_1089849_comb = p69_literal_1076349[p70_array_index_1089833_comb];
  assign p70_array_index_1089850_comb = p69_literal_1076351[p70_array_index_1089834_comb];
  assign p70_array_index_1089851_comb = p69_literal_1076353[p70_array_index_1089835_comb];
  assign p70_array_index_1089852_comb = p69_literal_1076355[p70_array_index_1089836_comb];
  assign p70_array_index_1089853_comb = p69_arr[p70_addedKey__64_comb[79:72]];
  assign p70_array_index_1089855_comb = p69_arr[p70_addedKey__64_comb[63:56]];
  assign p70_res7__368_comb = p70_array_index_1089847_comb ^ p70_array_index_1089848_comb ^ p70_array_index_1089849_comb ^ p70_array_index_1089850_comb ^ p70_array_index_1089851_comb ^ p70_array_index_1089852_comb ^ p70_array_index_1089853_comb ^ p69_literal_1076358[p70_array_index_1089838_comb] ^ p70_array_index_1089855_comb ^ p69_literal_1076355[p70_array_index_1089840_comb] ^ p69_literal_1076353[p70_array_index_1089841_comb] ^ p69_literal_1076351[p70_array_index_1089842_comb] ^ p69_literal_1076349[p70_array_index_1089843_comb] ^ p69_literal_1076347[p70_array_index_1089844_comb] ^ p69_literal_1076345[p70_array_index_1089845_comb] ^ p69_arr[p70_addedKey__64_comb[7:0]];
  assign p70_array_index_1089864_comb = p69_literal_1076345[p70_res7__368_comb];
  assign p70_array_index_1089865_comb = p69_literal_1076347[p70_array_index_1089831_comb];
  assign p70_array_index_1089866_comb = p69_literal_1076349[p70_array_index_1089832_comb];
  assign p70_array_index_1089867_comb = p69_literal_1076351[p70_array_index_1089833_comb];
  assign p70_array_index_1089868_comb = p69_literal_1076353[p70_array_index_1089834_comb];
  assign p70_array_index_1089869_comb = p69_literal_1076355[p70_array_index_1089835_comb];
  assign p70_res7__369_comb = p70_array_index_1089864_comb ^ p70_array_index_1089865_comb ^ p70_array_index_1089866_comb ^ p70_array_index_1089867_comb ^ p70_array_index_1089868_comb ^ p70_array_index_1089869_comb ^ p70_array_index_1089836_comb ^ p69_literal_1076358[p70_array_index_1089853_comb] ^ p70_array_index_1089838_comb ^ p69_literal_1076355[p70_array_index_1089855_comb] ^ p69_literal_1076353[p70_array_index_1089840_comb] ^ p69_literal_1076351[p70_array_index_1089841_comb] ^ p69_literal_1076349[p70_array_index_1089842_comb] ^ p69_literal_1076347[p70_array_index_1089843_comb] ^ p69_literal_1076345[p70_array_index_1089844_comb] ^ p70_array_index_1089845_comb;
  assign p70_array_index_1089879_comb = p69_literal_1076347[p70_res7__368_comb];
  assign p70_array_index_1089880_comb = p69_literal_1076349[p70_array_index_1089831_comb];
  assign p70_array_index_1089881_comb = p69_literal_1076351[p70_array_index_1089832_comb];
  assign p70_array_index_1089882_comb = p69_literal_1076353[p70_array_index_1089833_comb];
  assign p70_array_index_1089883_comb = p69_literal_1076355[p70_array_index_1089834_comb];
  assign p70_res7__370_comb = p69_literal_1076345[p70_res7__369_comb] ^ p70_array_index_1089879_comb ^ p70_array_index_1089880_comb ^ p70_array_index_1089881_comb ^ p70_array_index_1089882_comb ^ p70_array_index_1089883_comb ^ p70_array_index_1089835_comb ^ p69_literal_1076358[p70_array_index_1089836_comb] ^ p70_array_index_1089853_comb ^ p69_literal_1076355[p70_array_index_1089838_comb] ^ p69_literal_1076353[p70_array_index_1089855_comb] ^ p69_literal_1076351[p70_array_index_1089840_comb] ^ p69_literal_1076349[p70_array_index_1089841_comb] ^ p69_literal_1076347[p70_array_index_1089842_comb] ^ p69_literal_1076345[p70_array_index_1089843_comb] ^ p70_array_index_1089844_comb;
  assign p70_array_index_1089893_comb = p69_literal_1076347[p70_res7__369_comb];
  assign p70_array_index_1089894_comb = p69_literal_1076349[p70_res7__368_comb];
  assign p70_array_index_1089895_comb = p69_literal_1076351[p70_array_index_1089831_comb];
  assign p70_array_index_1089896_comb = p69_literal_1076353[p70_array_index_1089832_comb];
  assign p70_array_index_1089897_comb = p69_literal_1076355[p70_array_index_1089833_comb];
  assign p70_res7__371_comb = p69_literal_1076345[p70_res7__370_comb] ^ p70_array_index_1089893_comb ^ p70_array_index_1089894_comb ^ p70_array_index_1089895_comb ^ p70_array_index_1089896_comb ^ p70_array_index_1089897_comb ^ p70_array_index_1089834_comb ^ p69_literal_1076358[p70_array_index_1089835_comb] ^ p70_array_index_1089836_comb ^ p69_literal_1076355[p70_array_index_1089853_comb] ^ p69_literal_1076353[p70_array_index_1089838_comb] ^ p69_literal_1076351[p70_array_index_1089855_comb] ^ p69_literal_1076349[p70_array_index_1089840_comb] ^ p69_literal_1076347[p70_array_index_1089841_comb] ^ p69_literal_1076345[p70_array_index_1089842_comb] ^ p70_array_index_1089843_comb;
  assign p70_array_index_1089908_comb = p69_literal_1076349[p70_res7__369_comb];
  assign p70_array_index_1089909_comb = p69_literal_1076351[p70_res7__368_comb];
  assign p70_array_index_1089910_comb = p69_literal_1076353[p70_array_index_1089831_comb];
  assign p70_array_index_1089911_comb = p69_literal_1076355[p70_array_index_1089832_comb];
  assign p70_res7__372_comb = p69_literal_1076345[p70_res7__371_comb] ^ p69_literal_1076347[p70_res7__370_comb] ^ p70_array_index_1089908_comb ^ p70_array_index_1089909_comb ^ p70_array_index_1089910_comb ^ p70_array_index_1089911_comb ^ p70_array_index_1089833_comb ^ p69_literal_1076358[p70_array_index_1089834_comb] ^ p70_array_index_1089835_comb ^ p70_array_index_1089852_comb ^ p69_literal_1076353[p70_array_index_1089853_comb] ^ p69_literal_1076351[p70_array_index_1089838_comb] ^ p69_literal_1076349[p70_array_index_1089855_comb] ^ p69_literal_1076347[p70_array_index_1089840_comb] ^ p69_literal_1076345[p70_array_index_1089841_comb] ^ p70_array_index_1089842_comb;

  // Registers for pipe stage 70:
  reg [127:0] p70_xor_1089321;
  reg [127:0] p70_k7;
  reg [7:0] p70_array_index_1089831;
  reg [7:0] p70_array_index_1089832;
  reg [7:0] p70_array_index_1089833;
  reg [7:0] p70_array_index_1089834;
  reg [7:0] p70_array_index_1089835;
  reg [7:0] p70_array_index_1089836;
  reg [7:0] p70_array_index_1089838;
  reg [7:0] p70_array_index_1089840;
  reg [7:0] p70_array_index_1089841;
  reg [7:0] p70_array_index_1089847;
  reg [7:0] p70_array_index_1089848;
  reg [7:0] p70_array_index_1089849;
  reg [7:0] p70_array_index_1089850;
  reg [7:0] p70_array_index_1089851;
  reg [7:0] p70_array_index_1089853;
  reg [7:0] p70_array_index_1089855;
  reg [7:0] p70_res7__368;
  reg [7:0] p70_array_index_1089864;
  reg [7:0] p70_array_index_1089865;
  reg [7:0] p70_array_index_1089866;
  reg [7:0] p70_array_index_1089867;
  reg [7:0] p70_array_index_1089868;
  reg [7:0] p70_array_index_1089869;
  reg [7:0] p70_res7__369;
  reg [7:0] p70_array_index_1089879;
  reg [7:0] p70_array_index_1089880;
  reg [7:0] p70_array_index_1089881;
  reg [7:0] p70_array_index_1089882;
  reg [7:0] p70_array_index_1089883;
  reg [7:0] p70_res7__370;
  reg [7:0] p70_array_index_1089893;
  reg [7:0] p70_array_index_1089894;
  reg [7:0] p70_array_index_1089895;
  reg [7:0] p70_array_index_1089896;
  reg [7:0] p70_array_index_1089897;
  reg [7:0] p70_res7__371;
  reg [7:0] p70_array_index_1089908;
  reg [7:0] p70_array_index_1089909;
  reg [7:0] p70_array_index_1089910;
  reg [7:0] p70_array_index_1089911;
  reg [7:0] p70_res7__372;
  reg [127:0] p70_res__37;
  reg [7:0] p71_arr[256];
  reg [7:0] p71_literal_1076345[256];
  reg [7:0] p71_literal_1076347[256];
  reg [7:0] p71_literal_1076349[256];
  reg [7:0] p71_literal_1076351[256];
  reg [7:0] p71_literal_1076353[256];
  reg [7:0] p71_literal_1076355[256];
  reg [7:0] p71_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p70_xor_1089321 <= p69_xor_1089321;
    p70_k7 <= p69_k7;
    p70_array_index_1089831 <= p70_array_index_1089831_comb;
    p70_array_index_1089832 <= p70_array_index_1089832_comb;
    p70_array_index_1089833 <= p70_array_index_1089833_comb;
    p70_array_index_1089834 <= p70_array_index_1089834_comb;
    p70_array_index_1089835 <= p70_array_index_1089835_comb;
    p70_array_index_1089836 <= p70_array_index_1089836_comb;
    p70_array_index_1089838 <= p70_array_index_1089838_comb;
    p70_array_index_1089840 <= p70_array_index_1089840_comb;
    p70_array_index_1089841 <= p70_array_index_1089841_comb;
    p70_array_index_1089847 <= p70_array_index_1089847_comb;
    p70_array_index_1089848 <= p70_array_index_1089848_comb;
    p70_array_index_1089849 <= p70_array_index_1089849_comb;
    p70_array_index_1089850 <= p70_array_index_1089850_comb;
    p70_array_index_1089851 <= p70_array_index_1089851_comb;
    p70_array_index_1089853 <= p70_array_index_1089853_comb;
    p70_array_index_1089855 <= p70_array_index_1089855_comb;
    p70_res7__368 <= p70_res7__368_comb;
    p70_array_index_1089864 <= p70_array_index_1089864_comb;
    p70_array_index_1089865 <= p70_array_index_1089865_comb;
    p70_array_index_1089866 <= p70_array_index_1089866_comb;
    p70_array_index_1089867 <= p70_array_index_1089867_comb;
    p70_array_index_1089868 <= p70_array_index_1089868_comb;
    p70_array_index_1089869 <= p70_array_index_1089869_comb;
    p70_res7__369 <= p70_res7__369_comb;
    p70_array_index_1089879 <= p70_array_index_1089879_comb;
    p70_array_index_1089880 <= p70_array_index_1089880_comb;
    p70_array_index_1089881 <= p70_array_index_1089881_comb;
    p70_array_index_1089882 <= p70_array_index_1089882_comb;
    p70_array_index_1089883 <= p70_array_index_1089883_comb;
    p70_res7__370 <= p70_res7__370_comb;
    p70_array_index_1089893 <= p70_array_index_1089893_comb;
    p70_array_index_1089894 <= p70_array_index_1089894_comb;
    p70_array_index_1089895 <= p70_array_index_1089895_comb;
    p70_array_index_1089896 <= p70_array_index_1089896_comb;
    p70_array_index_1089897 <= p70_array_index_1089897_comb;
    p70_res7__371 <= p70_res7__371_comb;
    p70_array_index_1089908 <= p70_array_index_1089908_comb;
    p70_array_index_1089909 <= p70_array_index_1089909_comb;
    p70_array_index_1089910 <= p70_array_index_1089910_comb;
    p70_array_index_1089911 <= p70_array_index_1089911_comb;
    p70_res7__372 <= p70_res7__372_comb;
    p70_res__37 <= p69_res__37;
    p71_arr <= p70_arr;
    p71_literal_1076345 <= p70_literal_1076345;
    p71_literal_1076347 <= p70_literal_1076347;
    p71_literal_1076349 <= p70_literal_1076349;
    p71_literal_1076351 <= p70_literal_1076351;
    p71_literal_1076353 <= p70_literal_1076353;
    p71_literal_1076355 <= p70_literal_1076355;
    p71_literal_1076358 <= p70_literal_1076358;
  end

  // ===== Pipe stage 71:
  wire [7:0] p71_array_index_1090025_comb;
  wire [7:0] p71_array_index_1090026_comb;
  wire [7:0] p71_array_index_1090027_comb;
  wire [7:0] p71_array_index_1090028_comb;
  wire [7:0] p71_res7__373_comb;
  wire [7:0] p71_array_index_1090039_comb;
  wire [7:0] p71_array_index_1090040_comb;
  wire [7:0] p71_array_index_1090041_comb;
  wire [7:0] p71_res7__374_comb;
  wire [7:0] p71_array_index_1090051_comb;
  wire [7:0] p71_array_index_1090052_comb;
  wire [7:0] p71_array_index_1090053_comb;
  wire [7:0] p71_res7__375_comb;
  wire [7:0] p71_array_index_1090064_comb;
  wire [7:0] p71_array_index_1090065_comb;
  wire [7:0] p71_res7__376_comb;
  wire [7:0] p71_array_index_1090075_comb;
  wire [7:0] p71_array_index_1090076_comb;
  wire [7:0] p71_res7__377_comb;
  wire [7:0] p71_array_index_1090082_comb;
  wire [7:0] p71_array_index_1090083_comb;
  wire [7:0] p71_array_index_1090084_comb;
  wire [7:0] p71_array_index_1090085_comb;
  wire [7:0] p71_array_index_1090086_comb;
  wire [7:0] p71_array_index_1090087_comb;
  wire [7:0] p71_array_index_1090088_comb;
  wire [7:0] p71_array_index_1090089_comb;
  wire [7:0] p71_array_index_1090090_comb;
  assign p71_array_index_1090025_comb = p70_literal_1076349[p70_res7__370];
  assign p71_array_index_1090026_comb = p70_literal_1076351[p70_res7__369];
  assign p71_array_index_1090027_comb = p70_literal_1076353[p70_res7__368];
  assign p71_array_index_1090028_comb = p70_literal_1076355[p70_array_index_1089831];
  assign p71_res7__373_comb = p70_literal_1076345[p70_res7__372] ^ p70_literal_1076347[p70_res7__371] ^ p71_array_index_1090025_comb ^ p71_array_index_1090026_comb ^ p71_array_index_1090027_comb ^ p71_array_index_1090028_comb ^ p70_array_index_1089832 ^ p70_literal_1076358[p70_array_index_1089833] ^ p70_array_index_1089834 ^ p70_array_index_1089869 ^ p70_literal_1076353[p70_array_index_1089836] ^ p70_literal_1076351[p70_array_index_1089853] ^ p70_literal_1076349[p70_array_index_1089838] ^ p70_literal_1076347[p70_array_index_1089855] ^ p70_literal_1076345[p70_array_index_1089840] ^ p70_array_index_1089841;
  assign p71_array_index_1090039_comb = p70_literal_1076351[p70_res7__370];
  assign p71_array_index_1090040_comb = p70_literal_1076353[p70_res7__369];
  assign p71_array_index_1090041_comb = p70_literal_1076355[p70_res7__368];
  assign p71_res7__374_comb = p70_literal_1076345[p71_res7__373_comb] ^ p70_literal_1076347[p70_res7__372] ^ p70_literal_1076349[p70_res7__371] ^ p71_array_index_1090039_comb ^ p71_array_index_1090040_comb ^ p71_array_index_1090041_comb ^ p70_array_index_1089831 ^ p70_literal_1076358[p70_array_index_1089832] ^ p70_array_index_1089833 ^ p70_array_index_1089883 ^ p70_array_index_1089851 ^ p70_literal_1076351[p70_array_index_1089836] ^ p70_literal_1076349[p70_array_index_1089853] ^ p70_literal_1076347[p70_array_index_1089838] ^ p70_literal_1076345[p70_array_index_1089855] ^ p70_array_index_1089840;
  assign p71_array_index_1090051_comb = p70_literal_1076351[p70_res7__371];
  assign p71_array_index_1090052_comb = p70_literal_1076353[p70_res7__370];
  assign p71_array_index_1090053_comb = p70_literal_1076355[p70_res7__369];
  assign p71_res7__375_comb = p70_literal_1076345[p71_res7__374_comb] ^ p70_literal_1076347[p71_res7__373_comb] ^ p70_literal_1076349[p70_res7__372] ^ p71_array_index_1090051_comb ^ p71_array_index_1090052_comb ^ p71_array_index_1090053_comb ^ p70_res7__368 ^ p70_literal_1076358[p70_array_index_1089831] ^ p70_array_index_1089832 ^ p70_array_index_1089897 ^ p70_array_index_1089868 ^ p70_literal_1076351[p70_array_index_1089835] ^ p70_literal_1076349[p70_array_index_1089836] ^ p70_literal_1076347[p70_array_index_1089853] ^ p70_literal_1076345[p70_array_index_1089838] ^ p70_array_index_1089855;
  assign p71_array_index_1090064_comb = p70_literal_1076353[p70_res7__371];
  assign p71_array_index_1090065_comb = p70_literal_1076355[p70_res7__370];
  assign p71_res7__376_comb = p70_literal_1076345[p71_res7__375_comb] ^ p70_literal_1076347[p71_res7__374_comb] ^ p70_literal_1076349[p71_res7__373_comb] ^ p70_literal_1076351[p70_res7__372] ^ p71_array_index_1090064_comb ^ p71_array_index_1090065_comb ^ p70_res7__369 ^ p70_literal_1076358[p70_res7__368] ^ p70_array_index_1089831 ^ p70_array_index_1089911 ^ p70_array_index_1089882 ^ p70_array_index_1089850 ^ p70_literal_1076349[p70_array_index_1089835] ^ p70_literal_1076347[p70_array_index_1089836] ^ p70_literal_1076345[p70_array_index_1089853] ^ p70_array_index_1089838;
  assign p71_array_index_1090075_comb = p70_literal_1076353[p70_res7__372];
  assign p71_array_index_1090076_comb = p70_literal_1076355[p70_res7__371];
  assign p71_res7__377_comb = p70_literal_1076345[p71_res7__376_comb] ^ p70_literal_1076347[p71_res7__375_comb] ^ p70_literal_1076349[p71_res7__374_comb] ^ p70_literal_1076351[p71_res7__373_comb] ^ p71_array_index_1090075_comb ^ p71_array_index_1090076_comb ^ p70_res7__370 ^ p70_literal_1076358[p70_res7__369] ^ p70_res7__368 ^ p71_array_index_1090028_comb ^ p70_array_index_1089896 ^ p70_array_index_1089867 ^ p70_literal_1076349[p70_array_index_1089834] ^ p70_literal_1076347[p70_array_index_1089835] ^ p70_literal_1076345[p70_array_index_1089836] ^ p70_array_index_1089853;
  assign p71_array_index_1090082_comb = p70_literal_1076345[p71_res7__377_comb];
  assign p71_array_index_1090083_comb = p70_literal_1076347[p71_res7__376_comb];
  assign p71_array_index_1090084_comb = p70_literal_1076349[p71_res7__375_comb];
  assign p71_array_index_1090085_comb = p70_literal_1076351[p71_res7__374_comb];
  assign p71_array_index_1090086_comb = p70_literal_1076353[p71_res7__373_comb];
  assign p71_array_index_1090087_comb = p70_literal_1076355[p70_res7__372];
  assign p71_array_index_1090088_comb = p70_literal_1076358[p70_res7__370];
  assign p71_array_index_1090089_comb = p70_literal_1076347[p70_array_index_1089834];
  assign p71_array_index_1090090_comb = p70_literal_1076345[p70_array_index_1089835];

  // Registers for pipe stage 71:
  reg [127:0] p71_xor_1089321;
  reg [127:0] p71_k7;
  reg [7:0] p71_array_index_1089831;
  reg [7:0] p71_array_index_1089832;
  reg [7:0] p71_array_index_1089833;
  reg [7:0] p71_array_index_1089834;
  reg [7:0] p71_array_index_1089835;
  reg [7:0] p71_array_index_1089836;
  reg [7:0] p71_array_index_1089847;
  reg [7:0] p71_array_index_1089848;
  reg [7:0] p71_array_index_1089849;
  reg [7:0] p71_res7__368;
  reg [7:0] p71_array_index_1089864;
  reg [7:0] p71_array_index_1089865;
  reg [7:0] p71_array_index_1089866;
  reg [7:0] p71_res7__369;
  reg [7:0] p71_array_index_1089879;
  reg [7:0] p71_array_index_1089880;
  reg [7:0] p71_array_index_1089881;
  reg [7:0] p71_res7__370;
  reg [7:0] p71_array_index_1089893;
  reg [7:0] p71_array_index_1089894;
  reg [7:0] p71_array_index_1089895;
  reg [7:0] p71_res7__371;
  reg [7:0] p71_array_index_1089908;
  reg [7:0] p71_array_index_1089909;
  reg [7:0] p71_array_index_1089910;
  reg [7:0] p71_res7__372;
  reg [7:0] p71_array_index_1090025;
  reg [7:0] p71_array_index_1090026;
  reg [7:0] p71_array_index_1090027;
  reg [7:0] p71_res7__373;
  reg [7:0] p71_array_index_1090039;
  reg [7:0] p71_array_index_1090040;
  reg [7:0] p71_array_index_1090041;
  reg [7:0] p71_res7__374;
  reg [7:0] p71_array_index_1090051;
  reg [7:0] p71_array_index_1090052;
  reg [7:0] p71_array_index_1090053;
  reg [7:0] p71_res7__375;
  reg [7:0] p71_array_index_1090064;
  reg [7:0] p71_array_index_1090065;
  reg [7:0] p71_res7__376;
  reg [7:0] p71_array_index_1090075;
  reg [7:0] p71_array_index_1090076;
  reg [7:0] p71_res7__377;
  reg [7:0] p71_array_index_1090082;
  reg [7:0] p71_array_index_1090083;
  reg [7:0] p71_array_index_1090084;
  reg [7:0] p71_array_index_1090085;
  reg [7:0] p71_array_index_1090086;
  reg [7:0] p71_array_index_1090087;
  reg [7:0] p71_array_index_1090088;
  reg [7:0] p71_array_index_1090089;
  reg [7:0] p71_array_index_1090090;
  reg [127:0] p71_res__37;
  reg [7:0] p72_arr[256];
  reg [7:0] p72_literal_1076345[256];
  reg [7:0] p72_literal_1076347[256];
  reg [7:0] p72_literal_1076349[256];
  reg [7:0] p72_literal_1076351[256];
  reg [7:0] p72_literal_1076353[256];
  reg [7:0] p72_literal_1076355[256];
  reg [7:0] p72_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p71_xor_1089321 <= p70_xor_1089321;
    p71_k7 <= p70_k7;
    p71_array_index_1089831 <= p70_array_index_1089831;
    p71_array_index_1089832 <= p70_array_index_1089832;
    p71_array_index_1089833 <= p70_array_index_1089833;
    p71_array_index_1089834 <= p70_array_index_1089834;
    p71_array_index_1089835 <= p70_array_index_1089835;
    p71_array_index_1089836 <= p70_array_index_1089836;
    p71_array_index_1089847 <= p70_array_index_1089847;
    p71_array_index_1089848 <= p70_array_index_1089848;
    p71_array_index_1089849 <= p70_array_index_1089849;
    p71_res7__368 <= p70_res7__368;
    p71_array_index_1089864 <= p70_array_index_1089864;
    p71_array_index_1089865 <= p70_array_index_1089865;
    p71_array_index_1089866 <= p70_array_index_1089866;
    p71_res7__369 <= p70_res7__369;
    p71_array_index_1089879 <= p70_array_index_1089879;
    p71_array_index_1089880 <= p70_array_index_1089880;
    p71_array_index_1089881 <= p70_array_index_1089881;
    p71_res7__370 <= p70_res7__370;
    p71_array_index_1089893 <= p70_array_index_1089893;
    p71_array_index_1089894 <= p70_array_index_1089894;
    p71_array_index_1089895 <= p70_array_index_1089895;
    p71_res7__371 <= p70_res7__371;
    p71_array_index_1089908 <= p70_array_index_1089908;
    p71_array_index_1089909 <= p70_array_index_1089909;
    p71_array_index_1089910 <= p70_array_index_1089910;
    p71_res7__372 <= p70_res7__372;
    p71_array_index_1090025 <= p71_array_index_1090025_comb;
    p71_array_index_1090026 <= p71_array_index_1090026_comb;
    p71_array_index_1090027 <= p71_array_index_1090027_comb;
    p71_res7__373 <= p71_res7__373_comb;
    p71_array_index_1090039 <= p71_array_index_1090039_comb;
    p71_array_index_1090040 <= p71_array_index_1090040_comb;
    p71_array_index_1090041 <= p71_array_index_1090041_comb;
    p71_res7__374 <= p71_res7__374_comb;
    p71_array_index_1090051 <= p71_array_index_1090051_comb;
    p71_array_index_1090052 <= p71_array_index_1090052_comb;
    p71_array_index_1090053 <= p71_array_index_1090053_comb;
    p71_res7__375 <= p71_res7__375_comb;
    p71_array_index_1090064 <= p71_array_index_1090064_comb;
    p71_array_index_1090065 <= p71_array_index_1090065_comb;
    p71_res7__376 <= p71_res7__376_comb;
    p71_array_index_1090075 <= p71_array_index_1090075_comb;
    p71_array_index_1090076 <= p71_array_index_1090076_comb;
    p71_res7__377 <= p71_res7__377_comb;
    p71_array_index_1090082 <= p71_array_index_1090082_comb;
    p71_array_index_1090083 <= p71_array_index_1090083_comb;
    p71_array_index_1090084 <= p71_array_index_1090084_comb;
    p71_array_index_1090085 <= p71_array_index_1090085_comb;
    p71_array_index_1090086 <= p71_array_index_1090086_comb;
    p71_array_index_1090087 <= p71_array_index_1090087_comb;
    p71_array_index_1090088 <= p71_array_index_1090088_comb;
    p71_array_index_1090089 <= p71_array_index_1090089_comb;
    p71_array_index_1090090 <= p71_array_index_1090090_comb;
    p71_res__37 <= p70_res__37;
    p72_arr <= p71_arr;
    p72_literal_1076345 <= p71_literal_1076345;
    p72_literal_1076347 <= p71_literal_1076347;
    p72_literal_1076349 <= p71_literal_1076349;
    p72_literal_1076351 <= p71_literal_1076351;
    p72_literal_1076353 <= p71_literal_1076353;
    p72_literal_1076355 <= p71_literal_1076355;
    p72_literal_1076358 <= p71_literal_1076358;
  end

  // ===== Pipe stage 72:
  wire [7:0] p72_res7__378_comb;
  wire [7:0] p72_array_index_1090225_comb;
  wire [7:0] p72_res7__379_comb;
  wire [7:0] p72_res7__380_comb;
  wire [7:0] p72_res7__381_comb;
  wire [7:0] p72_res7__382_comb;
  wire [7:0] p72_res7__383_comb;
  wire [127:0] p72_res__23_comb;
  wire [127:0] p72_k6_comb;
  wire [127:0] p72_addedKey__38_comb;
  wire [7:0] p72_bit_slice_1090267_comb;
  wire [7:0] p72_bit_slice_1090268_comb;
  wire [7:0] p72_bit_slice_1090269_comb;
  wire [7:0] p72_bit_slice_1090270_comb;
  wire [7:0] p72_bit_slice_1090271_comb;
  wire [7:0] p72_bit_slice_1090272_comb;
  wire [7:0] p72_bit_slice_1090273_comb;
  wire [7:0] p72_bit_slice_1090274_comb;
  wire [7:0] p72_bit_slice_1090275_comb;
  wire [7:0] p72_bit_slice_1090276_comb;
  wire [7:0] p72_bit_slice_1090277_comb;
  wire [7:0] p72_bit_slice_1090278_comb;
  wire [7:0] p72_bit_slice_1090279_comb;
  wire [7:0] p72_bit_slice_1090280_comb;
  wire [7:0] p72_bit_slice_1090281_comb;
  wire [7:0] p72_bit_slice_1090282_comb;
  assign p72_res7__378_comb = p71_array_index_1090082 ^ p71_array_index_1090083 ^ p71_array_index_1090084 ^ p71_array_index_1090085 ^ p71_array_index_1090086 ^ p71_array_index_1090087 ^ p71_res7__371 ^ p71_array_index_1090088 ^ p71_res7__369 ^ p71_array_index_1090041 ^ p71_array_index_1089910 ^ p71_array_index_1089881 ^ p71_array_index_1089849 ^ p71_array_index_1090089 ^ p71_array_index_1090090 ^ p71_array_index_1089836;
  assign p72_array_index_1090225_comb = p71_literal_1076355[p71_res7__373];
  assign p72_res7__379_comb = p71_literal_1076345[p72_res7__378_comb] ^ p71_literal_1076347[p71_res7__377] ^ p71_literal_1076349[p71_res7__376] ^ p71_literal_1076351[p71_res7__375] ^ p71_literal_1076353[p71_res7__374] ^ p72_array_index_1090225_comb ^ p71_res7__372 ^ p71_literal_1076358[p71_res7__371] ^ p71_res7__370 ^ p71_array_index_1090053 ^ p71_array_index_1090027 ^ p71_array_index_1089895 ^ p71_array_index_1089866 ^ p71_literal_1076347[p71_array_index_1089833] ^ p71_literal_1076345[p71_array_index_1089834] ^ p71_array_index_1089835;
  assign p72_res7__380_comb = p71_literal_1076345[p72_res7__379_comb] ^ p71_literal_1076347[p72_res7__378_comb] ^ p71_literal_1076349[p71_res7__377] ^ p71_literal_1076351[p71_res7__376] ^ p71_literal_1076353[p71_res7__375] ^ p71_literal_1076355[p71_res7__374] ^ p71_res7__373 ^ p71_literal_1076358[p71_res7__372] ^ p71_res7__371 ^ p71_array_index_1090065 ^ p71_array_index_1090040 ^ p71_array_index_1089909 ^ p71_array_index_1089880 ^ p71_array_index_1089848 ^ p71_literal_1076345[p71_array_index_1089833] ^ p71_array_index_1089834;
  assign p72_res7__381_comb = p71_literal_1076345[p72_res7__380_comb] ^ p71_literal_1076347[p72_res7__379_comb] ^ p71_literal_1076349[p72_res7__378_comb] ^ p71_literal_1076351[p71_res7__377] ^ p71_literal_1076353[p71_res7__376] ^ p71_literal_1076355[p71_res7__375] ^ p71_res7__374 ^ p71_literal_1076358[p71_res7__373] ^ p71_res7__372 ^ p71_array_index_1090076 ^ p71_array_index_1090052 ^ p71_array_index_1090026 ^ p71_array_index_1089894 ^ p71_array_index_1089865 ^ p71_literal_1076345[p71_array_index_1089832] ^ p71_array_index_1089833;
  assign p72_res7__382_comb = p71_literal_1076345[p72_res7__381_comb] ^ p71_literal_1076347[p72_res7__380_comb] ^ p71_literal_1076349[p72_res7__379_comb] ^ p71_literal_1076351[p72_res7__378_comb] ^ p71_literal_1076353[p71_res7__377] ^ p71_literal_1076355[p71_res7__376] ^ p71_res7__375 ^ p71_literal_1076358[p71_res7__374] ^ p71_res7__373 ^ p71_array_index_1090087 ^ p71_array_index_1090064 ^ p71_array_index_1090039 ^ p71_array_index_1089908 ^ p71_array_index_1089879 ^ p71_array_index_1089847 ^ p71_array_index_1089832;
  assign p72_res7__383_comb = p71_literal_1076345[p72_res7__382_comb] ^ p71_literal_1076347[p72_res7__381_comb] ^ p71_literal_1076349[p72_res7__380_comb] ^ p71_literal_1076351[p72_res7__379_comb] ^ p71_literal_1076353[p72_res7__378_comb] ^ p71_literal_1076355[p71_res7__377] ^ p71_res7__376 ^ p71_literal_1076358[p71_res7__375] ^ p71_res7__374 ^ p72_array_index_1090225_comb ^ p71_array_index_1090075 ^ p71_array_index_1090051 ^ p71_array_index_1090025 ^ p71_array_index_1089893 ^ p71_array_index_1089864 ^ p71_array_index_1089831;
  assign p72_res__23_comb = {p72_res7__383_comb, p72_res7__382_comb, p72_res7__381_comb, p72_res7__380_comb, p72_res7__379_comb, p72_res7__378_comb, p71_res7__377, p71_res7__376, p71_res7__375, p71_res7__374, p71_res7__373, p71_res7__372, p71_res7__371, p71_res7__370, p71_res7__369, p71_res7__368};
  assign p72_k6_comb = p72_res__23_comb ^ p71_xor_1089321;
  assign p72_addedKey__38_comb = p72_k6_comb ^ p71_res__37;
  assign p72_bit_slice_1090267_comb = p72_addedKey__38_comb[127:120];
  assign p72_bit_slice_1090268_comb = p72_addedKey__38_comb[119:112];
  assign p72_bit_slice_1090269_comb = p72_addedKey__38_comb[111:104];
  assign p72_bit_slice_1090270_comb = p72_addedKey__38_comb[103:96];
  assign p72_bit_slice_1090271_comb = p72_addedKey__38_comb[95:88];
  assign p72_bit_slice_1090272_comb = p72_addedKey__38_comb[87:80];
  assign p72_bit_slice_1090273_comb = p72_addedKey__38_comb[71:64];
  assign p72_bit_slice_1090274_comb = p72_addedKey__38_comb[55:48];
  assign p72_bit_slice_1090275_comb = p72_addedKey__38_comb[47:40];
  assign p72_bit_slice_1090276_comb = p72_addedKey__38_comb[39:32];
  assign p72_bit_slice_1090277_comb = p72_addedKey__38_comb[31:24];
  assign p72_bit_slice_1090278_comb = p72_addedKey__38_comb[23:16];
  assign p72_bit_slice_1090279_comb = p72_addedKey__38_comb[15:8];
  assign p72_bit_slice_1090280_comb = p72_addedKey__38_comb[79:72];
  assign p72_bit_slice_1090281_comb = p72_addedKey__38_comb[63:56];
  assign p72_bit_slice_1090282_comb = p72_addedKey__38_comb[7:0];

  // Registers for pipe stage 72:
  reg [127:0] p72_k7;
  reg [127:0] p72_k6;
  reg [7:0] p72_bit_slice_1090267;
  reg [7:0] p72_bit_slice_1090268;
  reg [7:0] p72_bit_slice_1090269;
  reg [7:0] p72_bit_slice_1090270;
  reg [7:0] p72_bit_slice_1090271;
  reg [7:0] p72_bit_slice_1090272;
  reg [7:0] p72_bit_slice_1090273;
  reg [7:0] p72_bit_slice_1090274;
  reg [7:0] p72_bit_slice_1090275;
  reg [7:0] p72_bit_slice_1090276;
  reg [7:0] p72_bit_slice_1090277;
  reg [7:0] p72_bit_slice_1090278;
  reg [7:0] p72_bit_slice_1090279;
  reg [7:0] p72_bit_slice_1090280;
  reg [7:0] p72_bit_slice_1090281;
  reg [7:0] p72_bit_slice_1090282;
  reg [7:0] p73_arr[256];
  reg [7:0] p73_literal_1076345[256];
  reg [7:0] p73_literal_1076347[256];
  reg [7:0] p73_literal_1076349[256];
  reg [7:0] p73_literal_1076351[256];
  reg [7:0] p73_literal_1076353[256];
  reg [7:0] p73_literal_1076355[256];
  reg [7:0] p73_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p72_k7 <= p71_k7;
    p72_k6 <= p72_k6_comb;
    p72_bit_slice_1090267 <= p72_bit_slice_1090267_comb;
    p72_bit_slice_1090268 <= p72_bit_slice_1090268_comb;
    p72_bit_slice_1090269 <= p72_bit_slice_1090269_comb;
    p72_bit_slice_1090270 <= p72_bit_slice_1090270_comb;
    p72_bit_slice_1090271 <= p72_bit_slice_1090271_comb;
    p72_bit_slice_1090272 <= p72_bit_slice_1090272_comb;
    p72_bit_slice_1090273 <= p72_bit_slice_1090273_comb;
    p72_bit_slice_1090274 <= p72_bit_slice_1090274_comb;
    p72_bit_slice_1090275 <= p72_bit_slice_1090275_comb;
    p72_bit_slice_1090276 <= p72_bit_slice_1090276_comb;
    p72_bit_slice_1090277 <= p72_bit_slice_1090277_comb;
    p72_bit_slice_1090278 <= p72_bit_slice_1090278_comb;
    p72_bit_slice_1090279 <= p72_bit_slice_1090279_comb;
    p72_bit_slice_1090280 <= p72_bit_slice_1090280_comb;
    p72_bit_slice_1090281 <= p72_bit_slice_1090281_comb;
    p72_bit_slice_1090282 <= p72_bit_slice_1090282_comb;
    p73_arr <= p72_arr;
    p73_literal_1076345 <= p72_literal_1076345;
    p73_literal_1076347 <= p72_literal_1076347;
    p73_literal_1076349 <= p72_literal_1076349;
    p73_literal_1076351 <= p72_literal_1076351;
    p73_literal_1076353 <= p72_literal_1076353;
    p73_literal_1076355 <= p72_literal_1076355;
    p73_literal_1076358 <= p72_literal_1076358;
  end

  // ===== Pipe stage 73:
  wire [127:0] p73_addedKey__65_comb;
  wire [7:0] p73_array_index_1090350_comb;
  wire [7:0] p73_array_index_1090351_comb;
  wire [7:0] p73_array_index_1090352_comb;
  wire [7:0] p73_array_index_1090353_comb;
  wire [7:0] p73_array_index_1090354_comb;
  wire [7:0] p73_array_index_1090355_comb;
  wire [7:0] p73_array_index_1090357_comb;
  wire [7:0] p73_array_index_1090359_comb;
  wire [7:0] p73_array_index_1090360_comb;
  wire [7:0] p73_array_index_1090361_comb;
  wire [7:0] p73_array_index_1090362_comb;
  wire [7:0] p73_array_index_1090363_comb;
  wire [7:0] p73_array_index_1090364_comb;
  wire [7:0] p73_array_index_1090438_comb;
  wire [7:0] p73_array_index_1090439_comb;
  wire [7:0] p73_array_index_1090440_comb;
  wire [7:0] p73_array_index_1090441_comb;
  wire [7:0] p73_array_index_1090442_comb;
  wire [7:0] p73_array_index_1090443_comb;
  wire [7:0] p73_array_index_1090444_comb;
  wire [7:0] p73_array_index_1090445_comb;
  wire [7:0] p73_array_index_1090446_comb;
  wire [7:0] p73_array_index_1090447_comb;
  wire [7:0] p73_array_index_1090448_comb;
  wire [7:0] p73_array_index_1090449_comb;
  wire [7:0] p73_array_index_1090450_comb;
  wire [7:0] p73_array_index_1090366_comb;
  wire [7:0] p73_array_index_1090367_comb;
  wire [7:0] p73_array_index_1090368_comb;
  wire [7:0] p73_array_index_1090369_comb;
  wire [7:0] p73_array_index_1090370_comb;
  wire [7:0] p73_array_index_1090371_comb;
  wire [7:0] p73_array_index_1090372_comb;
  wire [7:0] p73_array_index_1090374_comb;
  wire [7:0] p73_array_index_1090451_comb;
  wire [7:0] p73_array_index_1090452_comb;
  wire [7:0] p73_array_index_1090453_comb;
  wire [7:0] p73_array_index_1090454_comb;
  wire [7:0] p73_array_index_1090455_comb;
  wire [7:0] p73_array_index_1090456_comb;
  wire [7:0] p73_array_index_1090457_comb;
  wire [7:0] p73_array_index_1090459_comb;
  wire [7:0] p73_res7__384_comb;
  wire [7:0] p73_res7__608_comb;
  wire [7:0] p73_array_index_1090383_comb;
  wire [7:0] p73_array_index_1090384_comb;
  wire [7:0] p73_array_index_1090385_comb;
  wire [7:0] p73_array_index_1090386_comb;
  wire [7:0] p73_array_index_1090387_comb;
  wire [7:0] p73_array_index_1090388_comb;
  wire [7:0] p73_array_index_1090468_comb;
  wire [7:0] p73_array_index_1090469_comb;
  wire [7:0] p73_array_index_1090470_comb;
  wire [7:0] p73_array_index_1090471_comb;
  wire [7:0] p73_array_index_1090472_comb;
  wire [7:0] p73_array_index_1090473_comb;
  wire [7:0] p73_res7__385_comb;
  wire [7:0] p73_res7__609_comb;
  wire [7:0] p73_array_index_1090398_comb;
  wire [7:0] p73_array_index_1090399_comb;
  wire [7:0] p73_array_index_1090400_comb;
  wire [7:0] p73_array_index_1090401_comb;
  wire [7:0] p73_array_index_1090402_comb;
  wire [7:0] p73_array_index_1090483_comb;
  wire [7:0] p73_array_index_1090484_comb;
  wire [7:0] p73_array_index_1090485_comb;
  wire [7:0] p73_array_index_1090486_comb;
  wire [7:0] p73_array_index_1090487_comb;
  wire [7:0] p73_res7__386_comb;
  wire [7:0] p73_res7__610_comb;
  wire [7:0] p73_array_index_1090412_comb;
  wire [7:0] p73_array_index_1090413_comb;
  wire [7:0] p73_array_index_1090414_comb;
  wire [7:0] p73_array_index_1090415_comb;
  wire [7:0] p73_array_index_1090416_comb;
  wire [7:0] p73_array_index_1090497_comb;
  wire [7:0] p73_array_index_1090498_comb;
  wire [7:0] p73_array_index_1090499_comb;
  wire [7:0] p73_array_index_1090500_comb;
  wire [7:0] p73_array_index_1090501_comb;
  wire [7:0] p73_res7__387_comb;
  wire [7:0] p73_res7__611_comb;
  wire [7:0] p73_array_index_1090427_comb;
  wire [7:0] p73_array_index_1090428_comb;
  wire [7:0] p73_array_index_1090429_comb;
  wire [7:0] p73_array_index_1090430_comb;
  wire [7:0] p73_array_index_1090512_comb;
  wire [7:0] p73_array_index_1090513_comb;
  wire [7:0] p73_array_index_1090514_comb;
  wire [7:0] p73_array_index_1090515_comb;
  wire [7:0] p73_res7__388_comb;
  wire [7:0] p73_res7__612_comb;
  assign p73_addedKey__65_comb = p72_k6 ^ 128'hb749_2c48_8547_80e0_69e9_9d53_b4b9_ea19;
  assign p73_array_index_1090350_comb = p72_arr[p73_addedKey__65_comb[127:120]];
  assign p73_array_index_1090351_comb = p72_arr[p73_addedKey__65_comb[119:112]];
  assign p73_array_index_1090352_comb = p72_arr[p73_addedKey__65_comb[111:104]];
  assign p73_array_index_1090353_comb = p72_arr[p73_addedKey__65_comb[103:96]];
  assign p73_array_index_1090354_comb = p72_arr[p73_addedKey__65_comb[95:88]];
  assign p73_array_index_1090355_comb = p72_arr[p73_addedKey__65_comb[87:80]];
  assign p73_array_index_1090357_comb = p72_arr[p73_addedKey__65_comb[71:64]];
  assign p73_array_index_1090359_comb = p72_arr[p73_addedKey__65_comb[55:48]];
  assign p73_array_index_1090360_comb = p72_arr[p73_addedKey__65_comb[47:40]];
  assign p73_array_index_1090361_comb = p72_arr[p73_addedKey__65_comb[39:32]];
  assign p73_array_index_1090362_comb = p72_arr[p73_addedKey__65_comb[31:24]];
  assign p73_array_index_1090363_comb = p72_arr[p73_addedKey__65_comb[23:16]];
  assign p73_array_index_1090364_comb = p72_arr[p73_addedKey__65_comb[15:8]];
  assign p73_array_index_1090438_comb = p72_arr[p72_bit_slice_1090267];
  assign p73_array_index_1090439_comb = p72_arr[p72_bit_slice_1090268];
  assign p73_array_index_1090440_comb = p72_arr[p72_bit_slice_1090269];
  assign p73_array_index_1090441_comb = p72_arr[p72_bit_slice_1090270];
  assign p73_array_index_1090442_comb = p72_arr[p72_bit_slice_1090271];
  assign p73_array_index_1090443_comb = p72_arr[p72_bit_slice_1090272];
  assign p73_array_index_1090444_comb = p72_arr[p72_bit_slice_1090273];
  assign p73_array_index_1090445_comb = p72_arr[p72_bit_slice_1090274];
  assign p73_array_index_1090446_comb = p72_arr[p72_bit_slice_1090275];
  assign p73_array_index_1090447_comb = p72_arr[p72_bit_slice_1090276];
  assign p73_array_index_1090448_comb = p72_arr[p72_bit_slice_1090277];
  assign p73_array_index_1090449_comb = p72_arr[p72_bit_slice_1090278];
  assign p73_array_index_1090450_comb = p72_arr[p72_bit_slice_1090279];
  assign p73_array_index_1090366_comb = p72_literal_1076345[p73_array_index_1090350_comb];
  assign p73_array_index_1090367_comb = p72_literal_1076347[p73_array_index_1090351_comb];
  assign p73_array_index_1090368_comb = p72_literal_1076349[p73_array_index_1090352_comb];
  assign p73_array_index_1090369_comb = p72_literal_1076351[p73_array_index_1090353_comb];
  assign p73_array_index_1090370_comb = p72_literal_1076353[p73_array_index_1090354_comb];
  assign p73_array_index_1090371_comb = p72_literal_1076355[p73_array_index_1090355_comb];
  assign p73_array_index_1090372_comb = p72_arr[p73_addedKey__65_comb[79:72]];
  assign p73_array_index_1090374_comb = p72_arr[p73_addedKey__65_comb[63:56]];
  assign p73_array_index_1090451_comb = p72_literal_1076345[p73_array_index_1090438_comb];
  assign p73_array_index_1090452_comb = p72_literal_1076347[p73_array_index_1090439_comb];
  assign p73_array_index_1090453_comb = p72_literal_1076349[p73_array_index_1090440_comb];
  assign p73_array_index_1090454_comb = p72_literal_1076351[p73_array_index_1090441_comb];
  assign p73_array_index_1090455_comb = p72_literal_1076353[p73_array_index_1090442_comb];
  assign p73_array_index_1090456_comb = p72_literal_1076355[p73_array_index_1090443_comb];
  assign p73_array_index_1090457_comb = p72_arr[p72_bit_slice_1090280];
  assign p73_array_index_1090459_comb = p72_arr[p72_bit_slice_1090281];
  assign p73_res7__384_comb = p73_array_index_1090366_comb ^ p73_array_index_1090367_comb ^ p73_array_index_1090368_comb ^ p73_array_index_1090369_comb ^ p73_array_index_1090370_comb ^ p73_array_index_1090371_comb ^ p73_array_index_1090372_comb ^ p72_literal_1076358[p73_array_index_1090357_comb] ^ p73_array_index_1090374_comb ^ p72_literal_1076355[p73_array_index_1090359_comb] ^ p72_literal_1076353[p73_array_index_1090360_comb] ^ p72_literal_1076351[p73_array_index_1090361_comb] ^ p72_literal_1076349[p73_array_index_1090362_comb] ^ p72_literal_1076347[p73_array_index_1090363_comb] ^ p72_literal_1076345[p73_array_index_1090364_comb] ^ p72_arr[p73_addedKey__65_comb[7:0]];
  assign p73_res7__608_comb = p73_array_index_1090451_comb ^ p73_array_index_1090452_comb ^ p73_array_index_1090453_comb ^ p73_array_index_1090454_comb ^ p73_array_index_1090455_comb ^ p73_array_index_1090456_comb ^ p73_array_index_1090457_comb ^ p72_literal_1076358[p73_array_index_1090444_comb] ^ p73_array_index_1090459_comb ^ p72_literal_1076355[p73_array_index_1090445_comb] ^ p72_literal_1076353[p73_array_index_1090446_comb] ^ p72_literal_1076351[p73_array_index_1090447_comb] ^ p72_literal_1076349[p73_array_index_1090448_comb] ^ p72_literal_1076347[p73_array_index_1090449_comb] ^ p72_literal_1076345[p73_array_index_1090450_comb] ^ p72_arr[p72_bit_slice_1090282];
  assign p73_array_index_1090383_comb = p72_literal_1076345[p73_res7__384_comb];
  assign p73_array_index_1090384_comb = p72_literal_1076347[p73_array_index_1090350_comb];
  assign p73_array_index_1090385_comb = p72_literal_1076349[p73_array_index_1090351_comb];
  assign p73_array_index_1090386_comb = p72_literal_1076351[p73_array_index_1090352_comb];
  assign p73_array_index_1090387_comb = p72_literal_1076353[p73_array_index_1090353_comb];
  assign p73_array_index_1090388_comb = p72_literal_1076355[p73_array_index_1090354_comb];
  assign p73_array_index_1090468_comb = p72_literal_1076345[p73_res7__608_comb];
  assign p73_array_index_1090469_comb = p72_literal_1076347[p73_array_index_1090438_comb];
  assign p73_array_index_1090470_comb = p72_literal_1076349[p73_array_index_1090439_comb];
  assign p73_array_index_1090471_comb = p72_literal_1076351[p73_array_index_1090440_comb];
  assign p73_array_index_1090472_comb = p72_literal_1076353[p73_array_index_1090441_comb];
  assign p73_array_index_1090473_comb = p72_literal_1076355[p73_array_index_1090442_comb];
  assign p73_res7__385_comb = p73_array_index_1090383_comb ^ p73_array_index_1090384_comb ^ p73_array_index_1090385_comb ^ p73_array_index_1090386_comb ^ p73_array_index_1090387_comb ^ p73_array_index_1090388_comb ^ p73_array_index_1090355_comb ^ p72_literal_1076358[p73_array_index_1090372_comb] ^ p73_array_index_1090357_comb ^ p72_literal_1076355[p73_array_index_1090374_comb] ^ p72_literal_1076353[p73_array_index_1090359_comb] ^ p72_literal_1076351[p73_array_index_1090360_comb] ^ p72_literal_1076349[p73_array_index_1090361_comb] ^ p72_literal_1076347[p73_array_index_1090362_comb] ^ p72_literal_1076345[p73_array_index_1090363_comb] ^ p73_array_index_1090364_comb;
  assign p73_res7__609_comb = p73_array_index_1090468_comb ^ p73_array_index_1090469_comb ^ p73_array_index_1090470_comb ^ p73_array_index_1090471_comb ^ p73_array_index_1090472_comb ^ p73_array_index_1090473_comb ^ p73_array_index_1090443_comb ^ p72_literal_1076358[p73_array_index_1090457_comb] ^ p73_array_index_1090444_comb ^ p72_literal_1076355[p73_array_index_1090459_comb] ^ p72_literal_1076353[p73_array_index_1090445_comb] ^ p72_literal_1076351[p73_array_index_1090446_comb] ^ p72_literal_1076349[p73_array_index_1090447_comb] ^ p72_literal_1076347[p73_array_index_1090448_comb] ^ p72_literal_1076345[p73_array_index_1090449_comb] ^ p73_array_index_1090450_comb;
  assign p73_array_index_1090398_comb = p72_literal_1076347[p73_res7__384_comb];
  assign p73_array_index_1090399_comb = p72_literal_1076349[p73_array_index_1090350_comb];
  assign p73_array_index_1090400_comb = p72_literal_1076351[p73_array_index_1090351_comb];
  assign p73_array_index_1090401_comb = p72_literal_1076353[p73_array_index_1090352_comb];
  assign p73_array_index_1090402_comb = p72_literal_1076355[p73_array_index_1090353_comb];
  assign p73_array_index_1090483_comb = p72_literal_1076347[p73_res7__608_comb];
  assign p73_array_index_1090484_comb = p72_literal_1076349[p73_array_index_1090438_comb];
  assign p73_array_index_1090485_comb = p72_literal_1076351[p73_array_index_1090439_comb];
  assign p73_array_index_1090486_comb = p72_literal_1076353[p73_array_index_1090440_comb];
  assign p73_array_index_1090487_comb = p72_literal_1076355[p73_array_index_1090441_comb];
  assign p73_res7__386_comb = p72_literal_1076345[p73_res7__385_comb] ^ p73_array_index_1090398_comb ^ p73_array_index_1090399_comb ^ p73_array_index_1090400_comb ^ p73_array_index_1090401_comb ^ p73_array_index_1090402_comb ^ p73_array_index_1090354_comb ^ p72_literal_1076358[p73_array_index_1090355_comb] ^ p73_array_index_1090372_comb ^ p72_literal_1076355[p73_array_index_1090357_comb] ^ p72_literal_1076353[p73_array_index_1090374_comb] ^ p72_literal_1076351[p73_array_index_1090359_comb] ^ p72_literal_1076349[p73_array_index_1090360_comb] ^ p72_literal_1076347[p73_array_index_1090361_comb] ^ p72_literal_1076345[p73_array_index_1090362_comb] ^ p73_array_index_1090363_comb;
  assign p73_res7__610_comb = p72_literal_1076345[p73_res7__609_comb] ^ p73_array_index_1090483_comb ^ p73_array_index_1090484_comb ^ p73_array_index_1090485_comb ^ p73_array_index_1090486_comb ^ p73_array_index_1090487_comb ^ p73_array_index_1090442_comb ^ p72_literal_1076358[p73_array_index_1090443_comb] ^ p73_array_index_1090457_comb ^ p72_literal_1076355[p73_array_index_1090444_comb] ^ p72_literal_1076353[p73_array_index_1090459_comb] ^ p72_literal_1076351[p73_array_index_1090445_comb] ^ p72_literal_1076349[p73_array_index_1090446_comb] ^ p72_literal_1076347[p73_array_index_1090447_comb] ^ p72_literal_1076345[p73_array_index_1090448_comb] ^ p73_array_index_1090449_comb;
  assign p73_array_index_1090412_comb = p72_literal_1076347[p73_res7__385_comb];
  assign p73_array_index_1090413_comb = p72_literal_1076349[p73_res7__384_comb];
  assign p73_array_index_1090414_comb = p72_literal_1076351[p73_array_index_1090350_comb];
  assign p73_array_index_1090415_comb = p72_literal_1076353[p73_array_index_1090351_comb];
  assign p73_array_index_1090416_comb = p72_literal_1076355[p73_array_index_1090352_comb];
  assign p73_array_index_1090497_comb = p72_literal_1076347[p73_res7__609_comb];
  assign p73_array_index_1090498_comb = p72_literal_1076349[p73_res7__608_comb];
  assign p73_array_index_1090499_comb = p72_literal_1076351[p73_array_index_1090438_comb];
  assign p73_array_index_1090500_comb = p72_literal_1076353[p73_array_index_1090439_comb];
  assign p73_array_index_1090501_comb = p72_literal_1076355[p73_array_index_1090440_comb];
  assign p73_res7__387_comb = p72_literal_1076345[p73_res7__386_comb] ^ p73_array_index_1090412_comb ^ p73_array_index_1090413_comb ^ p73_array_index_1090414_comb ^ p73_array_index_1090415_comb ^ p73_array_index_1090416_comb ^ p73_array_index_1090353_comb ^ p72_literal_1076358[p73_array_index_1090354_comb] ^ p73_array_index_1090355_comb ^ p72_literal_1076355[p73_array_index_1090372_comb] ^ p72_literal_1076353[p73_array_index_1090357_comb] ^ p72_literal_1076351[p73_array_index_1090374_comb] ^ p72_literal_1076349[p73_array_index_1090359_comb] ^ p72_literal_1076347[p73_array_index_1090360_comb] ^ p72_literal_1076345[p73_array_index_1090361_comb] ^ p73_array_index_1090362_comb;
  assign p73_res7__611_comb = p72_literal_1076345[p73_res7__610_comb] ^ p73_array_index_1090497_comb ^ p73_array_index_1090498_comb ^ p73_array_index_1090499_comb ^ p73_array_index_1090500_comb ^ p73_array_index_1090501_comb ^ p73_array_index_1090441_comb ^ p72_literal_1076358[p73_array_index_1090442_comb] ^ p73_array_index_1090443_comb ^ p72_literal_1076355[p73_array_index_1090457_comb] ^ p72_literal_1076353[p73_array_index_1090444_comb] ^ p72_literal_1076351[p73_array_index_1090459_comb] ^ p72_literal_1076349[p73_array_index_1090445_comb] ^ p72_literal_1076347[p73_array_index_1090446_comb] ^ p72_literal_1076345[p73_array_index_1090447_comb] ^ p73_array_index_1090448_comb;
  assign p73_array_index_1090427_comb = p72_literal_1076349[p73_res7__385_comb];
  assign p73_array_index_1090428_comb = p72_literal_1076351[p73_res7__384_comb];
  assign p73_array_index_1090429_comb = p72_literal_1076353[p73_array_index_1090350_comb];
  assign p73_array_index_1090430_comb = p72_literal_1076355[p73_array_index_1090351_comb];
  assign p73_array_index_1090512_comb = p72_literal_1076349[p73_res7__609_comb];
  assign p73_array_index_1090513_comb = p72_literal_1076351[p73_res7__608_comb];
  assign p73_array_index_1090514_comb = p72_literal_1076353[p73_array_index_1090438_comb];
  assign p73_array_index_1090515_comb = p72_literal_1076355[p73_array_index_1090439_comb];
  assign p73_res7__388_comb = p72_literal_1076345[p73_res7__387_comb] ^ p72_literal_1076347[p73_res7__386_comb] ^ p73_array_index_1090427_comb ^ p73_array_index_1090428_comb ^ p73_array_index_1090429_comb ^ p73_array_index_1090430_comb ^ p73_array_index_1090352_comb ^ p72_literal_1076358[p73_array_index_1090353_comb] ^ p73_array_index_1090354_comb ^ p73_array_index_1090371_comb ^ p72_literal_1076353[p73_array_index_1090372_comb] ^ p72_literal_1076351[p73_array_index_1090357_comb] ^ p72_literal_1076349[p73_array_index_1090374_comb] ^ p72_literal_1076347[p73_array_index_1090359_comb] ^ p72_literal_1076345[p73_array_index_1090360_comb] ^ p73_array_index_1090361_comb;
  assign p73_res7__612_comb = p72_literal_1076345[p73_res7__611_comb] ^ p72_literal_1076347[p73_res7__610_comb] ^ p73_array_index_1090512_comb ^ p73_array_index_1090513_comb ^ p73_array_index_1090514_comb ^ p73_array_index_1090515_comb ^ p73_array_index_1090440_comb ^ p72_literal_1076358[p73_array_index_1090441_comb] ^ p73_array_index_1090442_comb ^ p73_array_index_1090456_comb ^ p72_literal_1076353[p73_array_index_1090457_comb] ^ p72_literal_1076351[p73_array_index_1090444_comb] ^ p72_literal_1076349[p73_array_index_1090459_comb] ^ p72_literal_1076347[p73_array_index_1090445_comb] ^ p72_literal_1076345[p73_array_index_1090446_comb] ^ p73_array_index_1090447_comb;

  // Registers for pipe stage 73:
  reg [127:0] p73_k7;
  reg [127:0] p73_k6;
  reg [7:0] p73_array_index_1090350;
  reg [7:0] p73_array_index_1090351;
  reg [7:0] p73_array_index_1090352;
  reg [7:0] p73_array_index_1090353;
  reg [7:0] p73_array_index_1090354;
  reg [7:0] p73_array_index_1090355;
  reg [7:0] p73_array_index_1090357;
  reg [7:0] p73_array_index_1090359;
  reg [7:0] p73_array_index_1090360;
  reg [7:0] p73_array_index_1090366;
  reg [7:0] p73_array_index_1090367;
  reg [7:0] p73_array_index_1090368;
  reg [7:0] p73_array_index_1090369;
  reg [7:0] p73_array_index_1090370;
  reg [7:0] p73_array_index_1090372;
  reg [7:0] p73_array_index_1090374;
  reg [7:0] p73_res7__384;
  reg [7:0] p73_array_index_1090383;
  reg [7:0] p73_array_index_1090384;
  reg [7:0] p73_array_index_1090385;
  reg [7:0] p73_array_index_1090386;
  reg [7:0] p73_array_index_1090387;
  reg [7:0] p73_array_index_1090388;
  reg [7:0] p73_res7__385;
  reg [7:0] p73_array_index_1090398;
  reg [7:0] p73_array_index_1090399;
  reg [7:0] p73_array_index_1090400;
  reg [7:0] p73_array_index_1090401;
  reg [7:0] p73_array_index_1090402;
  reg [7:0] p73_res7__386;
  reg [7:0] p73_array_index_1090412;
  reg [7:0] p73_array_index_1090413;
  reg [7:0] p73_array_index_1090414;
  reg [7:0] p73_array_index_1090415;
  reg [7:0] p73_array_index_1090416;
  reg [7:0] p73_res7__387;
  reg [7:0] p73_array_index_1090427;
  reg [7:0] p73_array_index_1090428;
  reg [7:0] p73_array_index_1090429;
  reg [7:0] p73_array_index_1090430;
  reg [7:0] p73_res7__388;
  reg [7:0] p73_array_index_1090438;
  reg [7:0] p73_array_index_1090439;
  reg [7:0] p73_array_index_1090440;
  reg [7:0] p73_array_index_1090441;
  reg [7:0] p73_array_index_1090442;
  reg [7:0] p73_array_index_1090443;
  reg [7:0] p73_array_index_1090444;
  reg [7:0] p73_array_index_1090445;
  reg [7:0] p73_array_index_1090446;
  reg [7:0] p73_array_index_1090451;
  reg [7:0] p73_array_index_1090452;
  reg [7:0] p73_array_index_1090453;
  reg [7:0] p73_array_index_1090454;
  reg [7:0] p73_array_index_1090455;
  reg [7:0] p73_array_index_1090457;
  reg [7:0] p73_array_index_1090459;
  reg [7:0] p73_res7__608;
  reg [7:0] p73_array_index_1090468;
  reg [7:0] p73_array_index_1090469;
  reg [7:0] p73_array_index_1090470;
  reg [7:0] p73_array_index_1090471;
  reg [7:0] p73_array_index_1090472;
  reg [7:0] p73_array_index_1090473;
  reg [7:0] p73_res7__609;
  reg [7:0] p73_array_index_1090483;
  reg [7:0] p73_array_index_1090484;
  reg [7:0] p73_array_index_1090485;
  reg [7:0] p73_array_index_1090486;
  reg [7:0] p73_array_index_1090487;
  reg [7:0] p73_res7__610;
  reg [7:0] p73_array_index_1090497;
  reg [7:0] p73_array_index_1090498;
  reg [7:0] p73_array_index_1090499;
  reg [7:0] p73_array_index_1090500;
  reg [7:0] p73_array_index_1090501;
  reg [7:0] p73_res7__611;
  reg [7:0] p73_array_index_1090512;
  reg [7:0] p73_array_index_1090513;
  reg [7:0] p73_array_index_1090514;
  reg [7:0] p73_array_index_1090515;
  reg [7:0] p73_res7__612;
  reg [7:0] p74_arr[256];
  reg [7:0] p74_literal_1076345[256];
  reg [7:0] p74_literal_1076347[256];
  reg [7:0] p74_literal_1076349[256];
  reg [7:0] p74_literal_1076351[256];
  reg [7:0] p74_literal_1076353[256];
  reg [7:0] p74_literal_1076355[256];
  reg [7:0] p74_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p73_k7 <= p72_k7;
    p73_k6 <= p72_k6;
    p73_array_index_1090350 <= p73_array_index_1090350_comb;
    p73_array_index_1090351 <= p73_array_index_1090351_comb;
    p73_array_index_1090352 <= p73_array_index_1090352_comb;
    p73_array_index_1090353 <= p73_array_index_1090353_comb;
    p73_array_index_1090354 <= p73_array_index_1090354_comb;
    p73_array_index_1090355 <= p73_array_index_1090355_comb;
    p73_array_index_1090357 <= p73_array_index_1090357_comb;
    p73_array_index_1090359 <= p73_array_index_1090359_comb;
    p73_array_index_1090360 <= p73_array_index_1090360_comb;
    p73_array_index_1090366 <= p73_array_index_1090366_comb;
    p73_array_index_1090367 <= p73_array_index_1090367_comb;
    p73_array_index_1090368 <= p73_array_index_1090368_comb;
    p73_array_index_1090369 <= p73_array_index_1090369_comb;
    p73_array_index_1090370 <= p73_array_index_1090370_comb;
    p73_array_index_1090372 <= p73_array_index_1090372_comb;
    p73_array_index_1090374 <= p73_array_index_1090374_comb;
    p73_res7__384 <= p73_res7__384_comb;
    p73_array_index_1090383 <= p73_array_index_1090383_comb;
    p73_array_index_1090384 <= p73_array_index_1090384_comb;
    p73_array_index_1090385 <= p73_array_index_1090385_comb;
    p73_array_index_1090386 <= p73_array_index_1090386_comb;
    p73_array_index_1090387 <= p73_array_index_1090387_comb;
    p73_array_index_1090388 <= p73_array_index_1090388_comb;
    p73_res7__385 <= p73_res7__385_comb;
    p73_array_index_1090398 <= p73_array_index_1090398_comb;
    p73_array_index_1090399 <= p73_array_index_1090399_comb;
    p73_array_index_1090400 <= p73_array_index_1090400_comb;
    p73_array_index_1090401 <= p73_array_index_1090401_comb;
    p73_array_index_1090402 <= p73_array_index_1090402_comb;
    p73_res7__386 <= p73_res7__386_comb;
    p73_array_index_1090412 <= p73_array_index_1090412_comb;
    p73_array_index_1090413 <= p73_array_index_1090413_comb;
    p73_array_index_1090414 <= p73_array_index_1090414_comb;
    p73_array_index_1090415 <= p73_array_index_1090415_comb;
    p73_array_index_1090416 <= p73_array_index_1090416_comb;
    p73_res7__387 <= p73_res7__387_comb;
    p73_array_index_1090427 <= p73_array_index_1090427_comb;
    p73_array_index_1090428 <= p73_array_index_1090428_comb;
    p73_array_index_1090429 <= p73_array_index_1090429_comb;
    p73_array_index_1090430 <= p73_array_index_1090430_comb;
    p73_res7__388 <= p73_res7__388_comb;
    p73_array_index_1090438 <= p73_array_index_1090438_comb;
    p73_array_index_1090439 <= p73_array_index_1090439_comb;
    p73_array_index_1090440 <= p73_array_index_1090440_comb;
    p73_array_index_1090441 <= p73_array_index_1090441_comb;
    p73_array_index_1090442 <= p73_array_index_1090442_comb;
    p73_array_index_1090443 <= p73_array_index_1090443_comb;
    p73_array_index_1090444 <= p73_array_index_1090444_comb;
    p73_array_index_1090445 <= p73_array_index_1090445_comb;
    p73_array_index_1090446 <= p73_array_index_1090446_comb;
    p73_array_index_1090451 <= p73_array_index_1090451_comb;
    p73_array_index_1090452 <= p73_array_index_1090452_comb;
    p73_array_index_1090453 <= p73_array_index_1090453_comb;
    p73_array_index_1090454 <= p73_array_index_1090454_comb;
    p73_array_index_1090455 <= p73_array_index_1090455_comb;
    p73_array_index_1090457 <= p73_array_index_1090457_comb;
    p73_array_index_1090459 <= p73_array_index_1090459_comb;
    p73_res7__608 <= p73_res7__608_comb;
    p73_array_index_1090468 <= p73_array_index_1090468_comb;
    p73_array_index_1090469 <= p73_array_index_1090469_comb;
    p73_array_index_1090470 <= p73_array_index_1090470_comb;
    p73_array_index_1090471 <= p73_array_index_1090471_comb;
    p73_array_index_1090472 <= p73_array_index_1090472_comb;
    p73_array_index_1090473 <= p73_array_index_1090473_comb;
    p73_res7__609 <= p73_res7__609_comb;
    p73_array_index_1090483 <= p73_array_index_1090483_comb;
    p73_array_index_1090484 <= p73_array_index_1090484_comb;
    p73_array_index_1090485 <= p73_array_index_1090485_comb;
    p73_array_index_1090486 <= p73_array_index_1090486_comb;
    p73_array_index_1090487 <= p73_array_index_1090487_comb;
    p73_res7__610 <= p73_res7__610_comb;
    p73_array_index_1090497 <= p73_array_index_1090497_comb;
    p73_array_index_1090498 <= p73_array_index_1090498_comb;
    p73_array_index_1090499 <= p73_array_index_1090499_comb;
    p73_array_index_1090500 <= p73_array_index_1090500_comb;
    p73_array_index_1090501 <= p73_array_index_1090501_comb;
    p73_res7__611 <= p73_res7__611_comb;
    p73_array_index_1090512 <= p73_array_index_1090512_comb;
    p73_array_index_1090513 <= p73_array_index_1090513_comb;
    p73_array_index_1090514 <= p73_array_index_1090514_comb;
    p73_array_index_1090515 <= p73_array_index_1090515_comb;
    p73_res7__612 <= p73_res7__612_comb;
    p74_arr <= p73_arr;
    p74_literal_1076345 <= p73_literal_1076345;
    p74_literal_1076347 <= p73_literal_1076347;
    p74_literal_1076349 <= p73_literal_1076349;
    p74_literal_1076351 <= p73_literal_1076351;
    p74_literal_1076353 <= p73_literal_1076353;
    p74_literal_1076355 <= p73_literal_1076355;
    p74_literal_1076358 <= p73_literal_1076358;
  end

  // ===== Pipe stage 74:
  wire [7:0] p74_array_index_1090709_comb;
  wire [7:0] p74_array_index_1090710_comb;
  wire [7:0] p74_array_index_1090711_comb;
  wire [7:0] p74_array_index_1090712_comb;
  wire [7:0] p74_array_index_1090777_comb;
  wire [7:0] p74_array_index_1090778_comb;
  wire [7:0] p74_array_index_1090779_comb;
  wire [7:0] p74_array_index_1090780_comb;
  wire [7:0] p74_res7__389_comb;
  wire [7:0] p74_res7__613_comb;
  wire [7:0] p74_array_index_1090723_comb;
  wire [7:0] p74_array_index_1090724_comb;
  wire [7:0] p74_array_index_1090725_comb;
  wire [7:0] p74_array_index_1090791_comb;
  wire [7:0] p74_array_index_1090792_comb;
  wire [7:0] p74_array_index_1090793_comb;
  wire [7:0] p74_res7__390_comb;
  wire [7:0] p74_res7__614_comb;
  wire [7:0] p74_array_index_1090735_comb;
  wire [7:0] p74_array_index_1090736_comb;
  wire [7:0] p74_array_index_1090737_comb;
  wire [7:0] p74_array_index_1090803_comb;
  wire [7:0] p74_array_index_1090804_comb;
  wire [7:0] p74_array_index_1090805_comb;
  wire [7:0] p74_res7__391_comb;
  wire [7:0] p74_res7__615_comb;
  wire [7:0] p74_array_index_1090748_comb;
  wire [7:0] p74_array_index_1090749_comb;
  wire [7:0] p74_array_index_1090816_comb;
  wire [7:0] p74_array_index_1090817_comb;
  wire [7:0] p74_res7__392_comb;
  wire [7:0] p74_res7__616_comb;
  wire [7:0] p74_array_index_1090759_comb;
  wire [7:0] p74_array_index_1090760_comb;
  wire [7:0] p74_array_index_1090827_comb;
  wire [7:0] p74_array_index_1090828_comb;
  wire [7:0] p74_res7__393_comb;
  wire [7:0] p74_res7__617_comb;
  wire [7:0] p74_array_index_1090766_comb;
  wire [7:0] p74_array_index_1090767_comb;
  wire [7:0] p74_array_index_1090768_comb;
  wire [7:0] p74_array_index_1090769_comb;
  wire [7:0] p74_array_index_1090770_comb;
  wire [7:0] p74_array_index_1090771_comb;
  wire [7:0] p74_array_index_1090772_comb;
  wire [7:0] p74_array_index_1090773_comb;
  wire [7:0] p74_array_index_1090774_comb;
  wire [7:0] p74_array_index_1090834_comb;
  wire [7:0] p74_array_index_1090835_comb;
  wire [7:0] p74_array_index_1090836_comb;
  wire [7:0] p74_array_index_1090837_comb;
  wire [7:0] p74_array_index_1090838_comb;
  wire [7:0] p74_array_index_1090839_comb;
  wire [7:0] p74_array_index_1090840_comb;
  wire [7:0] p74_array_index_1090841_comb;
  wire [7:0] p74_array_index_1090842_comb;
  assign p74_array_index_1090709_comb = p73_literal_1076349[p73_res7__386];
  assign p74_array_index_1090710_comb = p73_literal_1076351[p73_res7__385];
  assign p74_array_index_1090711_comb = p73_literal_1076353[p73_res7__384];
  assign p74_array_index_1090712_comb = p73_literal_1076355[p73_array_index_1090350];
  assign p74_array_index_1090777_comb = p73_literal_1076349[p73_res7__610];
  assign p74_array_index_1090778_comb = p73_literal_1076351[p73_res7__609];
  assign p74_array_index_1090779_comb = p73_literal_1076353[p73_res7__608];
  assign p74_array_index_1090780_comb = p73_literal_1076355[p73_array_index_1090438];
  assign p74_res7__389_comb = p73_literal_1076345[p73_res7__388] ^ p73_literal_1076347[p73_res7__387] ^ p74_array_index_1090709_comb ^ p74_array_index_1090710_comb ^ p74_array_index_1090711_comb ^ p74_array_index_1090712_comb ^ p73_array_index_1090351 ^ p73_literal_1076358[p73_array_index_1090352] ^ p73_array_index_1090353 ^ p73_array_index_1090388 ^ p73_literal_1076353[p73_array_index_1090355] ^ p73_literal_1076351[p73_array_index_1090372] ^ p73_literal_1076349[p73_array_index_1090357] ^ p73_literal_1076347[p73_array_index_1090374] ^ p73_literal_1076345[p73_array_index_1090359] ^ p73_array_index_1090360;
  assign p74_res7__613_comb = p73_literal_1076345[p73_res7__612] ^ p73_literal_1076347[p73_res7__611] ^ p74_array_index_1090777_comb ^ p74_array_index_1090778_comb ^ p74_array_index_1090779_comb ^ p74_array_index_1090780_comb ^ p73_array_index_1090439 ^ p73_literal_1076358[p73_array_index_1090440] ^ p73_array_index_1090441 ^ p73_array_index_1090473 ^ p73_literal_1076353[p73_array_index_1090443] ^ p73_literal_1076351[p73_array_index_1090457] ^ p73_literal_1076349[p73_array_index_1090444] ^ p73_literal_1076347[p73_array_index_1090459] ^ p73_literal_1076345[p73_array_index_1090445] ^ p73_array_index_1090446;
  assign p74_array_index_1090723_comb = p73_literal_1076351[p73_res7__386];
  assign p74_array_index_1090724_comb = p73_literal_1076353[p73_res7__385];
  assign p74_array_index_1090725_comb = p73_literal_1076355[p73_res7__384];
  assign p74_array_index_1090791_comb = p73_literal_1076351[p73_res7__610];
  assign p74_array_index_1090792_comb = p73_literal_1076353[p73_res7__609];
  assign p74_array_index_1090793_comb = p73_literal_1076355[p73_res7__608];
  assign p74_res7__390_comb = p73_literal_1076345[p74_res7__389_comb] ^ p73_literal_1076347[p73_res7__388] ^ p73_literal_1076349[p73_res7__387] ^ p74_array_index_1090723_comb ^ p74_array_index_1090724_comb ^ p74_array_index_1090725_comb ^ p73_array_index_1090350 ^ p73_literal_1076358[p73_array_index_1090351] ^ p73_array_index_1090352 ^ p73_array_index_1090402 ^ p73_array_index_1090370 ^ p73_literal_1076351[p73_array_index_1090355] ^ p73_literal_1076349[p73_array_index_1090372] ^ p73_literal_1076347[p73_array_index_1090357] ^ p73_literal_1076345[p73_array_index_1090374] ^ p73_array_index_1090359;
  assign p74_res7__614_comb = p73_literal_1076345[p74_res7__613_comb] ^ p73_literal_1076347[p73_res7__612] ^ p73_literal_1076349[p73_res7__611] ^ p74_array_index_1090791_comb ^ p74_array_index_1090792_comb ^ p74_array_index_1090793_comb ^ p73_array_index_1090438 ^ p73_literal_1076358[p73_array_index_1090439] ^ p73_array_index_1090440 ^ p73_array_index_1090487 ^ p73_array_index_1090455 ^ p73_literal_1076351[p73_array_index_1090443] ^ p73_literal_1076349[p73_array_index_1090457] ^ p73_literal_1076347[p73_array_index_1090444] ^ p73_literal_1076345[p73_array_index_1090459] ^ p73_array_index_1090445;
  assign p74_array_index_1090735_comb = p73_literal_1076351[p73_res7__387];
  assign p74_array_index_1090736_comb = p73_literal_1076353[p73_res7__386];
  assign p74_array_index_1090737_comb = p73_literal_1076355[p73_res7__385];
  assign p74_array_index_1090803_comb = p73_literal_1076351[p73_res7__611];
  assign p74_array_index_1090804_comb = p73_literal_1076353[p73_res7__610];
  assign p74_array_index_1090805_comb = p73_literal_1076355[p73_res7__609];
  assign p74_res7__391_comb = p73_literal_1076345[p74_res7__390_comb] ^ p73_literal_1076347[p74_res7__389_comb] ^ p73_literal_1076349[p73_res7__388] ^ p74_array_index_1090735_comb ^ p74_array_index_1090736_comb ^ p74_array_index_1090737_comb ^ p73_res7__384 ^ p73_literal_1076358[p73_array_index_1090350] ^ p73_array_index_1090351 ^ p73_array_index_1090416 ^ p73_array_index_1090387 ^ p73_literal_1076351[p73_array_index_1090354] ^ p73_literal_1076349[p73_array_index_1090355] ^ p73_literal_1076347[p73_array_index_1090372] ^ p73_literal_1076345[p73_array_index_1090357] ^ p73_array_index_1090374;
  assign p74_res7__615_comb = p73_literal_1076345[p74_res7__614_comb] ^ p73_literal_1076347[p74_res7__613_comb] ^ p73_literal_1076349[p73_res7__612] ^ p74_array_index_1090803_comb ^ p74_array_index_1090804_comb ^ p74_array_index_1090805_comb ^ p73_res7__608 ^ p73_literal_1076358[p73_array_index_1090438] ^ p73_array_index_1090439 ^ p73_array_index_1090501 ^ p73_array_index_1090472 ^ p73_literal_1076351[p73_array_index_1090442] ^ p73_literal_1076349[p73_array_index_1090443] ^ p73_literal_1076347[p73_array_index_1090457] ^ p73_literal_1076345[p73_array_index_1090444] ^ p73_array_index_1090459;
  assign p74_array_index_1090748_comb = p73_literal_1076353[p73_res7__387];
  assign p74_array_index_1090749_comb = p73_literal_1076355[p73_res7__386];
  assign p74_array_index_1090816_comb = p73_literal_1076353[p73_res7__611];
  assign p74_array_index_1090817_comb = p73_literal_1076355[p73_res7__610];
  assign p74_res7__392_comb = p73_literal_1076345[p74_res7__391_comb] ^ p73_literal_1076347[p74_res7__390_comb] ^ p73_literal_1076349[p74_res7__389_comb] ^ p73_literal_1076351[p73_res7__388] ^ p74_array_index_1090748_comb ^ p74_array_index_1090749_comb ^ p73_res7__385 ^ p73_literal_1076358[p73_res7__384] ^ p73_array_index_1090350 ^ p73_array_index_1090430 ^ p73_array_index_1090401 ^ p73_array_index_1090369 ^ p73_literal_1076349[p73_array_index_1090354] ^ p73_literal_1076347[p73_array_index_1090355] ^ p73_literal_1076345[p73_array_index_1090372] ^ p73_array_index_1090357;
  assign p74_res7__616_comb = p73_literal_1076345[p74_res7__615_comb] ^ p73_literal_1076347[p74_res7__614_comb] ^ p73_literal_1076349[p74_res7__613_comb] ^ p73_literal_1076351[p73_res7__612] ^ p74_array_index_1090816_comb ^ p74_array_index_1090817_comb ^ p73_res7__609 ^ p73_literal_1076358[p73_res7__608] ^ p73_array_index_1090438 ^ p73_array_index_1090515 ^ p73_array_index_1090486 ^ p73_array_index_1090454 ^ p73_literal_1076349[p73_array_index_1090442] ^ p73_literal_1076347[p73_array_index_1090443] ^ p73_literal_1076345[p73_array_index_1090457] ^ p73_array_index_1090444;
  assign p74_array_index_1090759_comb = p73_literal_1076353[p73_res7__388];
  assign p74_array_index_1090760_comb = p73_literal_1076355[p73_res7__387];
  assign p74_array_index_1090827_comb = p73_literal_1076353[p73_res7__612];
  assign p74_array_index_1090828_comb = p73_literal_1076355[p73_res7__611];
  assign p74_res7__393_comb = p73_literal_1076345[p74_res7__392_comb] ^ p73_literal_1076347[p74_res7__391_comb] ^ p73_literal_1076349[p74_res7__390_comb] ^ p73_literal_1076351[p74_res7__389_comb] ^ p74_array_index_1090759_comb ^ p74_array_index_1090760_comb ^ p73_res7__386 ^ p73_literal_1076358[p73_res7__385] ^ p73_res7__384 ^ p74_array_index_1090712_comb ^ p73_array_index_1090415 ^ p73_array_index_1090386 ^ p73_literal_1076349[p73_array_index_1090353] ^ p73_literal_1076347[p73_array_index_1090354] ^ p73_literal_1076345[p73_array_index_1090355] ^ p73_array_index_1090372;
  assign p74_res7__617_comb = p73_literal_1076345[p74_res7__616_comb] ^ p73_literal_1076347[p74_res7__615_comb] ^ p73_literal_1076349[p74_res7__614_comb] ^ p73_literal_1076351[p74_res7__613_comb] ^ p74_array_index_1090827_comb ^ p74_array_index_1090828_comb ^ p73_res7__610 ^ p73_literal_1076358[p73_res7__609] ^ p73_res7__608 ^ p74_array_index_1090780_comb ^ p73_array_index_1090500 ^ p73_array_index_1090471 ^ p73_literal_1076349[p73_array_index_1090441] ^ p73_literal_1076347[p73_array_index_1090442] ^ p73_literal_1076345[p73_array_index_1090443] ^ p73_array_index_1090457;
  assign p74_array_index_1090766_comb = p73_literal_1076345[p74_res7__393_comb];
  assign p74_array_index_1090767_comb = p73_literal_1076347[p74_res7__392_comb];
  assign p74_array_index_1090768_comb = p73_literal_1076349[p74_res7__391_comb];
  assign p74_array_index_1090769_comb = p73_literal_1076351[p74_res7__390_comb];
  assign p74_array_index_1090770_comb = p73_literal_1076353[p74_res7__389_comb];
  assign p74_array_index_1090771_comb = p73_literal_1076355[p73_res7__388];
  assign p74_array_index_1090772_comb = p73_literal_1076358[p73_res7__386];
  assign p74_array_index_1090773_comb = p73_literal_1076347[p73_array_index_1090353];
  assign p74_array_index_1090774_comb = p73_literal_1076345[p73_array_index_1090354];
  assign p74_array_index_1090834_comb = p73_literal_1076345[p74_res7__617_comb];
  assign p74_array_index_1090835_comb = p73_literal_1076347[p74_res7__616_comb];
  assign p74_array_index_1090836_comb = p73_literal_1076349[p74_res7__615_comb];
  assign p74_array_index_1090837_comb = p73_literal_1076351[p74_res7__614_comb];
  assign p74_array_index_1090838_comb = p73_literal_1076353[p74_res7__613_comb];
  assign p74_array_index_1090839_comb = p73_literal_1076355[p73_res7__612];
  assign p74_array_index_1090840_comb = p73_literal_1076358[p73_res7__610];
  assign p74_array_index_1090841_comb = p73_literal_1076347[p73_array_index_1090441];
  assign p74_array_index_1090842_comb = p73_literal_1076345[p73_array_index_1090442];

  // Registers for pipe stage 74:
  reg [127:0] p74_k7;
  reg [127:0] p74_k6;
  reg [7:0] p74_array_index_1090350;
  reg [7:0] p74_array_index_1090351;
  reg [7:0] p74_array_index_1090352;
  reg [7:0] p74_array_index_1090353;
  reg [7:0] p74_array_index_1090354;
  reg [7:0] p74_array_index_1090355;
  reg [7:0] p74_array_index_1090366;
  reg [7:0] p74_array_index_1090367;
  reg [7:0] p74_array_index_1090368;
  reg [7:0] p74_res7__384;
  reg [7:0] p74_array_index_1090383;
  reg [7:0] p74_array_index_1090384;
  reg [7:0] p74_array_index_1090385;
  reg [7:0] p74_res7__385;
  reg [7:0] p74_array_index_1090398;
  reg [7:0] p74_array_index_1090399;
  reg [7:0] p74_array_index_1090400;
  reg [7:0] p74_res7__386;
  reg [7:0] p74_array_index_1090412;
  reg [7:0] p74_array_index_1090413;
  reg [7:0] p74_array_index_1090414;
  reg [7:0] p74_res7__387;
  reg [7:0] p74_array_index_1090427;
  reg [7:0] p74_array_index_1090428;
  reg [7:0] p74_array_index_1090429;
  reg [7:0] p74_res7__388;
  reg [7:0] p74_array_index_1090709;
  reg [7:0] p74_array_index_1090710;
  reg [7:0] p74_array_index_1090711;
  reg [7:0] p74_res7__389;
  reg [7:0] p74_array_index_1090723;
  reg [7:0] p74_array_index_1090724;
  reg [7:0] p74_array_index_1090725;
  reg [7:0] p74_res7__390;
  reg [7:0] p74_array_index_1090735;
  reg [7:0] p74_array_index_1090736;
  reg [7:0] p74_array_index_1090737;
  reg [7:0] p74_res7__391;
  reg [7:0] p74_array_index_1090748;
  reg [7:0] p74_array_index_1090749;
  reg [7:0] p74_res7__392;
  reg [7:0] p74_array_index_1090759;
  reg [7:0] p74_array_index_1090760;
  reg [7:0] p74_res7__393;
  reg [7:0] p74_array_index_1090766;
  reg [7:0] p74_array_index_1090767;
  reg [7:0] p74_array_index_1090768;
  reg [7:0] p74_array_index_1090769;
  reg [7:0] p74_array_index_1090770;
  reg [7:0] p74_array_index_1090771;
  reg [7:0] p74_array_index_1090772;
  reg [7:0] p74_array_index_1090773;
  reg [7:0] p74_array_index_1090774;
  reg [7:0] p74_array_index_1090438;
  reg [7:0] p74_array_index_1090439;
  reg [7:0] p74_array_index_1090440;
  reg [7:0] p74_array_index_1090441;
  reg [7:0] p74_array_index_1090442;
  reg [7:0] p74_array_index_1090443;
  reg [7:0] p74_array_index_1090451;
  reg [7:0] p74_array_index_1090452;
  reg [7:0] p74_array_index_1090453;
  reg [7:0] p74_res7__608;
  reg [7:0] p74_array_index_1090468;
  reg [7:0] p74_array_index_1090469;
  reg [7:0] p74_array_index_1090470;
  reg [7:0] p74_res7__609;
  reg [7:0] p74_array_index_1090483;
  reg [7:0] p74_array_index_1090484;
  reg [7:0] p74_array_index_1090485;
  reg [7:0] p74_res7__610;
  reg [7:0] p74_array_index_1090497;
  reg [7:0] p74_array_index_1090498;
  reg [7:0] p74_array_index_1090499;
  reg [7:0] p74_res7__611;
  reg [7:0] p74_array_index_1090512;
  reg [7:0] p74_array_index_1090513;
  reg [7:0] p74_array_index_1090514;
  reg [7:0] p74_res7__612;
  reg [7:0] p74_array_index_1090777;
  reg [7:0] p74_array_index_1090778;
  reg [7:0] p74_array_index_1090779;
  reg [7:0] p74_res7__613;
  reg [7:0] p74_array_index_1090791;
  reg [7:0] p74_array_index_1090792;
  reg [7:0] p74_array_index_1090793;
  reg [7:0] p74_res7__614;
  reg [7:0] p74_array_index_1090803;
  reg [7:0] p74_array_index_1090804;
  reg [7:0] p74_array_index_1090805;
  reg [7:0] p74_res7__615;
  reg [7:0] p74_array_index_1090816;
  reg [7:0] p74_array_index_1090817;
  reg [7:0] p74_res7__616;
  reg [7:0] p74_array_index_1090827;
  reg [7:0] p74_array_index_1090828;
  reg [7:0] p74_res7__617;
  reg [7:0] p74_array_index_1090834;
  reg [7:0] p74_array_index_1090835;
  reg [7:0] p74_array_index_1090836;
  reg [7:0] p74_array_index_1090837;
  reg [7:0] p74_array_index_1090838;
  reg [7:0] p74_array_index_1090839;
  reg [7:0] p74_array_index_1090840;
  reg [7:0] p74_array_index_1090841;
  reg [7:0] p74_array_index_1090842;
  reg [7:0] p75_arr[256];
  reg [7:0] p75_literal_1076345[256];
  reg [7:0] p75_literal_1076347[256];
  reg [7:0] p75_literal_1076349[256];
  reg [7:0] p75_literal_1076351[256];
  reg [7:0] p75_literal_1076353[256];
  reg [7:0] p75_literal_1076355[256];
  reg [7:0] p75_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p74_k7 <= p73_k7;
    p74_k6 <= p73_k6;
    p74_array_index_1090350 <= p73_array_index_1090350;
    p74_array_index_1090351 <= p73_array_index_1090351;
    p74_array_index_1090352 <= p73_array_index_1090352;
    p74_array_index_1090353 <= p73_array_index_1090353;
    p74_array_index_1090354 <= p73_array_index_1090354;
    p74_array_index_1090355 <= p73_array_index_1090355;
    p74_array_index_1090366 <= p73_array_index_1090366;
    p74_array_index_1090367 <= p73_array_index_1090367;
    p74_array_index_1090368 <= p73_array_index_1090368;
    p74_res7__384 <= p73_res7__384;
    p74_array_index_1090383 <= p73_array_index_1090383;
    p74_array_index_1090384 <= p73_array_index_1090384;
    p74_array_index_1090385 <= p73_array_index_1090385;
    p74_res7__385 <= p73_res7__385;
    p74_array_index_1090398 <= p73_array_index_1090398;
    p74_array_index_1090399 <= p73_array_index_1090399;
    p74_array_index_1090400 <= p73_array_index_1090400;
    p74_res7__386 <= p73_res7__386;
    p74_array_index_1090412 <= p73_array_index_1090412;
    p74_array_index_1090413 <= p73_array_index_1090413;
    p74_array_index_1090414 <= p73_array_index_1090414;
    p74_res7__387 <= p73_res7__387;
    p74_array_index_1090427 <= p73_array_index_1090427;
    p74_array_index_1090428 <= p73_array_index_1090428;
    p74_array_index_1090429 <= p73_array_index_1090429;
    p74_res7__388 <= p73_res7__388;
    p74_array_index_1090709 <= p74_array_index_1090709_comb;
    p74_array_index_1090710 <= p74_array_index_1090710_comb;
    p74_array_index_1090711 <= p74_array_index_1090711_comb;
    p74_res7__389 <= p74_res7__389_comb;
    p74_array_index_1090723 <= p74_array_index_1090723_comb;
    p74_array_index_1090724 <= p74_array_index_1090724_comb;
    p74_array_index_1090725 <= p74_array_index_1090725_comb;
    p74_res7__390 <= p74_res7__390_comb;
    p74_array_index_1090735 <= p74_array_index_1090735_comb;
    p74_array_index_1090736 <= p74_array_index_1090736_comb;
    p74_array_index_1090737 <= p74_array_index_1090737_comb;
    p74_res7__391 <= p74_res7__391_comb;
    p74_array_index_1090748 <= p74_array_index_1090748_comb;
    p74_array_index_1090749 <= p74_array_index_1090749_comb;
    p74_res7__392 <= p74_res7__392_comb;
    p74_array_index_1090759 <= p74_array_index_1090759_comb;
    p74_array_index_1090760 <= p74_array_index_1090760_comb;
    p74_res7__393 <= p74_res7__393_comb;
    p74_array_index_1090766 <= p74_array_index_1090766_comb;
    p74_array_index_1090767 <= p74_array_index_1090767_comb;
    p74_array_index_1090768 <= p74_array_index_1090768_comb;
    p74_array_index_1090769 <= p74_array_index_1090769_comb;
    p74_array_index_1090770 <= p74_array_index_1090770_comb;
    p74_array_index_1090771 <= p74_array_index_1090771_comb;
    p74_array_index_1090772 <= p74_array_index_1090772_comb;
    p74_array_index_1090773 <= p74_array_index_1090773_comb;
    p74_array_index_1090774 <= p74_array_index_1090774_comb;
    p74_array_index_1090438 <= p73_array_index_1090438;
    p74_array_index_1090439 <= p73_array_index_1090439;
    p74_array_index_1090440 <= p73_array_index_1090440;
    p74_array_index_1090441 <= p73_array_index_1090441;
    p74_array_index_1090442 <= p73_array_index_1090442;
    p74_array_index_1090443 <= p73_array_index_1090443;
    p74_array_index_1090451 <= p73_array_index_1090451;
    p74_array_index_1090452 <= p73_array_index_1090452;
    p74_array_index_1090453 <= p73_array_index_1090453;
    p74_res7__608 <= p73_res7__608;
    p74_array_index_1090468 <= p73_array_index_1090468;
    p74_array_index_1090469 <= p73_array_index_1090469;
    p74_array_index_1090470 <= p73_array_index_1090470;
    p74_res7__609 <= p73_res7__609;
    p74_array_index_1090483 <= p73_array_index_1090483;
    p74_array_index_1090484 <= p73_array_index_1090484;
    p74_array_index_1090485 <= p73_array_index_1090485;
    p74_res7__610 <= p73_res7__610;
    p74_array_index_1090497 <= p73_array_index_1090497;
    p74_array_index_1090498 <= p73_array_index_1090498;
    p74_array_index_1090499 <= p73_array_index_1090499;
    p74_res7__611 <= p73_res7__611;
    p74_array_index_1090512 <= p73_array_index_1090512;
    p74_array_index_1090513 <= p73_array_index_1090513;
    p74_array_index_1090514 <= p73_array_index_1090514;
    p74_res7__612 <= p73_res7__612;
    p74_array_index_1090777 <= p74_array_index_1090777_comb;
    p74_array_index_1090778 <= p74_array_index_1090778_comb;
    p74_array_index_1090779 <= p74_array_index_1090779_comb;
    p74_res7__613 <= p74_res7__613_comb;
    p74_array_index_1090791 <= p74_array_index_1090791_comb;
    p74_array_index_1090792 <= p74_array_index_1090792_comb;
    p74_array_index_1090793 <= p74_array_index_1090793_comb;
    p74_res7__614 <= p74_res7__614_comb;
    p74_array_index_1090803 <= p74_array_index_1090803_comb;
    p74_array_index_1090804 <= p74_array_index_1090804_comb;
    p74_array_index_1090805 <= p74_array_index_1090805_comb;
    p74_res7__615 <= p74_res7__615_comb;
    p74_array_index_1090816 <= p74_array_index_1090816_comb;
    p74_array_index_1090817 <= p74_array_index_1090817_comb;
    p74_res7__616 <= p74_res7__616_comb;
    p74_array_index_1090827 <= p74_array_index_1090827_comb;
    p74_array_index_1090828 <= p74_array_index_1090828_comb;
    p74_res7__617 <= p74_res7__617_comb;
    p74_array_index_1090834 <= p74_array_index_1090834_comb;
    p74_array_index_1090835 <= p74_array_index_1090835_comb;
    p74_array_index_1090836 <= p74_array_index_1090836_comb;
    p74_array_index_1090837 <= p74_array_index_1090837_comb;
    p74_array_index_1090838 <= p74_array_index_1090838_comb;
    p74_array_index_1090839 <= p74_array_index_1090839_comb;
    p74_array_index_1090840 <= p74_array_index_1090840_comb;
    p74_array_index_1090841 <= p74_array_index_1090841_comb;
    p74_array_index_1090842 <= p74_array_index_1090842_comb;
    p75_arr <= p74_arr;
    p75_literal_1076345 <= p74_literal_1076345;
    p75_literal_1076347 <= p74_literal_1076347;
    p75_literal_1076349 <= p74_literal_1076349;
    p75_literal_1076351 <= p74_literal_1076351;
    p75_literal_1076353 <= p74_literal_1076353;
    p75_literal_1076355 <= p74_literal_1076355;
    p75_literal_1076358 <= p74_literal_1076358;
  end

  // ===== Pipe stage 75:
  wire [7:0] p75_res7__618_comb;
  wire [7:0] p75_res7__394_comb;
  wire [7:0] p75_array_index_1091128_comb;
  wire [7:0] p75_array_index_1091081_comb;
  wire [7:0] p75_res7__619_comb;
  wire [7:0] p75_res7__395_comb;
  wire [7:0] p75_res7__620_comb;
  wire [7:0] p75_res7__396_comb;
  wire [7:0] p75_res7__621_comb;
  wire [7:0] p75_res7__397_comb;
  wire [7:0] p75_res7__622_comb;
  wire [7:0] p75_res7__398_comb;
  wire [7:0] p75_res7__623_comb;
  wire [7:0] p75_res7__399_comb;
  wire [127:0] p75_res__38_comb;
  wire [127:0] p75_res__24_comb;
  wire [127:0] p75_addedKey__39_comb;
  wire [127:0] p75_xor_1091121_comb;
  wire [7:0] p75_bit_slice_1091169_comb;
  wire [7:0] p75_bit_slice_1091170_comb;
  wire [7:0] p75_bit_slice_1091171_comb;
  wire [7:0] p75_bit_slice_1091172_comb;
  wire [7:0] p75_bit_slice_1091173_comb;
  wire [7:0] p75_bit_slice_1091174_comb;
  wire [7:0] p75_bit_slice_1091175_comb;
  wire [7:0] p75_bit_slice_1091176_comb;
  wire [7:0] p75_bit_slice_1091177_comb;
  wire [7:0] p75_bit_slice_1091178_comb;
  wire [7:0] p75_bit_slice_1091179_comb;
  wire [7:0] p75_bit_slice_1091180_comb;
  wire [7:0] p75_bit_slice_1091181_comb;
  wire [7:0] p75_bit_slice_1091182_comb;
  wire [7:0] p75_bit_slice_1091183_comb;
  wire [7:0] p75_bit_slice_1091184_comb;
  assign p75_res7__618_comb = p74_array_index_1090834 ^ p74_array_index_1090835 ^ p74_array_index_1090836 ^ p74_array_index_1090837 ^ p74_array_index_1090838 ^ p74_array_index_1090839 ^ p74_res7__611 ^ p74_array_index_1090840 ^ p74_res7__609 ^ p74_array_index_1090793 ^ p74_array_index_1090514 ^ p74_array_index_1090485 ^ p74_array_index_1090453 ^ p74_array_index_1090841 ^ p74_array_index_1090842 ^ p74_array_index_1090443;
  assign p75_res7__394_comb = p74_array_index_1090766 ^ p74_array_index_1090767 ^ p74_array_index_1090768 ^ p74_array_index_1090769 ^ p74_array_index_1090770 ^ p74_array_index_1090771 ^ p74_res7__387 ^ p74_array_index_1090772 ^ p74_res7__385 ^ p74_array_index_1090725 ^ p74_array_index_1090429 ^ p74_array_index_1090400 ^ p74_array_index_1090368 ^ p74_array_index_1090773 ^ p74_array_index_1090774 ^ p74_array_index_1090355;
  assign p75_array_index_1091128_comb = p74_literal_1076355[p74_res7__613];
  assign p75_array_index_1091081_comb = p74_literal_1076355[p74_res7__389];
  assign p75_res7__619_comb = p74_literal_1076345[p75_res7__618_comb] ^ p74_literal_1076347[p74_res7__617] ^ p74_literal_1076349[p74_res7__616] ^ p74_literal_1076351[p74_res7__615] ^ p74_literal_1076353[p74_res7__614] ^ p75_array_index_1091128_comb ^ p74_res7__612 ^ p74_literal_1076358[p74_res7__611] ^ p74_res7__610 ^ p74_array_index_1090805 ^ p74_array_index_1090779 ^ p74_array_index_1090499 ^ p74_array_index_1090470 ^ p74_literal_1076347[p74_array_index_1090440] ^ p74_literal_1076345[p74_array_index_1090441] ^ p74_array_index_1090442;
  assign p75_res7__395_comb = p74_literal_1076345[p75_res7__394_comb] ^ p74_literal_1076347[p74_res7__393] ^ p74_literal_1076349[p74_res7__392] ^ p74_literal_1076351[p74_res7__391] ^ p74_literal_1076353[p74_res7__390] ^ p75_array_index_1091081_comb ^ p74_res7__388 ^ p74_literal_1076358[p74_res7__387] ^ p74_res7__386 ^ p74_array_index_1090737 ^ p74_array_index_1090711 ^ p74_array_index_1090414 ^ p74_array_index_1090385 ^ p74_literal_1076347[p74_array_index_1090352] ^ p74_literal_1076345[p74_array_index_1090353] ^ p74_array_index_1090354;
  assign p75_res7__620_comb = p74_literal_1076345[p75_res7__619_comb] ^ p74_literal_1076347[p75_res7__618_comb] ^ p74_literal_1076349[p74_res7__617] ^ p74_literal_1076351[p74_res7__616] ^ p74_literal_1076353[p74_res7__615] ^ p74_literal_1076355[p74_res7__614] ^ p74_res7__613 ^ p74_literal_1076358[p74_res7__612] ^ p74_res7__611 ^ p74_array_index_1090817 ^ p74_array_index_1090792 ^ p74_array_index_1090513 ^ p74_array_index_1090484 ^ p74_array_index_1090452 ^ p74_literal_1076345[p74_array_index_1090440] ^ p74_array_index_1090441;
  assign p75_res7__396_comb = p74_literal_1076345[p75_res7__395_comb] ^ p74_literal_1076347[p75_res7__394_comb] ^ p74_literal_1076349[p74_res7__393] ^ p74_literal_1076351[p74_res7__392] ^ p74_literal_1076353[p74_res7__391] ^ p74_literal_1076355[p74_res7__390] ^ p74_res7__389 ^ p74_literal_1076358[p74_res7__388] ^ p74_res7__387 ^ p74_array_index_1090749 ^ p74_array_index_1090724 ^ p74_array_index_1090428 ^ p74_array_index_1090399 ^ p74_array_index_1090367 ^ p74_literal_1076345[p74_array_index_1090352] ^ p74_array_index_1090353;
  assign p75_res7__621_comb = p74_literal_1076345[p75_res7__620_comb] ^ p74_literal_1076347[p75_res7__619_comb] ^ p74_literal_1076349[p75_res7__618_comb] ^ p74_literal_1076351[p74_res7__617] ^ p74_literal_1076353[p74_res7__616] ^ p74_literal_1076355[p74_res7__615] ^ p74_res7__614 ^ p74_literal_1076358[p74_res7__613] ^ p74_res7__612 ^ p74_array_index_1090828 ^ p74_array_index_1090804 ^ p74_array_index_1090778 ^ p74_array_index_1090498 ^ p74_array_index_1090469 ^ p74_literal_1076345[p74_array_index_1090439] ^ p74_array_index_1090440;
  assign p75_res7__397_comb = p74_literal_1076345[p75_res7__396_comb] ^ p74_literal_1076347[p75_res7__395_comb] ^ p74_literal_1076349[p75_res7__394_comb] ^ p74_literal_1076351[p74_res7__393] ^ p74_literal_1076353[p74_res7__392] ^ p74_literal_1076355[p74_res7__391] ^ p74_res7__390 ^ p74_literal_1076358[p74_res7__389] ^ p74_res7__388 ^ p74_array_index_1090760 ^ p74_array_index_1090736 ^ p74_array_index_1090710 ^ p74_array_index_1090413 ^ p74_array_index_1090384 ^ p74_literal_1076345[p74_array_index_1090351] ^ p74_array_index_1090352;
  assign p75_res7__622_comb = p74_literal_1076345[p75_res7__621_comb] ^ p74_literal_1076347[p75_res7__620_comb] ^ p74_literal_1076349[p75_res7__619_comb] ^ p74_literal_1076351[p75_res7__618_comb] ^ p74_literal_1076353[p74_res7__617] ^ p74_literal_1076355[p74_res7__616] ^ p74_res7__615 ^ p74_literal_1076358[p74_res7__614] ^ p74_res7__613 ^ p74_array_index_1090839 ^ p74_array_index_1090816 ^ p74_array_index_1090791 ^ p74_array_index_1090512 ^ p74_array_index_1090483 ^ p74_array_index_1090451 ^ p74_array_index_1090439;
  assign p75_res7__398_comb = p74_literal_1076345[p75_res7__397_comb] ^ p74_literal_1076347[p75_res7__396_comb] ^ p74_literal_1076349[p75_res7__395_comb] ^ p74_literal_1076351[p75_res7__394_comb] ^ p74_literal_1076353[p74_res7__393] ^ p74_literal_1076355[p74_res7__392] ^ p74_res7__391 ^ p74_literal_1076358[p74_res7__390] ^ p74_res7__389 ^ p74_array_index_1090771 ^ p74_array_index_1090748 ^ p74_array_index_1090723 ^ p74_array_index_1090427 ^ p74_array_index_1090398 ^ p74_array_index_1090366 ^ p74_array_index_1090351;
  assign p75_res7__623_comb = p74_literal_1076345[p75_res7__622_comb] ^ p74_literal_1076347[p75_res7__621_comb] ^ p74_literal_1076349[p75_res7__620_comb] ^ p74_literal_1076351[p75_res7__619_comb] ^ p74_literal_1076353[p75_res7__618_comb] ^ p74_literal_1076355[p74_res7__617] ^ p74_res7__616 ^ p74_literal_1076358[p74_res7__615] ^ p74_res7__614 ^ p75_array_index_1091128_comb ^ p74_array_index_1090827 ^ p74_array_index_1090803 ^ p74_array_index_1090777 ^ p74_array_index_1090497 ^ p74_array_index_1090468 ^ p74_array_index_1090438;
  assign p75_res7__399_comb = p74_literal_1076345[p75_res7__398_comb] ^ p74_literal_1076347[p75_res7__397_comb] ^ p74_literal_1076349[p75_res7__396_comb] ^ p74_literal_1076351[p75_res7__395_comb] ^ p74_literal_1076353[p75_res7__394_comb] ^ p74_literal_1076355[p74_res7__393] ^ p74_res7__392 ^ p74_literal_1076358[p74_res7__391] ^ p74_res7__390 ^ p75_array_index_1091081_comb ^ p74_array_index_1090759 ^ p74_array_index_1090735 ^ p74_array_index_1090709 ^ p74_array_index_1090412 ^ p74_array_index_1090383 ^ p74_array_index_1090350;
  assign p75_res__38_comb = {p75_res7__623_comb, p75_res7__622_comb, p75_res7__621_comb, p75_res7__620_comb, p75_res7__619_comb, p75_res7__618_comb, p74_res7__617, p74_res7__616, p74_res7__615, p74_res7__614, p74_res7__613, p74_res7__612, p74_res7__611, p74_res7__610, p74_res7__609, p74_res7__608};
  assign p75_res__24_comb = {p75_res7__399_comb, p75_res7__398_comb, p75_res7__397_comb, p75_res7__396_comb, p75_res7__395_comb, p75_res7__394_comb, p74_res7__393, p74_res7__392, p74_res7__391, p74_res7__390, p74_res7__389, p74_res7__388, p74_res7__387, p74_res7__386, p74_res7__385, p74_res7__384};
  assign p75_addedKey__39_comb = p74_k7 ^ p75_res__38_comb;
  assign p75_xor_1091121_comb = p75_res__24_comb ^ p74_k7;
  assign p75_bit_slice_1091169_comb = p75_addedKey__39_comb[127:120];
  assign p75_bit_slice_1091170_comb = p75_addedKey__39_comb[119:112];
  assign p75_bit_slice_1091171_comb = p75_addedKey__39_comb[111:104];
  assign p75_bit_slice_1091172_comb = p75_addedKey__39_comb[103:96];
  assign p75_bit_slice_1091173_comb = p75_addedKey__39_comb[95:88];
  assign p75_bit_slice_1091174_comb = p75_addedKey__39_comb[87:80];
  assign p75_bit_slice_1091175_comb = p75_addedKey__39_comb[71:64];
  assign p75_bit_slice_1091176_comb = p75_addedKey__39_comb[55:48];
  assign p75_bit_slice_1091177_comb = p75_addedKey__39_comb[47:40];
  assign p75_bit_slice_1091178_comb = p75_addedKey__39_comb[39:32];
  assign p75_bit_slice_1091179_comb = p75_addedKey__39_comb[31:24];
  assign p75_bit_slice_1091180_comb = p75_addedKey__39_comb[23:16];
  assign p75_bit_slice_1091181_comb = p75_addedKey__39_comb[15:8];
  assign p75_bit_slice_1091182_comb = p75_addedKey__39_comb[79:72];
  assign p75_bit_slice_1091183_comb = p75_addedKey__39_comb[63:56];
  assign p75_bit_slice_1091184_comb = p75_addedKey__39_comb[7:0];

  // Registers for pipe stage 75:
  reg [127:0] p75_k6;
  reg [127:0] p75_xor_1091121;
  reg [7:0] p75_bit_slice_1091169;
  reg [7:0] p75_bit_slice_1091170;
  reg [7:0] p75_bit_slice_1091171;
  reg [7:0] p75_bit_slice_1091172;
  reg [7:0] p75_bit_slice_1091173;
  reg [7:0] p75_bit_slice_1091174;
  reg [7:0] p75_bit_slice_1091175;
  reg [7:0] p75_bit_slice_1091176;
  reg [7:0] p75_bit_slice_1091177;
  reg [7:0] p75_bit_slice_1091178;
  reg [7:0] p75_bit_slice_1091179;
  reg [7:0] p75_bit_slice_1091180;
  reg [7:0] p75_bit_slice_1091181;
  reg [7:0] p75_bit_slice_1091182;
  reg [7:0] p75_bit_slice_1091183;
  reg [7:0] p75_bit_slice_1091184;
  reg [7:0] p76_arr[256];
  reg [7:0] p76_literal_1076345[256];
  reg [7:0] p76_literal_1076347[256];
  reg [7:0] p76_literal_1076349[256];
  reg [7:0] p76_literal_1076351[256];
  reg [7:0] p76_literal_1076353[256];
  reg [7:0] p76_literal_1076355[256];
  reg [7:0] p76_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p75_k6 <= p74_k6;
    p75_xor_1091121 <= p75_xor_1091121_comb;
    p75_bit_slice_1091169 <= p75_bit_slice_1091169_comb;
    p75_bit_slice_1091170 <= p75_bit_slice_1091170_comb;
    p75_bit_slice_1091171 <= p75_bit_slice_1091171_comb;
    p75_bit_slice_1091172 <= p75_bit_slice_1091172_comb;
    p75_bit_slice_1091173 <= p75_bit_slice_1091173_comb;
    p75_bit_slice_1091174 <= p75_bit_slice_1091174_comb;
    p75_bit_slice_1091175 <= p75_bit_slice_1091175_comb;
    p75_bit_slice_1091176 <= p75_bit_slice_1091176_comb;
    p75_bit_slice_1091177 <= p75_bit_slice_1091177_comb;
    p75_bit_slice_1091178 <= p75_bit_slice_1091178_comb;
    p75_bit_slice_1091179 <= p75_bit_slice_1091179_comb;
    p75_bit_slice_1091180 <= p75_bit_slice_1091180_comb;
    p75_bit_slice_1091181 <= p75_bit_slice_1091181_comb;
    p75_bit_slice_1091182 <= p75_bit_slice_1091182_comb;
    p75_bit_slice_1091183 <= p75_bit_slice_1091183_comb;
    p75_bit_slice_1091184 <= p75_bit_slice_1091184_comb;
    p76_arr <= p75_arr;
    p76_literal_1076345 <= p75_literal_1076345;
    p76_literal_1076347 <= p75_literal_1076347;
    p76_literal_1076349 <= p75_literal_1076349;
    p76_literal_1076351 <= p75_literal_1076351;
    p76_literal_1076353 <= p75_literal_1076353;
    p76_literal_1076355 <= p75_literal_1076355;
    p76_literal_1076358 <= p75_literal_1076358;
  end

  // ===== Pipe stage 76:
  wire [127:0] p76_addedKey__66_comb;
  wire [7:0] p76_array_index_1091252_comb;
  wire [7:0] p76_array_index_1091253_comb;
  wire [7:0] p76_array_index_1091254_comb;
  wire [7:0] p76_array_index_1091255_comb;
  wire [7:0] p76_array_index_1091256_comb;
  wire [7:0] p76_array_index_1091257_comb;
  wire [7:0] p76_array_index_1091259_comb;
  wire [7:0] p76_array_index_1091261_comb;
  wire [7:0] p76_array_index_1091262_comb;
  wire [7:0] p76_array_index_1091263_comb;
  wire [7:0] p76_array_index_1091264_comb;
  wire [7:0] p76_array_index_1091265_comb;
  wire [7:0] p76_array_index_1091266_comb;
  wire [7:0] p76_array_index_1091340_comb;
  wire [7:0] p76_array_index_1091341_comb;
  wire [7:0] p76_array_index_1091342_comb;
  wire [7:0] p76_array_index_1091343_comb;
  wire [7:0] p76_array_index_1091344_comb;
  wire [7:0] p76_array_index_1091345_comb;
  wire [7:0] p76_array_index_1091346_comb;
  wire [7:0] p76_array_index_1091347_comb;
  wire [7:0] p76_array_index_1091348_comb;
  wire [7:0] p76_array_index_1091349_comb;
  wire [7:0] p76_array_index_1091350_comb;
  wire [7:0] p76_array_index_1091351_comb;
  wire [7:0] p76_array_index_1091352_comb;
  wire [7:0] p76_array_index_1091268_comb;
  wire [7:0] p76_array_index_1091269_comb;
  wire [7:0] p76_array_index_1091270_comb;
  wire [7:0] p76_array_index_1091271_comb;
  wire [7:0] p76_array_index_1091272_comb;
  wire [7:0] p76_array_index_1091273_comb;
  wire [7:0] p76_array_index_1091274_comb;
  wire [7:0] p76_array_index_1091276_comb;
  wire [7:0] p76_array_index_1091353_comb;
  wire [7:0] p76_array_index_1091354_comb;
  wire [7:0] p76_array_index_1091355_comb;
  wire [7:0] p76_array_index_1091356_comb;
  wire [7:0] p76_array_index_1091357_comb;
  wire [7:0] p76_array_index_1091358_comb;
  wire [7:0] p76_array_index_1091359_comb;
  wire [7:0] p76_array_index_1091361_comb;
  wire [7:0] p76_res7__400_comb;
  wire [7:0] p76_res7__624_comb;
  wire [7:0] p76_array_index_1091285_comb;
  wire [7:0] p76_array_index_1091286_comb;
  wire [7:0] p76_array_index_1091287_comb;
  wire [7:0] p76_array_index_1091288_comb;
  wire [7:0] p76_array_index_1091289_comb;
  wire [7:0] p76_array_index_1091290_comb;
  wire [7:0] p76_array_index_1091370_comb;
  wire [7:0] p76_array_index_1091371_comb;
  wire [7:0] p76_array_index_1091372_comb;
  wire [7:0] p76_array_index_1091373_comb;
  wire [7:0] p76_array_index_1091374_comb;
  wire [7:0] p76_array_index_1091375_comb;
  wire [7:0] p76_res7__401_comb;
  wire [7:0] p76_res7__625_comb;
  wire [7:0] p76_array_index_1091300_comb;
  wire [7:0] p76_array_index_1091301_comb;
  wire [7:0] p76_array_index_1091302_comb;
  wire [7:0] p76_array_index_1091303_comb;
  wire [7:0] p76_array_index_1091304_comb;
  wire [7:0] p76_array_index_1091385_comb;
  wire [7:0] p76_array_index_1091386_comb;
  wire [7:0] p76_array_index_1091387_comb;
  wire [7:0] p76_array_index_1091388_comb;
  wire [7:0] p76_array_index_1091389_comb;
  wire [7:0] p76_res7__402_comb;
  wire [7:0] p76_res7__626_comb;
  wire [7:0] p76_array_index_1091314_comb;
  wire [7:0] p76_array_index_1091315_comb;
  wire [7:0] p76_array_index_1091316_comb;
  wire [7:0] p76_array_index_1091317_comb;
  wire [7:0] p76_array_index_1091318_comb;
  wire [7:0] p76_array_index_1091399_comb;
  wire [7:0] p76_array_index_1091400_comb;
  wire [7:0] p76_array_index_1091401_comb;
  wire [7:0] p76_array_index_1091402_comb;
  wire [7:0] p76_array_index_1091403_comb;
  wire [7:0] p76_res7__403_comb;
  wire [7:0] p76_res7__627_comb;
  wire [7:0] p76_array_index_1091329_comb;
  wire [7:0] p76_array_index_1091330_comb;
  wire [7:0] p76_array_index_1091331_comb;
  wire [7:0] p76_array_index_1091332_comb;
  wire [7:0] p76_array_index_1091414_comb;
  wire [7:0] p76_array_index_1091415_comb;
  wire [7:0] p76_array_index_1091416_comb;
  wire [7:0] p76_array_index_1091417_comb;
  wire [7:0] p76_res7__404_comb;
  wire [7:0] p76_res7__628_comb;
  assign p76_addedKey__66_comb = p75_xor_1091121 ^ 128'h056c_b6de_319f_0eeb_8e80_9963_10f6_951a;
  assign p76_array_index_1091252_comb = p75_arr[p76_addedKey__66_comb[127:120]];
  assign p76_array_index_1091253_comb = p75_arr[p76_addedKey__66_comb[119:112]];
  assign p76_array_index_1091254_comb = p75_arr[p76_addedKey__66_comb[111:104]];
  assign p76_array_index_1091255_comb = p75_arr[p76_addedKey__66_comb[103:96]];
  assign p76_array_index_1091256_comb = p75_arr[p76_addedKey__66_comb[95:88]];
  assign p76_array_index_1091257_comb = p75_arr[p76_addedKey__66_comb[87:80]];
  assign p76_array_index_1091259_comb = p75_arr[p76_addedKey__66_comb[71:64]];
  assign p76_array_index_1091261_comb = p75_arr[p76_addedKey__66_comb[55:48]];
  assign p76_array_index_1091262_comb = p75_arr[p76_addedKey__66_comb[47:40]];
  assign p76_array_index_1091263_comb = p75_arr[p76_addedKey__66_comb[39:32]];
  assign p76_array_index_1091264_comb = p75_arr[p76_addedKey__66_comb[31:24]];
  assign p76_array_index_1091265_comb = p75_arr[p76_addedKey__66_comb[23:16]];
  assign p76_array_index_1091266_comb = p75_arr[p76_addedKey__66_comb[15:8]];
  assign p76_array_index_1091340_comb = p75_arr[p75_bit_slice_1091169];
  assign p76_array_index_1091341_comb = p75_arr[p75_bit_slice_1091170];
  assign p76_array_index_1091342_comb = p75_arr[p75_bit_slice_1091171];
  assign p76_array_index_1091343_comb = p75_arr[p75_bit_slice_1091172];
  assign p76_array_index_1091344_comb = p75_arr[p75_bit_slice_1091173];
  assign p76_array_index_1091345_comb = p75_arr[p75_bit_slice_1091174];
  assign p76_array_index_1091346_comb = p75_arr[p75_bit_slice_1091175];
  assign p76_array_index_1091347_comb = p75_arr[p75_bit_slice_1091176];
  assign p76_array_index_1091348_comb = p75_arr[p75_bit_slice_1091177];
  assign p76_array_index_1091349_comb = p75_arr[p75_bit_slice_1091178];
  assign p76_array_index_1091350_comb = p75_arr[p75_bit_slice_1091179];
  assign p76_array_index_1091351_comb = p75_arr[p75_bit_slice_1091180];
  assign p76_array_index_1091352_comb = p75_arr[p75_bit_slice_1091181];
  assign p76_array_index_1091268_comb = p75_literal_1076345[p76_array_index_1091252_comb];
  assign p76_array_index_1091269_comb = p75_literal_1076347[p76_array_index_1091253_comb];
  assign p76_array_index_1091270_comb = p75_literal_1076349[p76_array_index_1091254_comb];
  assign p76_array_index_1091271_comb = p75_literal_1076351[p76_array_index_1091255_comb];
  assign p76_array_index_1091272_comb = p75_literal_1076353[p76_array_index_1091256_comb];
  assign p76_array_index_1091273_comb = p75_literal_1076355[p76_array_index_1091257_comb];
  assign p76_array_index_1091274_comb = p75_arr[p76_addedKey__66_comb[79:72]];
  assign p76_array_index_1091276_comb = p75_arr[p76_addedKey__66_comb[63:56]];
  assign p76_array_index_1091353_comb = p75_literal_1076345[p76_array_index_1091340_comb];
  assign p76_array_index_1091354_comb = p75_literal_1076347[p76_array_index_1091341_comb];
  assign p76_array_index_1091355_comb = p75_literal_1076349[p76_array_index_1091342_comb];
  assign p76_array_index_1091356_comb = p75_literal_1076351[p76_array_index_1091343_comb];
  assign p76_array_index_1091357_comb = p75_literal_1076353[p76_array_index_1091344_comb];
  assign p76_array_index_1091358_comb = p75_literal_1076355[p76_array_index_1091345_comb];
  assign p76_array_index_1091359_comb = p75_arr[p75_bit_slice_1091182];
  assign p76_array_index_1091361_comb = p75_arr[p75_bit_slice_1091183];
  assign p76_res7__400_comb = p76_array_index_1091268_comb ^ p76_array_index_1091269_comb ^ p76_array_index_1091270_comb ^ p76_array_index_1091271_comb ^ p76_array_index_1091272_comb ^ p76_array_index_1091273_comb ^ p76_array_index_1091274_comb ^ p75_literal_1076358[p76_array_index_1091259_comb] ^ p76_array_index_1091276_comb ^ p75_literal_1076355[p76_array_index_1091261_comb] ^ p75_literal_1076353[p76_array_index_1091262_comb] ^ p75_literal_1076351[p76_array_index_1091263_comb] ^ p75_literal_1076349[p76_array_index_1091264_comb] ^ p75_literal_1076347[p76_array_index_1091265_comb] ^ p75_literal_1076345[p76_array_index_1091266_comb] ^ p75_arr[p76_addedKey__66_comb[7:0]];
  assign p76_res7__624_comb = p76_array_index_1091353_comb ^ p76_array_index_1091354_comb ^ p76_array_index_1091355_comb ^ p76_array_index_1091356_comb ^ p76_array_index_1091357_comb ^ p76_array_index_1091358_comb ^ p76_array_index_1091359_comb ^ p75_literal_1076358[p76_array_index_1091346_comb] ^ p76_array_index_1091361_comb ^ p75_literal_1076355[p76_array_index_1091347_comb] ^ p75_literal_1076353[p76_array_index_1091348_comb] ^ p75_literal_1076351[p76_array_index_1091349_comb] ^ p75_literal_1076349[p76_array_index_1091350_comb] ^ p75_literal_1076347[p76_array_index_1091351_comb] ^ p75_literal_1076345[p76_array_index_1091352_comb] ^ p75_arr[p75_bit_slice_1091184];
  assign p76_array_index_1091285_comb = p75_literal_1076345[p76_res7__400_comb];
  assign p76_array_index_1091286_comb = p75_literal_1076347[p76_array_index_1091252_comb];
  assign p76_array_index_1091287_comb = p75_literal_1076349[p76_array_index_1091253_comb];
  assign p76_array_index_1091288_comb = p75_literal_1076351[p76_array_index_1091254_comb];
  assign p76_array_index_1091289_comb = p75_literal_1076353[p76_array_index_1091255_comb];
  assign p76_array_index_1091290_comb = p75_literal_1076355[p76_array_index_1091256_comb];
  assign p76_array_index_1091370_comb = p75_literal_1076345[p76_res7__624_comb];
  assign p76_array_index_1091371_comb = p75_literal_1076347[p76_array_index_1091340_comb];
  assign p76_array_index_1091372_comb = p75_literal_1076349[p76_array_index_1091341_comb];
  assign p76_array_index_1091373_comb = p75_literal_1076351[p76_array_index_1091342_comb];
  assign p76_array_index_1091374_comb = p75_literal_1076353[p76_array_index_1091343_comb];
  assign p76_array_index_1091375_comb = p75_literal_1076355[p76_array_index_1091344_comb];
  assign p76_res7__401_comb = p76_array_index_1091285_comb ^ p76_array_index_1091286_comb ^ p76_array_index_1091287_comb ^ p76_array_index_1091288_comb ^ p76_array_index_1091289_comb ^ p76_array_index_1091290_comb ^ p76_array_index_1091257_comb ^ p75_literal_1076358[p76_array_index_1091274_comb] ^ p76_array_index_1091259_comb ^ p75_literal_1076355[p76_array_index_1091276_comb] ^ p75_literal_1076353[p76_array_index_1091261_comb] ^ p75_literal_1076351[p76_array_index_1091262_comb] ^ p75_literal_1076349[p76_array_index_1091263_comb] ^ p75_literal_1076347[p76_array_index_1091264_comb] ^ p75_literal_1076345[p76_array_index_1091265_comb] ^ p76_array_index_1091266_comb;
  assign p76_res7__625_comb = p76_array_index_1091370_comb ^ p76_array_index_1091371_comb ^ p76_array_index_1091372_comb ^ p76_array_index_1091373_comb ^ p76_array_index_1091374_comb ^ p76_array_index_1091375_comb ^ p76_array_index_1091345_comb ^ p75_literal_1076358[p76_array_index_1091359_comb] ^ p76_array_index_1091346_comb ^ p75_literal_1076355[p76_array_index_1091361_comb] ^ p75_literal_1076353[p76_array_index_1091347_comb] ^ p75_literal_1076351[p76_array_index_1091348_comb] ^ p75_literal_1076349[p76_array_index_1091349_comb] ^ p75_literal_1076347[p76_array_index_1091350_comb] ^ p75_literal_1076345[p76_array_index_1091351_comb] ^ p76_array_index_1091352_comb;
  assign p76_array_index_1091300_comb = p75_literal_1076347[p76_res7__400_comb];
  assign p76_array_index_1091301_comb = p75_literal_1076349[p76_array_index_1091252_comb];
  assign p76_array_index_1091302_comb = p75_literal_1076351[p76_array_index_1091253_comb];
  assign p76_array_index_1091303_comb = p75_literal_1076353[p76_array_index_1091254_comb];
  assign p76_array_index_1091304_comb = p75_literal_1076355[p76_array_index_1091255_comb];
  assign p76_array_index_1091385_comb = p75_literal_1076347[p76_res7__624_comb];
  assign p76_array_index_1091386_comb = p75_literal_1076349[p76_array_index_1091340_comb];
  assign p76_array_index_1091387_comb = p75_literal_1076351[p76_array_index_1091341_comb];
  assign p76_array_index_1091388_comb = p75_literal_1076353[p76_array_index_1091342_comb];
  assign p76_array_index_1091389_comb = p75_literal_1076355[p76_array_index_1091343_comb];
  assign p76_res7__402_comb = p75_literal_1076345[p76_res7__401_comb] ^ p76_array_index_1091300_comb ^ p76_array_index_1091301_comb ^ p76_array_index_1091302_comb ^ p76_array_index_1091303_comb ^ p76_array_index_1091304_comb ^ p76_array_index_1091256_comb ^ p75_literal_1076358[p76_array_index_1091257_comb] ^ p76_array_index_1091274_comb ^ p75_literal_1076355[p76_array_index_1091259_comb] ^ p75_literal_1076353[p76_array_index_1091276_comb] ^ p75_literal_1076351[p76_array_index_1091261_comb] ^ p75_literal_1076349[p76_array_index_1091262_comb] ^ p75_literal_1076347[p76_array_index_1091263_comb] ^ p75_literal_1076345[p76_array_index_1091264_comb] ^ p76_array_index_1091265_comb;
  assign p76_res7__626_comb = p75_literal_1076345[p76_res7__625_comb] ^ p76_array_index_1091385_comb ^ p76_array_index_1091386_comb ^ p76_array_index_1091387_comb ^ p76_array_index_1091388_comb ^ p76_array_index_1091389_comb ^ p76_array_index_1091344_comb ^ p75_literal_1076358[p76_array_index_1091345_comb] ^ p76_array_index_1091359_comb ^ p75_literal_1076355[p76_array_index_1091346_comb] ^ p75_literal_1076353[p76_array_index_1091361_comb] ^ p75_literal_1076351[p76_array_index_1091347_comb] ^ p75_literal_1076349[p76_array_index_1091348_comb] ^ p75_literal_1076347[p76_array_index_1091349_comb] ^ p75_literal_1076345[p76_array_index_1091350_comb] ^ p76_array_index_1091351_comb;
  assign p76_array_index_1091314_comb = p75_literal_1076347[p76_res7__401_comb];
  assign p76_array_index_1091315_comb = p75_literal_1076349[p76_res7__400_comb];
  assign p76_array_index_1091316_comb = p75_literal_1076351[p76_array_index_1091252_comb];
  assign p76_array_index_1091317_comb = p75_literal_1076353[p76_array_index_1091253_comb];
  assign p76_array_index_1091318_comb = p75_literal_1076355[p76_array_index_1091254_comb];
  assign p76_array_index_1091399_comb = p75_literal_1076347[p76_res7__625_comb];
  assign p76_array_index_1091400_comb = p75_literal_1076349[p76_res7__624_comb];
  assign p76_array_index_1091401_comb = p75_literal_1076351[p76_array_index_1091340_comb];
  assign p76_array_index_1091402_comb = p75_literal_1076353[p76_array_index_1091341_comb];
  assign p76_array_index_1091403_comb = p75_literal_1076355[p76_array_index_1091342_comb];
  assign p76_res7__403_comb = p75_literal_1076345[p76_res7__402_comb] ^ p76_array_index_1091314_comb ^ p76_array_index_1091315_comb ^ p76_array_index_1091316_comb ^ p76_array_index_1091317_comb ^ p76_array_index_1091318_comb ^ p76_array_index_1091255_comb ^ p75_literal_1076358[p76_array_index_1091256_comb] ^ p76_array_index_1091257_comb ^ p75_literal_1076355[p76_array_index_1091274_comb] ^ p75_literal_1076353[p76_array_index_1091259_comb] ^ p75_literal_1076351[p76_array_index_1091276_comb] ^ p75_literal_1076349[p76_array_index_1091261_comb] ^ p75_literal_1076347[p76_array_index_1091262_comb] ^ p75_literal_1076345[p76_array_index_1091263_comb] ^ p76_array_index_1091264_comb;
  assign p76_res7__627_comb = p75_literal_1076345[p76_res7__626_comb] ^ p76_array_index_1091399_comb ^ p76_array_index_1091400_comb ^ p76_array_index_1091401_comb ^ p76_array_index_1091402_comb ^ p76_array_index_1091403_comb ^ p76_array_index_1091343_comb ^ p75_literal_1076358[p76_array_index_1091344_comb] ^ p76_array_index_1091345_comb ^ p75_literal_1076355[p76_array_index_1091359_comb] ^ p75_literal_1076353[p76_array_index_1091346_comb] ^ p75_literal_1076351[p76_array_index_1091361_comb] ^ p75_literal_1076349[p76_array_index_1091347_comb] ^ p75_literal_1076347[p76_array_index_1091348_comb] ^ p75_literal_1076345[p76_array_index_1091349_comb] ^ p76_array_index_1091350_comb;
  assign p76_array_index_1091329_comb = p75_literal_1076349[p76_res7__401_comb];
  assign p76_array_index_1091330_comb = p75_literal_1076351[p76_res7__400_comb];
  assign p76_array_index_1091331_comb = p75_literal_1076353[p76_array_index_1091252_comb];
  assign p76_array_index_1091332_comb = p75_literal_1076355[p76_array_index_1091253_comb];
  assign p76_array_index_1091414_comb = p75_literal_1076349[p76_res7__625_comb];
  assign p76_array_index_1091415_comb = p75_literal_1076351[p76_res7__624_comb];
  assign p76_array_index_1091416_comb = p75_literal_1076353[p76_array_index_1091340_comb];
  assign p76_array_index_1091417_comb = p75_literal_1076355[p76_array_index_1091341_comb];
  assign p76_res7__404_comb = p75_literal_1076345[p76_res7__403_comb] ^ p75_literal_1076347[p76_res7__402_comb] ^ p76_array_index_1091329_comb ^ p76_array_index_1091330_comb ^ p76_array_index_1091331_comb ^ p76_array_index_1091332_comb ^ p76_array_index_1091254_comb ^ p75_literal_1076358[p76_array_index_1091255_comb] ^ p76_array_index_1091256_comb ^ p76_array_index_1091273_comb ^ p75_literal_1076353[p76_array_index_1091274_comb] ^ p75_literal_1076351[p76_array_index_1091259_comb] ^ p75_literal_1076349[p76_array_index_1091276_comb] ^ p75_literal_1076347[p76_array_index_1091261_comb] ^ p75_literal_1076345[p76_array_index_1091262_comb] ^ p76_array_index_1091263_comb;
  assign p76_res7__628_comb = p75_literal_1076345[p76_res7__627_comb] ^ p75_literal_1076347[p76_res7__626_comb] ^ p76_array_index_1091414_comb ^ p76_array_index_1091415_comb ^ p76_array_index_1091416_comb ^ p76_array_index_1091417_comb ^ p76_array_index_1091342_comb ^ p75_literal_1076358[p76_array_index_1091343_comb] ^ p76_array_index_1091344_comb ^ p76_array_index_1091358_comb ^ p75_literal_1076353[p76_array_index_1091359_comb] ^ p75_literal_1076351[p76_array_index_1091346_comb] ^ p75_literal_1076349[p76_array_index_1091361_comb] ^ p75_literal_1076347[p76_array_index_1091347_comb] ^ p75_literal_1076345[p76_array_index_1091348_comb] ^ p76_array_index_1091349_comb;

  // Registers for pipe stage 76:
  reg [127:0] p76_k6;
  reg [127:0] p76_xor_1091121;
  reg [7:0] p76_array_index_1091252;
  reg [7:0] p76_array_index_1091253;
  reg [7:0] p76_array_index_1091254;
  reg [7:0] p76_array_index_1091255;
  reg [7:0] p76_array_index_1091256;
  reg [7:0] p76_array_index_1091257;
  reg [7:0] p76_array_index_1091259;
  reg [7:0] p76_array_index_1091261;
  reg [7:0] p76_array_index_1091262;
  reg [7:0] p76_array_index_1091268;
  reg [7:0] p76_array_index_1091269;
  reg [7:0] p76_array_index_1091270;
  reg [7:0] p76_array_index_1091271;
  reg [7:0] p76_array_index_1091272;
  reg [7:0] p76_array_index_1091274;
  reg [7:0] p76_array_index_1091276;
  reg [7:0] p76_res7__400;
  reg [7:0] p76_array_index_1091285;
  reg [7:0] p76_array_index_1091286;
  reg [7:0] p76_array_index_1091287;
  reg [7:0] p76_array_index_1091288;
  reg [7:0] p76_array_index_1091289;
  reg [7:0] p76_array_index_1091290;
  reg [7:0] p76_res7__401;
  reg [7:0] p76_array_index_1091300;
  reg [7:0] p76_array_index_1091301;
  reg [7:0] p76_array_index_1091302;
  reg [7:0] p76_array_index_1091303;
  reg [7:0] p76_array_index_1091304;
  reg [7:0] p76_res7__402;
  reg [7:0] p76_array_index_1091314;
  reg [7:0] p76_array_index_1091315;
  reg [7:0] p76_array_index_1091316;
  reg [7:0] p76_array_index_1091317;
  reg [7:0] p76_array_index_1091318;
  reg [7:0] p76_res7__403;
  reg [7:0] p76_array_index_1091329;
  reg [7:0] p76_array_index_1091330;
  reg [7:0] p76_array_index_1091331;
  reg [7:0] p76_array_index_1091332;
  reg [7:0] p76_res7__404;
  reg [7:0] p76_array_index_1091340;
  reg [7:0] p76_array_index_1091341;
  reg [7:0] p76_array_index_1091342;
  reg [7:0] p76_array_index_1091343;
  reg [7:0] p76_array_index_1091344;
  reg [7:0] p76_array_index_1091345;
  reg [7:0] p76_array_index_1091346;
  reg [7:0] p76_array_index_1091347;
  reg [7:0] p76_array_index_1091348;
  reg [7:0] p76_array_index_1091353;
  reg [7:0] p76_array_index_1091354;
  reg [7:0] p76_array_index_1091355;
  reg [7:0] p76_array_index_1091356;
  reg [7:0] p76_array_index_1091357;
  reg [7:0] p76_array_index_1091359;
  reg [7:0] p76_array_index_1091361;
  reg [7:0] p76_res7__624;
  reg [7:0] p76_array_index_1091370;
  reg [7:0] p76_array_index_1091371;
  reg [7:0] p76_array_index_1091372;
  reg [7:0] p76_array_index_1091373;
  reg [7:0] p76_array_index_1091374;
  reg [7:0] p76_array_index_1091375;
  reg [7:0] p76_res7__625;
  reg [7:0] p76_array_index_1091385;
  reg [7:0] p76_array_index_1091386;
  reg [7:0] p76_array_index_1091387;
  reg [7:0] p76_array_index_1091388;
  reg [7:0] p76_array_index_1091389;
  reg [7:0] p76_res7__626;
  reg [7:0] p76_array_index_1091399;
  reg [7:0] p76_array_index_1091400;
  reg [7:0] p76_array_index_1091401;
  reg [7:0] p76_array_index_1091402;
  reg [7:0] p76_array_index_1091403;
  reg [7:0] p76_res7__627;
  reg [7:0] p76_array_index_1091414;
  reg [7:0] p76_array_index_1091415;
  reg [7:0] p76_array_index_1091416;
  reg [7:0] p76_array_index_1091417;
  reg [7:0] p76_res7__628;
  reg [7:0] p77_arr[256];
  reg [7:0] p77_literal_1076345[256];
  reg [7:0] p77_literal_1076347[256];
  reg [7:0] p77_literal_1076349[256];
  reg [7:0] p77_literal_1076351[256];
  reg [7:0] p77_literal_1076353[256];
  reg [7:0] p77_literal_1076355[256];
  reg [7:0] p77_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p76_k6 <= p75_k6;
    p76_xor_1091121 <= p75_xor_1091121;
    p76_array_index_1091252 <= p76_array_index_1091252_comb;
    p76_array_index_1091253 <= p76_array_index_1091253_comb;
    p76_array_index_1091254 <= p76_array_index_1091254_comb;
    p76_array_index_1091255 <= p76_array_index_1091255_comb;
    p76_array_index_1091256 <= p76_array_index_1091256_comb;
    p76_array_index_1091257 <= p76_array_index_1091257_comb;
    p76_array_index_1091259 <= p76_array_index_1091259_comb;
    p76_array_index_1091261 <= p76_array_index_1091261_comb;
    p76_array_index_1091262 <= p76_array_index_1091262_comb;
    p76_array_index_1091268 <= p76_array_index_1091268_comb;
    p76_array_index_1091269 <= p76_array_index_1091269_comb;
    p76_array_index_1091270 <= p76_array_index_1091270_comb;
    p76_array_index_1091271 <= p76_array_index_1091271_comb;
    p76_array_index_1091272 <= p76_array_index_1091272_comb;
    p76_array_index_1091274 <= p76_array_index_1091274_comb;
    p76_array_index_1091276 <= p76_array_index_1091276_comb;
    p76_res7__400 <= p76_res7__400_comb;
    p76_array_index_1091285 <= p76_array_index_1091285_comb;
    p76_array_index_1091286 <= p76_array_index_1091286_comb;
    p76_array_index_1091287 <= p76_array_index_1091287_comb;
    p76_array_index_1091288 <= p76_array_index_1091288_comb;
    p76_array_index_1091289 <= p76_array_index_1091289_comb;
    p76_array_index_1091290 <= p76_array_index_1091290_comb;
    p76_res7__401 <= p76_res7__401_comb;
    p76_array_index_1091300 <= p76_array_index_1091300_comb;
    p76_array_index_1091301 <= p76_array_index_1091301_comb;
    p76_array_index_1091302 <= p76_array_index_1091302_comb;
    p76_array_index_1091303 <= p76_array_index_1091303_comb;
    p76_array_index_1091304 <= p76_array_index_1091304_comb;
    p76_res7__402 <= p76_res7__402_comb;
    p76_array_index_1091314 <= p76_array_index_1091314_comb;
    p76_array_index_1091315 <= p76_array_index_1091315_comb;
    p76_array_index_1091316 <= p76_array_index_1091316_comb;
    p76_array_index_1091317 <= p76_array_index_1091317_comb;
    p76_array_index_1091318 <= p76_array_index_1091318_comb;
    p76_res7__403 <= p76_res7__403_comb;
    p76_array_index_1091329 <= p76_array_index_1091329_comb;
    p76_array_index_1091330 <= p76_array_index_1091330_comb;
    p76_array_index_1091331 <= p76_array_index_1091331_comb;
    p76_array_index_1091332 <= p76_array_index_1091332_comb;
    p76_res7__404 <= p76_res7__404_comb;
    p76_array_index_1091340 <= p76_array_index_1091340_comb;
    p76_array_index_1091341 <= p76_array_index_1091341_comb;
    p76_array_index_1091342 <= p76_array_index_1091342_comb;
    p76_array_index_1091343 <= p76_array_index_1091343_comb;
    p76_array_index_1091344 <= p76_array_index_1091344_comb;
    p76_array_index_1091345 <= p76_array_index_1091345_comb;
    p76_array_index_1091346 <= p76_array_index_1091346_comb;
    p76_array_index_1091347 <= p76_array_index_1091347_comb;
    p76_array_index_1091348 <= p76_array_index_1091348_comb;
    p76_array_index_1091353 <= p76_array_index_1091353_comb;
    p76_array_index_1091354 <= p76_array_index_1091354_comb;
    p76_array_index_1091355 <= p76_array_index_1091355_comb;
    p76_array_index_1091356 <= p76_array_index_1091356_comb;
    p76_array_index_1091357 <= p76_array_index_1091357_comb;
    p76_array_index_1091359 <= p76_array_index_1091359_comb;
    p76_array_index_1091361 <= p76_array_index_1091361_comb;
    p76_res7__624 <= p76_res7__624_comb;
    p76_array_index_1091370 <= p76_array_index_1091370_comb;
    p76_array_index_1091371 <= p76_array_index_1091371_comb;
    p76_array_index_1091372 <= p76_array_index_1091372_comb;
    p76_array_index_1091373 <= p76_array_index_1091373_comb;
    p76_array_index_1091374 <= p76_array_index_1091374_comb;
    p76_array_index_1091375 <= p76_array_index_1091375_comb;
    p76_res7__625 <= p76_res7__625_comb;
    p76_array_index_1091385 <= p76_array_index_1091385_comb;
    p76_array_index_1091386 <= p76_array_index_1091386_comb;
    p76_array_index_1091387 <= p76_array_index_1091387_comb;
    p76_array_index_1091388 <= p76_array_index_1091388_comb;
    p76_array_index_1091389 <= p76_array_index_1091389_comb;
    p76_res7__626 <= p76_res7__626_comb;
    p76_array_index_1091399 <= p76_array_index_1091399_comb;
    p76_array_index_1091400 <= p76_array_index_1091400_comb;
    p76_array_index_1091401 <= p76_array_index_1091401_comb;
    p76_array_index_1091402 <= p76_array_index_1091402_comb;
    p76_array_index_1091403 <= p76_array_index_1091403_comb;
    p76_res7__627 <= p76_res7__627_comb;
    p76_array_index_1091414 <= p76_array_index_1091414_comb;
    p76_array_index_1091415 <= p76_array_index_1091415_comb;
    p76_array_index_1091416 <= p76_array_index_1091416_comb;
    p76_array_index_1091417 <= p76_array_index_1091417_comb;
    p76_res7__628 <= p76_res7__628_comb;
    p77_arr <= p76_arr;
    p77_literal_1076345 <= p76_literal_1076345;
    p77_literal_1076347 <= p76_literal_1076347;
    p77_literal_1076349 <= p76_literal_1076349;
    p77_literal_1076351 <= p76_literal_1076351;
    p77_literal_1076353 <= p76_literal_1076353;
    p77_literal_1076355 <= p76_literal_1076355;
    p77_literal_1076358 <= p76_literal_1076358;
  end

  // ===== Pipe stage 77:
  wire [7:0] p77_array_index_1091611_comb;
  wire [7:0] p77_array_index_1091612_comb;
  wire [7:0] p77_array_index_1091613_comb;
  wire [7:0] p77_array_index_1091614_comb;
  wire [7:0] p77_res7__405_comb;
  wire [7:0] p77_array_index_1091679_comb;
  wire [7:0] p77_array_index_1091680_comb;
  wire [7:0] p77_array_index_1091681_comb;
  wire [7:0] p77_array_index_1091682_comb;
  wire [7:0] p77_array_index_1091625_comb;
  wire [7:0] p77_array_index_1091626_comb;
  wire [7:0] p77_array_index_1091627_comb;
  wire [7:0] p77_res7__629_comb;
  wire [7:0] p77_res7__406_comb;
  wire [7:0] p77_array_index_1091693_comb;
  wire [7:0] p77_array_index_1091694_comb;
  wire [7:0] p77_array_index_1091695_comb;
  wire [7:0] p77_array_index_1091637_comb;
  wire [7:0] p77_array_index_1091638_comb;
  wire [7:0] p77_array_index_1091639_comb;
  wire [7:0] p77_res7__630_comb;
  wire [7:0] p77_res7__407_comb;
  wire [7:0] p77_array_index_1091705_comb;
  wire [7:0] p77_array_index_1091706_comb;
  wire [7:0] p77_array_index_1091707_comb;
  wire [7:0] p77_array_index_1091650_comb;
  wire [7:0] p77_array_index_1091651_comb;
  wire [7:0] p77_res7__631_comb;
  wire [7:0] p77_res7__408_comb;
  wire [7:0] p77_array_index_1091718_comb;
  wire [7:0] p77_array_index_1091719_comb;
  wire [7:0] p77_array_index_1091661_comb;
  wire [7:0] p77_array_index_1091662_comb;
  wire [7:0] p77_res7__632_comb;
  wire [7:0] p77_res7__409_comb;
  wire [7:0] p77_array_index_1091729_comb;
  wire [7:0] p77_array_index_1091730_comb;
  wire [7:0] p77_array_index_1091668_comb;
  wire [7:0] p77_array_index_1091669_comb;
  wire [7:0] p77_array_index_1091670_comb;
  wire [7:0] p77_array_index_1091671_comb;
  wire [7:0] p77_array_index_1091672_comb;
  wire [7:0] p77_array_index_1091673_comb;
  wire [7:0] p77_array_index_1091674_comb;
  wire [7:0] p77_array_index_1091675_comb;
  wire [7:0] p77_array_index_1091676_comb;
  wire [7:0] p77_res7__633_comb;
  assign p77_array_index_1091611_comb = p76_literal_1076349[p76_res7__402];
  assign p77_array_index_1091612_comb = p76_literal_1076351[p76_res7__401];
  assign p77_array_index_1091613_comb = p76_literal_1076353[p76_res7__400];
  assign p77_array_index_1091614_comb = p76_literal_1076355[p76_array_index_1091252];
  assign p77_res7__405_comb = p76_literal_1076345[p76_res7__404] ^ p76_literal_1076347[p76_res7__403] ^ p77_array_index_1091611_comb ^ p77_array_index_1091612_comb ^ p77_array_index_1091613_comb ^ p77_array_index_1091614_comb ^ p76_array_index_1091253 ^ p76_literal_1076358[p76_array_index_1091254] ^ p76_array_index_1091255 ^ p76_array_index_1091290 ^ p76_literal_1076353[p76_array_index_1091257] ^ p76_literal_1076351[p76_array_index_1091274] ^ p76_literal_1076349[p76_array_index_1091259] ^ p76_literal_1076347[p76_array_index_1091276] ^ p76_literal_1076345[p76_array_index_1091261] ^ p76_array_index_1091262;
  assign p77_array_index_1091679_comb = p76_literal_1076349[p76_res7__626];
  assign p77_array_index_1091680_comb = p76_literal_1076351[p76_res7__625];
  assign p77_array_index_1091681_comb = p76_literal_1076353[p76_res7__624];
  assign p77_array_index_1091682_comb = p76_literal_1076355[p76_array_index_1091340];
  assign p77_array_index_1091625_comb = p76_literal_1076351[p76_res7__402];
  assign p77_array_index_1091626_comb = p76_literal_1076353[p76_res7__401];
  assign p77_array_index_1091627_comb = p76_literal_1076355[p76_res7__400];
  assign p77_res7__629_comb = p76_literal_1076345[p76_res7__628] ^ p76_literal_1076347[p76_res7__627] ^ p77_array_index_1091679_comb ^ p77_array_index_1091680_comb ^ p77_array_index_1091681_comb ^ p77_array_index_1091682_comb ^ p76_array_index_1091341 ^ p76_literal_1076358[p76_array_index_1091342] ^ p76_array_index_1091343 ^ p76_array_index_1091375 ^ p76_literal_1076353[p76_array_index_1091345] ^ p76_literal_1076351[p76_array_index_1091359] ^ p76_literal_1076349[p76_array_index_1091346] ^ p76_literal_1076347[p76_array_index_1091361] ^ p76_literal_1076345[p76_array_index_1091347] ^ p76_array_index_1091348;
  assign p77_res7__406_comb = p76_literal_1076345[p77_res7__405_comb] ^ p76_literal_1076347[p76_res7__404] ^ p76_literal_1076349[p76_res7__403] ^ p77_array_index_1091625_comb ^ p77_array_index_1091626_comb ^ p77_array_index_1091627_comb ^ p76_array_index_1091252 ^ p76_literal_1076358[p76_array_index_1091253] ^ p76_array_index_1091254 ^ p76_array_index_1091304 ^ p76_array_index_1091272 ^ p76_literal_1076351[p76_array_index_1091257] ^ p76_literal_1076349[p76_array_index_1091274] ^ p76_literal_1076347[p76_array_index_1091259] ^ p76_literal_1076345[p76_array_index_1091276] ^ p76_array_index_1091261;
  assign p77_array_index_1091693_comb = p76_literal_1076351[p76_res7__626];
  assign p77_array_index_1091694_comb = p76_literal_1076353[p76_res7__625];
  assign p77_array_index_1091695_comb = p76_literal_1076355[p76_res7__624];
  assign p77_array_index_1091637_comb = p76_literal_1076351[p76_res7__403];
  assign p77_array_index_1091638_comb = p76_literal_1076353[p76_res7__402];
  assign p77_array_index_1091639_comb = p76_literal_1076355[p76_res7__401];
  assign p77_res7__630_comb = p76_literal_1076345[p77_res7__629_comb] ^ p76_literal_1076347[p76_res7__628] ^ p76_literal_1076349[p76_res7__627] ^ p77_array_index_1091693_comb ^ p77_array_index_1091694_comb ^ p77_array_index_1091695_comb ^ p76_array_index_1091340 ^ p76_literal_1076358[p76_array_index_1091341] ^ p76_array_index_1091342 ^ p76_array_index_1091389 ^ p76_array_index_1091357 ^ p76_literal_1076351[p76_array_index_1091345] ^ p76_literal_1076349[p76_array_index_1091359] ^ p76_literal_1076347[p76_array_index_1091346] ^ p76_literal_1076345[p76_array_index_1091361] ^ p76_array_index_1091347;
  assign p77_res7__407_comb = p76_literal_1076345[p77_res7__406_comb] ^ p76_literal_1076347[p77_res7__405_comb] ^ p76_literal_1076349[p76_res7__404] ^ p77_array_index_1091637_comb ^ p77_array_index_1091638_comb ^ p77_array_index_1091639_comb ^ p76_res7__400 ^ p76_literal_1076358[p76_array_index_1091252] ^ p76_array_index_1091253 ^ p76_array_index_1091318 ^ p76_array_index_1091289 ^ p76_literal_1076351[p76_array_index_1091256] ^ p76_literal_1076349[p76_array_index_1091257] ^ p76_literal_1076347[p76_array_index_1091274] ^ p76_literal_1076345[p76_array_index_1091259] ^ p76_array_index_1091276;
  assign p77_array_index_1091705_comb = p76_literal_1076351[p76_res7__627];
  assign p77_array_index_1091706_comb = p76_literal_1076353[p76_res7__626];
  assign p77_array_index_1091707_comb = p76_literal_1076355[p76_res7__625];
  assign p77_array_index_1091650_comb = p76_literal_1076353[p76_res7__403];
  assign p77_array_index_1091651_comb = p76_literal_1076355[p76_res7__402];
  assign p77_res7__631_comb = p76_literal_1076345[p77_res7__630_comb] ^ p76_literal_1076347[p77_res7__629_comb] ^ p76_literal_1076349[p76_res7__628] ^ p77_array_index_1091705_comb ^ p77_array_index_1091706_comb ^ p77_array_index_1091707_comb ^ p76_res7__624 ^ p76_literal_1076358[p76_array_index_1091340] ^ p76_array_index_1091341 ^ p76_array_index_1091403 ^ p76_array_index_1091374 ^ p76_literal_1076351[p76_array_index_1091344] ^ p76_literal_1076349[p76_array_index_1091345] ^ p76_literal_1076347[p76_array_index_1091359] ^ p76_literal_1076345[p76_array_index_1091346] ^ p76_array_index_1091361;
  assign p77_res7__408_comb = p76_literal_1076345[p77_res7__407_comb] ^ p76_literal_1076347[p77_res7__406_comb] ^ p76_literal_1076349[p77_res7__405_comb] ^ p76_literal_1076351[p76_res7__404] ^ p77_array_index_1091650_comb ^ p77_array_index_1091651_comb ^ p76_res7__401 ^ p76_literal_1076358[p76_res7__400] ^ p76_array_index_1091252 ^ p76_array_index_1091332 ^ p76_array_index_1091303 ^ p76_array_index_1091271 ^ p76_literal_1076349[p76_array_index_1091256] ^ p76_literal_1076347[p76_array_index_1091257] ^ p76_literal_1076345[p76_array_index_1091274] ^ p76_array_index_1091259;
  assign p77_array_index_1091718_comb = p76_literal_1076353[p76_res7__627];
  assign p77_array_index_1091719_comb = p76_literal_1076355[p76_res7__626];
  assign p77_array_index_1091661_comb = p76_literal_1076353[p76_res7__404];
  assign p77_array_index_1091662_comb = p76_literal_1076355[p76_res7__403];
  assign p77_res7__632_comb = p76_literal_1076345[p77_res7__631_comb] ^ p76_literal_1076347[p77_res7__630_comb] ^ p76_literal_1076349[p77_res7__629_comb] ^ p76_literal_1076351[p76_res7__628] ^ p77_array_index_1091718_comb ^ p77_array_index_1091719_comb ^ p76_res7__625 ^ p76_literal_1076358[p76_res7__624] ^ p76_array_index_1091340 ^ p76_array_index_1091417 ^ p76_array_index_1091388 ^ p76_array_index_1091356 ^ p76_literal_1076349[p76_array_index_1091344] ^ p76_literal_1076347[p76_array_index_1091345] ^ p76_literal_1076345[p76_array_index_1091359] ^ p76_array_index_1091346;
  assign p77_res7__409_comb = p76_literal_1076345[p77_res7__408_comb] ^ p76_literal_1076347[p77_res7__407_comb] ^ p76_literal_1076349[p77_res7__406_comb] ^ p76_literal_1076351[p77_res7__405_comb] ^ p77_array_index_1091661_comb ^ p77_array_index_1091662_comb ^ p76_res7__402 ^ p76_literal_1076358[p76_res7__401] ^ p76_res7__400 ^ p77_array_index_1091614_comb ^ p76_array_index_1091317 ^ p76_array_index_1091288 ^ p76_literal_1076349[p76_array_index_1091255] ^ p76_literal_1076347[p76_array_index_1091256] ^ p76_literal_1076345[p76_array_index_1091257] ^ p76_array_index_1091274;
  assign p77_array_index_1091729_comb = p76_literal_1076353[p76_res7__628];
  assign p77_array_index_1091730_comb = p76_literal_1076355[p76_res7__627];
  assign p77_array_index_1091668_comb = p76_literal_1076345[p77_res7__409_comb];
  assign p77_array_index_1091669_comb = p76_literal_1076347[p77_res7__408_comb];
  assign p77_array_index_1091670_comb = p76_literal_1076349[p77_res7__407_comb];
  assign p77_array_index_1091671_comb = p76_literal_1076351[p77_res7__406_comb];
  assign p77_array_index_1091672_comb = p76_literal_1076353[p77_res7__405_comb];
  assign p77_array_index_1091673_comb = p76_literal_1076355[p76_res7__404];
  assign p77_array_index_1091674_comb = p76_literal_1076358[p76_res7__402];
  assign p77_array_index_1091675_comb = p76_literal_1076347[p76_array_index_1091255];
  assign p77_array_index_1091676_comb = p76_literal_1076345[p76_array_index_1091256];
  assign p77_res7__633_comb = p76_literal_1076345[p77_res7__632_comb] ^ p76_literal_1076347[p77_res7__631_comb] ^ p76_literal_1076349[p77_res7__630_comb] ^ p76_literal_1076351[p77_res7__629_comb] ^ p77_array_index_1091729_comb ^ p77_array_index_1091730_comb ^ p76_res7__626 ^ p76_literal_1076358[p76_res7__625] ^ p76_res7__624 ^ p77_array_index_1091682_comb ^ p76_array_index_1091402 ^ p76_array_index_1091373 ^ p76_literal_1076349[p76_array_index_1091343] ^ p76_literal_1076347[p76_array_index_1091344] ^ p76_literal_1076345[p76_array_index_1091345] ^ p76_array_index_1091359;

  // Registers for pipe stage 77:
  reg [127:0] p77_k6;
  reg [127:0] p77_xor_1091121;
  reg [7:0] p77_array_index_1091252;
  reg [7:0] p77_array_index_1091253;
  reg [7:0] p77_array_index_1091254;
  reg [7:0] p77_array_index_1091255;
  reg [7:0] p77_array_index_1091256;
  reg [7:0] p77_array_index_1091257;
  reg [7:0] p77_array_index_1091268;
  reg [7:0] p77_array_index_1091269;
  reg [7:0] p77_array_index_1091270;
  reg [7:0] p77_res7__400;
  reg [7:0] p77_array_index_1091285;
  reg [7:0] p77_array_index_1091286;
  reg [7:0] p77_array_index_1091287;
  reg [7:0] p77_res7__401;
  reg [7:0] p77_array_index_1091300;
  reg [7:0] p77_array_index_1091301;
  reg [7:0] p77_array_index_1091302;
  reg [7:0] p77_res7__402;
  reg [7:0] p77_array_index_1091314;
  reg [7:0] p77_array_index_1091315;
  reg [7:0] p77_array_index_1091316;
  reg [7:0] p77_res7__403;
  reg [7:0] p77_array_index_1091329;
  reg [7:0] p77_array_index_1091330;
  reg [7:0] p77_array_index_1091331;
  reg [7:0] p77_res7__404;
  reg [7:0] p77_array_index_1091611;
  reg [7:0] p77_array_index_1091612;
  reg [7:0] p77_array_index_1091613;
  reg [7:0] p77_res7__405;
  reg [7:0] p77_array_index_1091625;
  reg [7:0] p77_array_index_1091626;
  reg [7:0] p77_array_index_1091627;
  reg [7:0] p77_res7__406;
  reg [7:0] p77_array_index_1091637;
  reg [7:0] p77_array_index_1091638;
  reg [7:0] p77_array_index_1091639;
  reg [7:0] p77_res7__407;
  reg [7:0] p77_array_index_1091650;
  reg [7:0] p77_array_index_1091651;
  reg [7:0] p77_res7__408;
  reg [7:0] p77_array_index_1091661;
  reg [7:0] p77_array_index_1091662;
  reg [7:0] p77_res7__409;
  reg [7:0] p77_array_index_1091668;
  reg [7:0] p77_array_index_1091669;
  reg [7:0] p77_array_index_1091670;
  reg [7:0] p77_array_index_1091671;
  reg [7:0] p77_array_index_1091672;
  reg [7:0] p77_array_index_1091673;
  reg [7:0] p77_array_index_1091674;
  reg [7:0] p77_array_index_1091675;
  reg [7:0] p77_array_index_1091676;
  reg [7:0] p77_array_index_1091340;
  reg [7:0] p77_array_index_1091341;
  reg [7:0] p77_array_index_1091342;
  reg [7:0] p77_array_index_1091343;
  reg [7:0] p77_array_index_1091344;
  reg [7:0] p77_array_index_1091345;
  reg [7:0] p77_array_index_1091353;
  reg [7:0] p77_array_index_1091354;
  reg [7:0] p77_array_index_1091355;
  reg [7:0] p77_res7__624;
  reg [7:0] p77_array_index_1091370;
  reg [7:0] p77_array_index_1091371;
  reg [7:0] p77_array_index_1091372;
  reg [7:0] p77_res7__625;
  reg [7:0] p77_array_index_1091385;
  reg [7:0] p77_array_index_1091386;
  reg [7:0] p77_array_index_1091387;
  reg [7:0] p77_res7__626;
  reg [7:0] p77_array_index_1091399;
  reg [7:0] p77_array_index_1091400;
  reg [7:0] p77_array_index_1091401;
  reg [7:0] p77_res7__627;
  reg [7:0] p77_array_index_1091414;
  reg [7:0] p77_array_index_1091415;
  reg [7:0] p77_array_index_1091416;
  reg [7:0] p77_res7__628;
  reg [7:0] p77_array_index_1091679;
  reg [7:0] p77_array_index_1091680;
  reg [7:0] p77_array_index_1091681;
  reg [7:0] p77_res7__629;
  reg [7:0] p77_array_index_1091693;
  reg [7:0] p77_array_index_1091694;
  reg [7:0] p77_array_index_1091695;
  reg [7:0] p77_res7__630;
  reg [7:0] p77_array_index_1091705;
  reg [7:0] p77_array_index_1091706;
  reg [7:0] p77_array_index_1091707;
  reg [7:0] p77_res7__631;
  reg [7:0] p77_array_index_1091718;
  reg [7:0] p77_array_index_1091719;
  reg [7:0] p77_res7__632;
  reg [7:0] p77_array_index_1091729;
  reg [7:0] p77_array_index_1091730;
  reg [7:0] p77_res7__633;
  reg [7:0] p78_arr[256];
  reg [7:0] p78_literal_1076345[256];
  reg [7:0] p78_literal_1076347[256];
  reg [7:0] p78_literal_1076349[256];
  reg [7:0] p78_literal_1076351[256];
  reg [7:0] p78_literal_1076353[256];
  reg [7:0] p78_literal_1076355[256];
  reg [7:0] p78_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p77_k6 <= p76_k6;
    p77_xor_1091121 <= p76_xor_1091121;
    p77_array_index_1091252 <= p76_array_index_1091252;
    p77_array_index_1091253 <= p76_array_index_1091253;
    p77_array_index_1091254 <= p76_array_index_1091254;
    p77_array_index_1091255 <= p76_array_index_1091255;
    p77_array_index_1091256 <= p76_array_index_1091256;
    p77_array_index_1091257 <= p76_array_index_1091257;
    p77_array_index_1091268 <= p76_array_index_1091268;
    p77_array_index_1091269 <= p76_array_index_1091269;
    p77_array_index_1091270 <= p76_array_index_1091270;
    p77_res7__400 <= p76_res7__400;
    p77_array_index_1091285 <= p76_array_index_1091285;
    p77_array_index_1091286 <= p76_array_index_1091286;
    p77_array_index_1091287 <= p76_array_index_1091287;
    p77_res7__401 <= p76_res7__401;
    p77_array_index_1091300 <= p76_array_index_1091300;
    p77_array_index_1091301 <= p76_array_index_1091301;
    p77_array_index_1091302 <= p76_array_index_1091302;
    p77_res7__402 <= p76_res7__402;
    p77_array_index_1091314 <= p76_array_index_1091314;
    p77_array_index_1091315 <= p76_array_index_1091315;
    p77_array_index_1091316 <= p76_array_index_1091316;
    p77_res7__403 <= p76_res7__403;
    p77_array_index_1091329 <= p76_array_index_1091329;
    p77_array_index_1091330 <= p76_array_index_1091330;
    p77_array_index_1091331 <= p76_array_index_1091331;
    p77_res7__404 <= p76_res7__404;
    p77_array_index_1091611 <= p77_array_index_1091611_comb;
    p77_array_index_1091612 <= p77_array_index_1091612_comb;
    p77_array_index_1091613 <= p77_array_index_1091613_comb;
    p77_res7__405 <= p77_res7__405_comb;
    p77_array_index_1091625 <= p77_array_index_1091625_comb;
    p77_array_index_1091626 <= p77_array_index_1091626_comb;
    p77_array_index_1091627 <= p77_array_index_1091627_comb;
    p77_res7__406 <= p77_res7__406_comb;
    p77_array_index_1091637 <= p77_array_index_1091637_comb;
    p77_array_index_1091638 <= p77_array_index_1091638_comb;
    p77_array_index_1091639 <= p77_array_index_1091639_comb;
    p77_res7__407 <= p77_res7__407_comb;
    p77_array_index_1091650 <= p77_array_index_1091650_comb;
    p77_array_index_1091651 <= p77_array_index_1091651_comb;
    p77_res7__408 <= p77_res7__408_comb;
    p77_array_index_1091661 <= p77_array_index_1091661_comb;
    p77_array_index_1091662 <= p77_array_index_1091662_comb;
    p77_res7__409 <= p77_res7__409_comb;
    p77_array_index_1091668 <= p77_array_index_1091668_comb;
    p77_array_index_1091669 <= p77_array_index_1091669_comb;
    p77_array_index_1091670 <= p77_array_index_1091670_comb;
    p77_array_index_1091671 <= p77_array_index_1091671_comb;
    p77_array_index_1091672 <= p77_array_index_1091672_comb;
    p77_array_index_1091673 <= p77_array_index_1091673_comb;
    p77_array_index_1091674 <= p77_array_index_1091674_comb;
    p77_array_index_1091675 <= p77_array_index_1091675_comb;
    p77_array_index_1091676 <= p77_array_index_1091676_comb;
    p77_array_index_1091340 <= p76_array_index_1091340;
    p77_array_index_1091341 <= p76_array_index_1091341;
    p77_array_index_1091342 <= p76_array_index_1091342;
    p77_array_index_1091343 <= p76_array_index_1091343;
    p77_array_index_1091344 <= p76_array_index_1091344;
    p77_array_index_1091345 <= p76_array_index_1091345;
    p77_array_index_1091353 <= p76_array_index_1091353;
    p77_array_index_1091354 <= p76_array_index_1091354;
    p77_array_index_1091355 <= p76_array_index_1091355;
    p77_res7__624 <= p76_res7__624;
    p77_array_index_1091370 <= p76_array_index_1091370;
    p77_array_index_1091371 <= p76_array_index_1091371;
    p77_array_index_1091372 <= p76_array_index_1091372;
    p77_res7__625 <= p76_res7__625;
    p77_array_index_1091385 <= p76_array_index_1091385;
    p77_array_index_1091386 <= p76_array_index_1091386;
    p77_array_index_1091387 <= p76_array_index_1091387;
    p77_res7__626 <= p76_res7__626;
    p77_array_index_1091399 <= p76_array_index_1091399;
    p77_array_index_1091400 <= p76_array_index_1091400;
    p77_array_index_1091401 <= p76_array_index_1091401;
    p77_res7__627 <= p76_res7__627;
    p77_array_index_1091414 <= p76_array_index_1091414;
    p77_array_index_1091415 <= p76_array_index_1091415;
    p77_array_index_1091416 <= p76_array_index_1091416;
    p77_res7__628 <= p76_res7__628;
    p77_array_index_1091679 <= p77_array_index_1091679_comb;
    p77_array_index_1091680 <= p77_array_index_1091680_comb;
    p77_array_index_1091681 <= p77_array_index_1091681_comb;
    p77_res7__629 <= p77_res7__629_comb;
    p77_array_index_1091693 <= p77_array_index_1091693_comb;
    p77_array_index_1091694 <= p77_array_index_1091694_comb;
    p77_array_index_1091695 <= p77_array_index_1091695_comb;
    p77_res7__630 <= p77_res7__630_comb;
    p77_array_index_1091705 <= p77_array_index_1091705_comb;
    p77_array_index_1091706 <= p77_array_index_1091706_comb;
    p77_array_index_1091707 <= p77_array_index_1091707_comb;
    p77_res7__631 <= p77_res7__631_comb;
    p77_array_index_1091718 <= p77_array_index_1091718_comb;
    p77_array_index_1091719 <= p77_array_index_1091719_comb;
    p77_res7__632 <= p77_res7__632_comb;
    p77_array_index_1091729 <= p77_array_index_1091729_comb;
    p77_array_index_1091730 <= p77_array_index_1091730_comb;
    p77_res7__633 <= p77_res7__633_comb;
    p78_arr <= p77_arr;
    p78_literal_1076345 <= p77_literal_1076345;
    p78_literal_1076347 <= p77_literal_1076347;
    p78_literal_1076349 <= p77_literal_1076349;
    p78_literal_1076351 <= p77_literal_1076351;
    p78_literal_1076353 <= p77_literal_1076353;
    p78_literal_1076355 <= p77_literal_1076355;
    p78_literal_1076358 <= p77_literal_1076358;
  end

  // ===== Pipe stage 78:
  wire [7:0] p78_res7__410_comb;
  wire [7:0] p78_array_index_1091956_comb;
  wire [7:0] p78_res7__411_comb;
  wire [7:0] p78_array_index_1092002_comb;
  wire [7:0] p78_res7__412_comb;
  wire [7:0] p78_res7__634_comb;
  wire [7:0] p78_array_index_1092012_comb;
  wire [7:0] p78_res7__413_comb;
  wire [7:0] p78_res7__635_comb;
  wire [7:0] p78_res7__414_comb;
  wire [7:0] p78_res7__636_comb;
  wire [7:0] p78_res7__415_comb;
  wire [7:0] p78_res7__637_comb;
  wire [127:0] p78_res__25_comb;
  wire [127:0] p78_xor_1091996_comb;
  wire [7:0] p78_res7__638_comb;
  assign p78_res7__410_comb = p77_array_index_1091668 ^ p77_array_index_1091669 ^ p77_array_index_1091670 ^ p77_array_index_1091671 ^ p77_array_index_1091672 ^ p77_array_index_1091673 ^ p77_res7__403 ^ p77_array_index_1091674 ^ p77_res7__401 ^ p77_array_index_1091627 ^ p77_array_index_1091331 ^ p77_array_index_1091302 ^ p77_array_index_1091270 ^ p77_array_index_1091675 ^ p77_array_index_1091676 ^ p77_array_index_1091257;
  assign p78_array_index_1091956_comb = p77_literal_1076355[p77_res7__405];
  assign p78_res7__411_comb = p77_literal_1076345[p78_res7__410_comb] ^ p77_literal_1076347[p77_res7__409] ^ p77_literal_1076349[p77_res7__408] ^ p77_literal_1076351[p77_res7__407] ^ p77_literal_1076353[p77_res7__406] ^ p78_array_index_1091956_comb ^ p77_res7__404 ^ p77_literal_1076358[p77_res7__403] ^ p77_res7__402 ^ p77_array_index_1091639 ^ p77_array_index_1091613 ^ p77_array_index_1091316 ^ p77_array_index_1091287 ^ p77_literal_1076347[p77_array_index_1091254] ^ p77_literal_1076345[p77_array_index_1091255] ^ p77_array_index_1091256;
  assign p78_array_index_1092002_comb = p77_literal_1076355[p77_res7__628];
  assign p78_res7__412_comb = p77_literal_1076345[p78_res7__411_comb] ^ p77_literal_1076347[p78_res7__410_comb] ^ p77_literal_1076349[p77_res7__409] ^ p77_literal_1076351[p77_res7__408] ^ p77_literal_1076353[p77_res7__407] ^ p77_literal_1076355[p77_res7__406] ^ p77_res7__405 ^ p77_literal_1076358[p77_res7__404] ^ p77_res7__403 ^ p77_array_index_1091651 ^ p77_array_index_1091626 ^ p77_array_index_1091330 ^ p77_array_index_1091301 ^ p77_array_index_1091269 ^ p77_literal_1076345[p77_array_index_1091254] ^ p77_array_index_1091255;
  assign p78_res7__634_comb = p77_literal_1076345[p77_res7__633] ^ p77_literal_1076347[p77_res7__632] ^ p77_literal_1076349[p77_res7__631] ^ p77_literal_1076351[p77_res7__630] ^ p77_literal_1076353[p77_res7__629] ^ p78_array_index_1092002_comb ^ p77_res7__627 ^ p77_literal_1076358[p77_res7__626] ^ p77_res7__625 ^ p77_array_index_1091695 ^ p77_array_index_1091416 ^ p77_array_index_1091387 ^ p77_array_index_1091355 ^ p77_literal_1076347[p77_array_index_1091343] ^ p77_literal_1076345[p77_array_index_1091344] ^ p77_array_index_1091345;
  assign p78_array_index_1092012_comb = p77_literal_1076355[p77_res7__629];
  assign p78_res7__413_comb = p77_literal_1076345[p78_res7__412_comb] ^ p77_literal_1076347[p78_res7__411_comb] ^ p77_literal_1076349[p78_res7__410_comb] ^ p77_literal_1076351[p77_res7__409] ^ p77_literal_1076353[p77_res7__408] ^ p77_literal_1076355[p77_res7__407] ^ p77_res7__406 ^ p77_literal_1076358[p77_res7__405] ^ p77_res7__404 ^ p77_array_index_1091662 ^ p77_array_index_1091638 ^ p77_array_index_1091612 ^ p77_array_index_1091315 ^ p77_array_index_1091286 ^ p77_literal_1076345[p77_array_index_1091253] ^ p77_array_index_1091254;
  assign p78_res7__635_comb = p77_literal_1076345[p78_res7__634_comb] ^ p77_literal_1076347[p77_res7__633] ^ p77_literal_1076349[p77_res7__632] ^ p77_literal_1076351[p77_res7__631] ^ p77_literal_1076353[p77_res7__630] ^ p78_array_index_1092012_comb ^ p77_res7__628 ^ p77_literal_1076358[p77_res7__627] ^ p77_res7__626 ^ p77_array_index_1091707 ^ p77_array_index_1091681 ^ p77_array_index_1091401 ^ p77_array_index_1091372 ^ p77_literal_1076347[p77_array_index_1091342] ^ p77_literal_1076345[p77_array_index_1091343] ^ p77_array_index_1091344;
  assign p78_res7__414_comb = p77_literal_1076345[p78_res7__413_comb] ^ p77_literal_1076347[p78_res7__412_comb] ^ p77_literal_1076349[p78_res7__411_comb] ^ p77_literal_1076351[p78_res7__410_comb] ^ p77_literal_1076353[p77_res7__409] ^ p77_literal_1076355[p77_res7__408] ^ p77_res7__407 ^ p77_literal_1076358[p77_res7__406] ^ p77_res7__405 ^ p77_array_index_1091673 ^ p77_array_index_1091650 ^ p77_array_index_1091625 ^ p77_array_index_1091329 ^ p77_array_index_1091300 ^ p77_array_index_1091268 ^ p77_array_index_1091253;
  assign p78_res7__636_comb = p77_literal_1076345[p78_res7__635_comb] ^ p77_literal_1076347[p78_res7__634_comb] ^ p77_literal_1076349[p77_res7__633] ^ p77_literal_1076351[p77_res7__632] ^ p77_literal_1076353[p77_res7__631] ^ p77_literal_1076355[p77_res7__630] ^ p77_res7__629 ^ p77_literal_1076358[p77_res7__628] ^ p77_res7__627 ^ p77_array_index_1091719 ^ p77_array_index_1091694 ^ p77_array_index_1091415 ^ p77_array_index_1091386 ^ p77_array_index_1091354 ^ p77_literal_1076345[p77_array_index_1091342] ^ p77_array_index_1091343;
  assign p78_res7__415_comb = p77_literal_1076345[p78_res7__414_comb] ^ p77_literal_1076347[p78_res7__413_comb] ^ p77_literal_1076349[p78_res7__412_comb] ^ p77_literal_1076351[p78_res7__411_comb] ^ p77_literal_1076353[p78_res7__410_comb] ^ p77_literal_1076355[p77_res7__409] ^ p77_res7__408 ^ p77_literal_1076358[p77_res7__407] ^ p77_res7__406 ^ p78_array_index_1091956_comb ^ p77_array_index_1091661 ^ p77_array_index_1091637 ^ p77_array_index_1091611 ^ p77_array_index_1091314 ^ p77_array_index_1091285 ^ p77_array_index_1091252;
  assign p78_res7__637_comb = p77_literal_1076345[p78_res7__636_comb] ^ p77_literal_1076347[p78_res7__635_comb] ^ p77_literal_1076349[p78_res7__634_comb] ^ p77_literal_1076351[p77_res7__633] ^ p77_literal_1076353[p77_res7__632] ^ p77_literal_1076355[p77_res7__631] ^ p77_res7__630 ^ p77_literal_1076358[p77_res7__629] ^ p77_res7__628 ^ p77_array_index_1091730 ^ p77_array_index_1091706 ^ p77_array_index_1091680 ^ p77_array_index_1091400 ^ p77_array_index_1091371 ^ p77_literal_1076345[p77_array_index_1091341] ^ p77_array_index_1091342;
  assign p78_res__25_comb = {p78_res7__415_comb, p78_res7__414_comb, p78_res7__413_comb, p78_res7__412_comb, p78_res7__411_comb, p78_res7__410_comb, p77_res7__409, p77_res7__408, p77_res7__407, p77_res7__406, p77_res7__405, p77_res7__404, p77_res7__403, p77_res7__402, p77_res7__401, p77_res7__400};
  assign p78_xor_1091996_comb = p78_res__25_comb ^ p77_k6;
  assign p78_res7__638_comb = p77_literal_1076345[p78_res7__637_comb] ^ p77_literal_1076347[p78_res7__636_comb] ^ p77_literal_1076349[p78_res7__635_comb] ^ p77_literal_1076351[p78_res7__634_comb] ^ p77_literal_1076353[p77_res7__633] ^ p77_literal_1076355[p77_res7__632] ^ p77_res7__631 ^ p77_literal_1076358[p77_res7__630] ^ p77_res7__629 ^ p78_array_index_1092002_comb ^ p77_array_index_1091718 ^ p77_array_index_1091693 ^ p77_array_index_1091414 ^ p77_array_index_1091385 ^ p77_array_index_1091353 ^ p77_array_index_1091341;

  // Registers for pipe stage 78:
  reg [127:0] p78_xor_1091121;
  reg [127:0] p78_xor_1091996;
  reg [7:0] p78_array_index_1091340;
  reg [7:0] p78_res7__624;
  reg [7:0] p78_array_index_1091370;
  reg [7:0] p78_res7__625;
  reg [7:0] p78_res7__626;
  reg [7:0] p78_array_index_1091399;
  reg [7:0] p78_res7__627;
  reg [7:0] p78_res7__628;
  reg [7:0] p78_array_index_1091679;
  reg [7:0] p78_res7__629;
  reg [7:0] p78_res7__630;
  reg [7:0] p78_array_index_1091705;
  reg [7:0] p78_res7__631;
  reg [7:0] p78_res7__632;
  reg [7:0] p78_array_index_1091729;
  reg [7:0] p78_res7__633;
  reg [7:0] p78_res7__634;
  reg [7:0] p78_array_index_1092012;
  reg [7:0] p78_res7__635;
  reg [7:0] p78_res7__636;
  reg [7:0] p78_res7__637;
  reg [7:0] p78_res7__638;
  reg [7:0] p79_arr[256];
  reg [7:0] p79_literal_1076345[256];
  reg [7:0] p79_literal_1076347[256];
  reg [7:0] p79_literal_1076349[256];
  reg [7:0] p79_literal_1076351[256];
  reg [7:0] p79_literal_1076353[256];
  reg [7:0] p79_literal_1076355[256];
  reg [7:0] p79_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p78_xor_1091121 <= p77_xor_1091121;
    p78_xor_1091996 <= p78_xor_1091996_comb;
    p78_array_index_1091340 <= p77_array_index_1091340;
    p78_res7__624 <= p77_res7__624;
    p78_array_index_1091370 <= p77_array_index_1091370;
    p78_res7__625 <= p77_res7__625;
    p78_res7__626 <= p77_res7__626;
    p78_array_index_1091399 <= p77_array_index_1091399;
    p78_res7__627 <= p77_res7__627;
    p78_res7__628 <= p77_res7__628;
    p78_array_index_1091679 <= p77_array_index_1091679;
    p78_res7__629 <= p77_res7__629;
    p78_res7__630 <= p77_res7__630;
    p78_array_index_1091705 <= p77_array_index_1091705;
    p78_res7__631 <= p77_res7__631;
    p78_res7__632 <= p77_res7__632;
    p78_array_index_1091729 <= p77_array_index_1091729;
    p78_res7__633 <= p77_res7__633;
    p78_res7__634 <= p78_res7__634_comb;
    p78_array_index_1092012 <= p78_array_index_1092012_comb;
    p78_res7__635 <= p78_res7__635_comb;
    p78_res7__636 <= p78_res7__636_comb;
    p78_res7__637 <= p78_res7__637_comb;
    p78_res7__638 <= p78_res7__638_comb;
    p79_arr <= p78_arr;
    p79_literal_1076345 <= p78_literal_1076345;
    p79_literal_1076347 <= p78_literal_1076347;
    p79_literal_1076349 <= p78_literal_1076349;
    p79_literal_1076351 <= p78_literal_1076351;
    p79_literal_1076353 <= p78_literal_1076353;
    p79_literal_1076355 <= p78_literal_1076355;
    p79_literal_1076358 <= p78_literal_1076358;
  end

  // ===== Pipe stage 79:
  wire [127:0] p79_addedKey__67_comb;
  wire [7:0] p79_array_index_1092122_comb;
  wire [7:0] p79_array_index_1092123_comb;
  wire [7:0] p79_array_index_1092124_comb;
  wire [7:0] p79_array_index_1092125_comb;
  wire [7:0] p79_array_index_1092126_comb;
  wire [7:0] p79_array_index_1092127_comb;
  wire [7:0] p79_array_index_1092129_comb;
  wire [7:0] p79_array_index_1092131_comb;
  wire [7:0] p79_array_index_1092132_comb;
  wire [7:0] p79_array_index_1092133_comb;
  wire [7:0] p79_array_index_1092134_comb;
  wire [7:0] p79_array_index_1092135_comb;
  wire [7:0] p79_array_index_1092136_comb;
  wire [7:0] p79_array_index_1092138_comb;
  wire [7:0] p79_array_index_1092139_comb;
  wire [7:0] p79_array_index_1092140_comb;
  wire [7:0] p79_array_index_1092141_comb;
  wire [7:0] p79_array_index_1092142_comb;
  wire [7:0] p79_array_index_1092143_comb;
  wire [7:0] p79_array_index_1092144_comb;
  wire [7:0] p79_array_index_1092146_comb;
  wire [7:0] p79_res7__416_comb;
  wire [7:0] p79_array_index_1092155_comb;
  wire [7:0] p79_array_index_1092156_comb;
  wire [7:0] p79_array_index_1092157_comb;
  wire [7:0] p79_array_index_1092158_comb;
  wire [7:0] p79_array_index_1092159_comb;
  wire [7:0] p79_array_index_1092160_comb;
  wire [7:0] p79_res7__417_comb;
  wire [7:0] p79_array_index_1092170_comb;
  wire [7:0] p79_array_index_1092171_comb;
  wire [7:0] p79_array_index_1092172_comb;
  wire [7:0] p79_array_index_1092173_comb;
  wire [7:0] p79_array_index_1092174_comb;
  wire [7:0] p79_res7__418_comb;
  wire [7:0] p79_array_index_1092184_comb;
  wire [7:0] p79_array_index_1092185_comb;
  wire [7:0] p79_array_index_1092186_comb;
  wire [7:0] p79_array_index_1092187_comb;
  wire [7:0] p79_array_index_1092188_comb;
  wire [7:0] p79_res7__419_comb;
  wire [7:0] p79_array_index_1092199_comb;
  wire [7:0] p79_array_index_1092200_comb;
  wire [7:0] p79_array_index_1092201_comb;
  wire [7:0] p79_array_index_1092202_comb;
  wire [7:0] p79_res7__639_comb;
  wire [7:0] p79_res7__420_comb;
  wire [127:0] p79_res__39_comb;
  assign p79_addedKey__67_comb = p78_xor_1091996 ^ 128'h6bce_c0ac_5dd7_7453_d3a7_2473_cd72_011b;
  assign p79_array_index_1092122_comb = p78_arr[p79_addedKey__67_comb[127:120]];
  assign p79_array_index_1092123_comb = p78_arr[p79_addedKey__67_comb[119:112]];
  assign p79_array_index_1092124_comb = p78_arr[p79_addedKey__67_comb[111:104]];
  assign p79_array_index_1092125_comb = p78_arr[p79_addedKey__67_comb[103:96]];
  assign p79_array_index_1092126_comb = p78_arr[p79_addedKey__67_comb[95:88]];
  assign p79_array_index_1092127_comb = p78_arr[p79_addedKey__67_comb[87:80]];
  assign p79_array_index_1092129_comb = p78_arr[p79_addedKey__67_comb[71:64]];
  assign p79_array_index_1092131_comb = p78_arr[p79_addedKey__67_comb[55:48]];
  assign p79_array_index_1092132_comb = p78_arr[p79_addedKey__67_comb[47:40]];
  assign p79_array_index_1092133_comb = p78_arr[p79_addedKey__67_comb[39:32]];
  assign p79_array_index_1092134_comb = p78_arr[p79_addedKey__67_comb[31:24]];
  assign p79_array_index_1092135_comb = p78_arr[p79_addedKey__67_comb[23:16]];
  assign p79_array_index_1092136_comb = p78_arr[p79_addedKey__67_comb[15:8]];
  assign p79_array_index_1092138_comb = p78_literal_1076345[p79_array_index_1092122_comb];
  assign p79_array_index_1092139_comb = p78_literal_1076347[p79_array_index_1092123_comb];
  assign p79_array_index_1092140_comb = p78_literal_1076349[p79_array_index_1092124_comb];
  assign p79_array_index_1092141_comb = p78_literal_1076351[p79_array_index_1092125_comb];
  assign p79_array_index_1092142_comb = p78_literal_1076353[p79_array_index_1092126_comb];
  assign p79_array_index_1092143_comb = p78_literal_1076355[p79_array_index_1092127_comb];
  assign p79_array_index_1092144_comb = p78_arr[p79_addedKey__67_comb[79:72]];
  assign p79_array_index_1092146_comb = p78_arr[p79_addedKey__67_comb[63:56]];
  assign p79_res7__416_comb = p79_array_index_1092138_comb ^ p79_array_index_1092139_comb ^ p79_array_index_1092140_comb ^ p79_array_index_1092141_comb ^ p79_array_index_1092142_comb ^ p79_array_index_1092143_comb ^ p79_array_index_1092144_comb ^ p78_literal_1076358[p79_array_index_1092129_comb] ^ p79_array_index_1092146_comb ^ p78_literal_1076355[p79_array_index_1092131_comb] ^ p78_literal_1076353[p79_array_index_1092132_comb] ^ p78_literal_1076351[p79_array_index_1092133_comb] ^ p78_literal_1076349[p79_array_index_1092134_comb] ^ p78_literal_1076347[p79_array_index_1092135_comb] ^ p78_literal_1076345[p79_array_index_1092136_comb] ^ p78_arr[p79_addedKey__67_comb[7:0]];
  assign p79_array_index_1092155_comb = p78_literal_1076345[p79_res7__416_comb];
  assign p79_array_index_1092156_comb = p78_literal_1076347[p79_array_index_1092122_comb];
  assign p79_array_index_1092157_comb = p78_literal_1076349[p79_array_index_1092123_comb];
  assign p79_array_index_1092158_comb = p78_literal_1076351[p79_array_index_1092124_comb];
  assign p79_array_index_1092159_comb = p78_literal_1076353[p79_array_index_1092125_comb];
  assign p79_array_index_1092160_comb = p78_literal_1076355[p79_array_index_1092126_comb];
  assign p79_res7__417_comb = p79_array_index_1092155_comb ^ p79_array_index_1092156_comb ^ p79_array_index_1092157_comb ^ p79_array_index_1092158_comb ^ p79_array_index_1092159_comb ^ p79_array_index_1092160_comb ^ p79_array_index_1092127_comb ^ p78_literal_1076358[p79_array_index_1092144_comb] ^ p79_array_index_1092129_comb ^ p78_literal_1076355[p79_array_index_1092146_comb] ^ p78_literal_1076353[p79_array_index_1092131_comb] ^ p78_literal_1076351[p79_array_index_1092132_comb] ^ p78_literal_1076349[p79_array_index_1092133_comb] ^ p78_literal_1076347[p79_array_index_1092134_comb] ^ p78_literal_1076345[p79_array_index_1092135_comb] ^ p79_array_index_1092136_comb;
  assign p79_array_index_1092170_comb = p78_literal_1076347[p79_res7__416_comb];
  assign p79_array_index_1092171_comb = p78_literal_1076349[p79_array_index_1092122_comb];
  assign p79_array_index_1092172_comb = p78_literal_1076351[p79_array_index_1092123_comb];
  assign p79_array_index_1092173_comb = p78_literal_1076353[p79_array_index_1092124_comb];
  assign p79_array_index_1092174_comb = p78_literal_1076355[p79_array_index_1092125_comb];
  assign p79_res7__418_comb = p78_literal_1076345[p79_res7__417_comb] ^ p79_array_index_1092170_comb ^ p79_array_index_1092171_comb ^ p79_array_index_1092172_comb ^ p79_array_index_1092173_comb ^ p79_array_index_1092174_comb ^ p79_array_index_1092126_comb ^ p78_literal_1076358[p79_array_index_1092127_comb] ^ p79_array_index_1092144_comb ^ p78_literal_1076355[p79_array_index_1092129_comb] ^ p78_literal_1076353[p79_array_index_1092146_comb] ^ p78_literal_1076351[p79_array_index_1092131_comb] ^ p78_literal_1076349[p79_array_index_1092132_comb] ^ p78_literal_1076347[p79_array_index_1092133_comb] ^ p78_literal_1076345[p79_array_index_1092134_comb] ^ p79_array_index_1092135_comb;
  assign p79_array_index_1092184_comb = p78_literal_1076347[p79_res7__417_comb];
  assign p79_array_index_1092185_comb = p78_literal_1076349[p79_res7__416_comb];
  assign p79_array_index_1092186_comb = p78_literal_1076351[p79_array_index_1092122_comb];
  assign p79_array_index_1092187_comb = p78_literal_1076353[p79_array_index_1092123_comb];
  assign p79_array_index_1092188_comb = p78_literal_1076355[p79_array_index_1092124_comb];
  assign p79_res7__419_comb = p78_literal_1076345[p79_res7__418_comb] ^ p79_array_index_1092184_comb ^ p79_array_index_1092185_comb ^ p79_array_index_1092186_comb ^ p79_array_index_1092187_comb ^ p79_array_index_1092188_comb ^ p79_array_index_1092125_comb ^ p78_literal_1076358[p79_array_index_1092126_comb] ^ p79_array_index_1092127_comb ^ p78_literal_1076355[p79_array_index_1092144_comb] ^ p78_literal_1076353[p79_array_index_1092129_comb] ^ p78_literal_1076351[p79_array_index_1092146_comb] ^ p78_literal_1076349[p79_array_index_1092131_comb] ^ p78_literal_1076347[p79_array_index_1092132_comb] ^ p78_literal_1076345[p79_array_index_1092133_comb] ^ p79_array_index_1092134_comb;
  assign p79_array_index_1092199_comb = p78_literal_1076349[p79_res7__417_comb];
  assign p79_array_index_1092200_comb = p78_literal_1076351[p79_res7__416_comb];
  assign p79_array_index_1092201_comb = p78_literal_1076353[p79_array_index_1092122_comb];
  assign p79_array_index_1092202_comb = p78_literal_1076355[p79_array_index_1092123_comb];
  assign p79_res7__639_comb = p78_literal_1076345[p78_res7__638] ^ p78_literal_1076347[p78_res7__637] ^ p78_literal_1076349[p78_res7__636] ^ p78_literal_1076351[p78_res7__635] ^ p78_literal_1076353[p78_res7__634] ^ p78_literal_1076355[p78_res7__633] ^ p78_res7__632 ^ p78_literal_1076358[p78_res7__631] ^ p78_res7__630 ^ p78_array_index_1092012 ^ p78_array_index_1091729 ^ p78_array_index_1091705 ^ p78_array_index_1091679 ^ p78_array_index_1091399 ^ p78_array_index_1091370 ^ p78_array_index_1091340;
  assign p79_res7__420_comb = p78_literal_1076345[p79_res7__419_comb] ^ p78_literal_1076347[p79_res7__418_comb] ^ p79_array_index_1092199_comb ^ p79_array_index_1092200_comb ^ p79_array_index_1092201_comb ^ p79_array_index_1092202_comb ^ p79_array_index_1092124_comb ^ p78_literal_1076358[p79_array_index_1092125_comb] ^ p79_array_index_1092126_comb ^ p79_array_index_1092143_comb ^ p78_literal_1076353[p79_array_index_1092144_comb] ^ p78_literal_1076351[p79_array_index_1092129_comb] ^ p78_literal_1076349[p79_array_index_1092146_comb] ^ p78_literal_1076347[p79_array_index_1092131_comb] ^ p78_literal_1076345[p79_array_index_1092132_comb] ^ p79_array_index_1092133_comb;
  assign p79_res__39_comb = {p79_res7__639_comb, p78_res7__638, p78_res7__637, p78_res7__636, p78_res7__635, p78_res7__634, p78_res7__633, p78_res7__632, p78_res7__631, p78_res7__630, p78_res7__629, p78_res7__628, p78_res7__627, p78_res7__626, p78_res7__625, p78_res7__624};

  // Registers for pipe stage 79:
  reg [127:0] p79_xor_1091121;
  reg [127:0] p79_xor_1091996;
  reg [7:0] p79_array_index_1092122;
  reg [7:0] p79_array_index_1092123;
  reg [7:0] p79_array_index_1092124;
  reg [7:0] p79_array_index_1092125;
  reg [7:0] p79_array_index_1092126;
  reg [7:0] p79_array_index_1092127;
  reg [7:0] p79_array_index_1092129;
  reg [7:0] p79_array_index_1092131;
  reg [7:0] p79_array_index_1092132;
  reg [7:0] p79_array_index_1092138;
  reg [7:0] p79_array_index_1092139;
  reg [7:0] p79_array_index_1092140;
  reg [7:0] p79_array_index_1092141;
  reg [7:0] p79_array_index_1092142;
  reg [7:0] p79_array_index_1092144;
  reg [7:0] p79_array_index_1092146;
  reg [7:0] p79_res7__416;
  reg [7:0] p79_array_index_1092155;
  reg [7:0] p79_array_index_1092156;
  reg [7:0] p79_array_index_1092157;
  reg [7:0] p79_array_index_1092158;
  reg [7:0] p79_array_index_1092159;
  reg [7:0] p79_array_index_1092160;
  reg [7:0] p79_res7__417;
  reg [7:0] p79_array_index_1092170;
  reg [7:0] p79_array_index_1092171;
  reg [7:0] p79_array_index_1092172;
  reg [7:0] p79_array_index_1092173;
  reg [7:0] p79_array_index_1092174;
  reg [7:0] p79_res7__418;
  reg [7:0] p79_array_index_1092184;
  reg [7:0] p79_array_index_1092185;
  reg [7:0] p79_array_index_1092186;
  reg [7:0] p79_array_index_1092187;
  reg [7:0] p79_array_index_1092188;
  reg [7:0] p79_res7__419;
  reg [7:0] p79_array_index_1092199;
  reg [7:0] p79_array_index_1092200;
  reg [7:0] p79_array_index_1092201;
  reg [7:0] p79_array_index_1092202;
  reg [7:0] p79_res7__420;
  reg [127:0] p79_res__39;
  reg [7:0] p80_arr[256];
  reg [7:0] p80_literal_1076345[256];
  reg [7:0] p80_literal_1076347[256];
  reg [7:0] p80_literal_1076349[256];
  reg [7:0] p80_literal_1076351[256];
  reg [7:0] p80_literal_1076353[256];
  reg [7:0] p80_literal_1076355[256];
  reg [7:0] p80_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p79_xor_1091121 <= p78_xor_1091121;
    p79_xor_1091996 <= p78_xor_1091996;
    p79_array_index_1092122 <= p79_array_index_1092122_comb;
    p79_array_index_1092123 <= p79_array_index_1092123_comb;
    p79_array_index_1092124 <= p79_array_index_1092124_comb;
    p79_array_index_1092125 <= p79_array_index_1092125_comb;
    p79_array_index_1092126 <= p79_array_index_1092126_comb;
    p79_array_index_1092127 <= p79_array_index_1092127_comb;
    p79_array_index_1092129 <= p79_array_index_1092129_comb;
    p79_array_index_1092131 <= p79_array_index_1092131_comb;
    p79_array_index_1092132 <= p79_array_index_1092132_comb;
    p79_array_index_1092138 <= p79_array_index_1092138_comb;
    p79_array_index_1092139 <= p79_array_index_1092139_comb;
    p79_array_index_1092140 <= p79_array_index_1092140_comb;
    p79_array_index_1092141 <= p79_array_index_1092141_comb;
    p79_array_index_1092142 <= p79_array_index_1092142_comb;
    p79_array_index_1092144 <= p79_array_index_1092144_comb;
    p79_array_index_1092146 <= p79_array_index_1092146_comb;
    p79_res7__416 <= p79_res7__416_comb;
    p79_array_index_1092155 <= p79_array_index_1092155_comb;
    p79_array_index_1092156 <= p79_array_index_1092156_comb;
    p79_array_index_1092157 <= p79_array_index_1092157_comb;
    p79_array_index_1092158 <= p79_array_index_1092158_comb;
    p79_array_index_1092159 <= p79_array_index_1092159_comb;
    p79_array_index_1092160 <= p79_array_index_1092160_comb;
    p79_res7__417 <= p79_res7__417_comb;
    p79_array_index_1092170 <= p79_array_index_1092170_comb;
    p79_array_index_1092171 <= p79_array_index_1092171_comb;
    p79_array_index_1092172 <= p79_array_index_1092172_comb;
    p79_array_index_1092173 <= p79_array_index_1092173_comb;
    p79_array_index_1092174 <= p79_array_index_1092174_comb;
    p79_res7__418 <= p79_res7__418_comb;
    p79_array_index_1092184 <= p79_array_index_1092184_comb;
    p79_array_index_1092185 <= p79_array_index_1092185_comb;
    p79_array_index_1092186 <= p79_array_index_1092186_comb;
    p79_array_index_1092187 <= p79_array_index_1092187_comb;
    p79_array_index_1092188 <= p79_array_index_1092188_comb;
    p79_res7__419 <= p79_res7__419_comb;
    p79_array_index_1092199 <= p79_array_index_1092199_comb;
    p79_array_index_1092200 <= p79_array_index_1092200_comb;
    p79_array_index_1092201 <= p79_array_index_1092201_comb;
    p79_array_index_1092202 <= p79_array_index_1092202_comb;
    p79_res7__420 <= p79_res7__420_comb;
    p79_res__39 <= p79_res__39_comb;
    p80_arr <= p79_arr;
    p80_literal_1076345 <= p79_literal_1076345;
    p80_literal_1076347 <= p79_literal_1076347;
    p80_literal_1076349 <= p79_literal_1076349;
    p80_literal_1076351 <= p79_literal_1076351;
    p80_literal_1076353 <= p79_literal_1076353;
    p80_literal_1076355 <= p79_literal_1076355;
    p80_literal_1076358 <= p79_literal_1076358;
  end

  // ===== Pipe stage 80:
  wire [7:0] p80_array_index_1092325_comb;
  wire [7:0] p80_array_index_1092326_comb;
  wire [7:0] p80_array_index_1092327_comb;
  wire [7:0] p80_array_index_1092328_comb;
  wire [7:0] p80_res7__421_comb;
  wire [7:0] p80_array_index_1092339_comb;
  wire [7:0] p80_array_index_1092340_comb;
  wire [7:0] p80_array_index_1092341_comb;
  wire [7:0] p80_res7__422_comb;
  wire [7:0] p80_array_index_1092351_comb;
  wire [7:0] p80_array_index_1092352_comb;
  wire [7:0] p80_array_index_1092353_comb;
  wire [7:0] p80_res7__423_comb;
  wire [7:0] p80_array_index_1092364_comb;
  wire [7:0] p80_array_index_1092365_comb;
  wire [7:0] p80_res7__424_comb;
  wire [7:0] p80_array_index_1092375_comb;
  wire [7:0] p80_array_index_1092376_comb;
  wire [7:0] p80_res7__425_comb;
  wire [7:0] p80_array_index_1092382_comb;
  wire [7:0] p80_array_index_1092383_comb;
  wire [7:0] p80_array_index_1092384_comb;
  wire [7:0] p80_array_index_1092385_comb;
  wire [7:0] p80_array_index_1092386_comb;
  wire [7:0] p80_array_index_1092387_comb;
  wire [7:0] p80_array_index_1092388_comb;
  wire [7:0] p80_array_index_1092389_comb;
  wire [7:0] p80_array_index_1092390_comb;
  assign p80_array_index_1092325_comb = p79_literal_1076349[p79_res7__418];
  assign p80_array_index_1092326_comb = p79_literal_1076351[p79_res7__417];
  assign p80_array_index_1092327_comb = p79_literal_1076353[p79_res7__416];
  assign p80_array_index_1092328_comb = p79_literal_1076355[p79_array_index_1092122];
  assign p80_res7__421_comb = p79_literal_1076345[p79_res7__420] ^ p79_literal_1076347[p79_res7__419] ^ p80_array_index_1092325_comb ^ p80_array_index_1092326_comb ^ p80_array_index_1092327_comb ^ p80_array_index_1092328_comb ^ p79_array_index_1092123 ^ p79_literal_1076358[p79_array_index_1092124] ^ p79_array_index_1092125 ^ p79_array_index_1092160 ^ p79_literal_1076353[p79_array_index_1092127] ^ p79_literal_1076351[p79_array_index_1092144] ^ p79_literal_1076349[p79_array_index_1092129] ^ p79_literal_1076347[p79_array_index_1092146] ^ p79_literal_1076345[p79_array_index_1092131] ^ p79_array_index_1092132;
  assign p80_array_index_1092339_comb = p79_literal_1076351[p79_res7__418];
  assign p80_array_index_1092340_comb = p79_literal_1076353[p79_res7__417];
  assign p80_array_index_1092341_comb = p79_literal_1076355[p79_res7__416];
  assign p80_res7__422_comb = p79_literal_1076345[p80_res7__421_comb] ^ p79_literal_1076347[p79_res7__420] ^ p79_literal_1076349[p79_res7__419] ^ p80_array_index_1092339_comb ^ p80_array_index_1092340_comb ^ p80_array_index_1092341_comb ^ p79_array_index_1092122 ^ p79_literal_1076358[p79_array_index_1092123] ^ p79_array_index_1092124 ^ p79_array_index_1092174 ^ p79_array_index_1092142 ^ p79_literal_1076351[p79_array_index_1092127] ^ p79_literal_1076349[p79_array_index_1092144] ^ p79_literal_1076347[p79_array_index_1092129] ^ p79_literal_1076345[p79_array_index_1092146] ^ p79_array_index_1092131;
  assign p80_array_index_1092351_comb = p79_literal_1076351[p79_res7__419];
  assign p80_array_index_1092352_comb = p79_literal_1076353[p79_res7__418];
  assign p80_array_index_1092353_comb = p79_literal_1076355[p79_res7__417];
  assign p80_res7__423_comb = p79_literal_1076345[p80_res7__422_comb] ^ p79_literal_1076347[p80_res7__421_comb] ^ p79_literal_1076349[p79_res7__420] ^ p80_array_index_1092351_comb ^ p80_array_index_1092352_comb ^ p80_array_index_1092353_comb ^ p79_res7__416 ^ p79_literal_1076358[p79_array_index_1092122] ^ p79_array_index_1092123 ^ p79_array_index_1092188 ^ p79_array_index_1092159 ^ p79_literal_1076351[p79_array_index_1092126] ^ p79_literal_1076349[p79_array_index_1092127] ^ p79_literal_1076347[p79_array_index_1092144] ^ p79_literal_1076345[p79_array_index_1092129] ^ p79_array_index_1092146;
  assign p80_array_index_1092364_comb = p79_literal_1076353[p79_res7__419];
  assign p80_array_index_1092365_comb = p79_literal_1076355[p79_res7__418];
  assign p80_res7__424_comb = p79_literal_1076345[p80_res7__423_comb] ^ p79_literal_1076347[p80_res7__422_comb] ^ p79_literal_1076349[p80_res7__421_comb] ^ p79_literal_1076351[p79_res7__420] ^ p80_array_index_1092364_comb ^ p80_array_index_1092365_comb ^ p79_res7__417 ^ p79_literal_1076358[p79_res7__416] ^ p79_array_index_1092122 ^ p79_array_index_1092202 ^ p79_array_index_1092173 ^ p79_array_index_1092141 ^ p79_literal_1076349[p79_array_index_1092126] ^ p79_literal_1076347[p79_array_index_1092127] ^ p79_literal_1076345[p79_array_index_1092144] ^ p79_array_index_1092129;
  assign p80_array_index_1092375_comb = p79_literal_1076353[p79_res7__420];
  assign p80_array_index_1092376_comb = p79_literal_1076355[p79_res7__419];
  assign p80_res7__425_comb = p79_literal_1076345[p80_res7__424_comb] ^ p79_literal_1076347[p80_res7__423_comb] ^ p79_literal_1076349[p80_res7__422_comb] ^ p79_literal_1076351[p80_res7__421_comb] ^ p80_array_index_1092375_comb ^ p80_array_index_1092376_comb ^ p79_res7__418 ^ p79_literal_1076358[p79_res7__417] ^ p79_res7__416 ^ p80_array_index_1092328_comb ^ p79_array_index_1092187 ^ p79_array_index_1092158 ^ p79_literal_1076349[p79_array_index_1092125] ^ p79_literal_1076347[p79_array_index_1092126] ^ p79_literal_1076345[p79_array_index_1092127] ^ p79_array_index_1092144;
  assign p80_array_index_1092382_comb = p79_literal_1076345[p80_res7__425_comb];
  assign p80_array_index_1092383_comb = p79_literal_1076347[p80_res7__424_comb];
  assign p80_array_index_1092384_comb = p79_literal_1076349[p80_res7__423_comb];
  assign p80_array_index_1092385_comb = p79_literal_1076351[p80_res7__422_comb];
  assign p80_array_index_1092386_comb = p79_literal_1076353[p80_res7__421_comb];
  assign p80_array_index_1092387_comb = p79_literal_1076355[p79_res7__420];
  assign p80_array_index_1092388_comb = p79_literal_1076358[p79_res7__418];
  assign p80_array_index_1092389_comb = p79_literal_1076347[p79_array_index_1092125];
  assign p80_array_index_1092390_comb = p79_literal_1076345[p79_array_index_1092126];

  // Registers for pipe stage 80:
  reg [127:0] p80_xor_1091121;
  reg [127:0] p80_xor_1091996;
  reg [7:0] p80_array_index_1092122;
  reg [7:0] p80_array_index_1092123;
  reg [7:0] p80_array_index_1092124;
  reg [7:0] p80_array_index_1092125;
  reg [7:0] p80_array_index_1092126;
  reg [7:0] p80_array_index_1092127;
  reg [7:0] p80_array_index_1092138;
  reg [7:0] p80_array_index_1092139;
  reg [7:0] p80_array_index_1092140;
  reg [7:0] p80_res7__416;
  reg [7:0] p80_array_index_1092155;
  reg [7:0] p80_array_index_1092156;
  reg [7:0] p80_array_index_1092157;
  reg [7:0] p80_res7__417;
  reg [7:0] p80_array_index_1092170;
  reg [7:0] p80_array_index_1092171;
  reg [7:0] p80_array_index_1092172;
  reg [7:0] p80_res7__418;
  reg [7:0] p80_array_index_1092184;
  reg [7:0] p80_array_index_1092185;
  reg [7:0] p80_array_index_1092186;
  reg [7:0] p80_res7__419;
  reg [7:0] p80_array_index_1092199;
  reg [7:0] p80_array_index_1092200;
  reg [7:0] p80_array_index_1092201;
  reg [7:0] p80_res7__420;
  reg [7:0] p80_array_index_1092325;
  reg [7:0] p80_array_index_1092326;
  reg [7:0] p80_array_index_1092327;
  reg [7:0] p80_res7__421;
  reg [7:0] p80_array_index_1092339;
  reg [7:0] p80_array_index_1092340;
  reg [7:0] p80_array_index_1092341;
  reg [7:0] p80_res7__422;
  reg [7:0] p80_array_index_1092351;
  reg [7:0] p80_array_index_1092352;
  reg [7:0] p80_array_index_1092353;
  reg [7:0] p80_res7__423;
  reg [7:0] p80_array_index_1092364;
  reg [7:0] p80_array_index_1092365;
  reg [7:0] p80_res7__424;
  reg [7:0] p80_array_index_1092375;
  reg [7:0] p80_array_index_1092376;
  reg [7:0] p80_res7__425;
  reg [7:0] p80_array_index_1092382;
  reg [7:0] p80_array_index_1092383;
  reg [7:0] p80_array_index_1092384;
  reg [7:0] p80_array_index_1092385;
  reg [7:0] p80_array_index_1092386;
  reg [7:0] p80_array_index_1092387;
  reg [7:0] p80_array_index_1092388;
  reg [7:0] p80_array_index_1092389;
  reg [7:0] p80_array_index_1092390;
  reg [127:0] p80_res__39;
  reg [7:0] p81_arr[256];
  reg [7:0] p81_literal_1076345[256];
  reg [7:0] p81_literal_1076347[256];
  reg [7:0] p81_literal_1076349[256];
  reg [7:0] p81_literal_1076351[256];
  reg [7:0] p81_literal_1076353[256];
  reg [7:0] p81_literal_1076355[256];
  reg [7:0] p81_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p80_xor_1091121 <= p79_xor_1091121;
    p80_xor_1091996 <= p79_xor_1091996;
    p80_array_index_1092122 <= p79_array_index_1092122;
    p80_array_index_1092123 <= p79_array_index_1092123;
    p80_array_index_1092124 <= p79_array_index_1092124;
    p80_array_index_1092125 <= p79_array_index_1092125;
    p80_array_index_1092126 <= p79_array_index_1092126;
    p80_array_index_1092127 <= p79_array_index_1092127;
    p80_array_index_1092138 <= p79_array_index_1092138;
    p80_array_index_1092139 <= p79_array_index_1092139;
    p80_array_index_1092140 <= p79_array_index_1092140;
    p80_res7__416 <= p79_res7__416;
    p80_array_index_1092155 <= p79_array_index_1092155;
    p80_array_index_1092156 <= p79_array_index_1092156;
    p80_array_index_1092157 <= p79_array_index_1092157;
    p80_res7__417 <= p79_res7__417;
    p80_array_index_1092170 <= p79_array_index_1092170;
    p80_array_index_1092171 <= p79_array_index_1092171;
    p80_array_index_1092172 <= p79_array_index_1092172;
    p80_res7__418 <= p79_res7__418;
    p80_array_index_1092184 <= p79_array_index_1092184;
    p80_array_index_1092185 <= p79_array_index_1092185;
    p80_array_index_1092186 <= p79_array_index_1092186;
    p80_res7__419 <= p79_res7__419;
    p80_array_index_1092199 <= p79_array_index_1092199;
    p80_array_index_1092200 <= p79_array_index_1092200;
    p80_array_index_1092201 <= p79_array_index_1092201;
    p80_res7__420 <= p79_res7__420;
    p80_array_index_1092325 <= p80_array_index_1092325_comb;
    p80_array_index_1092326 <= p80_array_index_1092326_comb;
    p80_array_index_1092327 <= p80_array_index_1092327_comb;
    p80_res7__421 <= p80_res7__421_comb;
    p80_array_index_1092339 <= p80_array_index_1092339_comb;
    p80_array_index_1092340 <= p80_array_index_1092340_comb;
    p80_array_index_1092341 <= p80_array_index_1092341_comb;
    p80_res7__422 <= p80_res7__422_comb;
    p80_array_index_1092351 <= p80_array_index_1092351_comb;
    p80_array_index_1092352 <= p80_array_index_1092352_comb;
    p80_array_index_1092353 <= p80_array_index_1092353_comb;
    p80_res7__423 <= p80_res7__423_comb;
    p80_array_index_1092364 <= p80_array_index_1092364_comb;
    p80_array_index_1092365 <= p80_array_index_1092365_comb;
    p80_res7__424 <= p80_res7__424_comb;
    p80_array_index_1092375 <= p80_array_index_1092375_comb;
    p80_array_index_1092376 <= p80_array_index_1092376_comb;
    p80_res7__425 <= p80_res7__425_comb;
    p80_array_index_1092382 <= p80_array_index_1092382_comb;
    p80_array_index_1092383 <= p80_array_index_1092383_comb;
    p80_array_index_1092384 <= p80_array_index_1092384_comb;
    p80_array_index_1092385 <= p80_array_index_1092385_comb;
    p80_array_index_1092386 <= p80_array_index_1092386_comb;
    p80_array_index_1092387 <= p80_array_index_1092387_comb;
    p80_array_index_1092388 <= p80_array_index_1092388_comb;
    p80_array_index_1092389 <= p80_array_index_1092389_comb;
    p80_array_index_1092390 <= p80_array_index_1092390_comb;
    p80_res__39 <= p79_res__39;
    p81_arr <= p80_arr;
    p81_literal_1076345 <= p80_literal_1076345;
    p81_literal_1076347 <= p80_literal_1076347;
    p81_literal_1076349 <= p80_literal_1076349;
    p81_literal_1076351 <= p80_literal_1076351;
    p81_literal_1076353 <= p80_literal_1076353;
    p81_literal_1076355 <= p80_literal_1076355;
    p81_literal_1076358 <= p80_literal_1076358;
  end

  // ===== Pipe stage 81:
  wire [7:0] p81_res7__426_comb;
  wire [7:0] p81_array_index_1092525_comb;
  wire [7:0] p81_res7__427_comb;
  wire [7:0] p81_res7__428_comb;
  wire [7:0] p81_res7__429_comb;
  wire [7:0] p81_res7__430_comb;
  wire [7:0] p81_res7__431_comb;
  wire [127:0] p81_res__26_comb;
  wire [127:0] p81_xor_1092565_comb;
  assign p81_res7__426_comb = p80_array_index_1092382 ^ p80_array_index_1092383 ^ p80_array_index_1092384 ^ p80_array_index_1092385 ^ p80_array_index_1092386 ^ p80_array_index_1092387 ^ p80_res7__419 ^ p80_array_index_1092388 ^ p80_res7__417 ^ p80_array_index_1092341 ^ p80_array_index_1092201 ^ p80_array_index_1092172 ^ p80_array_index_1092140 ^ p80_array_index_1092389 ^ p80_array_index_1092390 ^ p80_array_index_1092127;
  assign p81_array_index_1092525_comb = p80_literal_1076355[p80_res7__421];
  assign p81_res7__427_comb = p80_literal_1076345[p81_res7__426_comb] ^ p80_literal_1076347[p80_res7__425] ^ p80_literal_1076349[p80_res7__424] ^ p80_literal_1076351[p80_res7__423] ^ p80_literal_1076353[p80_res7__422] ^ p81_array_index_1092525_comb ^ p80_res7__420 ^ p80_literal_1076358[p80_res7__419] ^ p80_res7__418 ^ p80_array_index_1092353 ^ p80_array_index_1092327 ^ p80_array_index_1092186 ^ p80_array_index_1092157 ^ p80_literal_1076347[p80_array_index_1092124] ^ p80_literal_1076345[p80_array_index_1092125] ^ p80_array_index_1092126;
  assign p81_res7__428_comb = p80_literal_1076345[p81_res7__427_comb] ^ p80_literal_1076347[p81_res7__426_comb] ^ p80_literal_1076349[p80_res7__425] ^ p80_literal_1076351[p80_res7__424] ^ p80_literal_1076353[p80_res7__423] ^ p80_literal_1076355[p80_res7__422] ^ p80_res7__421 ^ p80_literal_1076358[p80_res7__420] ^ p80_res7__419 ^ p80_array_index_1092365 ^ p80_array_index_1092340 ^ p80_array_index_1092200 ^ p80_array_index_1092171 ^ p80_array_index_1092139 ^ p80_literal_1076345[p80_array_index_1092124] ^ p80_array_index_1092125;
  assign p81_res7__429_comb = p80_literal_1076345[p81_res7__428_comb] ^ p80_literal_1076347[p81_res7__427_comb] ^ p80_literal_1076349[p81_res7__426_comb] ^ p80_literal_1076351[p80_res7__425] ^ p80_literal_1076353[p80_res7__424] ^ p80_literal_1076355[p80_res7__423] ^ p80_res7__422 ^ p80_literal_1076358[p80_res7__421] ^ p80_res7__420 ^ p80_array_index_1092376 ^ p80_array_index_1092352 ^ p80_array_index_1092326 ^ p80_array_index_1092185 ^ p80_array_index_1092156 ^ p80_literal_1076345[p80_array_index_1092123] ^ p80_array_index_1092124;
  assign p81_res7__430_comb = p80_literal_1076345[p81_res7__429_comb] ^ p80_literal_1076347[p81_res7__428_comb] ^ p80_literal_1076349[p81_res7__427_comb] ^ p80_literal_1076351[p81_res7__426_comb] ^ p80_literal_1076353[p80_res7__425] ^ p80_literal_1076355[p80_res7__424] ^ p80_res7__423 ^ p80_literal_1076358[p80_res7__422] ^ p80_res7__421 ^ p80_array_index_1092387 ^ p80_array_index_1092364 ^ p80_array_index_1092339 ^ p80_array_index_1092199 ^ p80_array_index_1092170 ^ p80_array_index_1092138 ^ p80_array_index_1092123;
  assign p81_res7__431_comb = p80_literal_1076345[p81_res7__430_comb] ^ p80_literal_1076347[p81_res7__429_comb] ^ p80_literal_1076349[p81_res7__428_comb] ^ p80_literal_1076351[p81_res7__427_comb] ^ p80_literal_1076353[p81_res7__426_comb] ^ p80_literal_1076355[p80_res7__425] ^ p80_res7__424 ^ p80_literal_1076358[p80_res7__423] ^ p80_res7__422 ^ p81_array_index_1092525_comb ^ p80_array_index_1092375 ^ p80_array_index_1092351 ^ p80_array_index_1092325 ^ p80_array_index_1092184 ^ p80_array_index_1092155 ^ p80_array_index_1092122;
  assign p81_res__26_comb = {p81_res7__431_comb, p81_res7__430_comb, p81_res7__429_comb, p81_res7__428_comb, p81_res7__427_comb, p81_res7__426_comb, p80_res7__425, p80_res7__424, p80_res7__423, p80_res7__422, p80_res7__421, p80_res7__420, p80_res7__419, p80_res7__418, p80_res7__417, p80_res7__416};
  assign p81_xor_1092565_comb = p81_res__26_comb ^ p80_xor_1091121;

  // Registers for pipe stage 81:
  reg [127:0] p81_xor_1091996;
  reg [127:0] p81_xor_1092565;
  reg [127:0] p81_res__39;
  reg [7:0] p82_arr[256];
  reg [7:0] p82_literal_1076345[256];
  reg [7:0] p82_literal_1076347[256];
  reg [7:0] p82_literal_1076349[256];
  reg [7:0] p82_literal_1076351[256];
  reg [7:0] p82_literal_1076353[256];
  reg [7:0] p82_literal_1076355[256];
  reg [7:0] p82_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p81_xor_1091996 <= p80_xor_1091996;
    p81_xor_1092565 <= p81_xor_1092565_comb;
    p81_res__39 <= p80_res__39;
    p82_arr <= p81_arr;
    p82_literal_1076345 <= p81_literal_1076345;
    p82_literal_1076347 <= p81_literal_1076347;
    p82_literal_1076349 <= p81_literal_1076349;
    p82_literal_1076351 <= p81_literal_1076351;
    p82_literal_1076353 <= p81_literal_1076353;
    p82_literal_1076355 <= p81_literal_1076355;
    p82_literal_1076358 <= p81_literal_1076358;
  end

  // ===== Pipe stage 82:
  wire [127:0] p82_addedKey__68_comb;
  wire [7:0] p82_array_index_1092603_comb;
  wire [7:0] p82_array_index_1092604_comb;
  wire [7:0] p82_array_index_1092605_comb;
  wire [7:0] p82_array_index_1092606_comb;
  wire [7:0] p82_array_index_1092607_comb;
  wire [7:0] p82_array_index_1092608_comb;
  wire [7:0] p82_array_index_1092610_comb;
  wire [7:0] p82_array_index_1092612_comb;
  wire [7:0] p82_array_index_1092613_comb;
  wire [7:0] p82_array_index_1092614_comb;
  wire [7:0] p82_array_index_1092615_comb;
  wire [7:0] p82_array_index_1092616_comb;
  wire [7:0] p82_array_index_1092617_comb;
  wire [7:0] p82_array_index_1092619_comb;
  wire [7:0] p82_array_index_1092620_comb;
  wire [7:0] p82_array_index_1092621_comb;
  wire [7:0] p82_array_index_1092622_comb;
  wire [7:0] p82_array_index_1092623_comb;
  wire [7:0] p82_array_index_1092624_comb;
  wire [7:0] p82_array_index_1092625_comb;
  wire [7:0] p82_array_index_1092627_comb;
  wire [7:0] p82_res7__432_comb;
  wire [7:0] p82_array_index_1092636_comb;
  wire [7:0] p82_array_index_1092637_comb;
  wire [7:0] p82_array_index_1092638_comb;
  wire [7:0] p82_array_index_1092639_comb;
  wire [7:0] p82_array_index_1092640_comb;
  wire [7:0] p82_array_index_1092641_comb;
  wire [7:0] p82_res7__433_comb;
  wire [7:0] p82_array_index_1092651_comb;
  wire [7:0] p82_array_index_1092652_comb;
  wire [7:0] p82_array_index_1092653_comb;
  wire [7:0] p82_array_index_1092654_comb;
  wire [7:0] p82_array_index_1092655_comb;
  wire [7:0] p82_res7__434_comb;
  wire [7:0] p82_array_index_1092665_comb;
  wire [7:0] p82_array_index_1092666_comb;
  wire [7:0] p82_array_index_1092667_comb;
  wire [7:0] p82_array_index_1092668_comb;
  wire [7:0] p82_array_index_1092669_comb;
  wire [7:0] p82_res7__435_comb;
  wire [7:0] p82_array_index_1092680_comb;
  wire [7:0] p82_array_index_1092681_comb;
  wire [7:0] p82_array_index_1092682_comb;
  wire [7:0] p82_array_index_1092683_comb;
  wire [7:0] p82_res7__436_comb;
  assign p82_addedKey__68_comb = p81_xor_1092565 ^ 128'ha226_4131_9aec_d1fd_8352_9103_9b68_6b1c;
  assign p82_array_index_1092603_comb = p81_arr[p82_addedKey__68_comb[127:120]];
  assign p82_array_index_1092604_comb = p81_arr[p82_addedKey__68_comb[119:112]];
  assign p82_array_index_1092605_comb = p81_arr[p82_addedKey__68_comb[111:104]];
  assign p82_array_index_1092606_comb = p81_arr[p82_addedKey__68_comb[103:96]];
  assign p82_array_index_1092607_comb = p81_arr[p82_addedKey__68_comb[95:88]];
  assign p82_array_index_1092608_comb = p81_arr[p82_addedKey__68_comb[87:80]];
  assign p82_array_index_1092610_comb = p81_arr[p82_addedKey__68_comb[71:64]];
  assign p82_array_index_1092612_comb = p81_arr[p82_addedKey__68_comb[55:48]];
  assign p82_array_index_1092613_comb = p81_arr[p82_addedKey__68_comb[47:40]];
  assign p82_array_index_1092614_comb = p81_arr[p82_addedKey__68_comb[39:32]];
  assign p82_array_index_1092615_comb = p81_arr[p82_addedKey__68_comb[31:24]];
  assign p82_array_index_1092616_comb = p81_arr[p82_addedKey__68_comb[23:16]];
  assign p82_array_index_1092617_comb = p81_arr[p82_addedKey__68_comb[15:8]];
  assign p82_array_index_1092619_comb = p81_literal_1076345[p82_array_index_1092603_comb];
  assign p82_array_index_1092620_comb = p81_literal_1076347[p82_array_index_1092604_comb];
  assign p82_array_index_1092621_comb = p81_literal_1076349[p82_array_index_1092605_comb];
  assign p82_array_index_1092622_comb = p81_literal_1076351[p82_array_index_1092606_comb];
  assign p82_array_index_1092623_comb = p81_literal_1076353[p82_array_index_1092607_comb];
  assign p82_array_index_1092624_comb = p81_literal_1076355[p82_array_index_1092608_comb];
  assign p82_array_index_1092625_comb = p81_arr[p82_addedKey__68_comb[79:72]];
  assign p82_array_index_1092627_comb = p81_arr[p82_addedKey__68_comb[63:56]];
  assign p82_res7__432_comb = p82_array_index_1092619_comb ^ p82_array_index_1092620_comb ^ p82_array_index_1092621_comb ^ p82_array_index_1092622_comb ^ p82_array_index_1092623_comb ^ p82_array_index_1092624_comb ^ p82_array_index_1092625_comb ^ p81_literal_1076358[p82_array_index_1092610_comb] ^ p82_array_index_1092627_comb ^ p81_literal_1076355[p82_array_index_1092612_comb] ^ p81_literal_1076353[p82_array_index_1092613_comb] ^ p81_literal_1076351[p82_array_index_1092614_comb] ^ p81_literal_1076349[p82_array_index_1092615_comb] ^ p81_literal_1076347[p82_array_index_1092616_comb] ^ p81_literal_1076345[p82_array_index_1092617_comb] ^ p81_arr[p82_addedKey__68_comb[7:0]];
  assign p82_array_index_1092636_comb = p81_literal_1076345[p82_res7__432_comb];
  assign p82_array_index_1092637_comb = p81_literal_1076347[p82_array_index_1092603_comb];
  assign p82_array_index_1092638_comb = p81_literal_1076349[p82_array_index_1092604_comb];
  assign p82_array_index_1092639_comb = p81_literal_1076351[p82_array_index_1092605_comb];
  assign p82_array_index_1092640_comb = p81_literal_1076353[p82_array_index_1092606_comb];
  assign p82_array_index_1092641_comb = p81_literal_1076355[p82_array_index_1092607_comb];
  assign p82_res7__433_comb = p82_array_index_1092636_comb ^ p82_array_index_1092637_comb ^ p82_array_index_1092638_comb ^ p82_array_index_1092639_comb ^ p82_array_index_1092640_comb ^ p82_array_index_1092641_comb ^ p82_array_index_1092608_comb ^ p81_literal_1076358[p82_array_index_1092625_comb] ^ p82_array_index_1092610_comb ^ p81_literal_1076355[p82_array_index_1092627_comb] ^ p81_literal_1076353[p82_array_index_1092612_comb] ^ p81_literal_1076351[p82_array_index_1092613_comb] ^ p81_literal_1076349[p82_array_index_1092614_comb] ^ p81_literal_1076347[p82_array_index_1092615_comb] ^ p81_literal_1076345[p82_array_index_1092616_comb] ^ p82_array_index_1092617_comb;
  assign p82_array_index_1092651_comb = p81_literal_1076347[p82_res7__432_comb];
  assign p82_array_index_1092652_comb = p81_literal_1076349[p82_array_index_1092603_comb];
  assign p82_array_index_1092653_comb = p81_literal_1076351[p82_array_index_1092604_comb];
  assign p82_array_index_1092654_comb = p81_literal_1076353[p82_array_index_1092605_comb];
  assign p82_array_index_1092655_comb = p81_literal_1076355[p82_array_index_1092606_comb];
  assign p82_res7__434_comb = p81_literal_1076345[p82_res7__433_comb] ^ p82_array_index_1092651_comb ^ p82_array_index_1092652_comb ^ p82_array_index_1092653_comb ^ p82_array_index_1092654_comb ^ p82_array_index_1092655_comb ^ p82_array_index_1092607_comb ^ p81_literal_1076358[p82_array_index_1092608_comb] ^ p82_array_index_1092625_comb ^ p81_literal_1076355[p82_array_index_1092610_comb] ^ p81_literal_1076353[p82_array_index_1092627_comb] ^ p81_literal_1076351[p82_array_index_1092612_comb] ^ p81_literal_1076349[p82_array_index_1092613_comb] ^ p81_literal_1076347[p82_array_index_1092614_comb] ^ p81_literal_1076345[p82_array_index_1092615_comb] ^ p82_array_index_1092616_comb;
  assign p82_array_index_1092665_comb = p81_literal_1076347[p82_res7__433_comb];
  assign p82_array_index_1092666_comb = p81_literal_1076349[p82_res7__432_comb];
  assign p82_array_index_1092667_comb = p81_literal_1076351[p82_array_index_1092603_comb];
  assign p82_array_index_1092668_comb = p81_literal_1076353[p82_array_index_1092604_comb];
  assign p82_array_index_1092669_comb = p81_literal_1076355[p82_array_index_1092605_comb];
  assign p82_res7__435_comb = p81_literal_1076345[p82_res7__434_comb] ^ p82_array_index_1092665_comb ^ p82_array_index_1092666_comb ^ p82_array_index_1092667_comb ^ p82_array_index_1092668_comb ^ p82_array_index_1092669_comb ^ p82_array_index_1092606_comb ^ p81_literal_1076358[p82_array_index_1092607_comb] ^ p82_array_index_1092608_comb ^ p81_literal_1076355[p82_array_index_1092625_comb] ^ p81_literal_1076353[p82_array_index_1092610_comb] ^ p81_literal_1076351[p82_array_index_1092627_comb] ^ p81_literal_1076349[p82_array_index_1092612_comb] ^ p81_literal_1076347[p82_array_index_1092613_comb] ^ p81_literal_1076345[p82_array_index_1092614_comb] ^ p82_array_index_1092615_comb;
  assign p82_array_index_1092680_comb = p81_literal_1076349[p82_res7__433_comb];
  assign p82_array_index_1092681_comb = p81_literal_1076351[p82_res7__432_comb];
  assign p82_array_index_1092682_comb = p81_literal_1076353[p82_array_index_1092603_comb];
  assign p82_array_index_1092683_comb = p81_literal_1076355[p82_array_index_1092604_comb];
  assign p82_res7__436_comb = p81_literal_1076345[p82_res7__435_comb] ^ p81_literal_1076347[p82_res7__434_comb] ^ p82_array_index_1092680_comb ^ p82_array_index_1092681_comb ^ p82_array_index_1092682_comb ^ p82_array_index_1092683_comb ^ p82_array_index_1092605_comb ^ p81_literal_1076358[p82_array_index_1092606_comb] ^ p82_array_index_1092607_comb ^ p82_array_index_1092624_comb ^ p81_literal_1076353[p82_array_index_1092625_comb] ^ p81_literal_1076351[p82_array_index_1092610_comb] ^ p81_literal_1076349[p82_array_index_1092627_comb] ^ p81_literal_1076347[p82_array_index_1092612_comb] ^ p81_literal_1076345[p82_array_index_1092613_comb] ^ p82_array_index_1092614_comb;

  // Registers for pipe stage 82:
  reg [127:0] p82_xor_1091996;
  reg [127:0] p82_xor_1092565;
  reg [7:0] p82_array_index_1092603;
  reg [7:0] p82_array_index_1092604;
  reg [7:0] p82_array_index_1092605;
  reg [7:0] p82_array_index_1092606;
  reg [7:0] p82_array_index_1092607;
  reg [7:0] p82_array_index_1092608;
  reg [7:0] p82_array_index_1092610;
  reg [7:0] p82_array_index_1092612;
  reg [7:0] p82_array_index_1092613;
  reg [7:0] p82_array_index_1092619;
  reg [7:0] p82_array_index_1092620;
  reg [7:0] p82_array_index_1092621;
  reg [7:0] p82_array_index_1092622;
  reg [7:0] p82_array_index_1092623;
  reg [7:0] p82_array_index_1092625;
  reg [7:0] p82_array_index_1092627;
  reg [7:0] p82_res7__432;
  reg [7:0] p82_array_index_1092636;
  reg [7:0] p82_array_index_1092637;
  reg [7:0] p82_array_index_1092638;
  reg [7:0] p82_array_index_1092639;
  reg [7:0] p82_array_index_1092640;
  reg [7:0] p82_array_index_1092641;
  reg [7:0] p82_res7__433;
  reg [7:0] p82_array_index_1092651;
  reg [7:0] p82_array_index_1092652;
  reg [7:0] p82_array_index_1092653;
  reg [7:0] p82_array_index_1092654;
  reg [7:0] p82_array_index_1092655;
  reg [7:0] p82_res7__434;
  reg [7:0] p82_array_index_1092665;
  reg [7:0] p82_array_index_1092666;
  reg [7:0] p82_array_index_1092667;
  reg [7:0] p82_array_index_1092668;
  reg [7:0] p82_array_index_1092669;
  reg [7:0] p82_res7__435;
  reg [7:0] p82_array_index_1092680;
  reg [7:0] p82_array_index_1092681;
  reg [7:0] p82_array_index_1092682;
  reg [7:0] p82_array_index_1092683;
  reg [7:0] p82_res7__436;
  reg [127:0] p82_res__39;
  reg [7:0] p83_arr[256];
  reg [7:0] p83_literal_1076345[256];
  reg [7:0] p83_literal_1076347[256];
  reg [7:0] p83_literal_1076349[256];
  reg [7:0] p83_literal_1076351[256];
  reg [7:0] p83_literal_1076353[256];
  reg [7:0] p83_literal_1076355[256];
  reg [7:0] p83_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p82_xor_1091996 <= p81_xor_1091996;
    p82_xor_1092565 <= p81_xor_1092565;
    p82_array_index_1092603 <= p82_array_index_1092603_comb;
    p82_array_index_1092604 <= p82_array_index_1092604_comb;
    p82_array_index_1092605 <= p82_array_index_1092605_comb;
    p82_array_index_1092606 <= p82_array_index_1092606_comb;
    p82_array_index_1092607 <= p82_array_index_1092607_comb;
    p82_array_index_1092608 <= p82_array_index_1092608_comb;
    p82_array_index_1092610 <= p82_array_index_1092610_comb;
    p82_array_index_1092612 <= p82_array_index_1092612_comb;
    p82_array_index_1092613 <= p82_array_index_1092613_comb;
    p82_array_index_1092619 <= p82_array_index_1092619_comb;
    p82_array_index_1092620 <= p82_array_index_1092620_comb;
    p82_array_index_1092621 <= p82_array_index_1092621_comb;
    p82_array_index_1092622 <= p82_array_index_1092622_comb;
    p82_array_index_1092623 <= p82_array_index_1092623_comb;
    p82_array_index_1092625 <= p82_array_index_1092625_comb;
    p82_array_index_1092627 <= p82_array_index_1092627_comb;
    p82_res7__432 <= p82_res7__432_comb;
    p82_array_index_1092636 <= p82_array_index_1092636_comb;
    p82_array_index_1092637 <= p82_array_index_1092637_comb;
    p82_array_index_1092638 <= p82_array_index_1092638_comb;
    p82_array_index_1092639 <= p82_array_index_1092639_comb;
    p82_array_index_1092640 <= p82_array_index_1092640_comb;
    p82_array_index_1092641 <= p82_array_index_1092641_comb;
    p82_res7__433 <= p82_res7__433_comb;
    p82_array_index_1092651 <= p82_array_index_1092651_comb;
    p82_array_index_1092652 <= p82_array_index_1092652_comb;
    p82_array_index_1092653 <= p82_array_index_1092653_comb;
    p82_array_index_1092654 <= p82_array_index_1092654_comb;
    p82_array_index_1092655 <= p82_array_index_1092655_comb;
    p82_res7__434 <= p82_res7__434_comb;
    p82_array_index_1092665 <= p82_array_index_1092665_comb;
    p82_array_index_1092666 <= p82_array_index_1092666_comb;
    p82_array_index_1092667 <= p82_array_index_1092667_comb;
    p82_array_index_1092668 <= p82_array_index_1092668_comb;
    p82_array_index_1092669 <= p82_array_index_1092669_comb;
    p82_res7__435 <= p82_res7__435_comb;
    p82_array_index_1092680 <= p82_array_index_1092680_comb;
    p82_array_index_1092681 <= p82_array_index_1092681_comb;
    p82_array_index_1092682 <= p82_array_index_1092682_comb;
    p82_array_index_1092683 <= p82_array_index_1092683_comb;
    p82_res7__436 <= p82_res7__436_comb;
    p82_res__39 <= p81_res__39;
    p83_arr <= p82_arr;
    p83_literal_1076345 <= p82_literal_1076345;
    p83_literal_1076347 <= p82_literal_1076347;
    p83_literal_1076349 <= p82_literal_1076349;
    p83_literal_1076351 <= p82_literal_1076351;
    p83_literal_1076353 <= p82_literal_1076353;
    p83_literal_1076355 <= p82_literal_1076355;
    p83_literal_1076358 <= p82_literal_1076358;
  end

  // ===== Pipe stage 83:
  wire [7:0] p83_array_index_1092797_comb;
  wire [7:0] p83_array_index_1092798_comb;
  wire [7:0] p83_array_index_1092799_comb;
  wire [7:0] p83_array_index_1092800_comb;
  wire [7:0] p83_res7__437_comb;
  wire [7:0] p83_array_index_1092811_comb;
  wire [7:0] p83_array_index_1092812_comb;
  wire [7:0] p83_array_index_1092813_comb;
  wire [7:0] p83_res7__438_comb;
  wire [7:0] p83_array_index_1092823_comb;
  wire [7:0] p83_array_index_1092824_comb;
  wire [7:0] p83_array_index_1092825_comb;
  wire [7:0] p83_res7__439_comb;
  wire [7:0] p83_array_index_1092836_comb;
  wire [7:0] p83_array_index_1092837_comb;
  wire [7:0] p83_res7__440_comb;
  wire [7:0] p83_array_index_1092847_comb;
  wire [7:0] p83_array_index_1092848_comb;
  wire [7:0] p83_res7__441_comb;
  wire [7:0] p83_array_index_1092854_comb;
  wire [7:0] p83_array_index_1092855_comb;
  wire [7:0] p83_array_index_1092856_comb;
  wire [7:0] p83_array_index_1092857_comb;
  wire [7:0] p83_array_index_1092858_comb;
  wire [7:0] p83_array_index_1092859_comb;
  wire [7:0] p83_array_index_1092860_comb;
  wire [7:0] p83_array_index_1092861_comb;
  wire [7:0] p83_array_index_1092862_comb;
  assign p83_array_index_1092797_comb = p82_literal_1076349[p82_res7__434];
  assign p83_array_index_1092798_comb = p82_literal_1076351[p82_res7__433];
  assign p83_array_index_1092799_comb = p82_literal_1076353[p82_res7__432];
  assign p83_array_index_1092800_comb = p82_literal_1076355[p82_array_index_1092603];
  assign p83_res7__437_comb = p82_literal_1076345[p82_res7__436] ^ p82_literal_1076347[p82_res7__435] ^ p83_array_index_1092797_comb ^ p83_array_index_1092798_comb ^ p83_array_index_1092799_comb ^ p83_array_index_1092800_comb ^ p82_array_index_1092604 ^ p82_literal_1076358[p82_array_index_1092605] ^ p82_array_index_1092606 ^ p82_array_index_1092641 ^ p82_literal_1076353[p82_array_index_1092608] ^ p82_literal_1076351[p82_array_index_1092625] ^ p82_literal_1076349[p82_array_index_1092610] ^ p82_literal_1076347[p82_array_index_1092627] ^ p82_literal_1076345[p82_array_index_1092612] ^ p82_array_index_1092613;
  assign p83_array_index_1092811_comb = p82_literal_1076351[p82_res7__434];
  assign p83_array_index_1092812_comb = p82_literal_1076353[p82_res7__433];
  assign p83_array_index_1092813_comb = p82_literal_1076355[p82_res7__432];
  assign p83_res7__438_comb = p82_literal_1076345[p83_res7__437_comb] ^ p82_literal_1076347[p82_res7__436] ^ p82_literal_1076349[p82_res7__435] ^ p83_array_index_1092811_comb ^ p83_array_index_1092812_comb ^ p83_array_index_1092813_comb ^ p82_array_index_1092603 ^ p82_literal_1076358[p82_array_index_1092604] ^ p82_array_index_1092605 ^ p82_array_index_1092655 ^ p82_array_index_1092623 ^ p82_literal_1076351[p82_array_index_1092608] ^ p82_literal_1076349[p82_array_index_1092625] ^ p82_literal_1076347[p82_array_index_1092610] ^ p82_literal_1076345[p82_array_index_1092627] ^ p82_array_index_1092612;
  assign p83_array_index_1092823_comb = p82_literal_1076351[p82_res7__435];
  assign p83_array_index_1092824_comb = p82_literal_1076353[p82_res7__434];
  assign p83_array_index_1092825_comb = p82_literal_1076355[p82_res7__433];
  assign p83_res7__439_comb = p82_literal_1076345[p83_res7__438_comb] ^ p82_literal_1076347[p83_res7__437_comb] ^ p82_literal_1076349[p82_res7__436] ^ p83_array_index_1092823_comb ^ p83_array_index_1092824_comb ^ p83_array_index_1092825_comb ^ p82_res7__432 ^ p82_literal_1076358[p82_array_index_1092603] ^ p82_array_index_1092604 ^ p82_array_index_1092669 ^ p82_array_index_1092640 ^ p82_literal_1076351[p82_array_index_1092607] ^ p82_literal_1076349[p82_array_index_1092608] ^ p82_literal_1076347[p82_array_index_1092625] ^ p82_literal_1076345[p82_array_index_1092610] ^ p82_array_index_1092627;
  assign p83_array_index_1092836_comb = p82_literal_1076353[p82_res7__435];
  assign p83_array_index_1092837_comb = p82_literal_1076355[p82_res7__434];
  assign p83_res7__440_comb = p82_literal_1076345[p83_res7__439_comb] ^ p82_literal_1076347[p83_res7__438_comb] ^ p82_literal_1076349[p83_res7__437_comb] ^ p82_literal_1076351[p82_res7__436] ^ p83_array_index_1092836_comb ^ p83_array_index_1092837_comb ^ p82_res7__433 ^ p82_literal_1076358[p82_res7__432] ^ p82_array_index_1092603 ^ p82_array_index_1092683 ^ p82_array_index_1092654 ^ p82_array_index_1092622 ^ p82_literal_1076349[p82_array_index_1092607] ^ p82_literal_1076347[p82_array_index_1092608] ^ p82_literal_1076345[p82_array_index_1092625] ^ p82_array_index_1092610;
  assign p83_array_index_1092847_comb = p82_literal_1076353[p82_res7__436];
  assign p83_array_index_1092848_comb = p82_literal_1076355[p82_res7__435];
  assign p83_res7__441_comb = p82_literal_1076345[p83_res7__440_comb] ^ p82_literal_1076347[p83_res7__439_comb] ^ p82_literal_1076349[p83_res7__438_comb] ^ p82_literal_1076351[p83_res7__437_comb] ^ p83_array_index_1092847_comb ^ p83_array_index_1092848_comb ^ p82_res7__434 ^ p82_literal_1076358[p82_res7__433] ^ p82_res7__432 ^ p83_array_index_1092800_comb ^ p82_array_index_1092668 ^ p82_array_index_1092639 ^ p82_literal_1076349[p82_array_index_1092606] ^ p82_literal_1076347[p82_array_index_1092607] ^ p82_literal_1076345[p82_array_index_1092608] ^ p82_array_index_1092625;
  assign p83_array_index_1092854_comb = p82_literal_1076345[p83_res7__441_comb];
  assign p83_array_index_1092855_comb = p82_literal_1076347[p83_res7__440_comb];
  assign p83_array_index_1092856_comb = p82_literal_1076349[p83_res7__439_comb];
  assign p83_array_index_1092857_comb = p82_literal_1076351[p83_res7__438_comb];
  assign p83_array_index_1092858_comb = p82_literal_1076353[p83_res7__437_comb];
  assign p83_array_index_1092859_comb = p82_literal_1076355[p82_res7__436];
  assign p83_array_index_1092860_comb = p82_literal_1076358[p82_res7__434];
  assign p83_array_index_1092861_comb = p82_literal_1076347[p82_array_index_1092606];
  assign p83_array_index_1092862_comb = p82_literal_1076345[p82_array_index_1092607];

  // Registers for pipe stage 83:
  reg [127:0] p83_xor_1091996;
  reg [127:0] p83_xor_1092565;
  reg [7:0] p83_array_index_1092603;
  reg [7:0] p83_array_index_1092604;
  reg [7:0] p83_array_index_1092605;
  reg [7:0] p83_array_index_1092606;
  reg [7:0] p83_array_index_1092607;
  reg [7:0] p83_array_index_1092608;
  reg [7:0] p83_array_index_1092619;
  reg [7:0] p83_array_index_1092620;
  reg [7:0] p83_array_index_1092621;
  reg [7:0] p83_res7__432;
  reg [7:0] p83_array_index_1092636;
  reg [7:0] p83_array_index_1092637;
  reg [7:0] p83_array_index_1092638;
  reg [7:0] p83_res7__433;
  reg [7:0] p83_array_index_1092651;
  reg [7:0] p83_array_index_1092652;
  reg [7:0] p83_array_index_1092653;
  reg [7:0] p83_res7__434;
  reg [7:0] p83_array_index_1092665;
  reg [7:0] p83_array_index_1092666;
  reg [7:0] p83_array_index_1092667;
  reg [7:0] p83_res7__435;
  reg [7:0] p83_array_index_1092680;
  reg [7:0] p83_array_index_1092681;
  reg [7:0] p83_array_index_1092682;
  reg [7:0] p83_res7__436;
  reg [7:0] p83_array_index_1092797;
  reg [7:0] p83_array_index_1092798;
  reg [7:0] p83_array_index_1092799;
  reg [7:0] p83_res7__437;
  reg [7:0] p83_array_index_1092811;
  reg [7:0] p83_array_index_1092812;
  reg [7:0] p83_array_index_1092813;
  reg [7:0] p83_res7__438;
  reg [7:0] p83_array_index_1092823;
  reg [7:0] p83_array_index_1092824;
  reg [7:0] p83_array_index_1092825;
  reg [7:0] p83_res7__439;
  reg [7:0] p83_array_index_1092836;
  reg [7:0] p83_array_index_1092837;
  reg [7:0] p83_res7__440;
  reg [7:0] p83_array_index_1092847;
  reg [7:0] p83_array_index_1092848;
  reg [7:0] p83_res7__441;
  reg [7:0] p83_array_index_1092854;
  reg [7:0] p83_array_index_1092855;
  reg [7:0] p83_array_index_1092856;
  reg [7:0] p83_array_index_1092857;
  reg [7:0] p83_array_index_1092858;
  reg [7:0] p83_array_index_1092859;
  reg [7:0] p83_array_index_1092860;
  reg [7:0] p83_array_index_1092861;
  reg [7:0] p83_array_index_1092862;
  reg [127:0] p83_res__39;
  reg [7:0] p84_arr[256];
  reg [7:0] p84_literal_1076345[256];
  reg [7:0] p84_literal_1076347[256];
  reg [7:0] p84_literal_1076349[256];
  reg [7:0] p84_literal_1076351[256];
  reg [7:0] p84_literal_1076353[256];
  reg [7:0] p84_literal_1076355[256];
  reg [7:0] p84_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p83_xor_1091996 <= p82_xor_1091996;
    p83_xor_1092565 <= p82_xor_1092565;
    p83_array_index_1092603 <= p82_array_index_1092603;
    p83_array_index_1092604 <= p82_array_index_1092604;
    p83_array_index_1092605 <= p82_array_index_1092605;
    p83_array_index_1092606 <= p82_array_index_1092606;
    p83_array_index_1092607 <= p82_array_index_1092607;
    p83_array_index_1092608 <= p82_array_index_1092608;
    p83_array_index_1092619 <= p82_array_index_1092619;
    p83_array_index_1092620 <= p82_array_index_1092620;
    p83_array_index_1092621 <= p82_array_index_1092621;
    p83_res7__432 <= p82_res7__432;
    p83_array_index_1092636 <= p82_array_index_1092636;
    p83_array_index_1092637 <= p82_array_index_1092637;
    p83_array_index_1092638 <= p82_array_index_1092638;
    p83_res7__433 <= p82_res7__433;
    p83_array_index_1092651 <= p82_array_index_1092651;
    p83_array_index_1092652 <= p82_array_index_1092652;
    p83_array_index_1092653 <= p82_array_index_1092653;
    p83_res7__434 <= p82_res7__434;
    p83_array_index_1092665 <= p82_array_index_1092665;
    p83_array_index_1092666 <= p82_array_index_1092666;
    p83_array_index_1092667 <= p82_array_index_1092667;
    p83_res7__435 <= p82_res7__435;
    p83_array_index_1092680 <= p82_array_index_1092680;
    p83_array_index_1092681 <= p82_array_index_1092681;
    p83_array_index_1092682 <= p82_array_index_1092682;
    p83_res7__436 <= p82_res7__436;
    p83_array_index_1092797 <= p83_array_index_1092797_comb;
    p83_array_index_1092798 <= p83_array_index_1092798_comb;
    p83_array_index_1092799 <= p83_array_index_1092799_comb;
    p83_res7__437 <= p83_res7__437_comb;
    p83_array_index_1092811 <= p83_array_index_1092811_comb;
    p83_array_index_1092812 <= p83_array_index_1092812_comb;
    p83_array_index_1092813 <= p83_array_index_1092813_comb;
    p83_res7__438 <= p83_res7__438_comb;
    p83_array_index_1092823 <= p83_array_index_1092823_comb;
    p83_array_index_1092824 <= p83_array_index_1092824_comb;
    p83_array_index_1092825 <= p83_array_index_1092825_comb;
    p83_res7__439 <= p83_res7__439_comb;
    p83_array_index_1092836 <= p83_array_index_1092836_comb;
    p83_array_index_1092837 <= p83_array_index_1092837_comb;
    p83_res7__440 <= p83_res7__440_comb;
    p83_array_index_1092847 <= p83_array_index_1092847_comb;
    p83_array_index_1092848 <= p83_array_index_1092848_comb;
    p83_res7__441 <= p83_res7__441_comb;
    p83_array_index_1092854 <= p83_array_index_1092854_comb;
    p83_array_index_1092855 <= p83_array_index_1092855_comb;
    p83_array_index_1092856 <= p83_array_index_1092856_comb;
    p83_array_index_1092857 <= p83_array_index_1092857_comb;
    p83_array_index_1092858 <= p83_array_index_1092858_comb;
    p83_array_index_1092859 <= p83_array_index_1092859_comb;
    p83_array_index_1092860 <= p83_array_index_1092860_comb;
    p83_array_index_1092861 <= p83_array_index_1092861_comb;
    p83_array_index_1092862 <= p83_array_index_1092862_comb;
    p83_res__39 <= p82_res__39;
    p84_arr <= p83_arr;
    p84_literal_1076345 <= p83_literal_1076345;
    p84_literal_1076347 <= p83_literal_1076347;
    p84_literal_1076349 <= p83_literal_1076349;
    p84_literal_1076351 <= p83_literal_1076351;
    p84_literal_1076353 <= p83_literal_1076353;
    p84_literal_1076355 <= p83_literal_1076355;
    p84_literal_1076358 <= p83_literal_1076358;
  end

  // ===== Pipe stage 84:
  wire [7:0] p84_res7__442_comb;
  wire [7:0] p84_array_index_1092997_comb;
  wire [7:0] p84_res7__443_comb;
  wire [7:0] p84_res7__444_comb;
  wire [7:0] p84_res7__445_comb;
  wire [7:0] p84_res7__446_comb;
  wire [7:0] p84_res7__447_comb;
  wire [127:0] p84_res__27_comb;
  wire [127:0] p84_xor_1093037_comb;
  assign p84_res7__442_comb = p83_array_index_1092854 ^ p83_array_index_1092855 ^ p83_array_index_1092856 ^ p83_array_index_1092857 ^ p83_array_index_1092858 ^ p83_array_index_1092859 ^ p83_res7__435 ^ p83_array_index_1092860 ^ p83_res7__433 ^ p83_array_index_1092813 ^ p83_array_index_1092682 ^ p83_array_index_1092653 ^ p83_array_index_1092621 ^ p83_array_index_1092861 ^ p83_array_index_1092862 ^ p83_array_index_1092608;
  assign p84_array_index_1092997_comb = p83_literal_1076355[p83_res7__437];
  assign p84_res7__443_comb = p83_literal_1076345[p84_res7__442_comb] ^ p83_literal_1076347[p83_res7__441] ^ p83_literal_1076349[p83_res7__440] ^ p83_literal_1076351[p83_res7__439] ^ p83_literal_1076353[p83_res7__438] ^ p84_array_index_1092997_comb ^ p83_res7__436 ^ p83_literal_1076358[p83_res7__435] ^ p83_res7__434 ^ p83_array_index_1092825 ^ p83_array_index_1092799 ^ p83_array_index_1092667 ^ p83_array_index_1092638 ^ p83_literal_1076347[p83_array_index_1092605] ^ p83_literal_1076345[p83_array_index_1092606] ^ p83_array_index_1092607;
  assign p84_res7__444_comb = p83_literal_1076345[p84_res7__443_comb] ^ p83_literal_1076347[p84_res7__442_comb] ^ p83_literal_1076349[p83_res7__441] ^ p83_literal_1076351[p83_res7__440] ^ p83_literal_1076353[p83_res7__439] ^ p83_literal_1076355[p83_res7__438] ^ p83_res7__437 ^ p83_literal_1076358[p83_res7__436] ^ p83_res7__435 ^ p83_array_index_1092837 ^ p83_array_index_1092812 ^ p83_array_index_1092681 ^ p83_array_index_1092652 ^ p83_array_index_1092620 ^ p83_literal_1076345[p83_array_index_1092605] ^ p83_array_index_1092606;
  assign p84_res7__445_comb = p83_literal_1076345[p84_res7__444_comb] ^ p83_literal_1076347[p84_res7__443_comb] ^ p83_literal_1076349[p84_res7__442_comb] ^ p83_literal_1076351[p83_res7__441] ^ p83_literal_1076353[p83_res7__440] ^ p83_literal_1076355[p83_res7__439] ^ p83_res7__438 ^ p83_literal_1076358[p83_res7__437] ^ p83_res7__436 ^ p83_array_index_1092848 ^ p83_array_index_1092824 ^ p83_array_index_1092798 ^ p83_array_index_1092666 ^ p83_array_index_1092637 ^ p83_literal_1076345[p83_array_index_1092604] ^ p83_array_index_1092605;
  assign p84_res7__446_comb = p83_literal_1076345[p84_res7__445_comb] ^ p83_literal_1076347[p84_res7__444_comb] ^ p83_literal_1076349[p84_res7__443_comb] ^ p83_literal_1076351[p84_res7__442_comb] ^ p83_literal_1076353[p83_res7__441] ^ p83_literal_1076355[p83_res7__440] ^ p83_res7__439 ^ p83_literal_1076358[p83_res7__438] ^ p83_res7__437 ^ p83_array_index_1092859 ^ p83_array_index_1092836 ^ p83_array_index_1092811 ^ p83_array_index_1092680 ^ p83_array_index_1092651 ^ p83_array_index_1092619 ^ p83_array_index_1092604;
  assign p84_res7__447_comb = p83_literal_1076345[p84_res7__446_comb] ^ p83_literal_1076347[p84_res7__445_comb] ^ p83_literal_1076349[p84_res7__444_comb] ^ p83_literal_1076351[p84_res7__443_comb] ^ p83_literal_1076353[p84_res7__442_comb] ^ p83_literal_1076355[p83_res7__441] ^ p83_res7__440 ^ p83_literal_1076358[p83_res7__439] ^ p83_res7__438 ^ p84_array_index_1092997_comb ^ p83_array_index_1092847 ^ p83_array_index_1092823 ^ p83_array_index_1092797 ^ p83_array_index_1092665 ^ p83_array_index_1092636 ^ p83_array_index_1092603;
  assign p84_res__27_comb = {p84_res7__447_comb, p84_res7__446_comb, p84_res7__445_comb, p84_res7__444_comb, p84_res7__443_comb, p84_res7__442_comb, p83_res7__441, p83_res7__440, p83_res7__439, p83_res7__438, p83_res7__437, p83_res7__436, p83_res7__435, p83_res7__434, p83_res7__433, p83_res7__432};
  assign p84_xor_1093037_comb = p84_res__27_comb ^ p83_xor_1091996;

  // Registers for pipe stage 84:
  reg [127:0] p84_xor_1092565;
  reg [127:0] p84_xor_1093037;
  reg [127:0] p84_res__39;
  reg [7:0] p85_arr[256];
  reg [7:0] p85_literal_1076345[256];
  reg [7:0] p85_literal_1076347[256];
  reg [7:0] p85_literal_1076349[256];
  reg [7:0] p85_literal_1076351[256];
  reg [7:0] p85_literal_1076353[256];
  reg [7:0] p85_literal_1076355[256];
  reg [7:0] p85_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p84_xor_1092565 <= p83_xor_1092565;
    p84_xor_1093037 <= p84_xor_1093037_comb;
    p84_res__39 <= p83_res__39;
    p85_arr <= p84_arr;
    p85_literal_1076345 <= p84_literal_1076345;
    p85_literal_1076347 <= p84_literal_1076347;
    p85_literal_1076349 <= p84_literal_1076349;
    p85_literal_1076351 <= p84_literal_1076351;
    p85_literal_1076353 <= p84_literal_1076353;
    p85_literal_1076355 <= p84_literal_1076355;
    p85_literal_1076358 <= p84_literal_1076358;
  end

  // ===== Pipe stage 85:
  wire [127:0] p85_addedKey__69_comb;
  wire [7:0] p85_array_index_1093075_comb;
  wire [7:0] p85_array_index_1093076_comb;
  wire [7:0] p85_array_index_1093077_comb;
  wire [7:0] p85_array_index_1093078_comb;
  wire [7:0] p85_array_index_1093079_comb;
  wire [7:0] p85_array_index_1093080_comb;
  wire [7:0] p85_array_index_1093082_comb;
  wire [7:0] p85_array_index_1093084_comb;
  wire [7:0] p85_array_index_1093085_comb;
  wire [7:0] p85_array_index_1093086_comb;
  wire [7:0] p85_array_index_1093087_comb;
  wire [7:0] p85_array_index_1093088_comb;
  wire [7:0] p85_array_index_1093089_comb;
  wire [7:0] p85_array_index_1093091_comb;
  wire [7:0] p85_array_index_1093092_comb;
  wire [7:0] p85_array_index_1093093_comb;
  wire [7:0] p85_array_index_1093094_comb;
  wire [7:0] p85_array_index_1093095_comb;
  wire [7:0] p85_array_index_1093096_comb;
  wire [7:0] p85_array_index_1093097_comb;
  wire [7:0] p85_array_index_1093099_comb;
  wire [7:0] p85_res7__448_comb;
  wire [7:0] p85_array_index_1093108_comb;
  wire [7:0] p85_array_index_1093109_comb;
  wire [7:0] p85_array_index_1093110_comb;
  wire [7:0] p85_array_index_1093111_comb;
  wire [7:0] p85_array_index_1093112_comb;
  wire [7:0] p85_array_index_1093113_comb;
  wire [7:0] p85_res7__449_comb;
  wire [7:0] p85_array_index_1093123_comb;
  wire [7:0] p85_array_index_1093124_comb;
  wire [7:0] p85_array_index_1093125_comb;
  wire [7:0] p85_array_index_1093126_comb;
  wire [7:0] p85_array_index_1093127_comb;
  wire [7:0] p85_res7__450_comb;
  wire [7:0] p85_array_index_1093137_comb;
  wire [7:0] p85_array_index_1093138_comb;
  wire [7:0] p85_array_index_1093139_comb;
  wire [7:0] p85_array_index_1093140_comb;
  wire [7:0] p85_array_index_1093141_comb;
  wire [7:0] p85_res7__451_comb;
  wire [7:0] p85_array_index_1093152_comb;
  wire [7:0] p85_array_index_1093153_comb;
  wire [7:0] p85_array_index_1093154_comb;
  wire [7:0] p85_array_index_1093155_comb;
  wire [7:0] p85_res7__452_comb;
  assign p85_addedKey__69_comb = p84_xor_1093037 ^ 128'hcc84_3743_f6a4_ab45_de75_2c13_46ec_ff1d;
  assign p85_array_index_1093075_comb = p84_arr[p85_addedKey__69_comb[127:120]];
  assign p85_array_index_1093076_comb = p84_arr[p85_addedKey__69_comb[119:112]];
  assign p85_array_index_1093077_comb = p84_arr[p85_addedKey__69_comb[111:104]];
  assign p85_array_index_1093078_comb = p84_arr[p85_addedKey__69_comb[103:96]];
  assign p85_array_index_1093079_comb = p84_arr[p85_addedKey__69_comb[95:88]];
  assign p85_array_index_1093080_comb = p84_arr[p85_addedKey__69_comb[87:80]];
  assign p85_array_index_1093082_comb = p84_arr[p85_addedKey__69_comb[71:64]];
  assign p85_array_index_1093084_comb = p84_arr[p85_addedKey__69_comb[55:48]];
  assign p85_array_index_1093085_comb = p84_arr[p85_addedKey__69_comb[47:40]];
  assign p85_array_index_1093086_comb = p84_arr[p85_addedKey__69_comb[39:32]];
  assign p85_array_index_1093087_comb = p84_arr[p85_addedKey__69_comb[31:24]];
  assign p85_array_index_1093088_comb = p84_arr[p85_addedKey__69_comb[23:16]];
  assign p85_array_index_1093089_comb = p84_arr[p85_addedKey__69_comb[15:8]];
  assign p85_array_index_1093091_comb = p84_literal_1076345[p85_array_index_1093075_comb];
  assign p85_array_index_1093092_comb = p84_literal_1076347[p85_array_index_1093076_comb];
  assign p85_array_index_1093093_comb = p84_literal_1076349[p85_array_index_1093077_comb];
  assign p85_array_index_1093094_comb = p84_literal_1076351[p85_array_index_1093078_comb];
  assign p85_array_index_1093095_comb = p84_literal_1076353[p85_array_index_1093079_comb];
  assign p85_array_index_1093096_comb = p84_literal_1076355[p85_array_index_1093080_comb];
  assign p85_array_index_1093097_comb = p84_arr[p85_addedKey__69_comb[79:72]];
  assign p85_array_index_1093099_comb = p84_arr[p85_addedKey__69_comb[63:56]];
  assign p85_res7__448_comb = p85_array_index_1093091_comb ^ p85_array_index_1093092_comb ^ p85_array_index_1093093_comb ^ p85_array_index_1093094_comb ^ p85_array_index_1093095_comb ^ p85_array_index_1093096_comb ^ p85_array_index_1093097_comb ^ p84_literal_1076358[p85_array_index_1093082_comb] ^ p85_array_index_1093099_comb ^ p84_literal_1076355[p85_array_index_1093084_comb] ^ p84_literal_1076353[p85_array_index_1093085_comb] ^ p84_literal_1076351[p85_array_index_1093086_comb] ^ p84_literal_1076349[p85_array_index_1093087_comb] ^ p84_literal_1076347[p85_array_index_1093088_comb] ^ p84_literal_1076345[p85_array_index_1093089_comb] ^ p84_arr[p85_addedKey__69_comb[7:0]];
  assign p85_array_index_1093108_comb = p84_literal_1076345[p85_res7__448_comb];
  assign p85_array_index_1093109_comb = p84_literal_1076347[p85_array_index_1093075_comb];
  assign p85_array_index_1093110_comb = p84_literal_1076349[p85_array_index_1093076_comb];
  assign p85_array_index_1093111_comb = p84_literal_1076351[p85_array_index_1093077_comb];
  assign p85_array_index_1093112_comb = p84_literal_1076353[p85_array_index_1093078_comb];
  assign p85_array_index_1093113_comb = p84_literal_1076355[p85_array_index_1093079_comb];
  assign p85_res7__449_comb = p85_array_index_1093108_comb ^ p85_array_index_1093109_comb ^ p85_array_index_1093110_comb ^ p85_array_index_1093111_comb ^ p85_array_index_1093112_comb ^ p85_array_index_1093113_comb ^ p85_array_index_1093080_comb ^ p84_literal_1076358[p85_array_index_1093097_comb] ^ p85_array_index_1093082_comb ^ p84_literal_1076355[p85_array_index_1093099_comb] ^ p84_literal_1076353[p85_array_index_1093084_comb] ^ p84_literal_1076351[p85_array_index_1093085_comb] ^ p84_literal_1076349[p85_array_index_1093086_comb] ^ p84_literal_1076347[p85_array_index_1093087_comb] ^ p84_literal_1076345[p85_array_index_1093088_comb] ^ p85_array_index_1093089_comb;
  assign p85_array_index_1093123_comb = p84_literal_1076347[p85_res7__448_comb];
  assign p85_array_index_1093124_comb = p84_literal_1076349[p85_array_index_1093075_comb];
  assign p85_array_index_1093125_comb = p84_literal_1076351[p85_array_index_1093076_comb];
  assign p85_array_index_1093126_comb = p84_literal_1076353[p85_array_index_1093077_comb];
  assign p85_array_index_1093127_comb = p84_literal_1076355[p85_array_index_1093078_comb];
  assign p85_res7__450_comb = p84_literal_1076345[p85_res7__449_comb] ^ p85_array_index_1093123_comb ^ p85_array_index_1093124_comb ^ p85_array_index_1093125_comb ^ p85_array_index_1093126_comb ^ p85_array_index_1093127_comb ^ p85_array_index_1093079_comb ^ p84_literal_1076358[p85_array_index_1093080_comb] ^ p85_array_index_1093097_comb ^ p84_literal_1076355[p85_array_index_1093082_comb] ^ p84_literal_1076353[p85_array_index_1093099_comb] ^ p84_literal_1076351[p85_array_index_1093084_comb] ^ p84_literal_1076349[p85_array_index_1093085_comb] ^ p84_literal_1076347[p85_array_index_1093086_comb] ^ p84_literal_1076345[p85_array_index_1093087_comb] ^ p85_array_index_1093088_comb;
  assign p85_array_index_1093137_comb = p84_literal_1076347[p85_res7__449_comb];
  assign p85_array_index_1093138_comb = p84_literal_1076349[p85_res7__448_comb];
  assign p85_array_index_1093139_comb = p84_literal_1076351[p85_array_index_1093075_comb];
  assign p85_array_index_1093140_comb = p84_literal_1076353[p85_array_index_1093076_comb];
  assign p85_array_index_1093141_comb = p84_literal_1076355[p85_array_index_1093077_comb];
  assign p85_res7__451_comb = p84_literal_1076345[p85_res7__450_comb] ^ p85_array_index_1093137_comb ^ p85_array_index_1093138_comb ^ p85_array_index_1093139_comb ^ p85_array_index_1093140_comb ^ p85_array_index_1093141_comb ^ p85_array_index_1093078_comb ^ p84_literal_1076358[p85_array_index_1093079_comb] ^ p85_array_index_1093080_comb ^ p84_literal_1076355[p85_array_index_1093097_comb] ^ p84_literal_1076353[p85_array_index_1093082_comb] ^ p84_literal_1076351[p85_array_index_1093099_comb] ^ p84_literal_1076349[p85_array_index_1093084_comb] ^ p84_literal_1076347[p85_array_index_1093085_comb] ^ p84_literal_1076345[p85_array_index_1093086_comb] ^ p85_array_index_1093087_comb;
  assign p85_array_index_1093152_comb = p84_literal_1076349[p85_res7__449_comb];
  assign p85_array_index_1093153_comb = p84_literal_1076351[p85_res7__448_comb];
  assign p85_array_index_1093154_comb = p84_literal_1076353[p85_array_index_1093075_comb];
  assign p85_array_index_1093155_comb = p84_literal_1076355[p85_array_index_1093076_comb];
  assign p85_res7__452_comb = p84_literal_1076345[p85_res7__451_comb] ^ p84_literal_1076347[p85_res7__450_comb] ^ p85_array_index_1093152_comb ^ p85_array_index_1093153_comb ^ p85_array_index_1093154_comb ^ p85_array_index_1093155_comb ^ p85_array_index_1093077_comb ^ p84_literal_1076358[p85_array_index_1093078_comb] ^ p85_array_index_1093079_comb ^ p85_array_index_1093096_comb ^ p84_literal_1076353[p85_array_index_1093097_comb] ^ p84_literal_1076351[p85_array_index_1093082_comb] ^ p84_literal_1076349[p85_array_index_1093099_comb] ^ p84_literal_1076347[p85_array_index_1093084_comb] ^ p84_literal_1076345[p85_array_index_1093085_comb] ^ p85_array_index_1093086_comb;

  // Registers for pipe stage 85:
  reg [127:0] p85_xor_1092565;
  reg [127:0] p85_xor_1093037;
  reg [7:0] p85_array_index_1093075;
  reg [7:0] p85_array_index_1093076;
  reg [7:0] p85_array_index_1093077;
  reg [7:0] p85_array_index_1093078;
  reg [7:0] p85_array_index_1093079;
  reg [7:0] p85_array_index_1093080;
  reg [7:0] p85_array_index_1093082;
  reg [7:0] p85_array_index_1093084;
  reg [7:0] p85_array_index_1093085;
  reg [7:0] p85_array_index_1093091;
  reg [7:0] p85_array_index_1093092;
  reg [7:0] p85_array_index_1093093;
  reg [7:0] p85_array_index_1093094;
  reg [7:0] p85_array_index_1093095;
  reg [7:0] p85_array_index_1093097;
  reg [7:0] p85_array_index_1093099;
  reg [7:0] p85_res7__448;
  reg [7:0] p85_array_index_1093108;
  reg [7:0] p85_array_index_1093109;
  reg [7:0] p85_array_index_1093110;
  reg [7:0] p85_array_index_1093111;
  reg [7:0] p85_array_index_1093112;
  reg [7:0] p85_array_index_1093113;
  reg [7:0] p85_res7__449;
  reg [7:0] p85_array_index_1093123;
  reg [7:0] p85_array_index_1093124;
  reg [7:0] p85_array_index_1093125;
  reg [7:0] p85_array_index_1093126;
  reg [7:0] p85_array_index_1093127;
  reg [7:0] p85_res7__450;
  reg [7:0] p85_array_index_1093137;
  reg [7:0] p85_array_index_1093138;
  reg [7:0] p85_array_index_1093139;
  reg [7:0] p85_array_index_1093140;
  reg [7:0] p85_array_index_1093141;
  reg [7:0] p85_res7__451;
  reg [7:0] p85_array_index_1093152;
  reg [7:0] p85_array_index_1093153;
  reg [7:0] p85_array_index_1093154;
  reg [7:0] p85_array_index_1093155;
  reg [7:0] p85_res7__452;
  reg [127:0] p85_res__39;
  reg [7:0] p86_arr[256];
  reg [7:0] p86_literal_1076345[256];
  reg [7:0] p86_literal_1076347[256];
  reg [7:0] p86_literal_1076349[256];
  reg [7:0] p86_literal_1076351[256];
  reg [7:0] p86_literal_1076353[256];
  reg [7:0] p86_literal_1076355[256];
  reg [7:0] p86_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p85_xor_1092565 <= p84_xor_1092565;
    p85_xor_1093037 <= p84_xor_1093037;
    p85_array_index_1093075 <= p85_array_index_1093075_comb;
    p85_array_index_1093076 <= p85_array_index_1093076_comb;
    p85_array_index_1093077 <= p85_array_index_1093077_comb;
    p85_array_index_1093078 <= p85_array_index_1093078_comb;
    p85_array_index_1093079 <= p85_array_index_1093079_comb;
    p85_array_index_1093080 <= p85_array_index_1093080_comb;
    p85_array_index_1093082 <= p85_array_index_1093082_comb;
    p85_array_index_1093084 <= p85_array_index_1093084_comb;
    p85_array_index_1093085 <= p85_array_index_1093085_comb;
    p85_array_index_1093091 <= p85_array_index_1093091_comb;
    p85_array_index_1093092 <= p85_array_index_1093092_comb;
    p85_array_index_1093093 <= p85_array_index_1093093_comb;
    p85_array_index_1093094 <= p85_array_index_1093094_comb;
    p85_array_index_1093095 <= p85_array_index_1093095_comb;
    p85_array_index_1093097 <= p85_array_index_1093097_comb;
    p85_array_index_1093099 <= p85_array_index_1093099_comb;
    p85_res7__448 <= p85_res7__448_comb;
    p85_array_index_1093108 <= p85_array_index_1093108_comb;
    p85_array_index_1093109 <= p85_array_index_1093109_comb;
    p85_array_index_1093110 <= p85_array_index_1093110_comb;
    p85_array_index_1093111 <= p85_array_index_1093111_comb;
    p85_array_index_1093112 <= p85_array_index_1093112_comb;
    p85_array_index_1093113 <= p85_array_index_1093113_comb;
    p85_res7__449 <= p85_res7__449_comb;
    p85_array_index_1093123 <= p85_array_index_1093123_comb;
    p85_array_index_1093124 <= p85_array_index_1093124_comb;
    p85_array_index_1093125 <= p85_array_index_1093125_comb;
    p85_array_index_1093126 <= p85_array_index_1093126_comb;
    p85_array_index_1093127 <= p85_array_index_1093127_comb;
    p85_res7__450 <= p85_res7__450_comb;
    p85_array_index_1093137 <= p85_array_index_1093137_comb;
    p85_array_index_1093138 <= p85_array_index_1093138_comb;
    p85_array_index_1093139 <= p85_array_index_1093139_comb;
    p85_array_index_1093140 <= p85_array_index_1093140_comb;
    p85_array_index_1093141 <= p85_array_index_1093141_comb;
    p85_res7__451 <= p85_res7__451_comb;
    p85_array_index_1093152 <= p85_array_index_1093152_comb;
    p85_array_index_1093153 <= p85_array_index_1093153_comb;
    p85_array_index_1093154 <= p85_array_index_1093154_comb;
    p85_array_index_1093155 <= p85_array_index_1093155_comb;
    p85_res7__452 <= p85_res7__452_comb;
    p85_res__39 <= p84_res__39;
    p86_arr <= p85_arr;
    p86_literal_1076345 <= p85_literal_1076345;
    p86_literal_1076347 <= p85_literal_1076347;
    p86_literal_1076349 <= p85_literal_1076349;
    p86_literal_1076351 <= p85_literal_1076351;
    p86_literal_1076353 <= p85_literal_1076353;
    p86_literal_1076355 <= p85_literal_1076355;
    p86_literal_1076358 <= p85_literal_1076358;
  end

  // ===== Pipe stage 86:
  wire [7:0] p86_array_index_1093269_comb;
  wire [7:0] p86_array_index_1093270_comb;
  wire [7:0] p86_array_index_1093271_comb;
  wire [7:0] p86_array_index_1093272_comb;
  wire [7:0] p86_res7__453_comb;
  wire [7:0] p86_array_index_1093283_comb;
  wire [7:0] p86_array_index_1093284_comb;
  wire [7:0] p86_array_index_1093285_comb;
  wire [7:0] p86_res7__454_comb;
  wire [7:0] p86_array_index_1093295_comb;
  wire [7:0] p86_array_index_1093296_comb;
  wire [7:0] p86_array_index_1093297_comb;
  wire [7:0] p86_res7__455_comb;
  wire [7:0] p86_array_index_1093308_comb;
  wire [7:0] p86_array_index_1093309_comb;
  wire [7:0] p86_res7__456_comb;
  wire [7:0] p86_array_index_1093319_comb;
  wire [7:0] p86_array_index_1093320_comb;
  wire [7:0] p86_res7__457_comb;
  wire [7:0] p86_array_index_1093326_comb;
  wire [7:0] p86_array_index_1093327_comb;
  wire [7:0] p86_array_index_1093328_comb;
  wire [7:0] p86_array_index_1093329_comb;
  wire [7:0] p86_array_index_1093330_comb;
  wire [7:0] p86_array_index_1093331_comb;
  wire [7:0] p86_array_index_1093332_comb;
  wire [7:0] p86_array_index_1093333_comb;
  wire [7:0] p86_array_index_1093334_comb;
  assign p86_array_index_1093269_comb = p85_literal_1076349[p85_res7__450];
  assign p86_array_index_1093270_comb = p85_literal_1076351[p85_res7__449];
  assign p86_array_index_1093271_comb = p85_literal_1076353[p85_res7__448];
  assign p86_array_index_1093272_comb = p85_literal_1076355[p85_array_index_1093075];
  assign p86_res7__453_comb = p85_literal_1076345[p85_res7__452] ^ p85_literal_1076347[p85_res7__451] ^ p86_array_index_1093269_comb ^ p86_array_index_1093270_comb ^ p86_array_index_1093271_comb ^ p86_array_index_1093272_comb ^ p85_array_index_1093076 ^ p85_literal_1076358[p85_array_index_1093077] ^ p85_array_index_1093078 ^ p85_array_index_1093113 ^ p85_literal_1076353[p85_array_index_1093080] ^ p85_literal_1076351[p85_array_index_1093097] ^ p85_literal_1076349[p85_array_index_1093082] ^ p85_literal_1076347[p85_array_index_1093099] ^ p85_literal_1076345[p85_array_index_1093084] ^ p85_array_index_1093085;
  assign p86_array_index_1093283_comb = p85_literal_1076351[p85_res7__450];
  assign p86_array_index_1093284_comb = p85_literal_1076353[p85_res7__449];
  assign p86_array_index_1093285_comb = p85_literal_1076355[p85_res7__448];
  assign p86_res7__454_comb = p85_literal_1076345[p86_res7__453_comb] ^ p85_literal_1076347[p85_res7__452] ^ p85_literal_1076349[p85_res7__451] ^ p86_array_index_1093283_comb ^ p86_array_index_1093284_comb ^ p86_array_index_1093285_comb ^ p85_array_index_1093075 ^ p85_literal_1076358[p85_array_index_1093076] ^ p85_array_index_1093077 ^ p85_array_index_1093127 ^ p85_array_index_1093095 ^ p85_literal_1076351[p85_array_index_1093080] ^ p85_literal_1076349[p85_array_index_1093097] ^ p85_literal_1076347[p85_array_index_1093082] ^ p85_literal_1076345[p85_array_index_1093099] ^ p85_array_index_1093084;
  assign p86_array_index_1093295_comb = p85_literal_1076351[p85_res7__451];
  assign p86_array_index_1093296_comb = p85_literal_1076353[p85_res7__450];
  assign p86_array_index_1093297_comb = p85_literal_1076355[p85_res7__449];
  assign p86_res7__455_comb = p85_literal_1076345[p86_res7__454_comb] ^ p85_literal_1076347[p86_res7__453_comb] ^ p85_literal_1076349[p85_res7__452] ^ p86_array_index_1093295_comb ^ p86_array_index_1093296_comb ^ p86_array_index_1093297_comb ^ p85_res7__448 ^ p85_literal_1076358[p85_array_index_1093075] ^ p85_array_index_1093076 ^ p85_array_index_1093141 ^ p85_array_index_1093112 ^ p85_literal_1076351[p85_array_index_1093079] ^ p85_literal_1076349[p85_array_index_1093080] ^ p85_literal_1076347[p85_array_index_1093097] ^ p85_literal_1076345[p85_array_index_1093082] ^ p85_array_index_1093099;
  assign p86_array_index_1093308_comb = p85_literal_1076353[p85_res7__451];
  assign p86_array_index_1093309_comb = p85_literal_1076355[p85_res7__450];
  assign p86_res7__456_comb = p85_literal_1076345[p86_res7__455_comb] ^ p85_literal_1076347[p86_res7__454_comb] ^ p85_literal_1076349[p86_res7__453_comb] ^ p85_literal_1076351[p85_res7__452] ^ p86_array_index_1093308_comb ^ p86_array_index_1093309_comb ^ p85_res7__449 ^ p85_literal_1076358[p85_res7__448] ^ p85_array_index_1093075 ^ p85_array_index_1093155 ^ p85_array_index_1093126 ^ p85_array_index_1093094 ^ p85_literal_1076349[p85_array_index_1093079] ^ p85_literal_1076347[p85_array_index_1093080] ^ p85_literal_1076345[p85_array_index_1093097] ^ p85_array_index_1093082;
  assign p86_array_index_1093319_comb = p85_literal_1076353[p85_res7__452];
  assign p86_array_index_1093320_comb = p85_literal_1076355[p85_res7__451];
  assign p86_res7__457_comb = p85_literal_1076345[p86_res7__456_comb] ^ p85_literal_1076347[p86_res7__455_comb] ^ p85_literal_1076349[p86_res7__454_comb] ^ p85_literal_1076351[p86_res7__453_comb] ^ p86_array_index_1093319_comb ^ p86_array_index_1093320_comb ^ p85_res7__450 ^ p85_literal_1076358[p85_res7__449] ^ p85_res7__448 ^ p86_array_index_1093272_comb ^ p85_array_index_1093140 ^ p85_array_index_1093111 ^ p85_literal_1076349[p85_array_index_1093078] ^ p85_literal_1076347[p85_array_index_1093079] ^ p85_literal_1076345[p85_array_index_1093080] ^ p85_array_index_1093097;
  assign p86_array_index_1093326_comb = p85_literal_1076345[p86_res7__457_comb];
  assign p86_array_index_1093327_comb = p85_literal_1076347[p86_res7__456_comb];
  assign p86_array_index_1093328_comb = p85_literal_1076349[p86_res7__455_comb];
  assign p86_array_index_1093329_comb = p85_literal_1076351[p86_res7__454_comb];
  assign p86_array_index_1093330_comb = p85_literal_1076353[p86_res7__453_comb];
  assign p86_array_index_1093331_comb = p85_literal_1076355[p85_res7__452];
  assign p86_array_index_1093332_comb = p85_literal_1076358[p85_res7__450];
  assign p86_array_index_1093333_comb = p85_literal_1076347[p85_array_index_1093078];
  assign p86_array_index_1093334_comb = p85_literal_1076345[p85_array_index_1093079];

  // Registers for pipe stage 86:
  reg [127:0] p86_xor_1092565;
  reg [127:0] p86_xor_1093037;
  reg [7:0] p86_array_index_1093075;
  reg [7:0] p86_array_index_1093076;
  reg [7:0] p86_array_index_1093077;
  reg [7:0] p86_array_index_1093078;
  reg [7:0] p86_array_index_1093079;
  reg [7:0] p86_array_index_1093080;
  reg [7:0] p86_array_index_1093091;
  reg [7:0] p86_array_index_1093092;
  reg [7:0] p86_array_index_1093093;
  reg [7:0] p86_res7__448;
  reg [7:0] p86_array_index_1093108;
  reg [7:0] p86_array_index_1093109;
  reg [7:0] p86_array_index_1093110;
  reg [7:0] p86_res7__449;
  reg [7:0] p86_array_index_1093123;
  reg [7:0] p86_array_index_1093124;
  reg [7:0] p86_array_index_1093125;
  reg [7:0] p86_res7__450;
  reg [7:0] p86_array_index_1093137;
  reg [7:0] p86_array_index_1093138;
  reg [7:0] p86_array_index_1093139;
  reg [7:0] p86_res7__451;
  reg [7:0] p86_array_index_1093152;
  reg [7:0] p86_array_index_1093153;
  reg [7:0] p86_array_index_1093154;
  reg [7:0] p86_res7__452;
  reg [7:0] p86_array_index_1093269;
  reg [7:0] p86_array_index_1093270;
  reg [7:0] p86_array_index_1093271;
  reg [7:0] p86_res7__453;
  reg [7:0] p86_array_index_1093283;
  reg [7:0] p86_array_index_1093284;
  reg [7:0] p86_array_index_1093285;
  reg [7:0] p86_res7__454;
  reg [7:0] p86_array_index_1093295;
  reg [7:0] p86_array_index_1093296;
  reg [7:0] p86_array_index_1093297;
  reg [7:0] p86_res7__455;
  reg [7:0] p86_array_index_1093308;
  reg [7:0] p86_array_index_1093309;
  reg [7:0] p86_res7__456;
  reg [7:0] p86_array_index_1093319;
  reg [7:0] p86_array_index_1093320;
  reg [7:0] p86_res7__457;
  reg [7:0] p86_array_index_1093326;
  reg [7:0] p86_array_index_1093327;
  reg [7:0] p86_array_index_1093328;
  reg [7:0] p86_array_index_1093329;
  reg [7:0] p86_array_index_1093330;
  reg [7:0] p86_array_index_1093331;
  reg [7:0] p86_array_index_1093332;
  reg [7:0] p86_array_index_1093333;
  reg [7:0] p86_array_index_1093334;
  reg [127:0] p86_res__39;
  reg [7:0] p87_arr[256];
  reg [7:0] p87_literal_1076345[256];
  reg [7:0] p87_literal_1076347[256];
  reg [7:0] p87_literal_1076349[256];
  reg [7:0] p87_literal_1076351[256];
  reg [7:0] p87_literal_1076353[256];
  reg [7:0] p87_literal_1076355[256];
  reg [7:0] p87_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p86_xor_1092565 <= p85_xor_1092565;
    p86_xor_1093037 <= p85_xor_1093037;
    p86_array_index_1093075 <= p85_array_index_1093075;
    p86_array_index_1093076 <= p85_array_index_1093076;
    p86_array_index_1093077 <= p85_array_index_1093077;
    p86_array_index_1093078 <= p85_array_index_1093078;
    p86_array_index_1093079 <= p85_array_index_1093079;
    p86_array_index_1093080 <= p85_array_index_1093080;
    p86_array_index_1093091 <= p85_array_index_1093091;
    p86_array_index_1093092 <= p85_array_index_1093092;
    p86_array_index_1093093 <= p85_array_index_1093093;
    p86_res7__448 <= p85_res7__448;
    p86_array_index_1093108 <= p85_array_index_1093108;
    p86_array_index_1093109 <= p85_array_index_1093109;
    p86_array_index_1093110 <= p85_array_index_1093110;
    p86_res7__449 <= p85_res7__449;
    p86_array_index_1093123 <= p85_array_index_1093123;
    p86_array_index_1093124 <= p85_array_index_1093124;
    p86_array_index_1093125 <= p85_array_index_1093125;
    p86_res7__450 <= p85_res7__450;
    p86_array_index_1093137 <= p85_array_index_1093137;
    p86_array_index_1093138 <= p85_array_index_1093138;
    p86_array_index_1093139 <= p85_array_index_1093139;
    p86_res7__451 <= p85_res7__451;
    p86_array_index_1093152 <= p85_array_index_1093152;
    p86_array_index_1093153 <= p85_array_index_1093153;
    p86_array_index_1093154 <= p85_array_index_1093154;
    p86_res7__452 <= p85_res7__452;
    p86_array_index_1093269 <= p86_array_index_1093269_comb;
    p86_array_index_1093270 <= p86_array_index_1093270_comb;
    p86_array_index_1093271 <= p86_array_index_1093271_comb;
    p86_res7__453 <= p86_res7__453_comb;
    p86_array_index_1093283 <= p86_array_index_1093283_comb;
    p86_array_index_1093284 <= p86_array_index_1093284_comb;
    p86_array_index_1093285 <= p86_array_index_1093285_comb;
    p86_res7__454 <= p86_res7__454_comb;
    p86_array_index_1093295 <= p86_array_index_1093295_comb;
    p86_array_index_1093296 <= p86_array_index_1093296_comb;
    p86_array_index_1093297 <= p86_array_index_1093297_comb;
    p86_res7__455 <= p86_res7__455_comb;
    p86_array_index_1093308 <= p86_array_index_1093308_comb;
    p86_array_index_1093309 <= p86_array_index_1093309_comb;
    p86_res7__456 <= p86_res7__456_comb;
    p86_array_index_1093319 <= p86_array_index_1093319_comb;
    p86_array_index_1093320 <= p86_array_index_1093320_comb;
    p86_res7__457 <= p86_res7__457_comb;
    p86_array_index_1093326 <= p86_array_index_1093326_comb;
    p86_array_index_1093327 <= p86_array_index_1093327_comb;
    p86_array_index_1093328 <= p86_array_index_1093328_comb;
    p86_array_index_1093329 <= p86_array_index_1093329_comb;
    p86_array_index_1093330 <= p86_array_index_1093330_comb;
    p86_array_index_1093331 <= p86_array_index_1093331_comb;
    p86_array_index_1093332 <= p86_array_index_1093332_comb;
    p86_array_index_1093333 <= p86_array_index_1093333_comb;
    p86_array_index_1093334 <= p86_array_index_1093334_comb;
    p86_res__39 <= p85_res__39;
    p87_arr <= p86_arr;
    p87_literal_1076345 <= p86_literal_1076345;
    p87_literal_1076347 <= p86_literal_1076347;
    p87_literal_1076349 <= p86_literal_1076349;
    p87_literal_1076351 <= p86_literal_1076351;
    p87_literal_1076353 <= p86_literal_1076353;
    p87_literal_1076355 <= p86_literal_1076355;
    p87_literal_1076358 <= p86_literal_1076358;
  end

  // ===== Pipe stage 87:
  wire [7:0] p87_res7__458_comb;
  wire [7:0] p87_array_index_1093469_comb;
  wire [7:0] p87_res7__459_comb;
  wire [7:0] p87_res7__460_comb;
  wire [7:0] p87_res7__461_comb;
  wire [7:0] p87_res7__462_comb;
  wire [7:0] p87_res7__463_comb;
  wire [127:0] p87_res__28_comb;
  wire [127:0] p87_xor_1093509_comb;
  assign p87_res7__458_comb = p86_array_index_1093326 ^ p86_array_index_1093327 ^ p86_array_index_1093328 ^ p86_array_index_1093329 ^ p86_array_index_1093330 ^ p86_array_index_1093331 ^ p86_res7__451 ^ p86_array_index_1093332 ^ p86_res7__449 ^ p86_array_index_1093285 ^ p86_array_index_1093154 ^ p86_array_index_1093125 ^ p86_array_index_1093093 ^ p86_array_index_1093333 ^ p86_array_index_1093334 ^ p86_array_index_1093080;
  assign p87_array_index_1093469_comb = p86_literal_1076355[p86_res7__453];
  assign p87_res7__459_comb = p86_literal_1076345[p87_res7__458_comb] ^ p86_literal_1076347[p86_res7__457] ^ p86_literal_1076349[p86_res7__456] ^ p86_literal_1076351[p86_res7__455] ^ p86_literal_1076353[p86_res7__454] ^ p87_array_index_1093469_comb ^ p86_res7__452 ^ p86_literal_1076358[p86_res7__451] ^ p86_res7__450 ^ p86_array_index_1093297 ^ p86_array_index_1093271 ^ p86_array_index_1093139 ^ p86_array_index_1093110 ^ p86_literal_1076347[p86_array_index_1093077] ^ p86_literal_1076345[p86_array_index_1093078] ^ p86_array_index_1093079;
  assign p87_res7__460_comb = p86_literal_1076345[p87_res7__459_comb] ^ p86_literal_1076347[p87_res7__458_comb] ^ p86_literal_1076349[p86_res7__457] ^ p86_literal_1076351[p86_res7__456] ^ p86_literal_1076353[p86_res7__455] ^ p86_literal_1076355[p86_res7__454] ^ p86_res7__453 ^ p86_literal_1076358[p86_res7__452] ^ p86_res7__451 ^ p86_array_index_1093309 ^ p86_array_index_1093284 ^ p86_array_index_1093153 ^ p86_array_index_1093124 ^ p86_array_index_1093092 ^ p86_literal_1076345[p86_array_index_1093077] ^ p86_array_index_1093078;
  assign p87_res7__461_comb = p86_literal_1076345[p87_res7__460_comb] ^ p86_literal_1076347[p87_res7__459_comb] ^ p86_literal_1076349[p87_res7__458_comb] ^ p86_literal_1076351[p86_res7__457] ^ p86_literal_1076353[p86_res7__456] ^ p86_literal_1076355[p86_res7__455] ^ p86_res7__454 ^ p86_literal_1076358[p86_res7__453] ^ p86_res7__452 ^ p86_array_index_1093320 ^ p86_array_index_1093296 ^ p86_array_index_1093270 ^ p86_array_index_1093138 ^ p86_array_index_1093109 ^ p86_literal_1076345[p86_array_index_1093076] ^ p86_array_index_1093077;
  assign p87_res7__462_comb = p86_literal_1076345[p87_res7__461_comb] ^ p86_literal_1076347[p87_res7__460_comb] ^ p86_literal_1076349[p87_res7__459_comb] ^ p86_literal_1076351[p87_res7__458_comb] ^ p86_literal_1076353[p86_res7__457] ^ p86_literal_1076355[p86_res7__456] ^ p86_res7__455 ^ p86_literal_1076358[p86_res7__454] ^ p86_res7__453 ^ p86_array_index_1093331 ^ p86_array_index_1093308 ^ p86_array_index_1093283 ^ p86_array_index_1093152 ^ p86_array_index_1093123 ^ p86_array_index_1093091 ^ p86_array_index_1093076;
  assign p87_res7__463_comb = p86_literal_1076345[p87_res7__462_comb] ^ p86_literal_1076347[p87_res7__461_comb] ^ p86_literal_1076349[p87_res7__460_comb] ^ p86_literal_1076351[p87_res7__459_comb] ^ p86_literal_1076353[p87_res7__458_comb] ^ p86_literal_1076355[p86_res7__457] ^ p86_res7__456 ^ p86_literal_1076358[p86_res7__455] ^ p86_res7__454 ^ p87_array_index_1093469_comb ^ p86_array_index_1093319 ^ p86_array_index_1093295 ^ p86_array_index_1093269 ^ p86_array_index_1093137 ^ p86_array_index_1093108 ^ p86_array_index_1093075;
  assign p87_res__28_comb = {p87_res7__463_comb, p87_res7__462_comb, p87_res7__461_comb, p87_res7__460_comb, p87_res7__459_comb, p87_res7__458_comb, p86_res7__457, p86_res7__456, p86_res7__455, p86_res7__454, p86_res7__453, p86_res7__452, p86_res7__451, p86_res7__450, p86_res7__449, p86_res7__448};
  assign p87_xor_1093509_comb = p87_res__28_comb ^ p86_xor_1092565;

  // Registers for pipe stage 87:
  reg [127:0] p87_xor_1093037;
  reg [127:0] p87_xor_1093509;
  reg [127:0] p87_res__39;
  reg [7:0] p88_arr[256];
  reg [7:0] p88_literal_1076345[256];
  reg [7:0] p88_literal_1076347[256];
  reg [7:0] p88_literal_1076349[256];
  reg [7:0] p88_literal_1076351[256];
  reg [7:0] p88_literal_1076353[256];
  reg [7:0] p88_literal_1076355[256];
  reg [7:0] p88_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p87_xor_1093037 <= p86_xor_1093037;
    p87_xor_1093509 <= p87_xor_1093509_comb;
    p87_res__39 <= p86_res__39;
    p88_arr <= p87_arr;
    p88_literal_1076345 <= p87_literal_1076345;
    p88_literal_1076347 <= p87_literal_1076347;
    p88_literal_1076349 <= p87_literal_1076349;
    p88_literal_1076351 <= p87_literal_1076351;
    p88_literal_1076353 <= p87_literal_1076353;
    p88_literal_1076355 <= p87_literal_1076355;
    p88_literal_1076358 <= p87_literal_1076358;
  end

  // ===== Pipe stage 88:
  wire [127:0] p88_addedKey__70_comb;
  wire [7:0] p88_array_index_1093547_comb;
  wire [7:0] p88_array_index_1093548_comb;
  wire [7:0] p88_array_index_1093549_comb;
  wire [7:0] p88_array_index_1093550_comb;
  wire [7:0] p88_array_index_1093551_comb;
  wire [7:0] p88_array_index_1093552_comb;
  wire [7:0] p88_array_index_1093554_comb;
  wire [7:0] p88_array_index_1093556_comb;
  wire [7:0] p88_array_index_1093557_comb;
  wire [7:0] p88_array_index_1093558_comb;
  wire [7:0] p88_array_index_1093559_comb;
  wire [7:0] p88_array_index_1093560_comb;
  wire [7:0] p88_array_index_1093561_comb;
  wire [7:0] p88_array_index_1093563_comb;
  wire [7:0] p88_array_index_1093564_comb;
  wire [7:0] p88_array_index_1093565_comb;
  wire [7:0] p88_array_index_1093566_comb;
  wire [7:0] p88_array_index_1093567_comb;
  wire [7:0] p88_array_index_1093568_comb;
  wire [7:0] p88_array_index_1093569_comb;
  wire [7:0] p88_array_index_1093571_comb;
  wire [7:0] p88_res7__464_comb;
  wire [7:0] p88_array_index_1093580_comb;
  wire [7:0] p88_array_index_1093581_comb;
  wire [7:0] p88_array_index_1093582_comb;
  wire [7:0] p88_array_index_1093583_comb;
  wire [7:0] p88_array_index_1093584_comb;
  wire [7:0] p88_array_index_1093585_comb;
  wire [7:0] p88_res7__465_comb;
  wire [7:0] p88_array_index_1093595_comb;
  wire [7:0] p88_array_index_1093596_comb;
  wire [7:0] p88_array_index_1093597_comb;
  wire [7:0] p88_array_index_1093598_comb;
  wire [7:0] p88_array_index_1093599_comb;
  wire [7:0] p88_res7__466_comb;
  wire [7:0] p88_array_index_1093609_comb;
  wire [7:0] p88_array_index_1093610_comb;
  wire [7:0] p88_array_index_1093611_comb;
  wire [7:0] p88_array_index_1093612_comb;
  wire [7:0] p88_array_index_1093613_comb;
  wire [7:0] p88_res7__467_comb;
  wire [7:0] p88_array_index_1093624_comb;
  wire [7:0] p88_array_index_1093625_comb;
  wire [7:0] p88_array_index_1093626_comb;
  wire [7:0] p88_array_index_1093627_comb;
  wire [7:0] p88_res7__468_comb;
  assign p88_addedKey__70_comb = p87_xor_1093509 ^ 128'h7ea1_add5_427c_254e_391c_2823_e2a3_801e;
  assign p88_array_index_1093547_comb = p87_arr[p88_addedKey__70_comb[127:120]];
  assign p88_array_index_1093548_comb = p87_arr[p88_addedKey__70_comb[119:112]];
  assign p88_array_index_1093549_comb = p87_arr[p88_addedKey__70_comb[111:104]];
  assign p88_array_index_1093550_comb = p87_arr[p88_addedKey__70_comb[103:96]];
  assign p88_array_index_1093551_comb = p87_arr[p88_addedKey__70_comb[95:88]];
  assign p88_array_index_1093552_comb = p87_arr[p88_addedKey__70_comb[87:80]];
  assign p88_array_index_1093554_comb = p87_arr[p88_addedKey__70_comb[71:64]];
  assign p88_array_index_1093556_comb = p87_arr[p88_addedKey__70_comb[55:48]];
  assign p88_array_index_1093557_comb = p87_arr[p88_addedKey__70_comb[47:40]];
  assign p88_array_index_1093558_comb = p87_arr[p88_addedKey__70_comb[39:32]];
  assign p88_array_index_1093559_comb = p87_arr[p88_addedKey__70_comb[31:24]];
  assign p88_array_index_1093560_comb = p87_arr[p88_addedKey__70_comb[23:16]];
  assign p88_array_index_1093561_comb = p87_arr[p88_addedKey__70_comb[15:8]];
  assign p88_array_index_1093563_comb = p87_literal_1076345[p88_array_index_1093547_comb];
  assign p88_array_index_1093564_comb = p87_literal_1076347[p88_array_index_1093548_comb];
  assign p88_array_index_1093565_comb = p87_literal_1076349[p88_array_index_1093549_comb];
  assign p88_array_index_1093566_comb = p87_literal_1076351[p88_array_index_1093550_comb];
  assign p88_array_index_1093567_comb = p87_literal_1076353[p88_array_index_1093551_comb];
  assign p88_array_index_1093568_comb = p87_literal_1076355[p88_array_index_1093552_comb];
  assign p88_array_index_1093569_comb = p87_arr[p88_addedKey__70_comb[79:72]];
  assign p88_array_index_1093571_comb = p87_arr[p88_addedKey__70_comb[63:56]];
  assign p88_res7__464_comb = p88_array_index_1093563_comb ^ p88_array_index_1093564_comb ^ p88_array_index_1093565_comb ^ p88_array_index_1093566_comb ^ p88_array_index_1093567_comb ^ p88_array_index_1093568_comb ^ p88_array_index_1093569_comb ^ p87_literal_1076358[p88_array_index_1093554_comb] ^ p88_array_index_1093571_comb ^ p87_literal_1076355[p88_array_index_1093556_comb] ^ p87_literal_1076353[p88_array_index_1093557_comb] ^ p87_literal_1076351[p88_array_index_1093558_comb] ^ p87_literal_1076349[p88_array_index_1093559_comb] ^ p87_literal_1076347[p88_array_index_1093560_comb] ^ p87_literal_1076345[p88_array_index_1093561_comb] ^ p87_arr[p88_addedKey__70_comb[7:0]];
  assign p88_array_index_1093580_comb = p87_literal_1076345[p88_res7__464_comb];
  assign p88_array_index_1093581_comb = p87_literal_1076347[p88_array_index_1093547_comb];
  assign p88_array_index_1093582_comb = p87_literal_1076349[p88_array_index_1093548_comb];
  assign p88_array_index_1093583_comb = p87_literal_1076351[p88_array_index_1093549_comb];
  assign p88_array_index_1093584_comb = p87_literal_1076353[p88_array_index_1093550_comb];
  assign p88_array_index_1093585_comb = p87_literal_1076355[p88_array_index_1093551_comb];
  assign p88_res7__465_comb = p88_array_index_1093580_comb ^ p88_array_index_1093581_comb ^ p88_array_index_1093582_comb ^ p88_array_index_1093583_comb ^ p88_array_index_1093584_comb ^ p88_array_index_1093585_comb ^ p88_array_index_1093552_comb ^ p87_literal_1076358[p88_array_index_1093569_comb] ^ p88_array_index_1093554_comb ^ p87_literal_1076355[p88_array_index_1093571_comb] ^ p87_literal_1076353[p88_array_index_1093556_comb] ^ p87_literal_1076351[p88_array_index_1093557_comb] ^ p87_literal_1076349[p88_array_index_1093558_comb] ^ p87_literal_1076347[p88_array_index_1093559_comb] ^ p87_literal_1076345[p88_array_index_1093560_comb] ^ p88_array_index_1093561_comb;
  assign p88_array_index_1093595_comb = p87_literal_1076347[p88_res7__464_comb];
  assign p88_array_index_1093596_comb = p87_literal_1076349[p88_array_index_1093547_comb];
  assign p88_array_index_1093597_comb = p87_literal_1076351[p88_array_index_1093548_comb];
  assign p88_array_index_1093598_comb = p87_literal_1076353[p88_array_index_1093549_comb];
  assign p88_array_index_1093599_comb = p87_literal_1076355[p88_array_index_1093550_comb];
  assign p88_res7__466_comb = p87_literal_1076345[p88_res7__465_comb] ^ p88_array_index_1093595_comb ^ p88_array_index_1093596_comb ^ p88_array_index_1093597_comb ^ p88_array_index_1093598_comb ^ p88_array_index_1093599_comb ^ p88_array_index_1093551_comb ^ p87_literal_1076358[p88_array_index_1093552_comb] ^ p88_array_index_1093569_comb ^ p87_literal_1076355[p88_array_index_1093554_comb] ^ p87_literal_1076353[p88_array_index_1093571_comb] ^ p87_literal_1076351[p88_array_index_1093556_comb] ^ p87_literal_1076349[p88_array_index_1093557_comb] ^ p87_literal_1076347[p88_array_index_1093558_comb] ^ p87_literal_1076345[p88_array_index_1093559_comb] ^ p88_array_index_1093560_comb;
  assign p88_array_index_1093609_comb = p87_literal_1076347[p88_res7__465_comb];
  assign p88_array_index_1093610_comb = p87_literal_1076349[p88_res7__464_comb];
  assign p88_array_index_1093611_comb = p87_literal_1076351[p88_array_index_1093547_comb];
  assign p88_array_index_1093612_comb = p87_literal_1076353[p88_array_index_1093548_comb];
  assign p88_array_index_1093613_comb = p87_literal_1076355[p88_array_index_1093549_comb];
  assign p88_res7__467_comb = p87_literal_1076345[p88_res7__466_comb] ^ p88_array_index_1093609_comb ^ p88_array_index_1093610_comb ^ p88_array_index_1093611_comb ^ p88_array_index_1093612_comb ^ p88_array_index_1093613_comb ^ p88_array_index_1093550_comb ^ p87_literal_1076358[p88_array_index_1093551_comb] ^ p88_array_index_1093552_comb ^ p87_literal_1076355[p88_array_index_1093569_comb] ^ p87_literal_1076353[p88_array_index_1093554_comb] ^ p87_literal_1076351[p88_array_index_1093571_comb] ^ p87_literal_1076349[p88_array_index_1093556_comb] ^ p87_literal_1076347[p88_array_index_1093557_comb] ^ p87_literal_1076345[p88_array_index_1093558_comb] ^ p88_array_index_1093559_comb;
  assign p88_array_index_1093624_comb = p87_literal_1076349[p88_res7__465_comb];
  assign p88_array_index_1093625_comb = p87_literal_1076351[p88_res7__464_comb];
  assign p88_array_index_1093626_comb = p87_literal_1076353[p88_array_index_1093547_comb];
  assign p88_array_index_1093627_comb = p87_literal_1076355[p88_array_index_1093548_comb];
  assign p88_res7__468_comb = p87_literal_1076345[p88_res7__467_comb] ^ p87_literal_1076347[p88_res7__466_comb] ^ p88_array_index_1093624_comb ^ p88_array_index_1093625_comb ^ p88_array_index_1093626_comb ^ p88_array_index_1093627_comb ^ p88_array_index_1093549_comb ^ p87_literal_1076358[p88_array_index_1093550_comb] ^ p88_array_index_1093551_comb ^ p88_array_index_1093568_comb ^ p87_literal_1076353[p88_array_index_1093569_comb] ^ p87_literal_1076351[p88_array_index_1093554_comb] ^ p87_literal_1076349[p88_array_index_1093571_comb] ^ p87_literal_1076347[p88_array_index_1093556_comb] ^ p87_literal_1076345[p88_array_index_1093557_comb] ^ p88_array_index_1093558_comb;

  // Registers for pipe stage 88:
  reg [127:0] p88_xor_1093037;
  reg [127:0] p88_xor_1093509;
  reg [7:0] p88_array_index_1093547;
  reg [7:0] p88_array_index_1093548;
  reg [7:0] p88_array_index_1093549;
  reg [7:0] p88_array_index_1093550;
  reg [7:0] p88_array_index_1093551;
  reg [7:0] p88_array_index_1093552;
  reg [7:0] p88_array_index_1093554;
  reg [7:0] p88_array_index_1093556;
  reg [7:0] p88_array_index_1093557;
  reg [7:0] p88_array_index_1093563;
  reg [7:0] p88_array_index_1093564;
  reg [7:0] p88_array_index_1093565;
  reg [7:0] p88_array_index_1093566;
  reg [7:0] p88_array_index_1093567;
  reg [7:0] p88_array_index_1093569;
  reg [7:0] p88_array_index_1093571;
  reg [7:0] p88_res7__464;
  reg [7:0] p88_array_index_1093580;
  reg [7:0] p88_array_index_1093581;
  reg [7:0] p88_array_index_1093582;
  reg [7:0] p88_array_index_1093583;
  reg [7:0] p88_array_index_1093584;
  reg [7:0] p88_array_index_1093585;
  reg [7:0] p88_res7__465;
  reg [7:0] p88_array_index_1093595;
  reg [7:0] p88_array_index_1093596;
  reg [7:0] p88_array_index_1093597;
  reg [7:0] p88_array_index_1093598;
  reg [7:0] p88_array_index_1093599;
  reg [7:0] p88_res7__466;
  reg [7:0] p88_array_index_1093609;
  reg [7:0] p88_array_index_1093610;
  reg [7:0] p88_array_index_1093611;
  reg [7:0] p88_array_index_1093612;
  reg [7:0] p88_array_index_1093613;
  reg [7:0] p88_res7__467;
  reg [7:0] p88_array_index_1093624;
  reg [7:0] p88_array_index_1093625;
  reg [7:0] p88_array_index_1093626;
  reg [7:0] p88_array_index_1093627;
  reg [7:0] p88_res7__468;
  reg [127:0] p88_res__39;
  reg [7:0] p89_arr[256];
  reg [7:0] p89_literal_1076345[256];
  reg [7:0] p89_literal_1076347[256];
  reg [7:0] p89_literal_1076349[256];
  reg [7:0] p89_literal_1076351[256];
  reg [7:0] p89_literal_1076353[256];
  reg [7:0] p89_literal_1076355[256];
  reg [7:0] p89_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p88_xor_1093037 <= p87_xor_1093037;
    p88_xor_1093509 <= p87_xor_1093509;
    p88_array_index_1093547 <= p88_array_index_1093547_comb;
    p88_array_index_1093548 <= p88_array_index_1093548_comb;
    p88_array_index_1093549 <= p88_array_index_1093549_comb;
    p88_array_index_1093550 <= p88_array_index_1093550_comb;
    p88_array_index_1093551 <= p88_array_index_1093551_comb;
    p88_array_index_1093552 <= p88_array_index_1093552_comb;
    p88_array_index_1093554 <= p88_array_index_1093554_comb;
    p88_array_index_1093556 <= p88_array_index_1093556_comb;
    p88_array_index_1093557 <= p88_array_index_1093557_comb;
    p88_array_index_1093563 <= p88_array_index_1093563_comb;
    p88_array_index_1093564 <= p88_array_index_1093564_comb;
    p88_array_index_1093565 <= p88_array_index_1093565_comb;
    p88_array_index_1093566 <= p88_array_index_1093566_comb;
    p88_array_index_1093567 <= p88_array_index_1093567_comb;
    p88_array_index_1093569 <= p88_array_index_1093569_comb;
    p88_array_index_1093571 <= p88_array_index_1093571_comb;
    p88_res7__464 <= p88_res7__464_comb;
    p88_array_index_1093580 <= p88_array_index_1093580_comb;
    p88_array_index_1093581 <= p88_array_index_1093581_comb;
    p88_array_index_1093582 <= p88_array_index_1093582_comb;
    p88_array_index_1093583 <= p88_array_index_1093583_comb;
    p88_array_index_1093584 <= p88_array_index_1093584_comb;
    p88_array_index_1093585 <= p88_array_index_1093585_comb;
    p88_res7__465 <= p88_res7__465_comb;
    p88_array_index_1093595 <= p88_array_index_1093595_comb;
    p88_array_index_1093596 <= p88_array_index_1093596_comb;
    p88_array_index_1093597 <= p88_array_index_1093597_comb;
    p88_array_index_1093598 <= p88_array_index_1093598_comb;
    p88_array_index_1093599 <= p88_array_index_1093599_comb;
    p88_res7__466 <= p88_res7__466_comb;
    p88_array_index_1093609 <= p88_array_index_1093609_comb;
    p88_array_index_1093610 <= p88_array_index_1093610_comb;
    p88_array_index_1093611 <= p88_array_index_1093611_comb;
    p88_array_index_1093612 <= p88_array_index_1093612_comb;
    p88_array_index_1093613 <= p88_array_index_1093613_comb;
    p88_res7__467 <= p88_res7__467_comb;
    p88_array_index_1093624 <= p88_array_index_1093624_comb;
    p88_array_index_1093625 <= p88_array_index_1093625_comb;
    p88_array_index_1093626 <= p88_array_index_1093626_comb;
    p88_array_index_1093627 <= p88_array_index_1093627_comb;
    p88_res7__468 <= p88_res7__468_comb;
    p88_res__39 <= p87_res__39;
    p89_arr <= p88_arr;
    p89_literal_1076345 <= p88_literal_1076345;
    p89_literal_1076347 <= p88_literal_1076347;
    p89_literal_1076349 <= p88_literal_1076349;
    p89_literal_1076351 <= p88_literal_1076351;
    p89_literal_1076353 <= p88_literal_1076353;
    p89_literal_1076355 <= p88_literal_1076355;
    p89_literal_1076358 <= p88_literal_1076358;
  end

  // ===== Pipe stage 89:
  wire [7:0] p89_array_index_1093741_comb;
  wire [7:0] p89_array_index_1093742_comb;
  wire [7:0] p89_array_index_1093743_comb;
  wire [7:0] p89_array_index_1093744_comb;
  wire [7:0] p89_res7__469_comb;
  wire [7:0] p89_array_index_1093755_comb;
  wire [7:0] p89_array_index_1093756_comb;
  wire [7:0] p89_array_index_1093757_comb;
  wire [7:0] p89_res7__470_comb;
  wire [7:0] p89_array_index_1093767_comb;
  wire [7:0] p89_array_index_1093768_comb;
  wire [7:0] p89_array_index_1093769_comb;
  wire [7:0] p89_res7__471_comb;
  wire [7:0] p89_array_index_1093780_comb;
  wire [7:0] p89_array_index_1093781_comb;
  wire [7:0] p89_res7__472_comb;
  wire [7:0] p89_array_index_1093791_comb;
  wire [7:0] p89_array_index_1093792_comb;
  wire [7:0] p89_res7__473_comb;
  wire [7:0] p89_array_index_1093798_comb;
  wire [7:0] p89_array_index_1093799_comb;
  wire [7:0] p89_array_index_1093800_comb;
  wire [7:0] p89_array_index_1093801_comb;
  wire [7:0] p89_array_index_1093802_comb;
  wire [7:0] p89_array_index_1093803_comb;
  wire [7:0] p89_array_index_1093804_comb;
  wire [7:0] p89_array_index_1093805_comb;
  wire [7:0] p89_array_index_1093806_comb;
  assign p89_array_index_1093741_comb = p88_literal_1076349[p88_res7__466];
  assign p89_array_index_1093742_comb = p88_literal_1076351[p88_res7__465];
  assign p89_array_index_1093743_comb = p88_literal_1076353[p88_res7__464];
  assign p89_array_index_1093744_comb = p88_literal_1076355[p88_array_index_1093547];
  assign p89_res7__469_comb = p88_literal_1076345[p88_res7__468] ^ p88_literal_1076347[p88_res7__467] ^ p89_array_index_1093741_comb ^ p89_array_index_1093742_comb ^ p89_array_index_1093743_comb ^ p89_array_index_1093744_comb ^ p88_array_index_1093548 ^ p88_literal_1076358[p88_array_index_1093549] ^ p88_array_index_1093550 ^ p88_array_index_1093585 ^ p88_literal_1076353[p88_array_index_1093552] ^ p88_literal_1076351[p88_array_index_1093569] ^ p88_literal_1076349[p88_array_index_1093554] ^ p88_literal_1076347[p88_array_index_1093571] ^ p88_literal_1076345[p88_array_index_1093556] ^ p88_array_index_1093557;
  assign p89_array_index_1093755_comb = p88_literal_1076351[p88_res7__466];
  assign p89_array_index_1093756_comb = p88_literal_1076353[p88_res7__465];
  assign p89_array_index_1093757_comb = p88_literal_1076355[p88_res7__464];
  assign p89_res7__470_comb = p88_literal_1076345[p89_res7__469_comb] ^ p88_literal_1076347[p88_res7__468] ^ p88_literal_1076349[p88_res7__467] ^ p89_array_index_1093755_comb ^ p89_array_index_1093756_comb ^ p89_array_index_1093757_comb ^ p88_array_index_1093547 ^ p88_literal_1076358[p88_array_index_1093548] ^ p88_array_index_1093549 ^ p88_array_index_1093599 ^ p88_array_index_1093567 ^ p88_literal_1076351[p88_array_index_1093552] ^ p88_literal_1076349[p88_array_index_1093569] ^ p88_literal_1076347[p88_array_index_1093554] ^ p88_literal_1076345[p88_array_index_1093571] ^ p88_array_index_1093556;
  assign p89_array_index_1093767_comb = p88_literal_1076351[p88_res7__467];
  assign p89_array_index_1093768_comb = p88_literal_1076353[p88_res7__466];
  assign p89_array_index_1093769_comb = p88_literal_1076355[p88_res7__465];
  assign p89_res7__471_comb = p88_literal_1076345[p89_res7__470_comb] ^ p88_literal_1076347[p89_res7__469_comb] ^ p88_literal_1076349[p88_res7__468] ^ p89_array_index_1093767_comb ^ p89_array_index_1093768_comb ^ p89_array_index_1093769_comb ^ p88_res7__464 ^ p88_literal_1076358[p88_array_index_1093547] ^ p88_array_index_1093548 ^ p88_array_index_1093613 ^ p88_array_index_1093584 ^ p88_literal_1076351[p88_array_index_1093551] ^ p88_literal_1076349[p88_array_index_1093552] ^ p88_literal_1076347[p88_array_index_1093569] ^ p88_literal_1076345[p88_array_index_1093554] ^ p88_array_index_1093571;
  assign p89_array_index_1093780_comb = p88_literal_1076353[p88_res7__467];
  assign p89_array_index_1093781_comb = p88_literal_1076355[p88_res7__466];
  assign p89_res7__472_comb = p88_literal_1076345[p89_res7__471_comb] ^ p88_literal_1076347[p89_res7__470_comb] ^ p88_literal_1076349[p89_res7__469_comb] ^ p88_literal_1076351[p88_res7__468] ^ p89_array_index_1093780_comb ^ p89_array_index_1093781_comb ^ p88_res7__465 ^ p88_literal_1076358[p88_res7__464] ^ p88_array_index_1093547 ^ p88_array_index_1093627 ^ p88_array_index_1093598 ^ p88_array_index_1093566 ^ p88_literal_1076349[p88_array_index_1093551] ^ p88_literal_1076347[p88_array_index_1093552] ^ p88_literal_1076345[p88_array_index_1093569] ^ p88_array_index_1093554;
  assign p89_array_index_1093791_comb = p88_literal_1076353[p88_res7__468];
  assign p89_array_index_1093792_comb = p88_literal_1076355[p88_res7__467];
  assign p89_res7__473_comb = p88_literal_1076345[p89_res7__472_comb] ^ p88_literal_1076347[p89_res7__471_comb] ^ p88_literal_1076349[p89_res7__470_comb] ^ p88_literal_1076351[p89_res7__469_comb] ^ p89_array_index_1093791_comb ^ p89_array_index_1093792_comb ^ p88_res7__466 ^ p88_literal_1076358[p88_res7__465] ^ p88_res7__464 ^ p89_array_index_1093744_comb ^ p88_array_index_1093612 ^ p88_array_index_1093583 ^ p88_literal_1076349[p88_array_index_1093550] ^ p88_literal_1076347[p88_array_index_1093551] ^ p88_literal_1076345[p88_array_index_1093552] ^ p88_array_index_1093569;
  assign p89_array_index_1093798_comb = p88_literal_1076345[p89_res7__473_comb];
  assign p89_array_index_1093799_comb = p88_literal_1076347[p89_res7__472_comb];
  assign p89_array_index_1093800_comb = p88_literal_1076349[p89_res7__471_comb];
  assign p89_array_index_1093801_comb = p88_literal_1076351[p89_res7__470_comb];
  assign p89_array_index_1093802_comb = p88_literal_1076353[p89_res7__469_comb];
  assign p89_array_index_1093803_comb = p88_literal_1076355[p88_res7__468];
  assign p89_array_index_1093804_comb = p88_literal_1076358[p88_res7__466];
  assign p89_array_index_1093805_comb = p88_literal_1076347[p88_array_index_1093550];
  assign p89_array_index_1093806_comb = p88_literal_1076345[p88_array_index_1093551];

  // Registers for pipe stage 89:
  reg [127:0] p89_xor_1093037;
  reg [127:0] p89_xor_1093509;
  reg [7:0] p89_array_index_1093547;
  reg [7:0] p89_array_index_1093548;
  reg [7:0] p89_array_index_1093549;
  reg [7:0] p89_array_index_1093550;
  reg [7:0] p89_array_index_1093551;
  reg [7:0] p89_array_index_1093552;
  reg [7:0] p89_array_index_1093563;
  reg [7:0] p89_array_index_1093564;
  reg [7:0] p89_array_index_1093565;
  reg [7:0] p89_res7__464;
  reg [7:0] p89_array_index_1093580;
  reg [7:0] p89_array_index_1093581;
  reg [7:0] p89_array_index_1093582;
  reg [7:0] p89_res7__465;
  reg [7:0] p89_array_index_1093595;
  reg [7:0] p89_array_index_1093596;
  reg [7:0] p89_array_index_1093597;
  reg [7:0] p89_res7__466;
  reg [7:0] p89_array_index_1093609;
  reg [7:0] p89_array_index_1093610;
  reg [7:0] p89_array_index_1093611;
  reg [7:0] p89_res7__467;
  reg [7:0] p89_array_index_1093624;
  reg [7:0] p89_array_index_1093625;
  reg [7:0] p89_array_index_1093626;
  reg [7:0] p89_res7__468;
  reg [7:0] p89_array_index_1093741;
  reg [7:0] p89_array_index_1093742;
  reg [7:0] p89_array_index_1093743;
  reg [7:0] p89_res7__469;
  reg [7:0] p89_array_index_1093755;
  reg [7:0] p89_array_index_1093756;
  reg [7:0] p89_array_index_1093757;
  reg [7:0] p89_res7__470;
  reg [7:0] p89_array_index_1093767;
  reg [7:0] p89_array_index_1093768;
  reg [7:0] p89_array_index_1093769;
  reg [7:0] p89_res7__471;
  reg [7:0] p89_array_index_1093780;
  reg [7:0] p89_array_index_1093781;
  reg [7:0] p89_res7__472;
  reg [7:0] p89_array_index_1093791;
  reg [7:0] p89_array_index_1093792;
  reg [7:0] p89_res7__473;
  reg [7:0] p89_array_index_1093798;
  reg [7:0] p89_array_index_1093799;
  reg [7:0] p89_array_index_1093800;
  reg [7:0] p89_array_index_1093801;
  reg [7:0] p89_array_index_1093802;
  reg [7:0] p89_array_index_1093803;
  reg [7:0] p89_array_index_1093804;
  reg [7:0] p89_array_index_1093805;
  reg [7:0] p89_array_index_1093806;
  reg [127:0] p89_res__39;
  reg [7:0] p90_arr[256];
  reg [7:0] p90_literal_1076345[256];
  reg [7:0] p90_literal_1076347[256];
  reg [7:0] p90_literal_1076349[256];
  reg [7:0] p90_literal_1076351[256];
  reg [7:0] p90_literal_1076353[256];
  reg [7:0] p90_literal_1076355[256];
  reg [7:0] p90_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p89_xor_1093037 <= p88_xor_1093037;
    p89_xor_1093509 <= p88_xor_1093509;
    p89_array_index_1093547 <= p88_array_index_1093547;
    p89_array_index_1093548 <= p88_array_index_1093548;
    p89_array_index_1093549 <= p88_array_index_1093549;
    p89_array_index_1093550 <= p88_array_index_1093550;
    p89_array_index_1093551 <= p88_array_index_1093551;
    p89_array_index_1093552 <= p88_array_index_1093552;
    p89_array_index_1093563 <= p88_array_index_1093563;
    p89_array_index_1093564 <= p88_array_index_1093564;
    p89_array_index_1093565 <= p88_array_index_1093565;
    p89_res7__464 <= p88_res7__464;
    p89_array_index_1093580 <= p88_array_index_1093580;
    p89_array_index_1093581 <= p88_array_index_1093581;
    p89_array_index_1093582 <= p88_array_index_1093582;
    p89_res7__465 <= p88_res7__465;
    p89_array_index_1093595 <= p88_array_index_1093595;
    p89_array_index_1093596 <= p88_array_index_1093596;
    p89_array_index_1093597 <= p88_array_index_1093597;
    p89_res7__466 <= p88_res7__466;
    p89_array_index_1093609 <= p88_array_index_1093609;
    p89_array_index_1093610 <= p88_array_index_1093610;
    p89_array_index_1093611 <= p88_array_index_1093611;
    p89_res7__467 <= p88_res7__467;
    p89_array_index_1093624 <= p88_array_index_1093624;
    p89_array_index_1093625 <= p88_array_index_1093625;
    p89_array_index_1093626 <= p88_array_index_1093626;
    p89_res7__468 <= p88_res7__468;
    p89_array_index_1093741 <= p89_array_index_1093741_comb;
    p89_array_index_1093742 <= p89_array_index_1093742_comb;
    p89_array_index_1093743 <= p89_array_index_1093743_comb;
    p89_res7__469 <= p89_res7__469_comb;
    p89_array_index_1093755 <= p89_array_index_1093755_comb;
    p89_array_index_1093756 <= p89_array_index_1093756_comb;
    p89_array_index_1093757 <= p89_array_index_1093757_comb;
    p89_res7__470 <= p89_res7__470_comb;
    p89_array_index_1093767 <= p89_array_index_1093767_comb;
    p89_array_index_1093768 <= p89_array_index_1093768_comb;
    p89_array_index_1093769 <= p89_array_index_1093769_comb;
    p89_res7__471 <= p89_res7__471_comb;
    p89_array_index_1093780 <= p89_array_index_1093780_comb;
    p89_array_index_1093781 <= p89_array_index_1093781_comb;
    p89_res7__472 <= p89_res7__472_comb;
    p89_array_index_1093791 <= p89_array_index_1093791_comb;
    p89_array_index_1093792 <= p89_array_index_1093792_comb;
    p89_res7__473 <= p89_res7__473_comb;
    p89_array_index_1093798 <= p89_array_index_1093798_comb;
    p89_array_index_1093799 <= p89_array_index_1093799_comb;
    p89_array_index_1093800 <= p89_array_index_1093800_comb;
    p89_array_index_1093801 <= p89_array_index_1093801_comb;
    p89_array_index_1093802 <= p89_array_index_1093802_comb;
    p89_array_index_1093803 <= p89_array_index_1093803_comb;
    p89_array_index_1093804 <= p89_array_index_1093804_comb;
    p89_array_index_1093805 <= p89_array_index_1093805_comb;
    p89_array_index_1093806 <= p89_array_index_1093806_comb;
    p89_res__39 <= p88_res__39;
    p90_arr <= p89_arr;
    p90_literal_1076345 <= p89_literal_1076345;
    p90_literal_1076347 <= p89_literal_1076347;
    p90_literal_1076349 <= p89_literal_1076349;
    p90_literal_1076351 <= p89_literal_1076351;
    p90_literal_1076353 <= p89_literal_1076353;
    p90_literal_1076355 <= p89_literal_1076355;
    p90_literal_1076358 <= p89_literal_1076358;
  end

  // ===== Pipe stage 90:
  wire [7:0] p90_res7__474_comb;
  wire [7:0] p90_array_index_1093941_comb;
  wire [7:0] p90_res7__475_comb;
  wire [7:0] p90_res7__476_comb;
  wire [7:0] p90_res7__477_comb;
  wire [7:0] p90_res7__478_comb;
  wire [7:0] p90_res7__479_comb;
  wire [127:0] p90_res__29_comb;
  wire [127:0] p90_xor_1093981_comb;
  assign p90_res7__474_comb = p89_array_index_1093798 ^ p89_array_index_1093799 ^ p89_array_index_1093800 ^ p89_array_index_1093801 ^ p89_array_index_1093802 ^ p89_array_index_1093803 ^ p89_res7__467 ^ p89_array_index_1093804 ^ p89_res7__465 ^ p89_array_index_1093757 ^ p89_array_index_1093626 ^ p89_array_index_1093597 ^ p89_array_index_1093565 ^ p89_array_index_1093805 ^ p89_array_index_1093806 ^ p89_array_index_1093552;
  assign p90_array_index_1093941_comb = p89_literal_1076355[p89_res7__469];
  assign p90_res7__475_comb = p89_literal_1076345[p90_res7__474_comb] ^ p89_literal_1076347[p89_res7__473] ^ p89_literal_1076349[p89_res7__472] ^ p89_literal_1076351[p89_res7__471] ^ p89_literal_1076353[p89_res7__470] ^ p90_array_index_1093941_comb ^ p89_res7__468 ^ p89_literal_1076358[p89_res7__467] ^ p89_res7__466 ^ p89_array_index_1093769 ^ p89_array_index_1093743 ^ p89_array_index_1093611 ^ p89_array_index_1093582 ^ p89_literal_1076347[p89_array_index_1093549] ^ p89_literal_1076345[p89_array_index_1093550] ^ p89_array_index_1093551;
  assign p90_res7__476_comb = p89_literal_1076345[p90_res7__475_comb] ^ p89_literal_1076347[p90_res7__474_comb] ^ p89_literal_1076349[p89_res7__473] ^ p89_literal_1076351[p89_res7__472] ^ p89_literal_1076353[p89_res7__471] ^ p89_literal_1076355[p89_res7__470] ^ p89_res7__469 ^ p89_literal_1076358[p89_res7__468] ^ p89_res7__467 ^ p89_array_index_1093781 ^ p89_array_index_1093756 ^ p89_array_index_1093625 ^ p89_array_index_1093596 ^ p89_array_index_1093564 ^ p89_literal_1076345[p89_array_index_1093549] ^ p89_array_index_1093550;
  assign p90_res7__477_comb = p89_literal_1076345[p90_res7__476_comb] ^ p89_literal_1076347[p90_res7__475_comb] ^ p89_literal_1076349[p90_res7__474_comb] ^ p89_literal_1076351[p89_res7__473] ^ p89_literal_1076353[p89_res7__472] ^ p89_literal_1076355[p89_res7__471] ^ p89_res7__470 ^ p89_literal_1076358[p89_res7__469] ^ p89_res7__468 ^ p89_array_index_1093792 ^ p89_array_index_1093768 ^ p89_array_index_1093742 ^ p89_array_index_1093610 ^ p89_array_index_1093581 ^ p89_literal_1076345[p89_array_index_1093548] ^ p89_array_index_1093549;
  assign p90_res7__478_comb = p89_literal_1076345[p90_res7__477_comb] ^ p89_literal_1076347[p90_res7__476_comb] ^ p89_literal_1076349[p90_res7__475_comb] ^ p89_literal_1076351[p90_res7__474_comb] ^ p89_literal_1076353[p89_res7__473] ^ p89_literal_1076355[p89_res7__472] ^ p89_res7__471 ^ p89_literal_1076358[p89_res7__470] ^ p89_res7__469 ^ p89_array_index_1093803 ^ p89_array_index_1093780 ^ p89_array_index_1093755 ^ p89_array_index_1093624 ^ p89_array_index_1093595 ^ p89_array_index_1093563 ^ p89_array_index_1093548;
  assign p90_res7__479_comb = p89_literal_1076345[p90_res7__478_comb] ^ p89_literal_1076347[p90_res7__477_comb] ^ p89_literal_1076349[p90_res7__476_comb] ^ p89_literal_1076351[p90_res7__475_comb] ^ p89_literal_1076353[p90_res7__474_comb] ^ p89_literal_1076355[p89_res7__473] ^ p89_res7__472 ^ p89_literal_1076358[p89_res7__471] ^ p89_res7__470 ^ p90_array_index_1093941_comb ^ p89_array_index_1093791 ^ p89_array_index_1093767 ^ p89_array_index_1093741 ^ p89_array_index_1093609 ^ p89_array_index_1093580 ^ p89_array_index_1093547;
  assign p90_res__29_comb = {p90_res7__479_comb, p90_res7__478_comb, p90_res7__477_comb, p90_res7__476_comb, p90_res7__475_comb, p90_res7__474_comb, p89_res7__473, p89_res7__472, p89_res7__471, p89_res7__470, p89_res7__469, p89_res7__468, p89_res7__467, p89_res7__466, p89_res7__465, p89_res7__464};
  assign p90_xor_1093981_comb = p90_res__29_comb ^ p89_xor_1093037;

  // Registers for pipe stage 90:
  reg [127:0] p90_xor_1093509;
  reg [127:0] p90_xor_1093981;
  reg [127:0] p90_res__39;
  reg [7:0] p91_arr[256];
  reg [7:0] p91_literal_1076345[256];
  reg [7:0] p91_literal_1076347[256];
  reg [7:0] p91_literal_1076349[256];
  reg [7:0] p91_literal_1076351[256];
  reg [7:0] p91_literal_1076353[256];
  reg [7:0] p91_literal_1076355[256];
  reg [7:0] p91_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p90_xor_1093509 <= p89_xor_1093509;
    p90_xor_1093981 <= p90_xor_1093981_comb;
    p90_res__39 <= p89_res__39;
    p91_arr <= p90_arr;
    p91_literal_1076345 <= p90_literal_1076345;
    p91_literal_1076347 <= p90_literal_1076347;
    p91_literal_1076349 <= p90_literal_1076349;
    p91_literal_1076351 <= p90_literal_1076351;
    p91_literal_1076353 <= p90_literal_1076353;
    p91_literal_1076355 <= p90_literal_1076355;
    p91_literal_1076358 <= p90_literal_1076358;
  end

  // ===== Pipe stage 91:
  wire [127:0] p91_addedKey__71_comb;
  wire [7:0] p91_array_index_1094019_comb;
  wire [7:0] p91_array_index_1094020_comb;
  wire [7:0] p91_array_index_1094021_comb;
  wire [7:0] p91_array_index_1094022_comb;
  wire [7:0] p91_array_index_1094023_comb;
  wire [7:0] p91_array_index_1094024_comb;
  wire [7:0] p91_array_index_1094026_comb;
  wire [7:0] p91_array_index_1094028_comb;
  wire [7:0] p91_array_index_1094029_comb;
  wire [7:0] p91_array_index_1094030_comb;
  wire [7:0] p91_array_index_1094031_comb;
  wire [7:0] p91_array_index_1094032_comb;
  wire [7:0] p91_array_index_1094033_comb;
  wire [7:0] p91_array_index_1094035_comb;
  wire [7:0] p91_array_index_1094036_comb;
  wire [7:0] p91_array_index_1094037_comb;
  wire [7:0] p91_array_index_1094038_comb;
  wire [7:0] p91_array_index_1094039_comb;
  wire [7:0] p91_array_index_1094040_comb;
  wire [7:0] p91_array_index_1094041_comb;
  wire [7:0] p91_array_index_1094043_comb;
  wire [7:0] p91_res7__480_comb;
  wire [7:0] p91_array_index_1094052_comb;
  wire [7:0] p91_array_index_1094053_comb;
  wire [7:0] p91_array_index_1094054_comb;
  wire [7:0] p91_array_index_1094055_comb;
  wire [7:0] p91_array_index_1094056_comb;
  wire [7:0] p91_array_index_1094057_comb;
  wire [7:0] p91_res7__481_comb;
  wire [7:0] p91_array_index_1094067_comb;
  wire [7:0] p91_array_index_1094068_comb;
  wire [7:0] p91_array_index_1094069_comb;
  wire [7:0] p91_array_index_1094070_comb;
  wire [7:0] p91_array_index_1094071_comb;
  wire [7:0] p91_res7__482_comb;
  wire [7:0] p91_array_index_1094081_comb;
  wire [7:0] p91_array_index_1094082_comb;
  wire [7:0] p91_array_index_1094083_comb;
  wire [7:0] p91_array_index_1094084_comb;
  wire [7:0] p91_array_index_1094085_comb;
  wire [7:0] p91_res7__483_comb;
  wire [7:0] p91_array_index_1094096_comb;
  wire [7:0] p91_array_index_1094097_comb;
  wire [7:0] p91_array_index_1094098_comb;
  wire [7:0] p91_array_index_1094099_comb;
  wire [7:0] p91_res7__484_comb;
  assign p91_addedKey__71_comb = p90_xor_1093981 ^ 128'h1003_dba7_2e34_5ff6_643b_9533_3f27_141f;
  assign p91_array_index_1094019_comb = p90_arr[p91_addedKey__71_comb[127:120]];
  assign p91_array_index_1094020_comb = p90_arr[p91_addedKey__71_comb[119:112]];
  assign p91_array_index_1094021_comb = p90_arr[p91_addedKey__71_comb[111:104]];
  assign p91_array_index_1094022_comb = p90_arr[p91_addedKey__71_comb[103:96]];
  assign p91_array_index_1094023_comb = p90_arr[p91_addedKey__71_comb[95:88]];
  assign p91_array_index_1094024_comb = p90_arr[p91_addedKey__71_comb[87:80]];
  assign p91_array_index_1094026_comb = p90_arr[p91_addedKey__71_comb[71:64]];
  assign p91_array_index_1094028_comb = p90_arr[p91_addedKey__71_comb[55:48]];
  assign p91_array_index_1094029_comb = p90_arr[p91_addedKey__71_comb[47:40]];
  assign p91_array_index_1094030_comb = p90_arr[p91_addedKey__71_comb[39:32]];
  assign p91_array_index_1094031_comb = p90_arr[p91_addedKey__71_comb[31:24]];
  assign p91_array_index_1094032_comb = p90_arr[p91_addedKey__71_comb[23:16]];
  assign p91_array_index_1094033_comb = p90_arr[p91_addedKey__71_comb[15:8]];
  assign p91_array_index_1094035_comb = p90_literal_1076345[p91_array_index_1094019_comb];
  assign p91_array_index_1094036_comb = p90_literal_1076347[p91_array_index_1094020_comb];
  assign p91_array_index_1094037_comb = p90_literal_1076349[p91_array_index_1094021_comb];
  assign p91_array_index_1094038_comb = p90_literal_1076351[p91_array_index_1094022_comb];
  assign p91_array_index_1094039_comb = p90_literal_1076353[p91_array_index_1094023_comb];
  assign p91_array_index_1094040_comb = p90_literal_1076355[p91_array_index_1094024_comb];
  assign p91_array_index_1094041_comb = p90_arr[p91_addedKey__71_comb[79:72]];
  assign p91_array_index_1094043_comb = p90_arr[p91_addedKey__71_comb[63:56]];
  assign p91_res7__480_comb = p91_array_index_1094035_comb ^ p91_array_index_1094036_comb ^ p91_array_index_1094037_comb ^ p91_array_index_1094038_comb ^ p91_array_index_1094039_comb ^ p91_array_index_1094040_comb ^ p91_array_index_1094041_comb ^ p90_literal_1076358[p91_array_index_1094026_comb] ^ p91_array_index_1094043_comb ^ p90_literal_1076355[p91_array_index_1094028_comb] ^ p90_literal_1076353[p91_array_index_1094029_comb] ^ p90_literal_1076351[p91_array_index_1094030_comb] ^ p90_literal_1076349[p91_array_index_1094031_comb] ^ p90_literal_1076347[p91_array_index_1094032_comb] ^ p90_literal_1076345[p91_array_index_1094033_comb] ^ p90_arr[p91_addedKey__71_comb[7:0]];
  assign p91_array_index_1094052_comb = p90_literal_1076345[p91_res7__480_comb];
  assign p91_array_index_1094053_comb = p90_literal_1076347[p91_array_index_1094019_comb];
  assign p91_array_index_1094054_comb = p90_literal_1076349[p91_array_index_1094020_comb];
  assign p91_array_index_1094055_comb = p90_literal_1076351[p91_array_index_1094021_comb];
  assign p91_array_index_1094056_comb = p90_literal_1076353[p91_array_index_1094022_comb];
  assign p91_array_index_1094057_comb = p90_literal_1076355[p91_array_index_1094023_comb];
  assign p91_res7__481_comb = p91_array_index_1094052_comb ^ p91_array_index_1094053_comb ^ p91_array_index_1094054_comb ^ p91_array_index_1094055_comb ^ p91_array_index_1094056_comb ^ p91_array_index_1094057_comb ^ p91_array_index_1094024_comb ^ p90_literal_1076358[p91_array_index_1094041_comb] ^ p91_array_index_1094026_comb ^ p90_literal_1076355[p91_array_index_1094043_comb] ^ p90_literal_1076353[p91_array_index_1094028_comb] ^ p90_literal_1076351[p91_array_index_1094029_comb] ^ p90_literal_1076349[p91_array_index_1094030_comb] ^ p90_literal_1076347[p91_array_index_1094031_comb] ^ p90_literal_1076345[p91_array_index_1094032_comb] ^ p91_array_index_1094033_comb;
  assign p91_array_index_1094067_comb = p90_literal_1076347[p91_res7__480_comb];
  assign p91_array_index_1094068_comb = p90_literal_1076349[p91_array_index_1094019_comb];
  assign p91_array_index_1094069_comb = p90_literal_1076351[p91_array_index_1094020_comb];
  assign p91_array_index_1094070_comb = p90_literal_1076353[p91_array_index_1094021_comb];
  assign p91_array_index_1094071_comb = p90_literal_1076355[p91_array_index_1094022_comb];
  assign p91_res7__482_comb = p90_literal_1076345[p91_res7__481_comb] ^ p91_array_index_1094067_comb ^ p91_array_index_1094068_comb ^ p91_array_index_1094069_comb ^ p91_array_index_1094070_comb ^ p91_array_index_1094071_comb ^ p91_array_index_1094023_comb ^ p90_literal_1076358[p91_array_index_1094024_comb] ^ p91_array_index_1094041_comb ^ p90_literal_1076355[p91_array_index_1094026_comb] ^ p90_literal_1076353[p91_array_index_1094043_comb] ^ p90_literal_1076351[p91_array_index_1094028_comb] ^ p90_literal_1076349[p91_array_index_1094029_comb] ^ p90_literal_1076347[p91_array_index_1094030_comb] ^ p90_literal_1076345[p91_array_index_1094031_comb] ^ p91_array_index_1094032_comb;
  assign p91_array_index_1094081_comb = p90_literal_1076347[p91_res7__481_comb];
  assign p91_array_index_1094082_comb = p90_literal_1076349[p91_res7__480_comb];
  assign p91_array_index_1094083_comb = p90_literal_1076351[p91_array_index_1094019_comb];
  assign p91_array_index_1094084_comb = p90_literal_1076353[p91_array_index_1094020_comb];
  assign p91_array_index_1094085_comb = p90_literal_1076355[p91_array_index_1094021_comb];
  assign p91_res7__483_comb = p90_literal_1076345[p91_res7__482_comb] ^ p91_array_index_1094081_comb ^ p91_array_index_1094082_comb ^ p91_array_index_1094083_comb ^ p91_array_index_1094084_comb ^ p91_array_index_1094085_comb ^ p91_array_index_1094022_comb ^ p90_literal_1076358[p91_array_index_1094023_comb] ^ p91_array_index_1094024_comb ^ p90_literal_1076355[p91_array_index_1094041_comb] ^ p90_literal_1076353[p91_array_index_1094026_comb] ^ p90_literal_1076351[p91_array_index_1094043_comb] ^ p90_literal_1076349[p91_array_index_1094028_comb] ^ p90_literal_1076347[p91_array_index_1094029_comb] ^ p90_literal_1076345[p91_array_index_1094030_comb] ^ p91_array_index_1094031_comb;
  assign p91_array_index_1094096_comb = p90_literal_1076349[p91_res7__481_comb];
  assign p91_array_index_1094097_comb = p90_literal_1076351[p91_res7__480_comb];
  assign p91_array_index_1094098_comb = p90_literal_1076353[p91_array_index_1094019_comb];
  assign p91_array_index_1094099_comb = p90_literal_1076355[p91_array_index_1094020_comb];
  assign p91_res7__484_comb = p90_literal_1076345[p91_res7__483_comb] ^ p90_literal_1076347[p91_res7__482_comb] ^ p91_array_index_1094096_comb ^ p91_array_index_1094097_comb ^ p91_array_index_1094098_comb ^ p91_array_index_1094099_comb ^ p91_array_index_1094021_comb ^ p90_literal_1076358[p91_array_index_1094022_comb] ^ p91_array_index_1094023_comb ^ p91_array_index_1094040_comb ^ p90_literal_1076353[p91_array_index_1094041_comb] ^ p90_literal_1076351[p91_array_index_1094026_comb] ^ p90_literal_1076349[p91_array_index_1094043_comb] ^ p90_literal_1076347[p91_array_index_1094028_comb] ^ p90_literal_1076345[p91_array_index_1094029_comb] ^ p91_array_index_1094030_comb;

  // Registers for pipe stage 91:
  reg [127:0] p91_xor_1093509;
  reg [127:0] p91_xor_1093981;
  reg [7:0] p91_array_index_1094019;
  reg [7:0] p91_array_index_1094020;
  reg [7:0] p91_array_index_1094021;
  reg [7:0] p91_array_index_1094022;
  reg [7:0] p91_array_index_1094023;
  reg [7:0] p91_array_index_1094024;
  reg [7:0] p91_array_index_1094026;
  reg [7:0] p91_array_index_1094028;
  reg [7:0] p91_array_index_1094029;
  reg [7:0] p91_array_index_1094035;
  reg [7:0] p91_array_index_1094036;
  reg [7:0] p91_array_index_1094037;
  reg [7:0] p91_array_index_1094038;
  reg [7:0] p91_array_index_1094039;
  reg [7:0] p91_array_index_1094041;
  reg [7:0] p91_array_index_1094043;
  reg [7:0] p91_res7__480;
  reg [7:0] p91_array_index_1094052;
  reg [7:0] p91_array_index_1094053;
  reg [7:0] p91_array_index_1094054;
  reg [7:0] p91_array_index_1094055;
  reg [7:0] p91_array_index_1094056;
  reg [7:0] p91_array_index_1094057;
  reg [7:0] p91_res7__481;
  reg [7:0] p91_array_index_1094067;
  reg [7:0] p91_array_index_1094068;
  reg [7:0] p91_array_index_1094069;
  reg [7:0] p91_array_index_1094070;
  reg [7:0] p91_array_index_1094071;
  reg [7:0] p91_res7__482;
  reg [7:0] p91_array_index_1094081;
  reg [7:0] p91_array_index_1094082;
  reg [7:0] p91_array_index_1094083;
  reg [7:0] p91_array_index_1094084;
  reg [7:0] p91_array_index_1094085;
  reg [7:0] p91_res7__483;
  reg [7:0] p91_array_index_1094096;
  reg [7:0] p91_array_index_1094097;
  reg [7:0] p91_array_index_1094098;
  reg [7:0] p91_array_index_1094099;
  reg [7:0] p91_res7__484;
  reg [127:0] p91_res__39;
  reg [7:0] p92_arr[256];
  reg [7:0] p92_literal_1076345[256];
  reg [7:0] p92_literal_1076347[256];
  reg [7:0] p92_literal_1076349[256];
  reg [7:0] p92_literal_1076351[256];
  reg [7:0] p92_literal_1076353[256];
  reg [7:0] p92_literal_1076355[256];
  reg [7:0] p92_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p91_xor_1093509 <= p90_xor_1093509;
    p91_xor_1093981 <= p90_xor_1093981;
    p91_array_index_1094019 <= p91_array_index_1094019_comb;
    p91_array_index_1094020 <= p91_array_index_1094020_comb;
    p91_array_index_1094021 <= p91_array_index_1094021_comb;
    p91_array_index_1094022 <= p91_array_index_1094022_comb;
    p91_array_index_1094023 <= p91_array_index_1094023_comb;
    p91_array_index_1094024 <= p91_array_index_1094024_comb;
    p91_array_index_1094026 <= p91_array_index_1094026_comb;
    p91_array_index_1094028 <= p91_array_index_1094028_comb;
    p91_array_index_1094029 <= p91_array_index_1094029_comb;
    p91_array_index_1094035 <= p91_array_index_1094035_comb;
    p91_array_index_1094036 <= p91_array_index_1094036_comb;
    p91_array_index_1094037 <= p91_array_index_1094037_comb;
    p91_array_index_1094038 <= p91_array_index_1094038_comb;
    p91_array_index_1094039 <= p91_array_index_1094039_comb;
    p91_array_index_1094041 <= p91_array_index_1094041_comb;
    p91_array_index_1094043 <= p91_array_index_1094043_comb;
    p91_res7__480 <= p91_res7__480_comb;
    p91_array_index_1094052 <= p91_array_index_1094052_comb;
    p91_array_index_1094053 <= p91_array_index_1094053_comb;
    p91_array_index_1094054 <= p91_array_index_1094054_comb;
    p91_array_index_1094055 <= p91_array_index_1094055_comb;
    p91_array_index_1094056 <= p91_array_index_1094056_comb;
    p91_array_index_1094057 <= p91_array_index_1094057_comb;
    p91_res7__481 <= p91_res7__481_comb;
    p91_array_index_1094067 <= p91_array_index_1094067_comb;
    p91_array_index_1094068 <= p91_array_index_1094068_comb;
    p91_array_index_1094069 <= p91_array_index_1094069_comb;
    p91_array_index_1094070 <= p91_array_index_1094070_comb;
    p91_array_index_1094071 <= p91_array_index_1094071_comb;
    p91_res7__482 <= p91_res7__482_comb;
    p91_array_index_1094081 <= p91_array_index_1094081_comb;
    p91_array_index_1094082 <= p91_array_index_1094082_comb;
    p91_array_index_1094083 <= p91_array_index_1094083_comb;
    p91_array_index_1094084 <= p91_array_index_1094084_comb;
    p91_array_index_1094085 <= p91_array_index_1094085_comb;
    p91_res7__483 <= p91_res7__483_comb;
    p91_array_index_1094096 <= p91_array_index_1094096_comb;
    p91_array_index_1094097 <= p91_array_index_1094097_comb;
    p91_array_index_1094098 <= p91_array_index_1094098_comb;
    p91_array_index_1094099 <= p91_array_index_1094099_comb;
    p91_res7__484 <= p91_res7__484_comb;
    p91_res__39 <= p90_res__39;
    p92_arr <= p91_arr;
    p92_literal_1076345 <= p91_literal_1076345;
    p92_literal_1076347 <= p91_literal_1076347;
    p92_literal_1076349 <= p91_literal_1076349;
    p92_literal_1076351 <= p91_literal_1076351;
    p92_literal_1076353 <= p91_literal_1076353;
    p92_literal_1076355 <= p91_literal_1076355;
    p92_literal_1076358 <= p91_literal_1076358;
  end

  // ===== Pipe stage 92:
  wire [7:0] p92_array_index_1094213_comb;
  wire [7:0] p92_array_index_1094214_comb;
  wire [7:0] p92_array_index_1094215_comb;
  wire [7:0] p92_array_index_1094216_comb;
  wire [7:0] p92_res7__485_comb;
  wire [7:0] p92_array_index_1094227_comb;
  wire [7:0] p92_array_index_1094228_comb;
  wire [7:0] p92_array_index_1094229_comb;
  wire [7:0] p92_res7__486_comb;
  wire [7:0] p92_array_index_1094239_comb;
  wire [7:0] p92_array_index_1094240_comb;
  wire [7:0] p92_array_index_1094241_comb;
  wire [7:0] p92_res7__487_comb;
  wire [7:0] p92_array_index_1094252_comb;
  wire [7:0] p92_array_index_1094253_comb;
  wire [7:0] p92_res7__488_comb;
  wire [7:0] p92_array_index_1094263_comb;
  wire [7:0] p92_array_index_1094264_comb;
  wire [7:0] p92_res7__489_comb;
  wire [7:0] p92_array_index_1094270_comb;
  wire [7:0] p92_array_index_1094271_comb;
  wire [7:0] p92_array_index_1094272_comb;
  wire [7:0] p92_array_index_1094273_comb;
  wire [7:0] p92_array_index_1094274_comb;
  wire [7:0] p92_array_index_1094275_comb;
  wire [7:0] p92_array_index_1094276_comb;
  wire [7:0] p92_array_index_1094277_comb;
  wire [7:0] p92_array_index_1094278_comb;
  assign p92_array_index_1094213_comb = p91_literal_1076349[p91_res7__482];
  assign p92_array_index_1094214_comb = p91_literal_1076351[p91_res7__481];
  assign p92_array_index_1094215_comb = p91_literal_1076353[p91_res7__480];
  assign p92_array_index_1094216_comb = p91_literal_1076355[p91_array_index_1094019];
  assign p92_res7__485_comb = p91_literal_1076345[p91_res7__484] ^ p91_literal_1076347[p91_res7__483] ^ p92_array_index_1094213_comb ^ p92_array_index_1094214_comb ^ p92_array_index_1094215_comb ^ p92_array_index_1094216_comb ^ p91_array_index_1094020 ^ p91_literal_1076358[p91_array_index_1094021] ^ p91_array_index_1094022 ^ p91_array_index_1094057 ^ p91_literal_1076353[p91_array_index_1094024] ^ p91_literal_1076351[p91_array_index_1094041] ^ p91_literal_1076349[p91_array_index_1094026] ^ p91_literal_1076347[p91_array_index_1094043] ^ p91_literal_1076345[p91_array_index_1094028] ^ p91_array_index_1094029;
  assign p92_array_index_1094227_comb = p91_literal_1076351[p91_res7__482];
  assign p92_array_index_1094228_comb = p91_literal_1076353[p91_res7__481];
  assign p92_array_index_1094229_comb = p91_literal_1076355[p91_res7__480];
  assign p92_res7__486_comb = p91_literal_1076345[p92_res7__485_comb] ^ p91_literal_1076347[p91_res7__484] ^ p91_literal_1076349[p91_res7__483] ^ p92_array_index_1094227_comb ^ p92_array_index_1094228_comb ^ p92_array_index_1094229_comb ^ p91_array_index_1094019 ^ p91_literal_1076358[p91_array_index_1094020] ^ p91_array_index_1094021 ^ p91_array_index_1094071 ^ p91_array_index_1094039 ^ p91_literal_1076351[p91_array_index_1094024] ^ p91_literal_1076349[p91_array_index_1094041] ^ p91_literal_1076347[p91_array_index_1094026] ^ p91_literal_1076345[p91_array_index_1094043] ^ p91_array_index_1094028;
  assign p92_array_index_1094239_comb = p91_literal_1076351[p91_res7__483];
  assign p92_array_index_1094240_comb = p91_literal_1076353[p91_res7__482];
  assign p92_array_index_1094241_comb = p91_literal_1076355[p91_res7__481];
  assign p92_res7__487_comb = p91_literal_1076345[p92_res7__486_comb] ^ p91_literal_1076347[p92_res7__485_comb] ^ p91_literal_1076349[p91_res7__484] ^ p92_array_index_1094239_comb ^ p92_array_index_1094240_comb ^ p92_array_index_1094241_comb ^ p91_res7__480 ^ p91_literal_1076358[p91_array_index_1094019] ^ p91_array_index_1094020 ^ p91_array_index_1094085 ^ p91_array_index_1094056 ^ p91_literal_1076351[p91_array_index_1094023] ^ p91_literal_1076349[p91_array_index_1094024] ^ p91_literal_1076347[p91_array_index_1094041] ^ p91_literal_1076345[p91_array_index_1094026] ^ p91_array_index_1094043;
  assign p92_array_index_1094252_comb = p91_literal_1076353[p91_res7__483];
  assign p92_array_index_1094253_comb = p91_literal_1076355[p91_res7__482];
  assign p92_res7__488_comb = p91_literal_1076345[p92_res7__487_comb] ^ p91_literal_1076347[p92_res7__486_comb] ^ p91_literal_1076349[p92_res7__485_comb] ^ p91_literal_1076351[p91_res7__484] ^ p92_array_index_1094252_comb ^ p92_array_index_1094253_comb ^ p91_res7__481 ^ p91_literal_1076358[p91_res7__480] ^ p91_array_index_1094019 ^ p91_array_index_1094099 ^ p91_array_index_1094070 ^ p91_array_index_1094038 ^ p91_literal_1076349[p91_array_index_1094023] ^ p91_literal_1076347[p91_array_index_1094024] ^ p91_literal_1076345[p91_array_index_1094041] ^ p91_array_index_1094026;
  assign p92_array_index_1094263_comb = p91_literal_1076353[p91_res7__484];
  assign p92_array_index_1094264_comb = p91_literal_1076355[p91_res7__483];
  assign p92_res7__489_comb = p91_literal_1076345[p92_res7__488_comb] ^ p91_literal_1076347[p92_res7__487_comb] ^ p91_literal_1076349[p92_res7__486_comb] ^ p91_literal_1076351[p92_res7__485_comb] ^ p92_array_index_1094263_comb ^ p92_array_index_1094264_comb ^ p91_res7__482 ^ p91_literal_1076358[p91_res7__481] ^ p91_res7__480 ^ p92_array_index_1094216_comb ^ p91_array_index_1094084 ^ p91_array_index_1094055 ^ p91_literal_1076349[p91_array_index_1094022] ^ p91_literal_1076347[p91_array_index_1094023] ^ p91_literal_1076345[p91_array_index_1094024] ^ p91_array_index_1094041;
  assign p92_array_index_1094270_comb = p91_literal_1076345[p92_res7__489_comb];
  assign p92_array_index_1094271_comb = p91_literal_1076347[p92_res7__488_comb];
  assign p92_array_index_1094272_comb = p91_literal_1076349[p92_res7__487_comb];
  assign p92_array_index_1094273_comb = p91_literal_1076351[p92_res7__486_comb];
  assign p92_array_index_1094274_comb = p91_literal_1076353[p92_res7__485_comb];
  assign p92_array_index_1094275_comb = p91_literal_1076355[p91_res7__484];
  assign p92_array_index_1094276_comb = p91_literal_1076358[p91_res7__482];
  assign p92_array_index_1094277_comb = p91_literal_1076347[p91_array_index_1094022];
  assign p92_array_index_1094278_comb = p91_literal_1076345[p91_array_index_1094023];

  // Registers for pipe stage 92:
  reg [127:0] p92_xor_1093509;
  reg [127:0] p92_xor_1093981;
  reg [7:0] p92_array_index_1094019;
  reg [7:0] p92_array_index_1094020;
  reg [7:0] p92_array_index_1094021;
  reg [7:0] p92_array_index_1094022;
  reg [7:0] p92_array_index_1094023;
  reg [7:0] p92_array_index_1094024;
  reg [7:0] p92_array_index_1094035;
  reg [7:0] p92_array_index_1094036;
  reg [7:0] p92_array_index_1094037;
  reg [7:0] p92_res7__480;
  reg [7:0] p92_array_index_1094052;
  reg [7:0] p92_array_index_1094053;
  reg [7:0] p92_array_index_1094054;
  reg [7:0] p92_res7__481;
  reg [7:0] p92_array_index_1094067;
  reg [7:0] p92_array_index_1094068;
  reg [7:0] p92_array_index_1094069;
  reg [7:0] p92_res7__482;
  reg [7:0] p92_array_index_1094081;
  reg [7:0] p92_array_index_1094082;
  reg [7:0] p92_array_index_1094083;
  reg [7:0] p92_res7__483;
  reg [7:0] p92_array_index_1094096;
  reg [7:0] p92_array_index_1094097;
  reg [7:0] p92_array_index_1094098;
  reg [7:0] p92_res7__484;
  reg [7:0] p92_array_index_1094213;
  reg [7:0] p92_array_index_1094214;
  reg [7:0] p92_array_index_1094215;
  reg [7:0] p92_res7__485;
  reg [7:0] p92_array_index_1094227;
  reg [7:0] p92_array_index_1094228;
  reg [7:0] p92_array_index_1094229;
  reg [7:0] p92_res7__486;
  reg [7:0] p92_array_index_1094239;
  reg [7:0] p92_array_index_1094240;
  reg [7:0] p92_array_index_1094241;
  reg [7:0] p92_res7__487;
  reg [7:0] p92_array_index_1094252;
  reg [7:0] p92_array_index_1094253;
  reg [7:0] p92_res7__488;
  reg [7:0] p92_array_index_1094263;
  reg [7:0] p92_array_index_1094264;
  reg [7:0] p92_res7__489;
  reg [7:0] p92_array_index_1094270;
  reg [7:0] p92_array_index_1094271;
  reg [7:0] p92_array_index_1094272;
  reg [7:0] p92_array_index_1094273;
  reg [7:0] p92_array_index_1094274;
  reg [7:0] p92_array_index_1094275;
  reg [7:0] p92_array_index_1094276;
  reg [7:0] p92_array_index_1094277;
  reg [7:0] p92_array_index_1094278;
  reg [127:0] p92_res__39;
  reg [7:0] p93_arr[256];
  reg [7:0] p93_literal_1076345[256];
  reg [7:0] p93_literal_1076347[256];
  reg [7:0] p93_literal_1076349[256];
  reg [7:0] p93_literal_1076351[256];
  reg [7:0] p93_literal_1076353[256];
  reg [7:0] p93_literal_1076355[256];
  reg [7:0] p93_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p92_xor_1093509 <= p91_xor_1093509;
    p92_xor_1093981 <= p91_xor_1093981;
    p92_array_index_1094019 <= p91_array_index_1094019;
    p92_array_index_1094020 <= p91_array_index_1094020;
    p92_array_index_1094021 <= p91_array_index_1094021;
    p92_array_index_1094022 <= p91_array_index_1094022;
    p92_array_index_1094023 <= p91_array_index_1094023;
    p92_array_index_1094024 <= p91_array_index_1094024;
    p92_array_index_1094035 <= p91_array_index_1094035;
    p92_array_index_1094036 <= p91_array_index_1094036;
    p92_array_index_1094037 <= p91_array_index_1094037;
    p92_res7__480 <= p91_res7__480;
    p92_array_index_1094052 <= p91_array_index_1094052;
    p92_array_index_1094053 <= p91_array_index_1094053;
    p92_array_index_1094054 <= p91_array_index_1094054;
    p92_res7__481 <= p91_res7__481;
    p92_array_index_1094067 <= p91_array_index_1094067;
    p92_array_index_1094068 <= p91_array_index_1094068;
    p92_array_index_1094069 <= p91_array_index_1094069;
    p92_res7__482 <= p91_res7__482;
    p92_array_index_1094081 <= p91_array_index_1094081;
    p92_array_index_1094082 <= p91_array_index_1094082;
    p92_array_index_1094083 <= p91_array_index_1094083;
    p92_res7__483 <= p91_res7__483;
    p92_array_index_1094096 <= p91_array_index_1094096;
    p92_array_index_1094097 <= p91_array_index_1094097;
    p92_array_index_1094098 <= p91_array_index_1094098;
    p92_res7__484 <= p91_res7__484;
    p92_array_index_1094213 <= p92_array_index_1094213_comb;
    p92_array_index_1094214 <= p92_array_index_1094214_comb;
    p92_array_index_1094215 <= p92_array_index_1094215_comb;
    p92_res7__485 <= p92_res7__485_comb;
    p92_array_index_1094227 <= p92_array_index_1094227_comb;
    p92_array_index_1094228 <= p92_array_index_1094228_comb;
    p92_array_index_1094229 <= p92_array_index_1094229_comb;
    p92_res7__486 <= p92_res7__486_comb;
    p92_array_index_1094239 <= p92_array_index_1094239_comb;
    p92_array_index_1094240 <= p92_array_index_1094240_comb;
    p92_array_index_1094241 <= p92_array_index_1094241_comb;
    p92_res7__487 <= p92_res7__487_comb;
    p92_array_index_1094252 <= p92_array_index_1094252_comb;
    p92_array_index_1094253 <= p92_array_index_1094253_comb;
    p92_res7__488 <= p92_res7__488_comb;
    p92_array_index_1094263 <= p92_array_index_1094263_comb;
    p92_array_index_1094264 <= p92_array_index_1094264_comb;
    p92_res7__489 <= p92_res7__489_comb;
    p92_array_index_1094270 <= p92_array_index_1094270_comb;
    p92_array_index_1094271 <= p92_array_index_1094271_comb;
    p92_array_index_1094272 <= p92_array_index_1094272_comb;
    p92_array_index_1094273 <= p92_array_index_1094273_comb;
    p92_array_index_1094274 <= p92_array_index_1094274_comb;
    p92_array_index_1094275 <= p92_array_index_1094275_comb;
    p92_array_index_1094276 <= p92_array_index_1094276_comb;
    p92_array_index_1094277 <= p92_array_index_1094277_comb;
    p92_array_index_1094278 <= p92_array_index_1094278_comb;
    p92_res__39 <= p91_res__39;
    p93_arr <= p92_arr;
    p93_literal_1076345 <= p92_literal_1076345;
    p93_literal_1076347 <= p92_literal_1076347;
    p93_literal_1076349 <= p92_literal_1076349;
    p93_literal_1076351 <= p92_literal_1076351;
    p93_literal_1076353 <= p92_literal_1076353;
    p93_literal_1076355 <= p92_literal_1076355;
    p93_literal_1076358 <= p92_literal_1076358;
  end

  // ===== Pipe stage 93:
  wire [7:0] p93_res7__490_comb;
  wire [7:0] p93_array_index_1094413_comb;
  wire [7:0] p93_res7__491_comb;
  wire [7:0] p93_res7__492_comb;
  wire [7:0] p93_res7__493_comb;
  wire [7:0] p93_res7__494_comb;
  wire [7:0] p93_res7__495_comb;
  wire [127:0] p93_res__30_comb;
  wire [127:0] p93_k9_comb;
  assign p93_res7__490_comb = p92_array_index_1094270 ^ p92_array_index_1094271 ^ p92_array_index_1094272 ^ p92_array_index_1094273 ^ p92_array_index_1094274 ^ p92_array_index_1094275 ^ p92_res7__483 ^ p92_array_index_1094276 ^ p92_res7__481 ^ p92_array_index_1094229 ^ p92_array_index_1094098 ^ p92_array_index_1094069 ^ p92_array_index_1094037 ^ p92_array_index_1094277 ^ p92_array_index_1094278 ^ p92_array_index_1094024;
  assign p93_array_index_1094413_comb = p92_literal_1076355[p92_res7__485];
  assign p93_res7__491_comb = p92_literal_1076345[p93_res7__490_comb] ^ p92_literal_1076347[p92_res7__489] ^ p92_literal_1076349[p92_res7__488] ^ p92_literal_1076351[p92_res7__487] ^ p92_literal_1076353[p92_res7__486] ^ p93_array_index_1094413_comb ^ p92_res7__484 ^ p92_literal_1076358[p92_res7__483] ^ p92_res7__482 ^ p92_array_index_1094241 ^ p92_array_index_1094215 ^ p92_array_index_1094083 ^ p92_array_index_1094054 ^ p92_literal_1076347[p92_array_index_1094021] ^ p92_literal_1076345[p92_array_index_1094022] ^ p92_array_index_1094023;
  assign p93_res7__492_comb = p92_literal_1076345[p93_res7__491_comb] ^ p92_literal_1076347[p93_res7__490_comb] ^ p92_literal_1076349[p92_res7__489] ^ p92_literal_1076351[p92_res7__488] ^ p92_literal_1076353[p92_res7__487] ^ p92_literal_1076355[p92_res7__486] ^ p92_res7__485 ^ p92_literal_1076358[p92_res7__484] ^ p92_res7__483 ^ p92_array_index_1094253 ^ p92_array_index_1094228 ^ p92_array_index_1094097 ^ p92_array_index_1094068 ^ p92_array_index_1094036 ^ p92_literal_1076345[p92_array_index_1094021] ^ p92_array_index_1094022;
  assign p93_res7__493_comb = p92_literal_1076345[p93_res7__492_comb] ^ p92_literal_1076347[p93_res7__491_comb] ^ p92_literal_1076349[p93_res7__490_comb] ^ p92_literal_1076351[p92_res7__489] ^ p92_literal_1076353[p92_res7__488] ^ p92_literal_1076355[p92_res7__487] ^ p92_res7__486 ^ p92_literal_1076358[p92_res7__485] ^ p92_res7__484 ^ p92_array_index_1094264 ^ p92_array_index_1094240 ^ p92_array_index_1094214 ^ p92_array_index_1094082 ^ p92_array_index_1094053 ^ p92_literal_1076345[p92_array_index_1094020] ^ p92_array_index_1094021;
  assign p93_res7__494_comb = p92_literal_1076345[p93_res7__493_comb] ^ p92_literal_1076347[p93_res7__492_comb] ^ p92_literal_1076349[p93_res7__491_comb] ^ p92_literal_1076351[p93_res7__490_comb] ^ p92_literal_1076353[p92_res7__489] ^ p92_literal_1076355[p92_res7__488] ^ p92_res7__487 ^ p92_literal_1076358[p92_res7__486] ^ p92_res7__485 ^ p92_array_index_1094275 ^ p92_array_index_1094252 ^ p92_array_index_1094227 ^ p92_array_index_1094096 ^ p92_array_index_1094067 ^ p92_array_index_1094035 ^ p92_array_index_1094020;
  assign p93_res7__495_comb = p92_literal_1076345[p93_res7__494_comb] ^ p92_literal_1076347[p93_res7__493_comb] ^ p92_literal_1076349[p93_res7__492_comb] ^ p92_literal_1076351[p93_res7__491_comb] ^ p92_literal_1076353[p93_res7__490_comb] ^ p92_literal_1076355[p92_res7__489] ^ p92_res7__488 ^ p92_literal_1076358[p92_res7__487] ^ p92_res7__486 ^ p93_array_index_1094413_comb ^ p92_array_index_1094263 ^ p92_array_index_1094239 ^ p92_array_index_1094213 ^ p92_array_index_1094081 ^ p92_array_index_1094052 ^ p92_array_index_1094019;
  assign p93_res__30_comb = {p93_res7__495_comb, p93_res7__494_comb, p93_res7__493_comb, p93_res7__492_comb, p93_res7__491_comb, p93_res7__490_comb, p92_res7__489, p92_res7__488, p92_res7__487, p92_res7__486, p92_res7__485, p92_res7__484, p92_res7__483, p92_res7__482, p92_res7__481, p92_res7__480};
  assign p93_k9_comb = p93_res__30_comb ^ p92_xor_1093509;

  // Registers for pipe stage 93:
  reg [127:0] p93_xor_1093981;
  reg [127:0] p93_k9;
  reg [127:0] p93_res__39;
  reg [7:0] p94_arr[256];
  reg [7:0] p94_literal_1076345[256];
  reg [7:0] p94_literal_1076347[256];
  reg [7:0] p94_literal_1076349[256];
  reg [7:0] p94_literal_1076351[256];
  reg [7:0] p94_literal_1076353[256];
  reg [7:0] p94_literal_1076355[256];
  reg [7:0] p94_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p93_xor_1093981 <= p92_xor_1093981;
    p93_k9 <= p93_k9_comb;
    p93_res__39 <= p92_res__39;
    p94_arr <= p93_arr;
    p94_literal_1076345 <= p93_literal_1076345;
    p94_literal_1076347 <= p93_literal_1076347;
    p94_literal_1076349 <= p93_literal_1076349;
    p94_literal_1076351 <= p93_literal_1076351;
    p94_literal_1076353 <= p93_literal_1076353;
    p94_literal_1076355 <= p93_literal_1076355;
    p94_literal_1076358 <= p93_literal_1076358;
  end

  // ===== Pipe stage 94:
  wire [127:0] p94_addedKey__72_comb;
  wire [7:0] p94_array_index_1094491_comb;
  wire [7:0] p94_array_index_1094492_comb;
  wire [7:0] p94_array_index_1094493_comb;
  wire [7:0] p94_array_index_1094494_comb;
  wire [7:0] p94_array_index_1094495_comb;
  wire [7:0] p94_array_index_1094496_comb;
  wire [7:0] p94_array_index_1094498_comb;
  wire [7:0] p94_array_index_1094500_comb;
  wire [7:0] p94_array_index_1094501_comb;
  wire [7:0] p94_array_index_1094502_comb;
  wire [7:0] p94_array_index_1094503_comb;
  wire [7:0] p94_array_index_1094504_comb;
  wire [7:0] p94_array_index_1094505_comb;
  wire [7:0] p94_array_index_1094507_comb;
  wire [7:0] p94_array_index_1094508_comb;
  wire [7:0] p94_array_index_1094509_comb;
  wire [7:0] p94_array_index_1094510_comb;
  wire [7:0] p94_array_index_1094511_comb;
  wire [7:0] p94_array_index_1094512_comb;
  wire [7:0] p94_array_index_1094513_comb;
  wire [7:0] p94_array_index_1094515_comb;
  wire [7:0] p94_res7__496_comb;
  wire [7:0] p94_array_index_1094524_comb;
  wire [7:0] p94_array_index_1094525_comb;
  wire [7:0] p94_array_index_1094526_comb;
  wire [7:0] p94_array_index_1094527_comb;
  wire [7:0] p94_array_index_1094528_comb;
  wire [7:0] p94_array_index_1094529_comb;
  wire [7:0] p94_res7__497_comb;
  wire [7:0] p94_array_index_1094539_comb;
  wire [7:0] p94_array_index_1094540_comb;
  wire [7:0] p94_array_index_1094541_comb;
  wire [7:0] p94_array_index_1094542_comb;
  wire [7:0] p94_array_index_1094543_comb;
  wire [7:0] p94_res7__498_comb;
  wire [7:0] p94_array_index_1094553_comb;
  wire [7:0] p94_array_index_1094554_comb;
  wire [7:0] p94_array_index_1094555_comb;
  wire [7:0] p94_array_index_1094556_comb;
  wire [7:0] p94_array_index_1094557_comb;
  wire [7:0] p94_res7__499_comb;
  wire [7:0] p94_array_index_1094568_comb;
  wire [7:0] p94_array_index_1094569_comb;
  wire [7:0] p94_array_index_1094570_comb;
  wire [7:0] p94_array_index_1094571_comb;
  wire [7:0] p94_res7__500_comb;
  assign p94_addedKey__72_comb = p93_k9 ^ 128'h5ea7_d858_1e14_9b61_f16a_c145_9ced_a820;
  assign p94_array_index_1094491_comb = p93_arr[p94_addedKey__72_comb[127:120]];
  assign p94_array_index_1094492_comb = p93_arr[p94_addedKey__72_comb[119:112]];
  assign p94_array_index_1094493_comb = p93_arr[p94_addedKey__72_comb[111:104]];
  assign p94_array_index_1094494_comb = p93_arr[p94_addedKey__72_comb[103:96]];
  assign p94_array_index_1094495_comb = p93_arr[p94_addedKey__72_comb[95:88]];
  assign p94_array_index_1094496_comb = p93_arr[p94_addedKey__72_comb[87:80]];
  assign p94_array_index_1094498_comb = p93_arr[p94_addedKey__72_comb[71:64]];
  assign p94_array_index_1094500_comb = p93_arr[p94_addedKey__72_comb[55:48]];
  assign p94_array_index_1094501_comb = p93_arr[p94_addedKey__72_comb[47:40]];
  assign p94_array_index_1094502_comb = p93_arr[p94_addedKey__72_comb[39:32]];
  assign p94_array_index_1094503_comb = p93_arr[p94_addedKey__72_comb[31:24]];
  assign p94_array_index_1094504_comb = p93_arr[p94_addedKey__72_comb[23:16]];
  assign p94_array_index_1094505_comb = p93_arr[p94_addedKey__72_comb[15:8]];
  assign p94_array_index_1094507_comb = p93_literal_1076345[p94_array_index_1094491_comb];
  assign p94_array_index_1094508_comb = p93_literal_1076347[p94_array_index_1094492_comb];
  assign p94_array_index_1094509_comb = p93_literal_1076349[p94_array_index_1094493_comb];
  assign p94_array_index_1094510_comb = p93_literal_1076351[p94_array_index_1094494_comb];
  assign p94_array_index_1094511_comb = p93_literal_1076353[p94_array_index_1094495_comb];
  assign p94_array_index_1094512_comb = p93_literal_1076355[p94_array_index_1094496_comb];
  assign p94_array_index_1094513_comb = p93_arr[p94_addedKey__72_comb[79:72]];
  assign p94_array_index_1094515_comb = p93_arr[p94_addedKey__72_comb[63:56]];
  assign p94_res7__496_comb = p94_array_index_1094507_comb ^ p94_array_index_1094508_comb ^ p94_array_index_1094509_comb ^ p94_array_index_1094510_comb ^ p94_array_index_1094511_comb ^ p94_array_index_1094512_comb ^ p94_array_index_1094513_comb ^ p93_literal_1076358[p94_array_index_1094498_comb] ^ p94_array_index_1094515_comb ^ p93_literal_1076355[p94_array_index_1094500_comb] ^ p93_literal_1076353[p94_array_index_1094501_comb] ^ p93_literal_1076351[p94_array_index_1094502_comb] ^ p93_literal_1076349[p94_array_index_1094503_comb] ^ p93_literal_1076347[p94_array_index_1094504_comb] ^ p93_literal_1076345[p94_array_index_1094505_comb] ^ p93_arr[p94_addedKey__72_comb[7:0]];
  assign p94_array_index_1094524_comb = p93_literal_1076345[p94_res7__496_comb];
  assign p94_array_index_1094525_comb = p93_literal_1076347[p94_array_index_1094491_comb];
  assign p94_array_index_1094526_comb = p93_literal_1076349[p94_array_index_1094492_comb];
  assign p94_array_index_1094527_comb = p93_literal_1076351[p94_array_index_1094493_comb];
  assign p94_array_index_1094528_comb = p93_literal_1076353[p94_array_index_1094494_comb];
  assign p94_array_index_1094529_comb = p93_literal_1076355[p94_array_index_1094495_comb];
  assign p94_res7__497_comb = p94_array_index_1094524_comb ^ p94_array_index_1094525_comb ^ p94_array_index_1094526_comb ^ p94_array_index_1094527_comb ^ p94_array_index_1094528_comb ^ p94_array_index_1094529_comb ^ p94_array_index_1094496_comb ^ p93_literal_1076358[p94_array_index_1094513_comb] ^ p94_array_index_1094498_comb ^ p93_literal_1076355[p94_array_index_1094515_comb] ^ p93_literal_1076353[p94_array_index_1094500_comb] ^ p93_literal_1076351[p94_array_index_1094501_comb] ^ p93_literal_1076349[p94_array_index_1094502_comb] ^ p93_literal_1076347[p94_array_index_1094503_comb] ^ p93_literal_1076345[p94_array_index_1094504_comb] ^ p94_array_index_1094505_comb;
  assign p94_array_index_1094539_comb = p93_literal_1076347[p94_res7__496_comb];
  assign p94_array_index_1094540_comb = p93_literal_1076349[p94_array_index_1094491_comb];
  assign p94_array_index_1094541_comb = p93_literal_1076351[p94_array_index_1094492_comb];
  assign p94_array_index_1094542_comb = p93_literal_1076353[p94_array_index_1094493_comb];
  assign p94_array_index_1094543_comb = p93_literal_1076355[p94_array_index_1094494_comb];
  assign p94_res7__498_comb = p93_literal_1076345[p94_res7__497_comb] ^ p94_array_index_1094539_comb ^ p94_array_index_1094540_comb ^ p94_array_index_1094541_comb ^ p94_array_index_1094542_comb ^ p94_array_index_1094543_comb ^ p94_array_index_1094495_comb ^ p93_literal_1076358[p94_array_index_1094496_comb] ^ p94_array_index_1094513_comb ^ p93_literal_1076355[p94_array_index_1094498_comb] ^ p93_literal_1076353[p94_array_index_1094515_comb] ^ p93_literal_1076351[p94_array_index_1094500_comb] ^ p93_literal_1076349[p94_array_index_1094501_comb] ^ p93_literal_1076347[p94_array_index_1094502_comb] ^ p93_literal_1076345[p94_array_index_1094503_comb] ^ p94_array_index_1094504_comb;
  assign p94_array_index_1094553_comb = p93_literal_1076347[p94_res7__497_comb];
  assign p94_array_index_1094554_comb = p93_literal_1076349[p94_res7__496_comb];
  assign p94_array_index_1094555_comb = p93_literal_1076351[p94_array_index_1094491_comb];
  assign p94_array_index_1094556_comb = p93_literal_1076353[p94_array_index_1094492_comb];
  assign p94_array_index_1094557_comb = p93_literal_1076355[p94_array_index_1094493_comb];
  assign p94_res7__499_comb = p93_literal_1076345[p94_res7__498_comb] ^ p94_array_index_1094553_comb ^ p94_array_index_1094554_comb ^ p94_array_index_1094555_comb ^ p94_array_index_1094556_comb ^ p94_array_index_1094557_comb ^ p94_array_index_1094494_comb ^ p93_literal_1076358[p94_array_index_1094495_comb] ^ p94_array_index_1094496_comb ^ p93_literal_1076355[p94_array_index_1094513_comb] ^ p93_literal_1076353[p94_array_index_1094498_comb] ^ p93_literal_1076351[p94_array_index_1094515_comb] ^ p93_literal_1076349[p94_array_index_1094500_comb] ^ p93_literal_1076347[p94_array_index_1094501_comb] ^ p93_literal_1076345[p94_array_index_1094502_comb] ^ p94_array_index_1094503_comb;
  assign p94_array_index_1094568_comb = p93_literal_1076349[p94_res7__497_comb];
  assign p94_array_index_1094569_comb = p93_literal_1076351[p94_res7__496_comb];
  assign p94_array_index_1094570_comb = p93_literal_1076353[p94_array_index_1094491_comb];
  assign p94_array_index_1094571_comb = p93_literal_1076355[p94_array_index_1094492_comb];
  assign p94_res7__500_comb = p93_literal_1076345[p94_res7__499_comb] ^ p93_literal_1076347[p94_res7__498_comb] ^ p94_array_index_1094568_comb ^ p94_array_index_1094569_comb ^ p94_array_index_1094570_comb ^ p94_array_index_1094571_comb ^ p94_array_index_1094493_comb ^ p93_literal_1076358[p94_array_index_1094494_comb] ^ p94_array_index_1094495_comb ^ p94_array_index_1094512_comb ^ p93_literal_1076353[p94_array_index_1094513_comb] ^ p93_literal_1076351[p94_array_index_1094498_comb] ^ p93_literal_1076349[p94_array_index_1094515_comb] ^ p93_literal_1076347[p94_array_index_1094500_comb] ^ p93_literal_1076345[p94_array_index_1094501_comb] ^ p94_array_index_1094502_comb;

  // Registers for pipe stage 94:
  reg [127:0] p94_xor_1093981;
  reg [127:0] p94_k9;
  reg [7:0] p94_array_index_1094491;
  reg [7:0] p94_array_index_1094492;
  reg [7:0] p94_array_index_1094493;
  reg [7:0] p94_array_index_1094494;
  reg [7:0] p94_array_index_1094495;
  reg [7:0] p94_array_index_1094496;
  reg [7:0] p94_array_index_1094498;
  reg [7:0] p94_array_index_1094500;
  reg [7:0] p94_array_index_1094501;
  reg [7:0] p94_array_index_1094507;
  reg [7:0] p94_array_index_1094508;
  reg [7:0] p94_array_index_1094509;
  reg [7:0] p94_array_index_1094510;
  reg [7:0] p94_array_index_1094511;
  reg [7:0] p94_array_index_1094513;
  reg [7:0] p94_array_index_1094515;
  reg [7:0] p94_res7__496;
  reg [7:0] p94_array_index_1094524;
  reg [7:0] p94_array_index_1094525;
  reg [7:0] p94_array_index_1094526;
  reg [7:0] p94_array_index_1094527;
  reg [7:0] p94_array_index_1094528;
  reg [7:0] p94_array_index_1094529;
  reg [7:0] p94_res7__497;
  reg [7:0] p94_array_index_1094539;
  reg [7:0] p94_array_index_1094540;
  reg [7:0] p94_array_index_1094541;
  reg [7:0] p94_array_index_1094542;
  reg [7:0] p94_array_index_1094543;
  reg [7:0] p94_res7__498;
  reg [7:0] p94_array_index_1094553;
  reg [7:0] p94_array_index_1094554;
  reg [7:0] p94_array_index_1094555;
  reg [7:0] p94_array_index_1094556;
  reg [7:0] p94_array_index_1094557;
  reg [7:0] p94_res7__499;
  reg [7:0] p94_array_index_1094568;
  reg [7:0] p94_array_index_1094569;
  reg [7:0] p94_array_index_1094570;
  reg [7:0] p94_array_index_1094571;
  reg [7:0] p94_res7__500;
  reg [127:0] p94_res__39;
  reg [7:0] p95_arr[256];
  reg [7:0] p95_literal_1076345[256];
  reg [7:0] p95_literal_1076347[256];
  reg [7:0] p95_literal_1076349[256];
  reg [7:0] p95_literal_1076351[256];
  reg [7:0] p95_literal_1076353[256];
  reg [7:0] p95_literal_1076355[256];
  reg [7:0] p95_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p94_xor_1093981 <= p93_xor_1093981;
    p94_k9 <= p93_k9;
    p94_array_index_1094491 <= p94_array_index_1094491_comb;
    p94_array_index_1094492 <= p94_array_index_1094492_comb;
    p94_array_index_1094493 <= p94_array_index_1094493_comb;
    p94_array_index_1094494 <= p94_array_index_1094494_comb;
    p94_array_index_1094495 <= p94_array_index_1094495_comb;
    p94_array_index_1094496 <= p94_array_index_1094496_comb;
    p94_array_index_1094498 <= p94_array_index_1094498_comb;
    p94_array_index_1094500 <= p94_array_index_1094500_comb;
    p94_array_index_1094501 <= p94_array_index_1094501_comb;
    p94_array_index_1094507 <= p94_array_index_1094507_comb;
    p94_array_index_1094508 <= p94_array_index_1094508_comb;
    p94_array_index_1094509 <= p94_array_index_1094509_comb;
    p94_array_index_1094510 <= p94_array_index_1094510_comb;
    p94_array_index_1094511 <= p94_array_index_1094511_comb;
    p94_array_index_1094513 <= p94_array_index_1094513_comb;
    p94_array_index_1094515 <= p94_array_index_1094515_comb;
    p94_res7__496 <= p94_res7__496_comb;
    p94_array_index_1094524 <= p94_array_index_1094524_comb;
    p94_array_index_1094525 <= p94_array_index_1094525_comb;
    p94_array_index_1094526 <= p94_array_index_1094526_comb;
    p94_array_index_1094527 <= p94_array_index_1094527_comb;
    p94_array_index_1094528 <= p94_array_index_1094528_comb;
    p94_array_index_1094529 <= p94_array_index_1094529_comb;
    p94_res7__497 <= p94_res7__497_comb;
    p94_array_index_1094539 <= p94_array_index_1094539_comb;
    p94_array_index_1094540 <= p94_array_index_1094540_comb;
    p94_array_index_1094541 <= p94_array_index_1094541_comb;
    p94_array_index_1094542 <= p94_array_index_1094542_comb;
    p94_array_index_1094543 <= p94_array_index_1094543_comb;
    p94_res7__498 <= p94_res7__498_comb;
    p94_array_index_1094553 <= p94_array_index_1094553_comb;
    p94_array_index_1094554 <= p94_array_index_1094554_comb;
    p94_array_index_1094555 <= p94_array_index_1094555_comb;
    p94_array_index_1094556 <= p94_array_index_1094556_comb;
    p94_array_index_1094557 <= p94_array_index_1094557_comb;
    p94_res7__499 <= p94_res7__499_comb;
    p94_array_index_1094568 <= p94_array_index_1094568_comb;
    p94_array_index_1094569 <= p94_array_index_1094569_comb;
    p94_array_index_1094570 <= p94_array_index_1094570_comb;
    p94_array_index_1094571 <= p94_array_index_1094571_comb;
    p94_res7__500 <= p94_res7__500_comb;
    p94_res__39 <= p93_res__39;
    p95_arr <= p94_arr;
    p95_literal_1076345 <= p94_literal_1076345;
    p95_literal_1076347 <= p94_literal_1076347;
    p95_literal_1076349 <= p94_literal_1076349;
    p95_literal_1076351 <= p94_literal_1076351;
    p95_literal_1076353 <= p94_literal_1076353;
    p95_literal_1076355 <= p94_literal_1076355;
    p95_literal_1076358 <= p94_literal_1076358;
  end

  // ===== Pipe stage 95:
  wire [7:0] p95_array_index_1094685_comb;
  wire [7:0] p95_array_index_1094686_comb;
  wire [7:0] p95_array_index_1094687_comb;
  wire [7:0] p95_array_index_1094688_comb;
  wire [7:0] p95_res7__501_comb;
  wire [7:0] p95_array_index_1094699_comb;
  wire [7:0] p95_array_index_1094700_comb;
  wire [7:0] p95_array_index_1094701_comb;
  wire [7:0] p95_res7__502_comb;
  wire [7:0] p95_array_index_1094711_comb;
  wire [7:0] p95_array_index_1094712_comb;
  wire [7:0] p95_array_index_1094713_comb;
  wire [7:0] p95_res7__503_comb;
  wire [7:0] p95_array_index_1094724_comb;
  wire [7:0] p95_array_index_1094725_comb;
  wire [7:0] p95_res7__504_comb;
  wire [7:0] p95_array_index_1094735_comb;
  wire [7:0] p95_array_index_1094736_comb;
  wire [7:0] p95_res7__505_comb;
  wire [7:0] p95_array_index_1094742_comb;
  wire [7:0] p95_array_index_1094743_comb;
  wire [7:0] p95_array_index_1094744_comb;
  wire [7:0] p95_array_index_1094745_comb;
  wire [7:0] p95_array_index_1094746_comb;
  wire [7:0] p95_array_index_1094747_comb;
  wire [7:0] p95_array_index_1094748_comb;
  wire [7:0] p95_array_index_1094749_comb;
  wire [7:0] p95_array_index_1094750_comb;
  assign p95_array_index_1094685_comb = p94_literal_1076349[p94_res7__498];
  assign p95_array_index_1094686_comb = p94_literal_1076351[p94_res7__497];
  assign p95_array_index_1094687_comb = p94_literal_1076353[p94_res7__496];
  assign p95_array_index_1094688_comb = p94_literal_1076355[p94_array_index_1094491];
  assign p95_res7__501_comb = p94_literal_1076345[p94_res7__500] ^ p94_literal_1076347[p94_res7__499] ^ p95_array_index_1094685_comb ^ p95_array_index_1094686_comb ^ p95_array_index_1094687_comb ^ p95_array_index_1094688_comb ^ p94_array_index_1094492 ^ p94_literal_1076358[p94_array_index_1094493] ^ p94_array_index_1094494 ^ p94_array_index_1094529 ^ p94_literal_1076353[p94_array_index_1094496] ^ p94_literal_1076351[p94_array_index_1094513] ^ p94_literal_1076349[p94_array_index_1094498] ^ p94_literal_1076347[p94_array_index_1094515] ^ p94_literal_1076345[p94_array_index_1094500] ^ p94_array_index_1094501;
  assign p95_array_index_1094699_comb = p94_literal_1076351[p94_res7__498];
  assign p95_array_index_1094700_comb = p94_literal_1076353[p94_res7__497];
  assign p95_array_index_1094701_comb = p94_literal_1076355[p94_res7__496];
  assign p95_res7__502_comb = p94_literal_1076345[p95_res7__501_comb] ^ p94_literal_1076347[p94_res7__500] ^ p94_literal_1076349[p94_res7__499] ^ p95_array_index_1094699_comb ^ p95_array_index_1094700_comb ^ p95_array_index_1094701_comb ^ p94_array_index_1094491 ^ p94_literal_1076358[p94_array_index_1094492] ^ p94_array_index_1094493 ^ p94_array_index_1094543 ^ p94_array_index_1094511 ^ p94_literal_1076351[p94_array_index_1094496] ^ p94_literal_1076349[p94_array_index_1094513] ^ p94_literal_1076347[p94_array_index_1094498] ^ p94_literal_1076345[p94_array_index_1094515] ^ p94_array_index_1094500;
  assign p95_array_index_1094711_comb = p94_literal_1076351[p94_res7__499];
  assign p95_array_index_1094712_comb = p94_literal_1076353[p94_res7__498];
  assign p95_array_index_1094713_comb = p94_literal_1076355[p94_res7__497];
  assign p95_res7__503_comb = p94_literal_1076345[p95_res7__502_comb] ^ p94_literal_1076347[p95_res7__501_comb] ^ p94_literal_1076349[p94_res7__500] ^ p95_array_index_1094711_comb ^ p95_array_index_1094712_comb ^ p95_array_index_1094713_comb ^ p94_res7__496 ^ p94_literal_1076358[p94_array_index_1094491] ^ p94_array_index_1094492 ^ p94_array_index_1094557 ^ p94_array_index_1094528 ^ p94_literal_1076351[p94_array_index_1094495] ^ p94_literal_1076349[p94_array_index_1094496] ^ p94_literal_1076347[p94_array_index_1094513] ^ p94_literal_1076345[p94_array_index_1094498] ^ p94_array_index_1094515;
  assign p95_array_index_1094724_comb = p94_literal_1076353[p94_res7__499];
  assign p95_array_index_1094725_comb = p94_literal_1076355[p94_res7__498];
  assign p95_res7__504_comb = p94_literal_1076345[p95_res7__503_comb] ^ p94_literal_1076347[p95_res7__502_comb] ^ p94_literal_1076349[p95_res7__501_comb] ^ p94_literal_1076351[p94_res7__500] ^ p95_array_index_1094724_comb ^ p95_array_index_1094725_comb ^ p94_res7__497 ^ p94_literal_1076358[p94_res7__496] ^ p94_array_index_1094491 ^ p94_array_index_1094571 ^ p94_array_index_1094542 ^ p94_array_index_1094510 ^ p94_literal_1076349[p94_array_index_1094495] ^ p94_literal_1076347[p94_array_index_1094496] ^ p94_literal_1076345[p94_array_index_1094513] ^ p94_array_index_1094498;
  assign p95_array_index_1094735_comb = p94_literal_1076353[p94_res7__500];
  assign p95_array_index_1094736_comb = p94_literal_1076355[p94_res7__499];
  assign p95_res7__505_comb = p94_literal_1076345[p95_res7__504_comb] ^ p94_literal_1076347[p95_res7__503_comb] ^ p94_literal_1076349[p95_res7__502_comb] ^ p94_literal_1076351[p95_res7__501_comb] ^ p95_array_index_1094735_comb ^ p95_array_index_1094736_comb ^ p94_res7__498 ^ p94_literal_1076358[p94_res7__497] ^ p94_res7__496 ^ p95_array_index_1094688_comb ^ p94_array_index_1094556 ^ p94_array_index_1094527 ^ p94_literal_1076349[p94_array_index_1094494] ^ p94_literal_1076347[p94_array_index_1094495] ^ p94_literal_1076345[p94_array_index_1094496] ^ p94_array_index_1094513;
  assign p95_array_index_1094742_comb = p94_literal_1076345[p95_res7__505_comb];
  assign p95_array_index_1094743_comb = p94_literal_1076347[p95_res7__504_comb];
  assign p95_array_index_1094744_comb = p94_literal_1076349[p95_res7__503_comb];
  assign p95_array_index_1094745_comb = p94_literal_1076351[p95_res7__502_comb];
  assign p95_array_index_1094746_comb = p94_literal_1076353[p95_res7__501_comb];
  assign p95_array_index_1094747_comb = p94_literal_1076355[p94_res7__500];
  assign p95_array_index_1094748_comb = p94_literal_1076358[p94_res7__498];
  assign p95_array_index_1094749_comb = p94_literal_1076347[p94_array_index_1094494];
  assign p95_array_index_1094750_comb = p94_literal_1076345[p94_array_index_1094495];

  // Registers for pipe stage 95:
  reg [127:0] p95_xor_1093981;
  reg [127:0] p95_k9;
  reg [7:0] p95_array_index_1094491;
  reg [7:0] p95_array_index_1094492;
  reg [7:0] p95_array_index_1094493;
  reg [7:0] p95_array_index_1094494;
  reg [7:0] p95_array_index_1094495;
  reg [7:0] p95_array_index_1094496;
  reg [7:0] p95_array_index_1094507;
  reg [7:0] p95_array_index_1094508;
  reg [7:0] p95_array_index_1094509;
  reg [7:0] p95_res7__496;
  reg [7:0] p95_array_index_1094524;
  reg [7:0] p95_array_index_1094525;
  reg [7:0] p95_array_index_1094526;
  reg [7:0] p95_res7__497;
  reg [7:0] p95_array_index_1094539;
  reg [7:0] p95_array_index_1094540;
  reg [7:0] p95_array_index_1094541;
  reg [7:0] p95_res7__498;
  reg [7:0] p95_array_index_1094553;
  reg [7:0] p95_array_index_1094554;
  reg [7:0] p95_array_index_1094555;
  reg [7:0] p95_res7__499;
  reg [7:0] p95_array_index_1094568;
  reg [7:0] p95_array_index_1094569;
  reg [7:0] p95_array_index_1094570;
  reg [7:0] p95_res7__500;
  reg [7:0] p95_array_index_1094685;
  reg [7:0] p95_array_index_1094686;
  reg [7:0] p95_array_index_1094687;
  reg [7:0] p95_res7__501;
  reg [7:0] p95_array_index_1094699;
  reg [7:0] p95_array_index_1094700;
  reg [7:0] p95_array_index_1094701;
  reg [7:0] p95_res7__502;
  reg [7:0] p95_array_index_1094711;
  reg [7:0] p95_array_index_1094712;
  reg [7:0] p95_array_index_1094713;
  reg [7:0] p95_res7__503;
  reg [7:0] p95_array_index_1094724;
  reg [7:0] p95_array_index_1094725;
  reg [7:0] p95_res7__504;
  reg [7:0] p95_array_index_1094735;
  reg [7:0] p95_array_index_1094736;
  reg [7:0] p95_res7__505;
  reg [7:0] p95_array_index_1094742;
  reg [7:0] p95_array_index_1094743;
  reg [7:0] p95_array_index_1094744;
  reg [7:0] p95_array_index_1094745;
  reg [7:0] p95_array_index_1094746;
  reg [7:0] p95_array_index_1094747;
  reg [7:0] p95_array_index_1094748;
  reg [7:0] p95_array_index_1094749;
  reg [7:0] p95_array_index_1094750;
  reg [127:0] p95_res__39;
  reg [7:0] p96_arr[256];
  reg [7:0] p96_literal_1076345[256];
  reg [7:0] p96_literal_1076347[256];
  reg [7:0] p96_literal_1076349[256];
  reg [7:0] p96_literal_1076351[256];
  reg [7:0] p96_literal_1076353[256];
  reg [7:0] p96_literal_1076355[256];
  reg [7:0] p96_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p95_xor_1093981 <= p94_xor_1093981;
    p95_k9 <= p94_k9;
    p95_array_index_1094491 <= p94_array_index_1094491;
    p95_array_index_1094492 <= p94_array_index_1094492;
    p95_array_index_1094493 <= p94_array_index_1094493;
    p95_array_index_1094494 <= p94_array_index_1094494;
    p95_array_index_1094495 <= p94_array_index_1094495;
    p95_array_index_1094496 <= p94_array_index_1094496;
    p95_array_index_1094507 <= p94_array_index_1094507;
    p95_array_index_1094508 <= p94_array_index_1094508;
    p95_array_index_1094509 <= p94_array_index_1094509;
    p95_res7__496 <= p94_res7__496;
    p95_array_index_1094524 <= p94_array_index_1094524;
    p95_array_index_1094525 <= p94_array_index_1094525;
    p95_array_index_1094526 <= p94_array_index_1094526;
    p95_res7__497 <= p94_res7__497;
    p95_array_index_1094539 <= p94_array_index_1094539;
    p95_array_index_1094540 <= p94_array_index_1094540;
    p95_array_index_1094541 <= p94_array_index_1094541;
    p95_res7__498 <= p94_res7__498;
    p95_array_index_1094553 <= p94_array_index_1094553;
    p95_array_index_1094554 <= p94_array_index_1094554;
    p95_array_index_1094555 <= p94_array_index_1094555;
    p95_res7__499 <= p94_res7__499;
    p95_array_index_1094568 <= p94_array_index_1094568;
    p95_array_index_1094569 <= p94_array_index_1094569;
    p95_array_index_1094570 <= p94_array_index_1094570;
    p95_res7__500 <= p94_res7__500;
    p95_array_index_1094685 <= p95_array_index_1094685_comb;
    p95_array_index_1094686 <= p95_array_index_1094686_comb;
    p95_array_index_1094687 <= p95_array_index_1094687_comb;
    p95_res7__501 <= p95_res7__501_comb;
    p95_array_index_1094699 <= p95_array_index_1094699_comb;
    p95_array_index_1094700 <= p95_array_index_1094700_comb;
    p95_array_index_1094701 <= p95_array_index_1094701_comb;
    p95_res7__502 <= p95_res7__502_comb;
    p95_array_index_1094711 <= p95_array_index_1094711_comb;
    p95_array_index_1094712 <= p95_array_index_1094712_comb;
    p95_array_index_1094713 <= p95_array_index_1094713_comb;
    p95_res7__503 <= p95_res7__503_comb;
    p95_array_index_1094724 <= p95_array_index_1094724_comb;
    p95_array_index_1094725 <= p95_array_index_1094725_comb;
    p95_res7__504 <= p95_res7__504_comb;
    p95_array_index_1094735 <= p95_array_index_1094735_comb;
    p95_array_index_1094736 <= p95_array_index_1094736_comb;
    p95_res7__505 <= p95_res7__505_comb;
    p95_array_index_1094742 <= p95_array_index_1094742_comb;
    p95_array_index_1094743 <= p95_array_index_1094743_comb;
    p95_array_index_1094744 <= p95_array_index_1094744_comb;
    p95_array_index_1094745 <= p95_array_index_1094745_comb;
    p95_array_index_1094746 <= p95_array_index_1094746_comb;
    p95_array_index_1094747 <= p95_array_index_1094747_comb;
    p95_array_index_1094748 <= p95_array_index_1094748_comb;
    p95_array_index_1094749 <= p95_array_index_1094749_comb;
    p95_array_index_1094750 <= p95_array_index_1094750_comb;
    p95_res__39 <= p94_res__39;
    p96_arr <= p95_arr;
    p96_literal_1076345 <= p95_literal_1076345;
    p96_literal_1076347 <= p95_literal_1076347;
    p96_literal_1076349 <= p95_literal_1076349;
    p96_literal_1076351 <= p95_literal_1076351;
    p96_literal_1076353 <= p95_literal_1076353;
    p96_literal_1076355 <= p95_literal_1076355;
    p96_literal_1076358 <= p95_literal_1076358;
  end

  // ===== Pipe stage 96:
  wire [7:0] p96_res7__506_comb;
  wire [7:0] p96_array_index_1094885_comb;
  wire [7:0] p96_res7__507_comb;
  wire [7:0] p96_res7__508_comb;
  wire [7:0] p96_res7__509_comb;
  wire [7:0] p96_res7__510_comb;
  wire [7:0] p96_res7__511_comb;
  wire [127:0] p96_res__31_comb;
  wire [127:0] p96_addedKey__40_comb;
  wire [7:0] p96_bit_slice_1094926_comb;
  wire [7:0] p96_bit_slice_1094927_comb;
  wire [7:0] p96_bit_slice_1094928_comb;
  wire [7:0] p96_bit_slice_1094929_comb;
  wire [7:0] p96_bit_slice_1094930_comb;
  wire [7:0] p96_bit_slice_1094931_comb;
  wire [7:0] p96_bit_slice_1094932_comb;
  wire [7:0] p96_bit_slice_1094933_comb;
  wire [7:0] p96_bit_slice_1094934_comb;
  wire [7:0] p96_bit_slice_1094935_comb;
  wire [7:0] p96_bit_slice_1094936_comb;
  wire [7:0] p96_bit_slice_1094937_comb;
  wire [7:0] p96_bit_slice_1094938_comb;
  wire [7:0] p96_bit_slice_1094939_comb;
  wire [7:0] p96_bit_slice_1094940_comb;
  wire [7:0] p96_bit_slice_1094941_comb;
  assign p96_res7__506_comb = p95_array_index_1094742 ^ p95_array_index_1094743 ^ p95_array_index_1094744 ^ p95_array_index_1094745 ^ p95_array_index_1094746 ^ p95_array_index_1094747 ^ p95_res7__499 ^ p95_array_index_1094748 ^ p95_res7__497 ^ p95_array_index_1094701 ^ p95_array_index_1094570 ^ p95_array_index_1094541 ^ p95_array_index_1094509 ^ p95_array_index_1094749 ^ p95_array_index_1094750 ^ p95_array_index_1094496;
  assign p96_array_index_1094885_comb = p95_literal_1076355[p95_res7__501];
  assign p96_res7__507_comb = p95_literal_1076345[p96_res7__506_comb] ^ p95_literal_1076347[p95_res7__505] ^ p95_literal_1076349[p95_res7__504] ^ p95_literal_1076351[p95_res7__503] ^ p95_literal_1076353[p95_res7__502] ^ p96_array_index_1094885_comb ^ p95_res7__500 ^ p95_literal_1076358[p95_res7__499] ^ p95_res7__498 ^ p95_array_index_1094713 ^ p95_array_index_1094687 ^ p95_array_index_1094555 ^ p95_array_index_1094526 ^ p95_literal_1076347[p95_array_index_1094493] ^ p95_literal_1076345[p95_array_index_1094494] ^ p95_array_index_1094495;
  assign p96_res7__508_comb = p95_literal_1076345[p96_res7__507_comb] ^ p95_literal_1076347[p96_res7__506_comb] ^ p95_literal_1076349[p95_res7__505] ^ p95_literal_1076351[p95_res7__504] ^ p95_literal_1076353[p95_res7__503] ^ p95_literal_1076355[p95_res7__502] ^ p95_res7__501 ^ p95_literal_1076358[p95_res7__500] ^ p95_res7__499 ^ p95_array_index_1094725 ^ p95_array_index_1094700 ^ p95_array_index_1094569 ^ p95_array_index_1094540 ^ p95_array_index_1094508 ^ p95_literal_1076345[p95_array_index_1094493] ^ p95_array_index_1094494;
  assign p96_res7__509_comb = p95_literal_1076345[p96_res7__508_comb] ^ p95_literal_1076347[p96_res7__507_comb] ^ p95_literal_1076349[p96_res7__506_comb] ^ p95_literal_1076351[p95_res7__505] ^ p95_literal_1076353[p95_res7__504] ^ p95_literal_1076355[p95_res7__503] ^ p95_res7__502 ^ p95_literal_1076358[p95_res7__501] ^ p95_res7__500 ^ p95_array_index_1094736 ^ p95_array_index_1094712 ^ p95_array_index_1094686 ^ p95_array_index_1094554 ^ p95_array_index_1094525 ^ p95_literal_1076345[p95_array_index_1094492] ^ p95_array_index_1094493;
  assign p96_res7__510_comb = p95_literal_1076345[p96_res7__509_comb] ^ p95_literal_1076347[p96_res7__508_comb] ^ p95_literal_1076349[p96_res7__507_comb] ^ p95_literal_1076351[p96_res7__506_comb] ^ p95_literal_1076353[p95_res7__505] ^ p95_literal_1076355[p95_res7__504] ^ p95_res7__503 ^ p95_literal_1076358[p95_res7__502] ^ p95_res7__501 ^ p95_array_index_1094747 ^ p95_array_index_1094724 ^ p95_array_index_1094699 ^ p95_array_index_1094568 ^ p95_array_index_1094539 ^ p95_array_index_1094507 ^ p95_array_index_1094492;
  assign p96_res7__511_comb = p95_literal_1076345[p96_res7__510_comb] ^ p95_literal_1076347[p96_res7__509_comb] ^ p95_literal_1076349[p96_res7__508_comb] ^ p95_literal_1076351[p96_res7__507_comb] ^ p95_literal_1076353[p96_res7__506_comb] ^ p95_literal_1076355[p95_res7__505] ^ p95_res7__504 ^ p95_literal_1076358[p95_res7__503] ^ p95_res7__502 ^ p96_array_index_1094885_comb ^ p95_array_index_1094735 ^ p95_array_index_1094711 ^ p95_array_index_1094685 ^ p95_array_index_1094553 ^ p95_array_index_1094524 ^ p95_array_index_1094491;
  assign p96_res__31_comb = {p96_res7__511_comb, p96_res7__510_comb, p96_res7__509_comb, p96_res7__508_comb, p96_res7__507_comb, p96_res7__506_comb, p95_res7__505, p95_res7__504, p95_res7__503, p95_res7__502, p95_res7__501, p95_res7__500, p95_res7__499, p95_res7__498, p95_res7__497, p95_res7__496};
  assign p96_addedKey__40_comb = p96_res__31_comb ^ p95_xor_1093981 ^ p95_res__39;
  assign p96_bit_slice_1094926_comb = p96_addedKey__40_comb[127:120];
  assign p96_bit_slice_1094927_comb = p96_addedKey__40_comb[119:112];
  assign p96_bit_slice_1094928_comb = p96_addedKey__40_comb[111:104];
  assign p96_bit_slice_1094929_comb = p96_addedKey__40_comb[103:96];
  assign p96_bit_slice_1094930_comb = p96_addedKey__40_comb[95:88];
  assign p96_bit_slice_1094931_comb = p96_addedKey__40_comb[87:80];
  assign p96_bit_slice_1094932_comb = p96_addedKey__40_comb[71:64];
  assign p96_bit_slice_1094933_comb = p96_addedKey__40_comb[55:48];
  assign p96_bit_slice_1094934_comb = p96_addedKey__40_comb[47:40];
  assign p96_bit_slice_1094935_comb = p96_addedKey__40_comb[39:32];
  assign p96_bit_slice_1094936_comb = p96_addedKey__40_comb[31:24];
  assign p96_bit_slice_1094937_comb = p96_addedKey__40_comb[23:16];
  assign p96_bit_slice_1094938_comb = p96_addedKey__40_comb[15:8];
  assign p96_bit_slice_1094939_comb = p96_addedKey__40_comb[79:72];
  assign p96_bit_slice_1094940_comb = p96_addedKey__40_comb[63:56];
  assign p96_bit_slice_1094941_comb = p96_addedKey__40_comb[7:0];

  // Registers for pipe stage 96:
  reg [127:0] p96_k9;
  reg [7:0] p96_bit_slice_1094926;
  reg [7:0] p96_bit_slice_1094927;
  reg [7:0] p96_bit_slice_1094928;
  reg [7:0] p96_bit_slice_1094929;
  reg [7:0] p96_bit_slice_1094930;
  reg [7:0] p96_bit_slice_1094931;
  reg [7:0] p96_bit_slice_1094932;
  reg [7:0] p96_bit_slice_1094933;
  reg [7:0] p96_bit_slice_1094934;
  reg [7:0] p96_bit_slice_1094935;
  reg [7:0] p96_bit_slice_1094936;
  reg [7:0] p96_bit_slice_1094937;
  reg [7:0] p96_bit_slice_1094938;
  reg [7:0] p96_bit_slice_1094939;
  reg [7:0] p96_bit_slice_1094940;
  reg [7:0] p96_bit_slice_1094941;
  reg [7:0] p97_literal_1076345[256];
  reg [7:0] p97_literal_1076347[256];
  reg [7:0] p97_literal_1076349[256];
  reg [7:0] p97_literal_1076351[256];
  reg [7:0] p97_literal_1076353[256];
  reg [7:0] p97_literal_1076355[256];
  reg [7:0] p97_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p96_k9 <= p95_k9;
    p96_bit_slice_1094926 <= p96_bit_slice_1094926_comb;
    p96_bit_slice_1094927 <= p96_bit_slice_1094927_comb;
    p96_bit_slice_1094928 <= p96_bit_slice_1094928_comb;
    p96_bit_slice_1094929 <= p96_bit_slice_1094929_comb;
    p96_bit_slice_1094930 <= p96_bit_slice_1094930_comb;
    p96_bit_slice_1094931 <= p96_bit_slice_1094931_comb;
    p96_bit_slice_1094932 <= p96_bit_slice_1094932_comb;
    p96_bit_slice_1094933 <= p96_bit_slice_1094933_comb;
    p96_bit_slice_1094934 <= p96_bit_slice_1094934_comb;
    p96_bit_slice_1094935 <= p96_bit_slice_1094935_comb;
    p96_bit_slice_1094936 <= p96_bit_slice_1094936_comb;
    p96_bit_slice_1094937 <= p96_bit_slice_1094937_comb;
    p96_bit_slice_1094938 <= p96_bit_slice_1094938_comb;
    p96_bit_slice_1094939 <= p96_bit_slice_1094939_comb;
    p96_bit_slice_1094940 <= p96_bit_slice_1094940_comb;
    p96_bit_slice_1094941 <= p96_bit_slice_1094941_comb;
    p97_literal_1076345 <= p96_literal_1076345;
    p97_literal_1076347 <= p96_literal_1076347;
    p97_literal_1076349 <= p96_literal_1076349;
    p97_literal_1076351 <= p96_literal_1076351;
    p97_literal_1076353 <= p96_literal_1076353;
    p97_literal_1076355 <= p96_literal_1076355;
    p97_literal_1076358 <= p96_literal_1076358;
  end

  // ===== Pipe stage 97:
  wire [7:0] p97_array_index_1094992_comb;
  wire [7:0] p97_array_index_1094993_comb;
  wire [7:0] p97_array_index_1094994_comb;
  wire [7:0] p97_array_index_1094995_comb;
  wire [7:0] p97_array_index_1094996_comb;
  wire [7:0] p97_array_index_1094997_comb;
  wire [7:0] p97_array_index_1094998_comb;
  wire [7:0] p97_array_index_1094999_comb;
  wire [7:0] p97_array_index_1095000_comb;
  wire [7:0] p97_array_index_1095001_comb;
  wire [7:0] p97_array_index_1095002_comb;
  wire [7:0] p97_array_index_1095003_comb;
  wire [7:0] p97_array_index_1095004_comb;
  wire [7:0] p97_array_index_1095005_comb;
  wire [7:0] p97_array_index_1095006_comb;
  wire [7:0] p97_array_index_1095007_comb;
  wire [7:0] p97_array_index_1095008_comb;
  wire [7:0] p97_array_index_1095009_comb;
  wire [7:0] p97_array_index_1095010_comb;
  wire [7:0] p97_array_index_1095011_comb;
  wire [7:0] p97_array_index_1095013_comb;
  wire [7:0] p97_res7__640_comb;
  wire [7:0] p97_array_index_1095022_comb;
  wire [7:0] p97_array_index_1095023_comb;
  wire [7:0] p97_array_index_1095024_comb;
  wire [7:0] p97_array_index_1095025_comb;
  wire [7:0] p97_array_index_1095026_comb;
  wire [7:0] p97_array_index_1095027_comb;
  wire [7:0] p97_res7__641_comb;
  wire [7:0] p97_array_index_1095037_comb;
  wire [7:0] p97_array_index_1095038_comb;
  wire [7:0] p97_array_index_1095039_comb;
  wire [7:0] p97_array_index_1095040_comb;
  wire [7:0] p97_array_index_1095041_comb;
  wire [7:0] p97_res7__642_comb;
  wire [7:0] p97_array_index_1095051_comb;
  wire [7:0] p97_array_index_1095052_comb;
  wire [7:0] p97_array_index_1095053_comb;
  wire [7:0] p97_array_index_1095054_comb;
  wire [7:0] p97_array_index_1095055_comb;
  wire [7:0] p97_res7__643_comb;
  wire [7:0] p97_array_index_1095066_comb;
  wire [7:0] p97_array_index_1095067_comb;
  wire [7:0] p97_array_index_1095068_comb;
  wire [7:0] p97_array_index_1095069_comb;
  wire [7:0] p97_res7__644_comb;
  assign p97_array_index_1094992_comb = p96_arr[p96_bit_slice_1094926];
  assign p97_array_index_1094993_comb = p96_arr[p96_bit_slice_1094927];
  assign p97_array_index_1094994_comb = p96_arr[p96_bit_slice_1094928];
  assign p97_array_index_1094995_comb = p96_arr[p96_bit_slice_1094929];
  assign p97_array_index_1094996_comb = p96_arr[p96_bit_slice_1094930];
  assign p97_array_index_1094997_comb = p96_arr[p96_bit_slice_1094931];
  assign p97_array_index_1094998_comb = p96_arr[p96_bit_slice_1094932];
  assign p97_array_index_1094999_comb = p96_arr[p96_bit_slice_1094933];
  assign p97_array_index_1095000_comb = p96_arr[p96_bit_slice_1094934];
  assign p97_array_index_1095001_comb = p96_arr[p96_bit_slice_1094935];
  assign p97_array_index_1095002_comb = p96_arr[p96_bit_slice_1094936];
  assign p97_array_index_1095003_comb = p96_arr[p96_bit_slice_1094937];
  assign p97_array_index_1095004_comb = p96_arr[p96_bit_slice_1094938];
  assign p97_array_index_1095005_comb = p96_literal_1076345[p97_array_index_1094992_comb];
  assign p97_array_index_1095006_comb = p96_literal_1076347[p97_array_index_1094993_comb];
  assign p97_array_index_1095007_comb = p96_literal_1076349[p97_array_index_1094994_comb];
  assign p97_array_index_1095008_comb = p96_literal_1076351[p97_array_index_1094995_comb];
  assign p97_array_index_1095009_comb = p96_literal_1076353[p97_array_index_1094996_comb];
  assign p97_array_index_1095010_comb = p96_literal_1076355[p97_array_index_1094997_comb];
  assign p97_array_index_1095011_comb = p96_arr[p96_bit_slice_1094939];
  assign p97_array_index_1095013_comb = p96_arr[p96_bit_slice_1094940];
  assign p97_res7__640_comb = p97_array_index_1095005_comb ^ p97_array_index_1095006_comb ^ p97_array_index_1095007_comb ^ p97_array_index_1095008_comb ^ p97_array_index_1095009_comb ^ p97_array_index_1095010_comb ^ p97_array_index_1095011_comb ^ p96_literal_1076358[p97_array_index_1094998_comb] ^ p97_array_index_1095013_comb ^ p96_literal_1076355[p97_array_index_1094999_comb] ^ p96_literal_1076353[p97_array_index_1095000_comb] ^ p96_literal_1076351[p97_array_index_1095001_comb] ^ p96_literal_1076349[p97_array_index_1095002_comb] ^ p96_literal_1076347[p97_array_index_1095003_comb] ^ p96_literal_1076345[p97_array_index_1095004_comb] ^ p96_arr[p96_bit_slice_1094941];
  assign p97_array_index_1095022_comb = p96_literal_1076345[p97_res7__640_comb];
  assign p97_array_index_1095023_comb = p96_literal_1076347[p97_array_index_1094992_comb];
  assign p97_array_index_1095024_comb = p96_literal_1076349[p97_array_index_1094993_comb];
  assign p97_array_index_1095025_comb = p96_literal_1076351[p97_array_index_1094994_comb];
  assign p97_array_index_1095026_comb = p96_literal_1076353[p97_array_index_1094995_comb];
  assign p97_array_index_1095027_comb = p96_literal_1076355[p97_array_index_1094996_comb];
  assign p97_res7__641_comb = p97_array_index_1095022_comb ^ p97_array_index_1095023_comb ^ p97_array_index_1095024_comb ^ p97_array_index_1095025_comb ^ p97_array_index_1095026_comb ^ p97_array_index_1095027_comb ^ p97_array_index_1094997_comb ^ p96_literal_1076358[p97_array_index_1095011_comb] ^ p97_array_index_1094998_comb ^ p96_literal_1076355[p97_array_index_1095013_comb] ^ p96_literal_1076353[p97_array_index_1094999_comb] ^ p96_literal_1076351[p97_array_index_1095000_comb] ^ p96_literal_1076349[p97_array_index_1095001_comb] ^ p96_literal_1076347[p97_array_index_1095002_comb] ^ p96_literal_1076345[p97_array_index_1095003_comb] ^ p97_array_index_1095004_comb;
  assign p97_array_index_1095037_comb = p96_literal_1076347[p97_res7__640_comb];
  assign p97_array_index_1095038_comb = p96_literal_1076349[p97_array_index_1094992_comb];
  assign p97_array_index_1095039_comb = p96_literal_1076351[p97_array_index_1094993_comb];
  assign p97_array_index_1095040_comb = p96_literal_1076353[p97_array_index_1094994_comb];
  assign p97_array_index_1095041_comb = p96_literal_1076355[p97_array_index_1094995_comb];
  assign p97_res7__642_comb = p96_literal_1076345[p97_res7__641_comb] ^ p97_array_index_1095037_comb ^ p97_array_index_1095038_comb ^ p97_array_index_1095039_comb ^ p97_array_index_1095040_comb ^ p97_array_index_1095041_comb ^ p97_array_index_1094996_comb ^ p96_literal_1076358[p97_array_index_1094997_comb] ^ p97_array_index_1095011_comb ^ p96_literal_1076355[p97_array_index_1094998_comb] ^ p96_literal_1076353[p97_array_index_1095013_comb] ^ p96_literal_1076351[p97_array_index_1094999_comb] ^ p96_literal_1076349[p97_array_index_1095000_comb] ^ p96_literal_1076347[p97_array_index_1095001_comb] ^ p96_literal_1076345[p97_array_index_1095002_comb] ^ p97_array_index_1095003_comb;
  assign p97_array_index_1095051_comb = p96_literal_1076347[p97_res7__641_comb];
  assign p97_array_index_1095052_comb = p96_literal_1076349[p97_res7__640_comb];
  assign p97_array_index_1095053_comb = p96_literal_1076351[p97_array_index_1094992_comb];
  assign p97_array_index_1095054_comb = p96_literal_1076353[p97_array_index_1094993_comb];
  assign p97_array_index_1095055_comb = p96_literal_1076355[p97_array_index_1094994_comb];
  assign p97_res7__643_comb = p96_literal_1076345[p97_res7__642_comb] ^ p97_array_index_1095051_comb ^ p97_array_index_1095052_comb ^ p97_array_index_1095053_comb ^ p97_array_index_1095054_comb ^ p97_array_index_1095055_comb ^ p97_array_index_1094995_comb ^ p96_literal_1076358[p97_array_index_1094996_comb] ^ p97_array_index_1094997_comb ^ p96_literal_1076355[p97_array_index_1095011_comb] ^ p96_literal_1076353[p97_array_index_1094998_comb] ^ p96_literal_1076351[p97_array_index_1095013_comb] ^ p96_literal_1076349[p97_array_index_1094999_comb] ^ p96_literal_1076347[p97_array_index_1095000_comb] ^ p96_literal_1076345[p97_array_index_1095001_comb] ^ p97_array_index_1095002_comb;
  assign p97_array_index_1095066_comb = p96_literal_1076349[p97_res7__641_comb];
  assign p97_array_index_1095067_comb = p96_literal_1076351[p97_res7__640_comb];
  assign p97_array_index_1095068_comb = p96_literal_1076353[p97_array_index_1094992_comb];
  assign p97_array_index_1095069_comb = p96_literal_1076355[p97_array_index_1094993_comb];
  assign p97_res7__644_comb = p96_literal_1076345[p97_res7__643_comb] ^ p96_literal_1076347[p97_res7__642_comb] ^ p97_array_index_1095066_comb ^ p97_array_index_1095067_comb ^ p97_array_index_1095068_comb ^ p97_array_index_1095069_comb ^ p97_array_index_1094994_comb ^ p96_literal_1076358[p97_array_index_1094995_comb] ^ p97_array_index_1094996_comb ^ p97_array_index_1095010_comb ^ p96_literal_1076353[p97_array_index_1095011_comb] ^ p96_literal_1076351[p97_array_index_1094998_comb] ^ p96_literal_1076349[p97_array_index_1095013_comb] ^ p96_literal_1076347[p97_array_index_1094999_comb] ^ p96_literal_1076345[p97_array_index_1095000_comb] ^ p97_array_index_1095001_comb;

  // Registers for pipe stage 97:
  reg [127:0] p97_k9;
  reg [7:0] p97_array_index_1094992;
  reg [7:0] p97_array_index_1094993;
  reg [7:0] p97_array_index_1094994;
  reg [7:0] p97_array_index_1094995;
  reg [7:0] p97_array_index_1094996;
  reg [7:0] p97_array_index_1094997;
  reg [7:0] p97_array_index_1094998;
  reg [7:0] p97_array_index_1094999;
  reg [7:0] p97_array_index_1095000;
  reg [7:0] p97_array_index_1095005;
  reg [7:0] p97_array_index_1095006;
  reg [7:0] p97_array_index_1095007;
  reg [7:0] p97_array_index_1095008;
  reg [7:0] p97_array_index_1095009;
  reg [7:0] p97_array_index_1095011;
  reg [7:0] p97_array_index_1095013;
  reg [7:0] p97_res7__640;
  reg [7:0] p97_array_index_1095022;
  reg [7:0] p97_array_index_1095023;
  reg [7:0] p97_array_index_1095024;
  reg [7:0] p97_array_index_1095025;
  reg [7:0] p97_array_index_1095026;
  reg [7:0] p97_array_index_1095027;
  reg [7:0] p97_res7__641;
  reg [7:0] p97_array_index_1095037;
  reg [7:0] p97_array_index_1095038;
  reg [7:0] p97_array_index_1095039;
  reg [7:0] p97_array_index_1095040;
  reg [7:0] p97_array_index_1095041;
  reg [7:0] p97_res7__642;
  reg [7:0] p97_array_index_1095051;
  reg [7:0] p97_array_index_1095052;
  reg [7:0] p97_array_index_1095053;
  reg [7:0] p97_array_index_1095054;
  reg [7:0] p97_array_index_1095055;
  reg [7:0] p97_res7__643;
  reg [7:0] p97_array_index_1095066;
  reg [7:0] p97_array_index_1095067;
  reg [7:0] p97_array_index_1095068;
  reg [7:0] p97_array_index_1095069;
  reg [7:0] p97_res7__644;
  reg [7:0] p98_literal_1076345[256];
  reg [7:0] p98_literal_1076347[256];
  reg [7:0] p98_literal_1076349[256];
  reg [7:0] p98_literal_1076351[256];
  reg [7:0] p98_literal_1076353[256];
  always_ff @ (posedge clk) begin
    p97_k9 <= p96_k9;
    p97_array_index_1094992 <= p97_array_index_1094992_comb;
    p97_array_index_1094993 <= p97_array_index_1094993_comb;
    p97_array_index_1094994 <= p97_array_index_1094994_comb;
    p97_array_index_1094995 <= p97_array_index_1094995_comb;
    p97_array_index_1094996 <= p97_array_index_1094996_comb;
    p97_array_index_1094997 <= p97_array_index_1094997_comb;
    p97_array_index_1094998 <= p97_array_index_1094998_comb;
    p97_array_index_1094999 <= p97_array_index_1094999_comb;
    p97_array_index_1095000 <= p97_array_index_1095000_comb;
    p97_array_index_1095005 <= p97_array_index_1095005_comb;
    p97_array_index_1095006 <= p97_array_index_1095006_comb;
    p97_array_index_1095007 <= p97_array_index_1095007_comb;
    p97_array_index_1095008 <= p97_array_index_1095008_comb;
    p97_array_index_1095009 <= p97_array_index_1095009_comb;
    p97_array_index_1095011 <= p97_array_index_1095011_comb;
    p97_array_index_1095013 <= p97_array_index_1095013_comb;
    p97_res7__640 <= p97_res7__640_comb;
    p97_array_index_1095022 <= p97_array_index_1095022_comb;
    p97_array_index_1095023 <= p97_array_index_1095023_comb;
    p97_array_index_1095024 <= p97_array_index_1095024_comb;
    p97_array_index_1095025 <= p97_array_index_1095025_comb;
    p97_array_index_1095026 <= p97_array_index_1095026_comb;
    p97_array_index_1095027 <= p97_array_index_1095027_comb;
    p97_res7__641 <= p97_res7__641_comb;
    p97_array_index_1095037 <= p97_array_index_1095037_comb;
    p97_array_index_1095038 <= p97_array_index_1095038_comb;
    p97_array_index_1095039 <= p97_array_index_1095039_comb;
    p97_array_index_1095040 <= p97_array_index_1095040_comb;
    p97_array_index_1095041 <= p97_array_index_1095041_comb;
    p97_res7__642 <= p97_res7__642_comb;
    p97_array_index_1095051 <= p97_array_index_1095051_comb;
    p97_array_index_1095052 <= p97_array_index_1095052_comb;
    p97_array_index_1095053 <= p97_array_index_1095053_comb;
    p97_array_index_1095054 <= p97_array_index_1095054_comb;
    p97_array_index_1095055 <= p97_array_index_1095055_comb;
    p97_res7__643 <= p97_res7__643_comb;
    p97_array_index_1095066 <= p97_array_index_1095066_comb;
    p97_array_index_1095067 <= p97_array_index_1095067_comb;
    p97_array_index_1095068 <= p97_array_index_1095068_comb;
    p97_array_index_1095069 <= p97_array_index_1095069_comb;
    p97_res7__644 <= p97_res7__644_comb;
    p98_literal_1076345 <= p97_literal_1076345;
    p98_literal_1076347 <= p97_literal_1076347;
    p98_literal_1076349 <= p97_literal_1076349;
    p98_literal_1076351 <= p97_literal_1076351;
    p98_literal_1076353 <= p97_literal_1076353;
  end

  // ===== Pipe stage 98:
  wire [7:0] p98_array_index_1095177_comb;
  wire [7:0] p98_array_index_1095178_comb;
  wire [7:0] p98_array_index_1095179_comb;
  wire [7:0] p98_array_index_1095180_comb;
  wire [7:0] p98_res7__645_comb;
  wire [7:0] p98_array_index_1095191_comb;
  wire [7:0] p98_array_index_1095192_comb;
  wire [7:0] p98_array_index_1095193_comb;
  wire [7:0] p98_res7__646_comb;
  wire [7:0] p98_array_index_1095203_comb;
  wire [7:0] p98_array_index_1095204_comb;
  wire [7:0] p98_array_index_1095205_comb;
  wire [7:0] p98_res7__647_comb;
  wire [7:0] p98_array_index_1095216_comb;
  wire [7:0] p98_array_index_1095217_comb;
  wire [7:0] p98_res7__648_comb;
  wire [7:0] p98_array_index_1095227_comb;
  wire [7:0] p98_array_index_1095228_comb;
  wire [7:0] p98_res7__649_comb;
  wire [7:0] p98_array_index_1095234_comb;
  wire [7:0] p98_array_index_1095235_comb;
  wire [7:0] p98_array_index_1095236_comb;
  wire [7:0] p98_array_index_1095237_comb;
  wire [7:0] p98_array_index_1095238_comb;
  wire [7:0] p98_array_index_1095239_comb;
  wire [7:0] p98_array_index_1095240_comb;
  wire [7:0] p98_array_index_1095241_comb;
  wire [7:0] p98_array_index_1095242_comb;
  wire [7:0] p98_array_index_1095243_comb;
  wire [7:0] p98_array_index_1095244_comb;
  wire [7:0] p98_array_index_1095245_comb;
  wire [7:0] p98_array_index_1095246_comb;
  wire [7:0] p98_array_index_1095247_comb;
  wire [7:0] p98_array_index_1095248_comb;
  wire [7:0] p98_array_index_1095249_comb;
  wire [7:0] p98_array_index_1095250_comb;
  wire [7:0] p98_array_index_1095251_comb;
  wire [7:0] p98_array_index_1095252_comb;
  assign p98_array_index_1095177_comb = p97_literal_1076349[p97_res7__642];
  assign p98_array_index_1095178_comb = p97_literal_1076351[p97_res7__641];
  assign p98_array_index_1095179_comb = p97_literal_1076353[p97_res7__640];
  assign p98_array_index_1095180_comb = p97_literal_1076355[p97_array_index_1094992];
  assign p98_res7__645_comb = p97_literal_1076345[p97_res7__644] ^ p97_literal_1076347[p97_res7__643] ^ p98_array_index_1095177_comb ^ p98_array_index_1095178_comb ^ p98_array_index_1095179_comb ^ p98_array_index_1095180_comb ^ p97_array_index_1094993 ^ p97_literal_1076358[p97_array_index_1094994] ^ p97_array_index_1094995 ^ p97_array_index_1095027 ^ p97_literal_1076353[p97_array_index_1094997] ^ p97_literal_1076351[p97_array_index_1095011] ^ p97_literal_1076349[p97_array_index_1094998] ^ p97_literal_1076347[p97_array_index_1095013] ^ p97_literal_1076345[p97_array_index_1094999] ^ p97_array_index_1095000;
  assign p98_array_index_1095191_comb = p97_literal_1076351[p97_res7__642];
  assign p98_array_index_1095192_comb = p97_literal_1076353[p97_res7__641];
  assign p98_array_index_1095193_comb = p97_literal_1076355[p97_res7__640];
  assign p98_res7__646_comb = p97_literal_1076345[p98_res7__645_comb] ^ p97_literal_1076347[p97_res7__644] ^ p97_literal_1076349[p97_res7__643] ^ p98_array_index_1095191_comb ^ p98_array_index_1095192_comb ^ p98_array_index_1095193_comb ^ p97_array_index_1094992 ^ p97_literal_1076358[p97_array_index_1094993] ^ p97_array_index_1094994 ^ p97_array_index_1095041 ^ p97_array_index_1095009 ^ p97_literal_1076351[p97_array_index_1094997] ^ p97_literal_1076349[p97_array_index_1095011] ^ p97_literal_1076347[p97_array_index_1094998] ^ p97_literal_1076345[p97_array_index_1095013] ^ p97_array_index_1094999;
  assign p98_array_index_1095203_comb = p97_literal_1076351[p97_res7__643];
  assign p98_array_index_1095204_comb = p97_literal_1076353[p97_res7__642];
  assign p98_array_index_1095205_comb = p97_literal_1076355[p97_res7__641];
  assign p98_res7__647_comb = p97_literal_1076345[p98_res7__646_comb] ^ p97_literal_1076347[p98_res7__645_comb] ^ p97_literal_1076349[p97_res7__644] ^ p98_array_index_1095203_comb ^ p98_array_index_1095204_comb ^ p98_array_index_1095205_comb ^ p97_res7__640 ^ p97_literal_1076358[p97_array_index_1094992] ^ p97_array_index_1094993 ^ p97_array_index_1095055 ^ p97_array_index_1095026 ^ p97_literal_1076351[p97_array_index_1094996] ^ p97_literal_1076349[p97_array_index_1094997] ^ p97_literal_1076347[p97_array_index_1095011] ^ p97_literal_1076345[p97_array_index_1094998] ^ p97_array_index_1095013;
  assign p98_array_index_1095216_comb = p97_literal_1076353[p97_res7__643];
  assign p98_array_index_1095217_comb = p97_literal_1076355[p97_res7__642];
  assign p98_res7__648_comb = p97_literal_1076345[p98_res7__647_comb] ^ p97_literal_1076347[p98_res7__646_comb] ^ p97_literal_1076349[p98_res7__645_comb] ^ p97_literal_1076351[p97_res7__644] ^ p98_array_index_1095216_comb ^ p98_array_index_1095217_comb ^ p97_res7__641 ^ p97_literal_1076358[p97_res7__640] ^ p97_array_index_1094992 ^ p97_array_index_1095069 ^ p97_array_index_1095040 ^ p97_array_index_1095008 ^ p97_literal_1076349[p97_array_index_1094996] ^ p97_literal_1076347[p97_array_index_1094997] ^ p97_literal_1076345[p97_array_index_1095011] ^ p97_array_index_1094998;
  assign p98_array_index_1095227_comb = p97_literal_1076353[p97_res7__644];
  assign p98_array_index_1095228_comb = p97_literal_1076355[p97_res7__643];
  assign p98_res7__649_comb = p97_literal_1076345[p98_res7__648_comb] ^ p97_literal_1076347[p98_res7__647_comb] ^ p97_literal_1076349[p98_res7__646_comb] ^ p97_literal_1076351[p98_res7__645_comb] ^ p98_array_index_1095227_comb ^ p98_array_index_1095228_comb ^ p97_res7__642 ^ p97_literal_1076358[p97_res7__641] ^ p97_res7__640 ^ p98_array_index_1095180_comb ^ p97_array_index_1095054 ^ p97_array_index_1095025 ^ p97_literal_1076349[p97_array_index_1094995] ^ p97_literal_1076347[p97_array_index_1094996] ^ p97_literal_1076345[p97_array_index_1094997] ^ p97_array_index_1095011;
  assign p98_array_index_1095234_comb = p97_literal_1076345[p98_res7__649_comb];
  assign p98_array_index_1095235_comb = p97_literal_1076347[p98_res7__648_comb];
  assign p98_array_index_1095236_comb = p97_literal_1076349[p98_res7__647_comb];
  assign p98_array_index_1095237_comb = p97_literal_1076351[p98_res7__646_comb];
  assign p98_array_index_1095238_comb = p97_literal_1076353[p98_res7__645_comb];
  assign p98_array_index_1095239_comb = p97_literal_1076355[p97_res7__644];
  assign p98_array_index_1095240_comb = p97_literal_1076358[p97_res7__642];
  assign p98_array_index_1095241_comb = p97_literal_1076347[p97_array_index_1094995];
  assign p98_array_index_1095242_comb = p97_literal_1076345[p97_array_index_1094996];
  assign p98_array_index_1095243_comb = p97_literal_1076355[p98_res7__645_comb];
  assign p98_array_index_1095244_comb = p97_literal_1076358[p97_res7__643];
  assign p98_array_index_1095245_comb = p97_literal_1076355[p98_res7__646_comb];
  assign p98_array_index_1095246_comb = p97_literal_1076358[p97_res7__644];
  assign p98_array_index_1095247_comb = p97_literal_1076355[p98_res7__647_comb];
  assign p98_array_index_1095248_comb = p97_literal_1076358[p98_res7__645_comb];
  assign p98_array_index_1095249_comb = p97_literal_1076355[p98_res7__648_comb];
  assign p98_array_index_1095250_comb = p97_literal_1076358[p98_res7__646_comb];
  assign p98_array_index_1095251_comb = p97_literal_1076355[p98_res7__649_comb];
  assign p98_array_index_1095252_comb = p97_literal_1076358[p98_res7__647_comb];

  // Registers for pipe stage 98:
  reg [127:0] p98_k9;
  reg [7:0] p98_array_index_1094992;
  reg [7:0] p98_array_index_1094993;
  reg [7:0] p98_array_index_1094994;
  reg [7:0] p98_array_index_1094995;
  reg [7:0] p98_array_index_1094996;
  reg [7:0] p98_array_index_1094997;
  reg [7:0] p98_array_index_1095005;
  reg [7:0] p98_array_index_1095006;
  reg [7:0] p98_array_index_1095007;
  reg [7:0] p98_res7__640;
  reg [7:0] p98_array_index_1095022;
  reg [7:0] p98_array_index_1095023;
  reg [7:0] p98_array_index_1095024;
  reg [7:0] p98_res7__641;
  reg [7:0] p98_array_index_1095037;
  reg [7:0] p98_array_index_1095038;
  reg [7:0] p98_array_index_1095039;
  reg [7:0] p98_res7__642;
  reg [7:0] p98_array_index_1095051;
  reg [7:0] p98_array_index_1095052;
  reg [7:0] p98_array_index_1095053;
  reg [7:0] p98_res7__643;
  reg [7:0] p98_array_index_1095066;
  reg [7:0] p98_array_index_1095067;
  reg [7:0] p98_array_index_1095068;
  reg [7:0] p98_res7__644;
  reg [7:0] p98_array_index_1095177;
  reg [7:0] p98_array_index_1095178;
  reg [7:0] p98_array_index_1095179;
  reg [7:0] p98_res7__645;
  reg [7:0] p98_array_index_1095191;
  reg [7:0] p98_array_index_1095192;
  reg [7:0] p98_array_index_1095193;
  reg [7:0] p98_res7__646;
  reg [7:0] p98_array_index_1095203;
  reg [7:0] p98_array_index_1095204;
  reg [7:0] p98_array_index_1095205;
  reg [7:0] p98_res7__647;
  reg [7:0] p98_array_index_1095216;
  reg [7:0] p98_array_index_1095217;
  reg [7:0] p98_res7__648;
  reg [7:0] p98_array_index_1095227;
  reg [7:0] p98_array_index_1095228;
  reg [7:0] p98_res7__649;
  reg [7:0] p98_array_index_1095234;
  reg [7:0] p98_array_index_1095235;
  reg [7:0] p98_array_index_1095236;
  reg [7:0] p98_array_index_1095237;
  reg [7:0] p98_array_index_1095238;
  reg [7:0] p98_array_index_1095239;
  reg [7:0] p98_array_index_1095240;
  reg [7:0] p98_array_index_1095241;
  reg [7:0] p98_array_index_1095242;
  reg [7:0] p98_array_index_1095243;
  reg [7:0] p98_array_index_1095244;
  reg [7:0] p98_array_index_1095245;
  reg [7:0] p98_array_index_1095246;
  reg [7:0] p98_array_index_1095247;
  reg [7:0] p98_array_index_1095248;
  reg [7:0] p98_array_index_1095249;
  reg [7:0] p98_array_index_1095250;
  reg [7:0] p98_array_index_1095251;
  reg [7:0] p98_array_index_1095252;
  always_ff @ (posedge clk) begin
    p98_k9 <= p97_k9;
    p98_array_index_1094992 <= p97_array_index_1094992;
    p98_array_index_1094993 <= p97_array_index_1094993;
    p98_array_index_1094994 <= p97_array_index_1094994;
    p98_array_index_1094995 <= p97_array_index_1094995;
    p98_array_index_1094996 <= p97_array_index_1094996;
    p98_array_index_1094997 <= p97_array_index_1094997;
    p98_array_index_1095005 <= p97_array_index_1095005;
    p98_array_index_1095006 <= p97_array_index_1095006;
    p98_array_index_1095007 <= p97_array_index_1095007;
    p98_res7__640 <= p97_res7__640;
    p98_array_index_1095022 <= p97_array_index_1095022;
    p98_array_index_1095023 <= p97_array_index_1095023;
    p98_array_index_1095024 <= p97_array_index_1095024;
    p98_res7__641 <= p97_res7__641;
    p98_array_index_1095037 <= p97_array_index_1095037;
    p98_array_index_1095038 <= p97_array_index_1095038;
    p98_array_index_1095039 <= p97_array_index_1095039;
    p98_res7__642 <= p97_res7__642;
    p98_array_index_1095051 <= p97_array_index_1095051;
    p98_array_index_1095052 <= p97_array_index_1095052;
    p98_array_index_1095053 <= p97_array_index_1095053;
    p98_res7__643 <= p97_res7__643;
    p98_array_index_1095066 <= p97_array_index_1095066;
    p98_array_index_1095067 <= p97_array_index_1095067;
    p98_array_index_1095068 <= p97_array_index_1095068;
    p98_res7__644 <= p97_res7__644;
    p98_array_index_1095177 <= p98_array_index_1095177_comb;
    p98_array_index_1095178 <= p98_array_index_1095178_comb;
    p98_array_index_1095179 <= p98_array_index_1095179_comb;
    p98_res7__645 <= p98_res7__645_comb;
    p98_array_index_1095191 <= p98_array_index_1095191_comb;
    p98_array_index_1095192 <= p98_array_index_1095192_comb;
    p98_array_index_1095193 <= p98_array_index_1095193_comb;
    p98_res7__646 <= p98_res7__646_comb;
    p98_array_index_1095203 <= p98_array_index_1095203_comb;
    p98_array_index_1095204 <= p98_array_index_1095204_comb;
    p98_array_index_1095205 <= p98_array_index_1095205_comb;
    p98_res7__647 <= p98_res7__647_comb;
    p98_array_index_1095216 <= p98_array_index_1095216_comb;
    p98_array_index_1095217 <= p98_array_index_1095217_comb;
    p98_res7__648 <= p98_res7__648_comb;
    p98_array_index_1095227 <= p98_array_index_1095227_comb;
    p98_array_index_1095228 <= p98_array_index_1095228_comb;
    p98_res7__649 <= p98_res7__649_comb;
    p98_array_index_1095234 <= p98_array_index_1095234_comb;
    p98_array_index_1095235 <= p98_array_index_1095235_comb;
    p98_array_index_1095236 <= p98_array_index_1095236_comb;
    p98_array_index_1095237 <= p98_array_index_1095237_comb;
    p98_array_index_1095238 <= p98_array_index_1095238_comb;
    p98_array_index_1095239 <= p98_array_index_1095239_comb;
    p98_array_index_1095240 <= p98_array_index_1095240_comb;
    p98_array_index_1095241 <= p98_array_index_1095241_comb;
    p98_array_index_1095242 <= p98_array_index_1095242_comb;
    p98_array_index_1095243 <= p98_array_index_1095243_comb;
    p98_array_index_1095244 <= p98_array_index_1095244_comb;
    p98_array_index_1095245 <= p98_array_index_1095245_comb;
    p98_array_index_1095246 <= p98_array_index_1095246_comb;
    p98_array_index_1095247 <= p98_array_index_1095247_comb;
    p98_array_index_1095248 <= p98_array_index_1095248_comb;
    p98_array_index_1095249 <= p98_array_index_1095249_comb;
    p98_array_index_1095250 <= p98_array_index_1095250_comb;
    p98_array_index_1095251 <= p98_array_index_1095251_comb;
    p98_array_index_1095252 <= p98_array_index_1095252_comb;
  end

  // ===== Pipe stage 99:
  wire [7:0] p99_res7__650_comb;
  wire [7:0] p99_res7__651_comb;
  wire [7:0] p99_res7__652_comb;
  wire [7:0] p99_res7__653_comb;
  wire [7:0] p99_res7__654_comb;
  wire [7:0] p99_res7__655_comb;
  wire [127:0] p99_newValue_comb;
  wire [127:0] p99_xor_1095427_comb;
  assign p99_res7__650_comb = p98_array_index_1095234 ^ p98_array_index_1095235 ^ p98_array_index_1095236 ^ p98_array_index_1095237 ^ p98_array_index_1095238 ^ p98_array_index_1095239 ^ p98_res7__643 ^ p98_array_index_1095240 ^ p98_res7__641 ^ p98_array_index_1095193 ^ p98_array_index_1095068 ^ p98_array_index_1095039 ^ p98_array_index_1095007 ^ p98_array_index_1095241 ^ p98_array_index_1095242 ^ p98_array_index_1094997;
  assign p99_res7__651_comb = p98_literal_1076345[p99_res7__650_comb] ^ p98_literal_1076347[p98_res7__649] ^ p98_literal_1076349[p98_res7__648] ^ p98_literal_1076351[p98_res7__647] ^ p98_literal_1076353[p98_res7__646] ^ p98_array_index_1095243 ^ p98_res7__644 ^ p98_array_index_1095244 ^ p98_res7__642 ^ p98_array_index_1095205 ^ p98_array_index_1095179 ^ p98_array_index_1095053 ^ p98_array_index_1095024 ^ p98_literal_1076347[p98_array_index_1094994] ^ p98_literal_1076345[p98_array_index_1094995] ^ p98_array_index_1094996;
  assign p99_res7__652_comb = p98_literal_1076345[p99_res7__651_comb] ^ p98_literal_1076347[p99_res7__650_comb] ^ p98_literal_1076349[p98_res7__649] ^ p98_literal_1076351[p98_res7__648] ^ p98_literal_1076353[p98_res7__647] ^ p98_array_index_1095245 ^ p98_res7__645 ^ p98_array_index_1095246 ^ p98_res7__643 ^ p98_array_index_1095217 ^ p98_array_index_1095192 ^ p98_array_index_1095067 ^ p98_array_index_1095038 ^ p98_array_index_1095006 ^ p98_literal_1076345[p98_array_index_1094994] ^ p98_array_index_1094995;
  assign p99_res7__653_comb = p98_literal_1076345[p99_res7__652_comb] ^ p98_literal_1076347[p99_res7__651_comb] ^ p98_literal_1076349[p99_res7__650_comb] ^ p98_literal_1076351[p98_res7__649] ^ p98_literal_1076353[p98_res7__648] ^ p98_array_index_1095247 ^ p98_res7__646 ^ p98_array_index_1095248 ^ p98_res7__644 ^ p98_array_index_1095228 ^ p98_array_index_1095204 ^ p98_array_index_1095178 ^ p98_array_index_1095052 ^ p98_array_index_1095023 ^ p98_literal_1076345[p98_array_index_1094993] ^ p98_array_index_1094994;
  assign p99_res7__654_comb = p98_literal_1076345[p99_res7__653_comb] ^ p98_literal_1076347[p99_res7__652_comb] ^ p98_literal_1076349[p99_res7__651_comb] ^ p98_literal_1076351[p99_res7__650_comb] ^ p98_literal_1076353[p98_res7__649] ^ p98_array_index_1095249 ^ p98_res7__647 ^ p98_array_index_1095250 ^ p98_res7__645 ^ p98_array_index_1095239 ^ p98_array_index_1095216 ^ p98_array_index_1095191 ^ p98_array_index_1095066 ^ p98_array_index_1095037 ^ p98_array_index_1095005 ^ p98_array_index_1094993;
  assign p99_res7__655_comb = p98_literal_1076345[p99_res7__654_comb] ^ p98_literal_1076347[p99_res7__653_comb] ^ p98_literal_1076349[p99_res7__652_comb] ^ p98_literal_1076351[p99_res7__651_comb] ^ p98_literal_1076353[p99_res7__650_comb] ^ p98_array_index_1095251 ^ p98_res7__648 ^ p98_array_index_1095252 ^ p98_res7__646 ^ p98_array_index_1095243 ^ p98_array_index_1095227 ^ p98_array_index_1095203 ^ p98_array_index_1095177 ^ p98_array_index_1095051 ^ p98_array_index_1095022 ^ p98_array_index_1094992;
  assign p99_newValue_comb = {p99_res7__655_comb, p99_res7__654_comb, p99_res7__653_comb, p99_res7__652_comb, p99_res7__651_comb, p99_res7__650_comb, p98_res7__649, p98_res7__648, p98_res7__647, p98_res7__646, p98_res7__645, p98_res7__644, p98_res7__643, p98_res7__642, p98_res7__641, p98_res7__640};
  assign p99_xor_1095427_comb = p99_newValue_comb ^ p98_k9;

  // Registers for pipe stage 99:
  reg [127:0] p99_xor_1095427;
  always_ff @ (posedge clk) begin
    p99_xor_1095427 <= p99_xor_1095427_comb;
  end
  assign out = p99_xor_1095427;
endmodule
