// IWLS benchmark module "MultiplierA_32" printed on Wed May 29 22:12:33 2002
module MultiplierA_32(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \30 , \31 , \32 , \33 , \34 , \68 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ;
output
  \68 ;
reg
  \2 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ;
wire
  \[59] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \166 ,
  \167 ,
  \168 ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \197 ,
  \198 ,
  \199 ,
  \[33] ,
  \[34] ,
  \[35] ,
  \200 ,
  \201 ,
  \202 ,
  \203 ,
  \207 ,
  \209 ,
  \[36] ,
  \211 ,
  \213 ,
  \215 ,
  \217 ,
  \219 ,
  \[37] ,
  \221 ,
  \223 ,
  \225 ,
  \227 ,
  \229 ,
  \[38] ,
  \231 ,
  \233 ,
  \235 ,
  \237 ,
  \239 ,
  \[39] ,
  \241 ,
  \243 ,
  \245 ,
  \247 ,
  \249 ,
  \251 ,
  \253 ,
  \255 ,
  \257 ,
  \259 ,
  \261 ,
  \263 ,
  \265 ,
  \268 ,
  \269 ,
  \272 ,
  \274 ,
  \275 ,
  \276 ,
  \277 ,
  \278 ,
  \280 ,
  \282 ,
  \284 ,
  \286 ,
  \288 ,
  \290 ,
  \292 ,
  \294 ,
  \296 ,
  \298 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \300 ,
  \302 ,
  \304 ,
  \306 ,
  \308 ,
  \[46] ,
  \310 ,
  \312 ,
  \314 ,
  \316 ,
  \318 ,
  \[47] ,
  \320 ,
  \322 ,
  \324 ,
  \326 ,
  \328 ,
  \[48] ,
  \330 ,
  \332 ,
  \334 ,
  \336 ,
  \338 ,
  \[49] ,
  \340 ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ;
assign
  \[59]  = \193 ,
  \[60]  = \194 ,
  \[61]  = \195 ,
  \[62]  = \196 ,
  \[63]  = \197 ,
  \[64]  = \198 ,
  \166  = (\280  & \265 ) | ((\280  & \66 ) | (\265  & \66 )),
  \167  = (~\340  & \36 ) | (\340  & ~\36 ),
  \168  = (~\338  & (~\207  & \37 )) | ((~\338  & (\207  & ~\37 )) | ((\338  & (~\207  & ~\37 )) | (\338  & (\207  & \37 )))),
  \169  = (~\336  & (~\209  & \38 )) | ((~\336  & (\209  & ~\38 )) | ((\336  & (~\209  & ~\38 )) | (\336  & (\209  & \38 )))),
  \170  = (~\334  & (~\211  & \39 )) | ((~\334  & (\211  & ~\39 )) | ((\334  & (~\211  & ~\39 )) | (\334  & (\211  & \39 )))),
  \171  = (~\332  & (~\213  & \40 )) | ((~\332  & (\213  & ~\40 )) | ((\332  & (~\213  & ~\40 )) | (\332  & (\213  & \40 )))),
  \172  = (~\330  & (~\215  & \41 )) | ((~\330  & (\215  & ~\41 )) | ((\330  & (~\215  & ~\41 )) | (\330  & (\215  & \41 )))),
  \173  = (~\328  & (~\217  & \42 )) | ((~\328  & (\217  & ~\42 )) | ((\328  & (~\217  & ~\42 )) | (\328  & (\217  & \42 )))),
  \174  = (~\326  & (~\219  & \43 )) | ((~\326  & (\219  & ~\43 )) | ((\326  & (~\219  & ~\43 )) | (\326  & (\219  & \43 )))),
  \175  = (~\324  & (~\221  & \44 )) | ((~\324  & (\221  & ~\44 )) | ((\324  & (~\221  & ~\44 )) | (\324  & (\221  & \44 )))),
  \176  = (~\322  & (~\223  & \45 )) | ((~\322  & (\223  & ~\45 )) | ((\322  & (~\223  & ~\45 )) | (\322  & (\223  & \45 )))),
  \177  = (~\320  & (~\225  & \46 )) | ((~\320  & (\225  & ~\46 )) | ((\320  & (~\225  & ~\46 )) | (\320  & (\225  & \46 )))),
  \178  = (~\318  & (~\227  & \47 )) | ((~\318  & (\227  & ~\47 )) | ((\318  & (~\227  & ~\47 )) | (\318  & (\227  & \47 )))),
  \179  = (~\316  & (~\229  & \48 )) | ((~\316  & (\229  & ~\48 )) | ((\316  & (~\229  & ~\48 )) | (\316  & (\229  & \48 )))),
  \180  = (~\314  & (~\231  & \49 )) | ((~\314  & (\231  & ~\49 )) | ((\314  & (~\231  & ~\49 )) | (\314  & (\231  & \49 )))),
  \181  = (~\312  & (~\233  & \50 )) | ((~\312  & (\233  & ~\50 )) | ((\312  & (~\233  & ~\50 )) | (\312  & (\233  & \50 )))),
  \182  = (~\310  & (~\235  & \51 )) | ((~\310  & (\235  & ~\51 )) | ((\310  & (~\235  & ~\51 )) | (\310  & (\235  & \51 )))),
  \183  = (~\308  & (~\237  & \52 )) | ((~\308  & (\237  & ~\52 )) | ((\308  & (~\237  & ~\52 )) | (\308  & (\237  & \52 )))),
  \184  = (~\306  & (~\239  & \53 )) | ((~\306  & (\239  & ~\53 )) | ((\306  & (~\239  & ~\53 )) | (\306  & (\239  & \53 )))),
  \185  = (~\304  & (~\241  & \54 )) | ((~\304  & (\241  & ~\54 )) | ((\304  & (~\241  & ~\54 )) | (\304  & (\241  & \54 )))),
  \186  = (~\302  & (~\243  & \55 )) | ((~\302  & (\243  & ~\55 )) | ((\302  & (~\243  & ~\55 )) | (\302  & (\243  & \55 )))),
  \187  = (~\300  & (~\245  & \56 )) | ((~\300  & (\245  & ~\56 )) | ((\300  & (~\245  & ~\56 )) | (\300  & (\245  & \56 )))),
  \188  = (~\298  & (~\247  & \57 )) | ((~\298  & (\247  & ~\57 )) | ((\298  & (~\247  & ~\57 )) | (\298  & (\247  & \57 )))),
  \189  = (~\296  & (~\249  & \58 )) | ((~\296  & (\249  & ~\58 )) | ((\296  & (~\249  & ~\58 )) | (\296  & (\249  & \58 )))),
  \190  = (~\294  & (~\251  & \59 )) | ((~\294  & (\251  & ~\59 )) | ((\294  & (~\251  & ~\59 )) | (\294  & (\251  & \59 )))),
  \191  = (~\292  & (~\253  & \60 )) | ((~\292  & (\253  & ~\60 )) | ((\292  & (~\253  & ~\60 )) | (\292  & (\253  & \60 )))),
  \192  = (~\290  & (~\255  & \61 )) | ((~\290  & (\255  & ~\61 )) | ((\290  & (~\255  & ~\61 )) | (\290  & (\255  & \61 )))),
  \193  = (~\288  & (~\257  & \62 )) | ((~\288  & (\257  & ~\62 )) | ((\288  & (~\257  & ~\62 )) | (\288  & (\257  & \62 )))),
  \194  = (~\286  & (~\259  & \63 )) | ((~\286  & (\259  & ~\63 )) | ((\286  & (~\259  & ~\63 )) | (\286  & (\259  & \63 )))),
  \195  = (~\284  & (~\261  & \64 )) | ((~\284  & (\261  & ~\64 )) | ((\284  & (~\261  & ~\64 )) | (\284  & (\261  & \64 )))),
  \196  = (~\282  & (~\263  & \65 )) | ((~\282  & (\263  & ~\65 )) | ((\282  & (~\263  & ~\65 )) | (\282  & (\263  & \65 )))),
  \197  = (~\280  & (~\265  & \66 )) | ((~\280  & (\265  & ~\66 )) | ((\280  & (~\265  & ~\66 )) | (\280  & (\265  & \66 )))),
  \198  = (~\268  & \2 ) | (\268  & ~\2 ),
  \199  = \269  & ~\166 ,
  \[33]  = \203 ,
  \[34]  = \168 ,
  \[35]  = \169 ,
  \200  = \272  & \166 ,
  \201  = \274  & \166 ,
  \202  = \275  & \166 ,
  \203  = \277  | \276 ,
  \207  = \340  & \36 ,
  \209  = (\338  & \207 ) | ((\338  & \37 ) | (\207  & \37 )),
  \[36]  = \170 ,
  \211  = (\336  & \209 ) | ((\336  & \38 ) | (\209  & \38 )),
  \213  = (\334  & \211 ) | ((\334  & \39 ) | (\211  & \39 )),
  \215  = (\332  & \213 ) | ((\332  & \40 ) | (\213  & \40 )),
  \217  = (\330  & \215 ) | ((\330  & \41 ) | (\215  & \41 )),
  \219  = (\328  & \217 ) | ((\328  & \42 ) | (\217  & \42 )),
  \[37]  = \171 ,
  \221  = (\326  & \219 ) | ((\326  & \43 ) | (\219  & \43 )),
  \223  = (\324  & \221 ) | ((\324  & \44 ) | (\221  & \44 )),
  \225  = (\322  & \223 ) | ((\322  & \45 ) | (\223  & \45 )),
  \227  = (\320  & \225 ) | ((\320  & \46 ) | (\225  & \46 )),
  \229  = (\318  & \227 ) | ((\318  & \47 ) | (\227  & \47 )),
  \[38]  = \172 ,
  \231  = (\316  & \229 ) | ((\316  & \48 ) | (\229  & \48 )),
  \233  = (\314  & \231 ) | ((\314  & \49 ) | (\231  & \49 )),
  \235  = (\312  & \233 ) | ((\312  & \50 ) | (\233  & \50 )),
  \237  = (\310  & \235 ) | ((\310  & \51 ) | (\235  & \51 )),
  \239  = (\308  & \237 ) | ((\308  & \52 ) | (\237  & \52 )),
  \[39]  = \173 ,
  \241  = (\306  & \239 ) | ((\306  & \53 ) | (\239  & \53 )),
  \243  = (\304  & \241 ) | ((\304  & \54 ) | (\241  & \54 )),
  \245  = (\302  & \243 ) | ((\302  & \55 ) | (\243  & \55 )),
  \247  = (\300  & \245 ) | ((\300  & \56 ) | (\245  & \56 )),
  \249  = (\298  & \247 ) | ((\298  & \57 ) | (\247  & \57 )),
  \251  = (\296  & \249 ) | ((\296  & \58 ) | (\249  & \58 )),
  \253  = (\294  & \251 ) | ((\294  & \59 ) | (\251  & \59 )),
  \255  = (\292  & \253 ) | ((\292  & \60 ) | (\253  & \60 )),
  \257  = (\290  & \255 ) | ((\290  & \61 ) | (\255  & \61 )),
  \259  = (\288  & \257 ) | ((\288  & \62 ) | (\257  & \62 )),
  \261  = (\286  & \259 ) | ((\286  & \63 ) | (\259  & \63 )),
  \263  = (\284  & \261 ) | ((\284  & \64 ) | (\261  & \64 )),
  \265  = (\282  & \263 ) | ((\282  & \65 ) | (\263  & \65 )),
  \268  = (~\278  & \166 ) | (\278  & ~\166 ),
  \269  = \278  & \2 ,
  \272  = ~\278  & \2 ,
  \274  = \278  & ~\2 ,
  \275  = \278  & \2 ,
  \276  = \200  | \199 ,
  \277  = \202  | \201 ,
  \278  = \34  & \1 ,
  \280  = \33  & \1 ,
  \282  = \32  & \1 ,
  \284  = \31  & \1 ,
  \286  = \30  & \1 ,
  \288  = \29  & \1 ,
  \290  = \28  & \1 ,
  \292  = \27  & \1 ,
  \294  = \26  & \1 ,
  \296  = \25  & \1 ,
  \298  = \24  & \1 ,
  \[40]  = \174 ,
  \[41]  = \175 ,
  \[42]  = \176 ,
  \[43]  = \177 ,
  \[44]  = \178 ,
  \[45]  = \179 ,
  \300  = \23  & \1 ,
  \302  = \22  & \1 ,
  \304  = \21  & \1 ,
  \306  = \20  & \1 ,
  \308  = \19  & \1 ,
  \[46]  = \180 ,
  \310  = \18  & \1 ,
  \312  = \17  & \1 ,
  \314  = \16  & \1 ,
  \316  = \15  & \1 ,
  \318  = \14  & \1 ,
  \[47]  = \181 ,
  \320  = \13  & \1 ,
  \322  = \12  & \1 ,
  \324  = \11  & \1 ,
  \326  = \10  & \1 ,
  \328  = \9  & \1 ,
  \[48]  = \182 ,
  \330  = \8  & \1 ,
  \332  = \7  & \1 ,
  \334  = \6  & \1 ,
  \336  = \5  & \1 ,
  \338  = \4  & \1 ,
  \[49]  = \183 ,
  \340  = \3  & \1 ,
  \68  = \167 ,
  \[50]  = \184 ,
  \[51]  = \185 ,
  \[52]  = \186 ,
  \[53]  = \187 ,
  \[54]  = \188 ,
  \[55]  = \189 ,
  \[56]  = \190 ,
  \[57]  = \191 ,
  \[58]  = \192 ;
always begin
  \2  = \[33] ;
  \36  = \[34] ;
  \37  = \[35] ;
  \38  = \[36] ;
  \39  = \[37] ;
  \40  = \[38] ;
  \41  = \[39] ;
  \42  = \[40] ;
  \43  = \[41] ;
  \44  = \[42] ;
  \45  = \[43] ;
  \46  = \[44] ;
  \47  = \[45] ;
  \48  = \[46] ;
  \49  = \[47] ;
  \50  = \[48] ;
  \51  = \[49] ;
  \52  = \[50] ;
  \53  = \[51] ;
  \54  = \[52] ;
  \55  = \[53] ;
  \56  = \[54] ;
  \57  = \[55] ;
  \58  = \[56] ;
  \59  = \[57] ;
  \60  = \[58] ;
  \61  = \[59] ;
  \62  = \[60] ;
  \63  = \[61] ;
  \64  = \[62] ;
  \65  = \[63] ;
  \66  = \[64] ;
end
initial begin
  \2  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
  \49  = 0;
  \50  = 0;
  \51  = 0;
  \52  = 0;
  \53  = 0;
  \54  = 0;
  \55  = 0;
  \56  = 0;
  \57  = 0;
  \58  = 0;
  \59  = 0;
  \60  = 0;
  \61  = 0;
  \62  = 0;
  \63  = 0;
  \64  = 0;
  \65  = 0;
  \66  = 0;
end
endmodule

