module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
output n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
 n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
 n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
 n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
 n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
 n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
 n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
 n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
 n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
 n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
 n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
 n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
 n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
wire n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
 n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
 n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
 n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
 n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
 n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
 n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
 n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
 n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
 n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
 n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
 n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
 n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
 n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
 n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
 n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
 n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
 n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
 n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
 n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
 n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , 
 n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
 n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , 
 n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , 
 n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , 
 n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , 
 n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , 
 n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , 
 n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , 
 n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , 
 n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , 
 n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , 
 n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , 
 n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , 
 n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , 
 n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , 
 n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , 
 n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , 
 n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
 n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , 
 n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
 n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , 
 n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , 
 n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , 
 n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
 n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
 n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
 n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , 
 n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , 
 n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , 
 n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
 n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , 
 n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , 
 n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , 
 n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
 n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
 n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
 n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , 
 n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , 
 n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
 n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , 
 n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , 
 n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , 
 n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
 n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
 n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , 
 n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
 n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
 n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , 
 n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , 
 n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , 
 n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , 
 n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , 
 n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , 
 n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , 
 n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
 n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , 
 n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , 
 n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , 
 n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , 
 n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , 
 n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , 
 n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , 
 n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , 
 n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , 
 n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , 
 n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
 n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , 
 n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , 
 n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , 
 n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
 n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
 n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , 
 n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , 
 n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , 
 n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , 
 n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , 
 n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , 
 n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , 
 n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , 
 n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , 
 n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , 
 n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , 
 n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
 n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
 n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
 n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
 n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
 n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
 n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , 
 n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , 
 n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , 
 n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
 n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
 n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
 n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
 n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
 n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
 n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
 n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
 n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
 n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
 n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
 n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
 n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
 n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , 
 n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , 
 n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , 
 n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , 
 n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , 
 n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
 n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , 
 n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , 
 n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , 
 n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , 
 n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
 n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
 n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
 n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , 
 n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , 
 n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , 
 n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , 
 n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
 n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , 
 n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , 
 n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , 
 n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , 
 n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , 
 n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , 
 n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , 
 n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , 
 n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , 
 n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , 
 n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , 
 n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
 n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , 
 n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , 
 n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , 
 n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , 
 n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , 
 n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , 
 n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , 
 n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , 
 n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , 
 n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , 
 n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , 
 n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , 
 n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , 
 n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , 
 n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
 n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , 
 n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
 n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , 
 n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , 
 n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , 
 n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , 
 n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
 n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , 
 n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , 
 n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , 
 n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , 
 n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , 
 n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , 
 n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
 n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
 n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , 
 n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , 
 n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , 
 n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , 
 n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , 
 n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
 n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , 
 n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , 
 n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , 
 n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , 
 n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , 
 n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , 
 n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , 
 n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , 
 n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , 
 n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
 n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
 n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , 
 n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , 
 n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , 
 n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , 
 n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , 
 n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , 
 n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , 
 n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , 
 n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
 n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
 n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , 
 n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , 
 n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
 n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
 n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
 n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
 n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , 
 n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , 
 n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , 
 n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , 
 n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , 
 n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , 
 n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , 
 n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , 
 n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , 
 n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , 
 n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , 
 n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , 
 n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , 
 n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , 
 n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , 
 n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , 
 n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , 
 n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , 
 n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , 
 n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , 
 n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , 
 n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , 
 n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , 
 n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , 
 n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , 
 n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , 
 n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , 
 n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , 
 n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , 
 n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , 
 n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , 
 n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , 
 n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , 
 n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , 
 n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , 
 n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , 
 n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , 
 n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , 
 n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , 
 n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , 
 n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , 
 n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , 
 n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , 
 n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , 
 n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
 n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
 n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , 
 n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , 
 n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , 
 n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , 
 n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , 
 n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , 
 n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , 
 n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , 
 n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , 
 n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , 
 n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , 
 n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , 
 n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , 
 n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , 
 n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , 
 n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , 
 n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , 
 n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , 
 n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , 
 n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , 
 n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , 
 n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , 
 n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , 
 n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , 
 n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , 
 n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , 
 n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , 
 n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
 n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , 
 n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
 n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
 n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
 n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
 n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , 
 n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
 n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , 
 n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
 n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , 
 n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , 
 n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , 
 n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , 
 n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , 
 n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , 
 n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , 
 n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , 
 n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , 
 n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , 
 n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , 
 n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , 
 n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , 
 n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , 
 n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , 
 n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
 n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
 n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
 n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , 
 n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , 
 n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , 
 n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , 
 n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , 
 n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , 
 n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , 
 n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
 n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , 
 n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
 n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
 n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
 n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
 n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
 n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
 n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
 n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , 
 n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , 
 n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
 n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , 
 n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
 n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
 n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
 n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
 n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
 n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , 
 n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , 
 n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , 
 n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , 
 n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , 
 n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
 n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , 
 n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , 
 n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , 
 n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , 
 n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , 
 n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , 
 n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , 
 n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , 
 n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , 
 n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
 n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , 
 n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , 
 n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , 
 n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , 
 n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , 
 n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , 
 n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , 
 n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , 
 n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , 
 n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , 
 n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , 
 n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , 
 n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , 
 n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , 
 n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , 
 n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , 
 n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , 
 n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , 
 n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , 
 n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , 
 n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , 
 n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , 
 n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , 
 n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , 
 n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , 
 n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , 
 n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , 
 n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , 
 n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , 
 n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , 
 n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , 
 n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , 
 n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , 
 n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , 
 n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , 
 n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , 
 n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , 
 n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , 
 n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , 
 n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , 
 n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , 
 n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , 
 n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , 
 n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , 
 n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , 
 n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , 
 n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , 
 n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , 
 n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , 
 n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , 
 n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , 
 n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , 
 n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , 
 n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , 
 n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , 
 n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , 
 n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , 
 n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , 
 n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , 
 n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , 
 n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , 
 n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , 
 n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , 
 n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , 
 n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , 
 n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , 
 n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
 n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , 
 n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , 
 n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , 
 n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , 
 n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , 
 n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , 
 n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
 n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , 
 n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , 
 n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
 n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
 n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , 
 n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , 
 n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , 
 n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , 
 n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , 
 n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , 
 n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , 
 n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , 
 n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , 
 n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , 
 n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , 
 n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
 n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , 
 n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , 
 n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , 
 n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , 
 n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , 
 n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , 
 n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , 
 n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , 
 n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , 
 n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , 
 n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , 
 n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , 
 n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , 
 n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , 
 n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , 
 n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , 
 n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , 
 n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , 
 n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , 
 n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , 
 n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , 
 n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , 
 n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , 
 n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , 
 n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , 
 n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , 
 n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , 
 n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , 
 n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , 
 n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , 
 n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , 
 n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , 
 n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , 
 n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , 
 n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , 
 n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , 
 n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , 
 n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , 
 n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , 
 n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , 
 n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , 
 n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , 
 n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , 
 n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , 
 n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , 
 n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , 
 n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , 
 n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , 
 n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , 
 n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , 
 n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , 
 n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , 
 n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , 
 n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , 
 n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , 
 n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , 
 n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , 
 n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , 
 n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , 
 n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , 
 n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , 
 n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , 
 n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , 
 n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , 
 n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , 
 n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , 
 n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , 
 n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , 
 n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , 
 n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , 
 n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
 n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
 n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , 
 n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , 
 n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , 
 n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , 
 n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , 
 n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , 
 n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , 
 n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , 
 n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , 
 n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , 
 n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , 
 n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , 
 n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , 
 n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , 
 n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , 
 n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , 
 n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , 
 n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , 
 n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , 
 n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , 
 n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , 
 n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , 
 n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , 
 n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , 
 n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , 
 n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , 
 n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , 
 n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , 
 n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , 
 n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , 
 n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , 
 n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , 
 n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , 
 n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , 
 n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , 
 n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , 
 n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , 
 n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , 
 n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , 
 n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , 
 n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , 
 n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , 
 n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , 
 n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , 
 n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , 
 n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , 
 n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , 
 n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , 
 n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , 
 n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , 
 n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , 
 n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , 
 n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , 
 n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , 
 n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , 
 n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , 
 n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , 
 n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , 
 n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , 
 n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , 
 n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , 
 n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , 
 n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , 
 n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , 
 n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , 
 n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , 
 n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , 
 n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
 n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , 
 n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , 
 n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , 
 n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , 
 n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , 
 n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , 
 n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , 
 n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , 
 n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
 n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
 n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
 n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
 n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
 n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , 
 n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , 
 n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , 
 n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , 
 n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , 
 n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , 
 n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , 
 n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , 
 n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , 
 n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , 
 n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , 
 n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , 
 n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , 
 n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , 
 n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , 
 n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , 
 n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
 n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
 n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , 
 n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , 
 n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , 
 n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , 
 n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , 
 n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , 
 n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , 
 n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , 
 n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , 
 n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , 
 n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , 
 n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , 
 n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , 
 n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , 
 n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , 
 n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , 
 n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , 
 n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , 
 n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , 
 n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , 
 n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , 
 n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , 
 n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , 
 n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , 
 n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , 
 n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , 
 n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , 
 n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , 
 n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , 
 n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , 
 n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , 
 n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , 
 n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , 
 n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , 
 n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , 
 n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , 
 n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
 n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
 n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
 n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , 
 n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , 
 n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , 
 n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , 
 n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , 
 n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , 
 n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , 
 n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , 
 n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , 
 n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , 
 n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , 
 n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , 
 n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , 
 n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
 n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , 
 n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , 
 n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , 
 n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , 
 n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , 
 n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , 
 n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , 
 n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
 n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
 n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
 n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
 n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , 
 n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , 
 n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
 n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
 n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
 n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
 n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
 n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
 n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
 n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
 n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
 n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
 n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , 
 n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , 
 n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , 
 n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , 
 n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , 
 n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , 
 n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , 
 n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , 
 n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , 
 n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , 
 n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , 
 n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , 
 n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , 
 n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , 
 n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , 
 n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , 
 n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , 
 n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , 
 n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , 
 n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , 
 n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , 
 n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , 
 n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , 
 n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , 
 n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , 
 n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , 
 n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , 
 n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , 
 n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , 
 n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , 
 n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , 
 n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , 
 n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , 
 n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , 
 n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , 
 n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , 
 n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , 
 n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , 
 n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , 
 n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , 
 n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , 
 n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , 
 n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , 
 n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , 
 n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , 
 n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , 
 n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , 
 n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , 
 n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , 
 n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , 
 n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
 n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , 
 n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , 
 n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , 
 n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , 
 n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , 
 n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , 
 n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , 
 n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , 
 n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , 
 n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , 
 n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , 
 n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , 
 n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , 
 n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , 
 n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , 
 n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , 
 n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , 
 n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , 
 n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , 
 n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , 
 n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , 
 n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , 
 n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , 
 n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , 
 n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , 
 n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , 
 n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , 
 n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , 
 n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , 
 n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , 
 n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , 
 n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , 
 n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , 
 n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , 
 n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , 
 n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , 
 n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , 
 n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , 
 n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , 
 n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , 
 n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , 
 n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , 
 n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , 
 n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , 
 n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , 
 n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , 
 n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , 
 n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , 
 n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , 
 n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , 
 n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , 
 n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , 
 n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , 
 n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , 
 n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , 
 n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , 
 n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , 
 n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , 
 n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , 
 n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , 
 n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , 
 n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , 
 n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , 
 n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , 
 n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , 
 n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , 
 n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , 
 n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , 
 n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , 
 n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , 
 n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , 
 n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , 
 n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , 
 n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , 
 n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , 
 n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , 
 n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , 
 n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , 
 n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , 
 n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , 
 n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , 
 n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , 
 n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , 
 n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , 
 n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , 
 n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , 
 n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , 
 n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , 
 n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , 
 n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , 
 n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , 
 n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , 
 n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , 
 n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , 
 n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , 
 n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , 
 n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , 
 n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , 
 n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , 
 n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , 
 n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , 
 n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , 
 n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , 
 n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , 
 n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , 
 n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , 
 n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , 
 n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , 
 n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , 
 n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , 
 n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , 
 n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , 
 n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , 
 n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , 
 n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , 
 n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , 
 n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , 
 n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , 
 n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , 
 n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , 
 n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , 
 n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , 
 n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , 
 n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , 
 n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , 
 n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , 
 n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , 
 n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , 
 n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , 
 n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , 
 n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , 
 n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , 
 n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , 
 n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , 
 n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , 
 n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , 
 n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , 
 n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , 
 n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , 
 n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , 
 n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , 
 n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , 
 n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , 
 n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , 
 n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , 
 n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
 n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , 
 n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , 
 n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , 
 n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
 n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , 
 n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
 n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
 n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , 
 n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , 
 n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , 
 n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , 
 n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , 
 n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , 
 n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , 
 n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , 
 n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , 
 n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , 
 n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , 
 n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , 
 n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , 
 n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , 
 n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , 
 n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , 
 n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , 
 n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , 
 n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , 
 n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , 
 n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , 
 n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , 
 n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , 
 n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , 
 n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , 
 n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , 
 n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , 
 n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , 
 n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , 
 n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , 
 n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , 
 n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , 
 n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , 
 n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , 
 n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , 
 n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , 
 n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , 
 n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , 
 n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , 
 n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , 
 n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , 
 n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , 
 n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , 
 n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , 
 n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , 
 n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , 
 n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , 
 n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , 
 n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , 
 n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , 
 n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , 
 n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , 
 n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , 
 n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , 
 n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , 
 n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , 
 n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , 
 n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , 
 n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , 
 n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , 
 n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , 
 n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , 
 n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , 
 n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , 
 n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , 
 n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , 
 n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , 
 n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , 
 n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , 
 n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , 
 n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , 
 n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , 
 n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , 
 n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , 
 n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , 
 n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , 
 n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , 
 n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , 
 n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , 
 n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , 
 n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , 
 n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , 
 n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , 
 n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , 
 n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , 
 n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , 
 n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , 
 n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , 
 n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , 
 n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , 
 n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , 
 n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , 
 n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , 
 n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , 
 n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , 
 n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , 
 n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , 
 n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , 
 n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , 
 n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , 
 n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , 
 n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , 
 n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , 
 n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , 
 n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , 
 n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , 
 n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , 
 n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , 
 n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , 
 n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , 
 n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , 
 n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , 
 n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , 
 n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , 
 n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , 
 n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , 
 n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , 
 n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , 
 n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , 
 n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , 
 n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , 
 n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , 
 n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , 
 n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , 
 n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , 
 n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , 
 n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , 
 n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , 
 n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , 
 n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , 
 n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , 
 n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , 
 n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , 
 n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , 
 n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , 
 n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , 
 n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , 
 n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , 
 n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , 
 n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , 
 n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , 
 n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , 
 n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , 
 n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , 
 n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , 
 n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , 
 n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , 
 n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , 
 n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , 
 n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , 
 n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , 
 n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , 
 n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , 
 n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , 
 n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , 
 n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , 
 n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , 
 n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , 
 n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , 
 n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , 
 n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , 
 n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , 
 n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , 
 n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , 
 n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , 
 n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , 
 n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , 
 n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , 
 n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , 
 n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , 
 n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , 
 n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , 
 n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , 
 n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , 
 n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , 
 n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , 
 n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , 
 n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , 
 n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , 
 n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , 
 n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , 
 n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , 
 n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , 
 n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , 
 n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , 
 n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , 
 n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , 
 n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , 
 n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , 
 n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , 
 n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , 
 n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , 
 n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , 
 n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , 
 n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , 
 n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , 
 n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , 
 n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , 
 n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , 
 n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , 
 n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , 
 n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , 
 n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , 
 n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , 
 n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , 
 n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , 
 n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , 
 n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , 
 n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , 
 n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , 
 n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , 
 n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , 
 n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , 
 n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , 
 n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , 
 n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , 
 n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , 
 n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , 
 n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , 
 n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , 
 n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , 
 n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , 
 n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , 
 n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , 
 n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , 
 n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , 
 n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , 
 n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , 
 n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , 
 n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , 
 n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , 
 n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , 
 n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , 
 n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , 
 n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , 
 n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , 
 n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , 
 n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , 
 n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , 
 n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , 
 n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , 
 n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , 
 n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , 
 n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , 
 n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , 
 n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , 
 n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , 
 n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , 
 n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , 
 n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , 
 n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , 
 n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , 
 n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , 
 n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , 
 n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , 
 n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , 
 n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , 
 n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , 
 n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , 
 n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , 
 n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , 
 n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , 
 n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , 
 n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , 
 n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , 
 n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , 
 n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , 
 n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , 
 n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , 
 n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , 
 n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , 
 n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , 
 n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , 
 n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , 
 n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , 
 n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , 
 n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , 
 n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , 
 n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , 
 n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , 
 n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , 
 n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , 
 n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , 
 n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , 
 n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , 
 n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , 
 n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , 
 n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , 
 n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , 
 n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , 
 n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , 
 n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , 
 n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , 
 n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , 
 n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , 
 n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , 
 n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , 
 n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , 
 n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , 
 n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , 
 n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , 
 n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , 
 n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , 
 n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , 
 n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , 
 n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , 
 n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , 
 n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , 
 n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , 
 n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , 
 n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , 
 n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , 
 n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , 
 n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , 
 n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , 
 n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , 
 n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , 
 n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , 
 n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , 
 n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , 
 n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , 
 n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , 
 n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , 
 n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , 
 n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , 
 n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , 
 n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , 
 n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , 
 n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , 
 n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , 
 n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , 
 n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , 
 n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , 
 n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , 
 n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , 
 n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , 
 n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , 
 n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , 
 n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , 
 n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , 
 n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , 
 n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , 
 n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , 
 n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , 
 n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , 
 n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , 
 n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , 
 n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , 
 n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
 n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , 
 n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , 
 n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , 
 n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , 
 n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , 
 n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , 
 n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , 
 n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , 
 n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , 
 n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , 
 n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , 
 n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , 
 n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , 
 n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , 
 n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , 
 n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , 
 n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , 
 n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , 
 n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , 
 n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , 
 n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , 
 n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , 
 n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , 
 n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , 
 n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , 
 n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , 
 n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , 
 n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , 
 n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , 
 n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , 
 n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , 
 n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , 
 n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , 
 n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , 
 n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , 
 n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , 
 n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , 
 n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , 
 n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , 
 n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , 
 n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , 
 n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , 
 n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , 
 n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , 
 n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , 
 n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , 
 n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , 
 n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , 
 n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , 
 n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , 
 n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , 
 n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , 
 n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , 
 n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , 
 n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , 
 n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , 
 n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , 
 n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , 
 n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , 
 n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , 
 n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , 
 n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , 
 n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , 
 n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , 
 n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , 
 n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , 
 n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , 
 n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , 
 n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , 
 n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , 
 n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , 
 n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , 
 n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , 
 n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , 
 n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , 
 n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , 
 n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , 
 n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , 
 n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , 
 n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , 
 n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , 
 n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , 
 n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , 
 n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , 
 n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , 
 n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , 
 n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , 
 n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , 
 n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , 
 n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , 
 n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , 
 n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , 
 n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , 
 n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , 
 n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , 
 n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , 
 n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , 
 n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , 
 n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , 
 n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , 
 n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , 
 n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , 
 n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , 
 n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , 
 n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , 
 n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , 
 n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , 
 n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , 
 n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , 
 n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , 
 n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , 
 n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , 
 n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , 
 n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , 
 n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , 
 n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , 
 n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , 
 n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , 
 n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , 
 n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , 
 n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , 
 n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , 
 n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , 
 n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , 
 n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , 
 n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , 
 n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , 
 n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , 
 n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , 
 n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , 
 n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , 
 n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , 
 n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , 
 n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , 
 n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , 
 n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , 
 n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , 
 n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , 
 n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , 
 n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , 
 n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , 
 n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , 
 n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , 
 n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , 
 n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , 
 n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , 
 n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , 
 n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , 
 n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , 
 n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , 
 n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , 
 n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , 
 n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , 
 n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , 
 n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , 
 n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , 
 n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , 
 n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , 
 n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , 
 n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , 
 n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , 
 n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , 
 n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , 
 n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , 
 n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , 
 n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , 
 n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , 
 n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , 
 n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , 
 n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , 
 n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , 
 n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , 
 n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , 
 n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , 
 n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , 
 n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , 
 n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , 
 n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , 
 n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , 
 n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , 
 n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , 
 n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , 
 n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , 
 n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , 
 n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , 
 n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , 
 n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , 
 n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , 
 n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , 
 n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , 
 n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , 
 n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , 
 n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , 
 n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , 
 n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , 
 n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , 
 n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , 
 n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , 
 n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , 
 n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , 
 n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , 
 n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , 
 n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , 
 n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , 
 n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , 
 n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , 
 n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , 
 n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , 
 n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , 
 n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , 
 n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , 
 n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , 
 n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , 
 n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , 
 n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , 
 n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , 
 n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , 
 n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , 
 n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , 
 n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , 
 n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , 
 n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , 
 n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , 
 n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , 
 n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , 
 n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , 
 n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , 
 n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , 
 n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , 
 n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , 
 n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , 
 n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , 
 n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , 
 n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , 
 n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , 
 n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , 
 n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , 
 n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , 
 n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , 
 n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , 
 n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , 
 n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , 
 n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , 
 n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , 
 n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , 
 n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , 
 n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , 
 n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , 
 n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , 
 n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , 
 n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , 
 n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , 
 n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , 
 n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , 
 n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , 
 n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , 
 n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , 
 n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , 
 n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , 
 n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , 
 n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , 
 n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , 
 n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , 
 n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , 
 n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , 
 n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , 
 n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , 
 n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , 
 n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , 
 n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , 
 n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , 
 n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , 
 n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , 
 n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , 
 n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , 
 n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , 
 n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , 
 n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , 
 n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , 
 n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , 
 n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , 
 n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , 
 n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , 
 n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , 
 n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , 
 n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , 
 n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , 
 n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , 
 n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , 
 n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , 
 n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , 
 n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , 
 n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , 
 n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , 
 n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , 
 n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , 
 n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , 
 n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , 
 n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , 
 n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , 
 n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , 
 n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , 
 n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , 
 n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , 
 n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , 
 n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , 
 n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , 
 n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , 
 n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , 
 n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , 
 n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , 
 n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , 
 n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , 
 n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , 
 n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , 
 n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , 
 n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , 
 n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , 
 n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , 
 n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , 
 n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , 
 n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , 
 n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , 
 n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , 
 n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , 
 n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , 
 n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , 
 n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , 
 n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , 
 n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , 
 n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , 
 n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , 
 n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , 
 n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , 
 n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , 
 n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , 
 n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , 
 n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , 
 n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , 
 n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , 
 n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , 
 n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , 
 n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , 
 n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , 
 n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , 
 n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , 
 n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , 
 n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , 
 n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , 
 n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , 
 n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , 
 n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , 
 n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , 
 n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , 
 n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , 
 n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , 
 n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , 
 n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , 
 n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , 
 n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , 
 n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , 
 n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , 
 n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , 
 n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , 
 n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , 
 n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , 
 n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , 
 n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , 
 n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , 
 n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , 
 n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , 
 n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , 
 n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , 
 n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , 
 n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , 
 n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , 
 n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , 
 n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , 
 n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , 
 n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , 
 n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , 
 n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , 
 n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , 
 n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , 
 n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , 
 n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , 
 n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , 
 n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , 
 n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , 
 n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , 
 n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , 
 n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , 
 n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , 
 n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , 
 n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , 
 n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , 
 n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , 
 n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , 
 n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , 
 n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , 
 n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , 
 n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , 
 n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , 
 n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , 
 n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , 
 n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , 
 n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , 
 n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , 
 n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , 
 n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , 
 n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , 
 n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , 
 n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , 
 n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , 
 n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , 
 n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , 
 n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , 
 n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , 
 n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , 
 n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , 
 n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , 
 n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , 
 n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , 
 n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , 
 n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , 
 n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , 
 n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , 
 n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , 
 n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , 
 n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , 
 n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , 
 n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , 
 n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , 
 n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , 
 n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , 
 n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , 
 n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , 
 n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , 
 n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , 
 n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , 
 n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , 
 n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , 
 n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , 
 n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , 
 n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , 
 n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , 
 n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , 
 n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , 
 n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , 
 n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , 
 n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , 
 n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , 
 n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , 
 n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , 
 n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , 
 n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , 
 n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , 
 n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , 
 n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , 
 n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , 
 n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , 
 n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , 
 n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , 
 n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , 
 n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , 
 n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , 
 n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , 
 n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , 
 n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , 
 n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , 
 n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , 
 n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , 
 n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , 
 n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , 
 n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , 
 n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , 
 n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , 
 n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , 
 n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , 
 n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , 
 n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , 
 n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , 
 n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , 
 n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , 
 n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , 
 n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , 
 n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , 
 n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , 
 n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , 
 n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , 
 n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , 
 n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , 
 n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , 
 n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , 
 n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , 
 n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , 
 n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , 
 n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , 
 n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , 
 n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , 
 n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , 
 n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , 
 n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , 
 n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , 
 n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , 
 n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , 
 n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , 
 n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , 
 n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , 
 n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , 
 n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , 
 n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , 
 n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , 
 n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , 
 n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , 
 n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , 
 n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , 
 n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , 
 n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , 
 n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , 
 n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , 
 n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , 
 n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , 
 n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , 
 n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , 
 n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , 
 n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , 
 n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , 
 n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , 
 n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , 
 n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , 
 n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , 
 n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , 
 n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , 
 n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , 
 n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , 
 n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , 
 n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , 
 n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , 
 n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , 
 n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , 
 n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , 
 n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , 
 n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , 
 n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , 
 n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , 
 n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , 
 n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , 
 n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , 
 n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , 
 n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , 
 n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , 
 n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , 
 n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , 
 n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , 
 n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , 
 n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , 
 n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , 
 n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , 
 n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , 
 n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , 
 n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , 
 n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , 
 n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , 
 n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , 
 n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , 
 n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , 
 n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , 
 n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , 
 n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , 
 n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , 
 n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , 
 n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , 
 n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , 
 n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , 
 n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , 
 n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , 
 n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , 
 n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , 
 n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , 
 n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , 
 n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , 
 n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , 
 n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , 
 n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , 
 n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , 
 n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , 
 n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , 
 n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , 
 n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , 
 n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , 
 n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , 
 n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , 
 n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , 
 n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , 
 n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , 
 n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , 
 n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , 
 n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , 
 n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , 
 n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , 
 n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , 
 n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , 
 n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , 
 n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , 
 n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , 
 n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , 
 n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , 
 n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , 
 n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , 
 n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , 
 n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , 
 n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , 
 n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , 
 n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , 
 n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , 
 n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , 
 n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , 
 n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , 
 n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , 
 n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , 
 n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , 
 n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , 
 n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , 
 n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , 
 n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , 
 n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , 
 n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , 
 n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , 
 n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , 
 n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , 
 n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , 
 n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , 
 n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , 
 n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , 
 n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , 
 n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , 
 n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , 
 n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , 
 n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , 
 n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , 
 n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , 
 n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , 
 n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , 
 n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , 
 n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , 
 n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , 
 n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , 
 n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , 
 n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , 
 n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , 
 n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , 
 n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , 
 n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , 
 n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , 
 n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , 
 n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , 
 n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , 
 n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , 
 n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , 
 n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , 
 n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , 
 n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , 
 n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , 
 n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , 
 n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , 
 n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , 
 n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , 
 n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , 
 n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , 
 n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , 
 n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , 
 n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , 
 n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , 
 n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , 
 n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , 
 n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , 
 n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , 
 n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , 
 n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , 
 n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , 
 n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , 
 n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , 
 n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , 
 n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , 
 n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , 
 n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , 
 n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , 
 n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , 
 n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , 
 n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , 
 n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , 
 n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , 
 n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , 
 n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , 
 n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , 
 n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , 
 n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , 
 n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , 
 n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , 
 n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , 
 n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , 
 n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , 
 n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , 
 n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , 
 n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , 
 n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , 
 n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , 
 n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , 
 n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , 
 n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , 
 n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , 
 n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , 
 n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , 
 n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , 
 n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , 
 n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , 
 n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , 
 n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , 
 n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , 
 n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , 
 n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , 
 n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , 
 n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , 
 n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , 
 n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , 
 n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , 
 n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , 
 n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , 
 n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , 
 n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , 
 n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , 
 n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , 
 n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , 
 n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , 
 n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , 
 n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , 
 n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , 
 n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , 
 n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , 
 n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , 
 n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , 
 n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , 
 n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , 
 n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , 
 n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , 
 n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , 
 n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , 
 n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , 
 n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , 
 n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , 
 n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , 
 n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , 
 n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , 
 n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , 
 n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , 
 n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , 
 n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , 
 n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , 
 n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , 
 n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , 
 n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , 
 n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , 
 n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , 
 n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , 
 n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , 
 n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , 
 n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , 
 n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , 
 n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , 
 n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , 
 n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , 
 n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , 
 n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , 
 n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , 
 n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , 
 n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , 
 n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , 
 n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , 
 n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , 
 n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , 
 n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , 
 n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , 
 n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , 
 n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , 
 n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , 
 n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , 
 n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , 
 n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , 
 n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , 
 n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , 
 n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , 
 n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , 
 n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , 
 n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , 
 n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , 
 n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , 
 n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , 
 n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , 
 n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , 
 n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , 
 n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , 
 n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , 
 n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , 
 n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , 
 n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , 
 n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , 
 n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , 
 n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , 
 n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , 
 n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , 
 n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , 
 n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , 
 n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , 
 n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , 
 n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , 
 n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , 
 n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , 
 n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , 
 n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , 
 n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , 
 n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , 
 n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , 
 n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , 
 n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , 
 n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , 
 n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , 
 n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , 
 n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , 
 n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , 
 n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , 
 n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , 
 n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , 
 n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , 
 n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , 
 n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , 
 n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , 
 n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , 
 n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , 
 n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , 
 n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , 
 n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , 
 n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , 
 n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , 
 n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , 
 n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , 
 n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , 
 n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , 
 n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , 
 n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , 
 n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , 
 n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , 
 n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , 
 n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , 
 n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , 
 n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , 
 n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , 
 n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , 
 n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , 
 n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , 
 n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , 
 n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , 
 n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , 
 n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , 
 n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , 
 n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , 
 n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , 
 n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , 
 n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , 
 n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , 
 n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , 
 n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , 
 n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , 
 n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , 
 n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , 
 n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , 
 n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , 
 n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , 
 n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , 
 n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , 
 n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , 
 n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , 
 n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , 
 n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , 
 n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , 
 n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , 
 n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , 
 n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , 
 n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , 
 n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , 
 n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , 
 n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , 
 n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , 
 n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , 
 n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , 
 n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , 
 n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , 
 n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , 
 n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , 
 n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , 
 n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , 
 n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , 
 n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , 
 n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , 
 n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , 
 n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , 
 n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , 
 n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , 
 n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , 
 n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , 
 n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , 
 n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , 
 n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , 
 n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , 
 n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , 
 n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , 
 n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , 
 n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , 
 n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , 
 n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , 
 n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , 
 n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , 
 n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , 
 n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , 
 n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , 
 n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , 
 n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , 
 n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , 
 n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , 
 n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , 
 n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , 
 n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , 
 n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , 
 n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , 
 n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , 
 n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , 
 n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , 
 n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , 
 n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , 
 n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , 
 n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , 
 n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , 
 n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , 
 n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , 
 n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , 
 n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , 
 n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , 
 n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , 
 n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , 
 n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , 
 n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , 
 n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , 
 n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , 
 n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , 
 n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , 
 n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , 
 n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , 
 n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , 
 n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , 
 n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , 
 n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , 
 n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , 
 n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , 
 n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , 
 n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , 
 n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , 
 n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , 
 n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , 
 n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , 
 n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , 
 n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , 
 n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , 
 n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , 
 n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , 
 n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , 
 n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , 
 n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , 
 n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , 
 n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , 
 n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , 
 n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , 
 n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , 
 n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , 
 n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , 
 n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , 
 n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , 
 n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , 
 n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , 
 n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , 
 n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , 
 n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , 
 n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , 
 n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , 
 n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , 
 n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , 
 n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , 
 n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , 
 n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , 
 n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , 
 n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , 
 n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , 
 n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , 
 n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , 
 n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , 
 n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , 
 n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , 
 n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , 
 n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , 
 n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , 
 n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , 
 n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , 
 n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , 
 n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , 
 n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , 
 n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , 
 n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , 
 n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , 
 n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , 
 n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , 
 n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , 
 n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , 
 n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , 
 n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , 
 n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , 
 n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , 
 n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , 
 n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , 
 n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , 
 n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , 
 n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , 
 n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , 
 n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , 
 n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , 
 n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , 
 n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , 
 n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , 
 n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , 
 n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , 
 n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , 
 n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , 
 n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , 
 n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , 
 n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , 
 n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , 
 n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , 
 n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , 
 n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , 
 n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , 
 n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , 
 n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , 
 n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , 
 n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , 
 n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , 
 n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , 
 n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , 
 n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , 
 n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , 
 n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , 
 n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , 
 n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , 
 n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , 
 n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , 
 n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , 
 n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , 
 n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , 
 n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , 
 n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , 
 n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , 
 n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , 
 n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , 
 n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , 
 n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , 
 n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , 
 n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , 
 n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , 
 n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , 
 n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , 
 n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , 
 n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , 
 n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , 
 n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , 
 n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , 
 n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , 
 n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , 
 n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , 
 n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , 
 n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , 
 n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , 
 n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , 
 n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , 
 n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , 
 n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , 
 n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , 
 n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , 
 n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , 
 n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , 
 n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , 
 n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , 
 n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , 
 n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , 
 n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , 
 n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , 
 n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , 
 n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , 
 n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , 
 n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , 
 n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , 
 n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , 
 n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , 
 n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , 
 n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , 
 n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , 
 n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , 
 n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , 
 n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , 
 n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , 
 n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , 
 n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , 
 n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , 
 n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , 
 n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , 
 n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , 
 n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , 
 n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , 
 n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , 
 n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , 
 n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , 
 n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , 
 n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , 
 n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , 
 n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , 
 n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , 
 n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , 
 n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , 
 n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , 
 n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , 
 n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , 
 n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , 
 n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , 
 n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , 
 n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , 
 n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , 
 n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , 
 n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , 
 n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , 
 n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , 
 n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , 
 n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , 
 n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , 
 n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , 
 n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , 
 n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , 
 n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , 
 n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , 
 n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , 
 n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , 
 n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , 
 n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , 
 n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , 
 n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , 
 n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , 
 n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , 
 n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , 
 n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , 
 n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , 
 n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , 
 n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , 
 n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , 
 n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , 
 n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , 
 n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , 
 n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , 
 n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , 
 n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , 
 n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , 
 n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , 
 n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , 
 n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , 
 n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , 
 n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , 
 n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , 
 n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , 
 n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , 
 n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , 
 n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , 
 n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , 
 n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , 
 n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , 
 n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , 
 n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , 
 n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , 
 n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , 
 n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , 
 n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , 
 n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , 
 n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , 
 n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , 
 n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , 
 n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , 
 n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , 
 n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , 
 n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , 
 n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , 
 n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , 
 n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , 
 n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , 
 n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , 
 n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , 
 n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , 
 n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , 
 n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , 
 n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , 
 n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , 
 n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , 
 n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , 
 n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , 
 n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , 
 n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , 
 n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , 
 n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , 
 n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , 
 n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , 
 n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , 
 n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , 
 n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , 
 n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , 
 n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , 
 n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , 
 n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , 
 n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , 
 n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , 
 n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , 
 n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , 
 n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , 
 n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , 
 n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , 
 n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , 
 n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , 
 n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , 
 n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , 
 n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , 
 n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , 
 n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , 
 n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , 
 n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , 
 n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , 
 n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , 
 n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , 
 n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , 
 n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , 
 n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , 
 n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
 n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
 n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
 n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
 n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
 n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
 n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
 n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
 n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , 
 n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , 
 n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , 
 n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , 
 n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , 
 n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , 
 n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , 
 n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , 
 n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , 
 n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , 
 n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , 
 n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
 n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , 
 n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , 
 n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , 
 n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , 
 n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , 
 n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , 
 n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , 
 n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , 
 n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , 
 n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , 
 n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , 
 n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , 
 n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , 
 n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , 
 n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , 
 n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , 
 n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , 
 n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , 
 n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , 
 n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , 
 n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , 
 n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , 
 n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , 
 n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , 
 n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , 
 n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , 
 n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , 
 n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , 
 n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , 
 n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , 
 n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , 
 n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , 
 n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , 
 n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , 
 n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , 
 n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , 
 n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , 
 n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , 
 n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , 
 n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , 
 n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , 
 n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , 
 n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , 
 n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , 
 n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , 
 n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , 
 n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , 
 n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , 
 n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , 
 n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , 
 n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , 
 n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , 
 n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , 
 n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , 
 n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , 
 n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , 
 n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , 
 n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , 
 n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , 
 n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , 
 n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , 
 n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , 
 n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , 
 n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , 
 n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , 
 n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , 
 n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , 
 n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , 
 n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , 
 n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , 
 n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , 
 n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , 
 n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , 
 n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , 
 n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , 
 n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , 
 n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , 
 n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , 
 n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , 
 n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , 
 n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , 
 n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , 
 n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , 
 n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , 
 n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , 
 n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , 
 n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , 
 n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , 
 n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , 
 n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , 
 n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , 
 n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , 
 n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , 
 n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , 
 n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , 
 n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , 
 n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , 
 n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , 
 n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , 
 n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , 
 n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , 
 n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , 
 n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , 
 n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , 
 n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , 
 n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , 
 n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , 
 n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , 
 n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , 
 n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , 
 n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , 
 n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , 
 n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , 
 n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , 
 n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , 
 n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , 
 n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , 
 n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , 
 n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , 
 n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , 
 n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , 
 n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , 
 n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , 
 n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , 
 n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , 
 n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , 
 n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , 
 n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , 
 n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , 
 n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , 
 n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , 
 n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , 
 n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , 
 n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , 
 n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , 
 n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , 
 n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , 
 n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , 
 n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , 
 n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , 
 n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , 
 n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , 
 n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , 
 n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , 
 n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , 
 n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , 
 n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , 
 n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , 
 n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , 
 n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , 
 n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , 
 n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , 
 n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , 
 n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , 
 n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , 
 n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , 
 n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , 
 n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , 
 n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , 
 n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , 
 n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , 
 n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , 
 n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , 
 n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , 
 n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , 
 n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , 
 n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , 
 n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , 
 n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , 
 n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , 
 n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , 
 n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , 
 n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , 
 n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , 
 n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , 
 n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , 
 n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , 
 n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , 
 n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , 
 n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , 
 n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , 
 n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , 
 n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , 
 n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , 
 n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , 
 n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , 
 n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , 
 n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , 
 n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , 
 n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , 
 n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , 
 n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , 
 n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , 
 n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , 
 n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , 
 n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , 
 n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , 
 n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , 
 n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , 
 n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , 
 n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , 
 n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , 
 n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , 
 n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , 
 n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , 
 n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , 
 n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , 
 n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , 
 n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , 
 n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , 
 n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , 
 n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , 
 n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , 
 n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , 
 n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , 
 n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , 
 n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , 
 n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , 
 n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , 
 n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , 
 n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , 
 n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , 
 n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , 
 n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , 
 n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , 
 n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , 
 n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , 
 n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , 
 n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , 
 n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , 
 n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , 
 n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , 
 n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , 
 n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , 
 n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , 
 n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , 
 n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , 
 n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , 
 n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , 
 n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , 
 n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , 
 n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , 
 n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , 
 n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , 
 n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , 
 n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , 
 n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , 
 n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , 
 n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , 
 n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , 
 n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , 
 n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , 
 n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , 
 n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , 
 n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , 
 n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , 
 n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , 
 n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , 
 n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , 
 n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , 
 n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , 
 n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , 
 n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , 
 n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , 
 n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , 
 n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , 
 n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , 
 n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , 
 n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , 
 n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , 
 n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , 
 n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , 
 n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , 
 n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , 
 n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , 
 n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , 
 n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , 
 n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , 
 n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , 
 n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , 
 n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , 
 n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , 
 n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , 
 n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , 
 n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , 
 n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , 
 n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , 
 n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , 
 n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , 
 n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , 
 n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , 
 n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , 
 n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , 
 n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , 
 n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , 
 n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , 
 n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , 
 n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , 
 n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , 
 n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , 
 n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , 
 n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
 n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , 
 n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , 
 n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , 
 n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , 
 n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , 
 n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , 
 n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , 
 n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , 
 n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , 
 n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , 
 n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , 
 n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , 
 n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , 
 n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , 
 n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , 
 n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , 
 n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , 
 n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , 
 n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , 
 n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , 
 n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , 
 n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , 
 n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , 
 n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , 
 n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , 
 n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , 
 n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , 
 n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , 
 n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , 
 n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , 
 n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , 
 n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , 
 n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , 
 n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , 
 n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , 
 n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , 
 n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , 
 n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , 
 n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , 
 n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , 
 n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , 
 C0n , C0 , C1n , C1 ;
buf ( n454 , n0 );
buf ( n455 , n1 );
buf ( n456 , n2 );
buf ( n457 , n3 );
buf ( n458 , n4 );
buf ( n459 , n5 );
buf ( n460 , n6 );
buf ( n461 , n7 );
buf ( n462 , n8 );
buf ( n463 , n9 );
buf ( n464 , n10 );
buf ( n465 , n11 );
buf ( n466 , n12 );
buf ( n467 , n13 );
buf ( n468 , n14 );
buf ( n469 , n15 );
buf ( n470 , n16 );
buf ( n471 , n17 );
buf ( n472 , n18 );
buf ( n473 , n19 );
buf ( n474 , n20 );
buf ( n475 , n21 );
buf ( n476 , n22 );
buf ( n477 , n23 );
buf ( n478 , n24 );
buf ( n479 , n25 );
buf ( n480 , n26 );
buf ( n481 , n27 );
buf ( n482 , n28 );
buf ( n483 , n29 );
buf ( n484 , n30 );
buf ( n485 , n31 );
buf ( n486 , n32 );
buf ( n487 , n33 );
buf ( n488 , n34 );
buf ( n489 , n35 );
buf ( n490 , n36 );
buf ( n491 , n37 );
buf ( n492 , n38 );
buf ( n493 , n39 );
buf ( n494 , n40 );
buf ( n495 , n41 );
buf ( n496 , n42 );
buf ( n497 , n43 );
buf ( n498 , n44 );
buf ( n499 , n45 );
buf ( n500 , n46 );
buf ( n501 , n47 );
buf ( n502 , n48 );
buf ( n503 , n49 );
buf ( n504 , n50 );
buf ( n505 , n51 );
buf ( n506 , n52 );
buf ( n507 , n53 );
buf ( n508 , n54 );
buf ( n509 , n55 );
buf ( n510 , n56 );
buf ( n511 , n57 );
buf ( n512 , n58 );
buf ( n513 , n59 );
buf ( n514 , n60 );
buf ( n515 , n61 );
buf ( n516 , n62 );
buf ( n517 , n63 );
buf ( n518 , n64 );
buf ( n519 , n65 );
buf ( n520 , n66 );
buf ( n521 , n67 );
buf ( n522 , n68 );
buf ( n523 , n69 );
buf ( n524 , n70 );
buf ( n525 , n71 );
buf ( n526 , n72 );
buf ( n527 , n73 );
buf ( n528 , n74 );
buf ( n529 , n75 );
buf ( n530 , n76 );
buf ( n531 , n77 );
buf ( n532 , n78 );
buf ( n533 , n79 );
buf ( n534 , n80 );
buf ( n535 , n81 );
buf ( n536 , n82 );
buf ( n537 , n83 );
buf ( n538 , n84 );
buf ( n539 , n85 );
buf ( n540 , n86 );
buf ( n541 , n87 );
buf ( n542 , n88 );
buf ( n543 , n89 );
buf ( n544 , n90 );
buf ( n545 , n91 );
buf ( n546 , n92 );
buf ( n547 , n93 );
buf ( n548 , n94 );
buf ( n549 , n95 );
buf ( n550 , n96 );
buf ( n551 , n97 );
buf ( n552 , n98 );
buf ( n99 , n553 );
buf ( n100 , n554 );
buf ( n101 , n555 );
buf ( n102 , n556 );
buf ( n103 , n557 );
buf ( n104 , n558 );
buf ( n105 , n559 );
buf ( n106 , n560 );
buf ( n107 , n561 );
buf ( n108 , n562 );
buf ( n109 , n563 );
buf ( n110 , n564 );
buf ( n111 , n565 );
buf ( n112 , n566 );
buf ( n113 , n567 );
buf ( n114 , n568 );
buf ( n115 , n569 );
buf ( n116 , n570 );
buf ( n117 , n571 );
buf ( n118 , n572 );
buf ( n119 , n573 );
buf ( n120 , n574 );
buf ( n121 , n575 );
buf ( n122 , n576 );
buf ( n123 , n577 );
buf ( n124 , n578 );
buf ( n125 , n579 );
buf ( n126 , n580 );
buf ( n127 , n581 );
buf ( n128 , n582 );
buf ( n129 , n583 );
buf ( n130 , n584 );
buf ( n131 , n585 );
buf ( n132 , n586 );
buf ( n133 , n587 );
buf ( n134 , n588 );
buf ( n135 , n589 );
buf ( n136 , n590 );
buf ( n137 , n591 );
buf ( n138 , n592 );
buf ( n139 , n593 );
buf ( n140 , n594 );
buf ( n141 , n595 );
buf ( n142 , n596 );
buf ( n143 , n597 );
buf ( n144 , n598 );
buf ( n145 , n599 );
buf ( n146 , n600 );
buf ( n147 , n601 );
buf ( n148 , n602 );
buf ( n149 , n603 );
buf ( n150 , n604 );
buf ( n151 , n605 );
buf ( n152 , n606 );
buf ( n153 , n607 );
buf ( n154 , n608 );
buf ( n155 , n609 );
buf ( n156 , n610 );
buf ( n157 , n611 );
buf ( n158 , n612 );
buf ( n159 , n613 );
buf ( n160 , n614 );
buf ( n161 , n615 );
buf ( n162 , n616 );
buf ( n163 , n617 );
buf ( n164 , n618 );
buf ( n165 , n619 );
buf ( n166 , n620 );
buf ( n167 , n621 );
buf ( n168 , n622 );
buf ( n169 , n623 );
buf ( n170 , n624 );
buf ( n171 , n625 );
buf ( n172 , n626 );
buf ( n173 , n627 );
buf ( n174 , n628 );
buf ( n175 , n629 );
buf ( n176 , n630 );
buf ( n177 , n631 );
buf ( n178 , n632 );
buf ( n179 , n633 );
buf ( n180 , n634 );
buf ( n181 , n635 );
buf ( n182 , n636 );
buf ( n183 , n637 );
buf ( n184 , n638 );
buf ( n185 , n639 );
buf ( n186 , n640 );
buf ( n187 , n641 );
buf ( n188 , n642 );
buf ( n189 , n643 );
buf ( n190 , n644 );
buf ( n191 , n645 );
buf ( n192 , n646 );
buf ( n193 , n647 );
buf ( n194 , n648 );
buf ( n195 , n649 );
buf ( n196 , n650 );
buf ( n197 , n651 );
buf ( n198 , n652 );
buf ( n199 , n653 );
buf ( n200 , n654 );
buf ( n201 , n655 );
buf ( n202 , n656 );
buf ( n203 , n657 );
buf ( n204 , n658 );
buf ( n205 , n659 );
buf ( n206 , n660 );
buf ( n207 , n661 );
buf ( n208 , n662 );
buf ( n209 , n663 );
buf ( n210 , n664 );
buf ( n211 , n665 );
buf ( n212 , n666 );
buf ( n213 , n667 );
buf ( n214 , n668 );
buf ( n215 , n669 );
buf ( n216 , n670 );
buf ( n217 , n671 );
buf ( n218 , n672 );
buf ( n219 , n673 );
buf ( n220 , n674 );
buf ( n221 , n675 );
buf ( n222 , n676 );
buf ( n223 , n677 );
buf ( n224 , n678 );
buf ( n225 , n679 );
buf ( n226 , n680 );
buf ( n553 , C0 );
buf ( n554 , C0 );
buf ( n555 , C0 );
buf ( n556 , C0 );
buf ( n557 , C0 );
buf ( n558 , C0 );
buf ( n559 , C0 );
buf ( n560 , C0 );
buf ( n561 , C0 );
buf ( n562 , C0 );
buf ( n563 , C0 );
buf ( n564 , C0 );
buf ( n565 , C0 );
buf ( n566 , C0 );
buf ( n567 , C0 );
buf ( n568 , C0 );
buf ( n569 , n28762 );
buf ( n570 , n28774 );
buf ( n571 , n28764 );
buf ( n572 , n28631 );
buf ( n573 , n27609 );
buf ( n574 , n28549 );
buf ( n575 , n28496 );
buf ( n576 , n28457 );
buf ( n577 , n25261 );
buf ( n578 , n25395 );
buf ( n579 , n25436 );
buf ( n580 , n25296 );
buf ( n581 , n25469 );
buf ( n582 , n25465 );
buf ( n583 , n25498 );
buf ( n584 , n29314 );
buf ( n585 , n16710 );
buf ( n586 , n16718 );
buf ( n587 , n15982 );
buf ( n588 , n16057 );
buf ( n589 , n16072 );
buf ( n590 , n16019 );
buf ( n591 , n16758 );
buf ( n592 , n17474 );
buf ( n593 , n17447 );
buf ( n594 , n17453 );
buf ( n595 , n17484 );
buf ( n596 , n16880 );
buf ( n597 , n16786 );
buf ( n598 , n16835 );
buf ( n599 , n16846 );
buf ( n600 , n16817 );
buf ( n601 , n16895 );
buf ( n602 , n16936 );
buf ( n603 , n16977 );
buf ( n604 , n17014 );
buf ( n605 , n17049 );
buf ( n606 , n17086 );
buf ( n607 , n17123 );
buf ( n608 , n17161 );
buf ( n609 , n17196 );
buf ( n610 , n17228 );
buf ( n611 , n17247 );
buf ( n612 , n29186 );
buf ( n613 , n29196 );
buf ( n614 , n29298 );
buf ( n615 , n29200 );
buf ( n616 , n27310 );
buf ( n617 , C0 );
buf ( n618 , C0 );
buf ( n619 , C0 );
buf ( n620 , C0 );
buf ( n621 , C0 );
buf ( n622 , C0 );
buf ( n623 , C0 );
buf ( n624 , C0 );
buf ( n625 , C0 );
buf ( n626 , C0 );
buf ( n627 , C0 );
buf ( n628 , C0 );
buf ( n629 , C0 );
buf ( n630 , C0 );
buf ( n631 , C0 );
buf ( n632 , C0 );
buf ( n633 , n29241 );
buf ( n634 , n29071 );
buf ( n635 , n29062 );
buf ( n636 , n29117 );
buf ( n637 , n29283 );
buf ( n638 , n29050 );
buf ( n639 , n29164 );
buf ( n640 , n29114 );
buf ( n641 , n29088 );
buf ( n642 , n29133 );
buf ( n643 , n29028 );
buf ( n644 , n29151 );
buf ( n645 , n27022 );
buf ( n646 , n28986 );
buf ( n647 , n27083 );
buf ( n648 , n29003 );
buf ( n649 , n28976 );
buf ( n650 , n27150 );
buf ( n651 , n28959 );
buf ( n652 , n27182 );
buf ( n653 , n23839 );
buf ( n654 , n29292 );
buf ( n655 , n29313 );
buf ( n656 , n23883 );
buf ( n657 , n23894 );
buf ( n658 , n23906 );
buf ( n659 , n29234 );
buf ( n660 , n23933 );
buf ( n661 , n29224 );
buf ( n662 , n23950 );
buf ( n663 , n27040 );
buf ( n664 , n27047 );
buf ( n665 , n27066 );
buf ( n666 , n27095 );
buf ( n667 , n29266 );
buf ( n668 , n27109 );
buf ( n669 , n29180 );
buf ( n670 , n29246 );
buf ( n671 , n27121 );
buf ( n672 , n27132 );
buf ( n673 , n27157 );
buf ( n674 , n29251 );
buf ( n675 , n27325 );
buf ( n676 , n29309 );
buf ( n677 , n29205 );
buf ( n678 , n29271 );
buf ( n679 , n29297 );
buf ( n680 , n29192 );
not ( n681 , n504 );
nand ( n682 , n681 , n503 );
not ( n683 , n682 );
xor ( n684 , n503 , n520 );
and ( n685 , n683 , n684 );
not ( n686 , n685 );
not ( n687 , n502 );
not ( n688 , n503 );
not ( n689 , n688 );
or ( n690 , n687 , n689 );
not ( n691 , n502 );
nand ( n692 , n691 , n503 );
nand ( n693 , n690 , n692 );
buf ( n694 , n693 );
nand ( n695 , n520 , n694 );
nand ( n696 , n686 , n695 );
xor ( n697 , n503 , n519 );
not ( n698 , n697 );
nand ( n699 , n503 , n504 );
nor ( n700 , n698 , n699 , n520 );
or ( n701 , n696 , n700 );
not ( n702 , n697 );
not ( n703 , n683 );
or ( n704 , n702 , n703 );
xor ( n705 , n518 , n503 );
nand ( n706 , n705 , n504 );
nand ( n707 , n704 , n706 );
nand ( n708 , n701 , n707 );
nand ( n709 , C1 , n708 );
not ( n710 , n709 );
not ( n711 , n504 );
xor ( n712 , n503 , n517 );
not ( n713 , n712 );
or ( n714 , n711 , n713 );
nand ( n715 , n705 , n683 );
nand ( n716 , n714 , n715 );
or ( n717 , n520 , n502 );
nand ( n718 , n717 , n503 );
nand ( n719 , n520 , n502 );
and ( n720 , n718 , n719 , n501 );
and ( n721 , n716 , n720 );
not ( n722 , n716 );
not ( n723 , n720 );
and ( n724 , n722 , n723 );
nor ( n725 , n721 , n724 );
xor ( n726 , n501 , n520 );
not ( n727 , n726 );
and ( n728 , n502 , n503 );
not ( n729 , n502 );
not ( n730 , n503 );
and ( n731 , n729 , n730 );
nor ( n732 , n728 , n731 );
not ( n733 , n732 );
xor ( n734 , n501 , n502 );
nand ( n735 , n733 , n734 );
not ( n736 , n735 );
not ( n737 , n736 );
or ( n738 , n727 , n737 );
xor ( n739 , n519 , n501 );
nand ( n740 , n739 , n694 );
nand ( n741 , n738 , n740 );
nor ( n742 , n725 , n741 );
not ( n743 , n742 );
not ( n744 , n743 );
or ( n745 , n710 , n744 );
nand ( n746 , n741 , n725 );
nand ( n747 , n745 , n746 );
not ( n748 , n747 );
xor ( n749 , n500 , n501 );
and ( n750 , n749 , n520 );
not ( n751 , n750 );
nand ( n752 , n734 , n739 );
or ( n753 , n752 , n694 );
not ( n754 , n518 );
not ( n755 , n501 );
not ( n756 , n755 );
or ( n757 , n754 , n756 );
not ( n758 , n518 );
nand ( n759 , n758 , n501 );
nand ( n760 , n757 , n759 );
xor ( n761 , n502 , n503 );
nand ( n762 , n760 , n761 );
nand ( n763 , n753 , n762 );
not ( n764 , n763 );
not ( n765 , n764 );
or ( n766 , n751 , n765 );
not ( n767 , n750 );
nand ( n768 , n767 , n763 );
nand ( n769 , n766 , n768 );
not ( n770 , n504 );
xor ( n771 , n503 , n516 );
not ( n772 , n771 );
or ( n773 , n770 , n772 );
nand ( n774 , n712 , n683 );
nand ( n775 , n773 , n774 );
not ( n776 , n775 );
and ( n777 , n769 , n776 );
not ( n778 , n769 );
and ( n779 , n778 , n775 );
nor ( n780 , n777 , n779 );
and ( n781 , n716 , n720 );
and ( n782 , n780 , n781 );
nand ( n783 , n748 , n782 );
not ( n784 , n781 );
nand ( n785 , n780 , n784 );
not ( n786 , n785 );
nor ( n787 , n780 , n784 );
or ( n788 , n786 , n787 );
nand ( n789 , n788 , n747 );
nor ( n790 , n780 , n781 );
nand ( n791 , n748 , n790 );
nand ( n792 , n783 , n789 , n791 );
not ( n793 , n455 );
nand ( n794 , n792 , n793 );
not ( n795 , n761 );
xor ( n796 , n513 , n501 );
not ( n797 , n796 );
or ( n798 , n795 , n797 );
xor ( n799 , n501 , n514 );
not ( n800 , n503 );
nand ( n801 , n800 , n502 );
nand ( n802 , n503 , n691 );
nand ( n803 , n734 , n799 , n801 , n802 );
nand ( n804 , n798 , n803 );
not ( n805 , n497 );
or ( n806 , n520 , n496 );
not ( n807 , n806 );
or ( n808 , n805 , n807 );
nand ( n809 , n520 , n496 );
and ( n810 , n809 , n495 );
nand ( n811 , n808 , n810 );
not ( n812 , n811 );
and ( n813 , n804 , n812 );
xor ( n814 , n494 , n495 );
nand ( n815 , n814 , n520 );
and ( n816 , n517 , n497 );
not ( n817 , n517 );
not ( n818 , n497 );
and ( n819 , n817 , n818 );
nor ( n820 , n816 , n819 );
not ( n821 , n820 );
xor ( n822 , n498 , n499 );
not ( n823 , n822 );
not ( n824 , n497 );
not ( n825 , n498 );
not ( n826 , n825 );
or ( n827 , n824 , n826 );
not ( n828 , n497 );
nand ( n829 , n828 , n498 );
nand ( n830 , n827 , n829 );
nand ( n831 , n823 , n830 );
not ( n832 , n831 );
not ( n833 , n832 );
or ( n834 , n821 , n833 );
xor ( n835 , n516 , n497 );
buf ( n836 , n822 );
nand ( n837 , n835 , n836 );
nand ( n838 , n834 , n837 );
xor ( n839 , n815 , n838 );
and ( n840 , n796 , n734 );
not ( n841 , n840 );
not ( n842 , n694 );
not ( n843 , n842 );
or ( n844 , n841 , n843 );
not ( n845 , n733 );
xor ( n846 , n512 , n501 );
nand ( n847 , n845 , n846 );
nand ( n848 , n844 , n847 );
xnor ( n849 , n839 , n848 );
xor ( n850 , n813 , n849 );
xor ( n851 , n520 , n495 );
not ( n852 , n851 );
not ( n853 , n497 );
nor ( n854 , n853 , n496 );
not ( n855 , n854 );
nand ( n856 , n818 , n496 );
xor ( n857 , n496 , n495 );
nand ( n858 , n855 , n856 , n857 );
not ( n859 , n858 );
not ( n860 , n859 );
or ( n861 , n852 , n860 );
and ( n862 , n496 , n497 );
not ( n863 , n496 );
not ( n864 , n497 );
and ( n865 , n863 , n864 );
nor ( n866 , n862 , n865 );
buf ( n867 , n866 );
xor ( n868 , n519 , n495 );
nand ( n869 , n867 , n868 );
nand ( n870 , n861 , n869 );
not ( n871 , n870 );
and ( n872 , n503 , n512 );
not ( n873 , n503 );
not ( n874 , n512 );
and ( n875 , n873 , n874 );
nor ( n876 , n872 , n875 );
not ( n877 , n876 );
not ( n878 , n683 );
or ( n879 , n877 , n878 );
xor ( n880 , n511 , n503 );
nand ( n881 , n880 , n504 );
nand ( n882 , n879 , n881 );
not ( n883 , n882 );
or ( n884 , n871 , n883 );
nor ( n885 , n882 , n870 );
xor ( n886 , n518 , n497 );
not ( n887 , n886 );
and ( n888 , n823 , n830 );
not ( n889 , n888 );
or ( n890 , n887 , n889 );
nand ( n891 , n836 , n820 );
nand ( n892 , n890 , n891 );
not ( n893 , n892 );
or ( n894 , n885 , n893 );
nand ( n895 , n884 , n894 );
xor ( n896 , n850 , n895 );
not ( n897 , n504 );
xor ( n898 , n503 , n510 );
not ( n899 , n898 );
or ( n900 , n897 , n899 );
nand ( n901 , n880 , n683 );
nand ( n902 , n900 , n901 );
not ( n903 , n902 );
not ( n904 , n903 );
not ( n905 , n868 );
not ( n906 , n828 );
not ( n907 , n496 );
not ( n908 , n907 );
or ( n909 , n906 , n908 );
nand ( n910 , n496 , n497 );
nand ( n911 , n909 , n910 );
and ( n912 , n911 , n857 );
not ( n913 , n912 );
or ( n914 , n905 , n913 );
and ( n915 , n518 , n495 );
not ( n916 , n518 );
not ( n917 , n495 );
and ( n918 , n916 , n917 );
nor ( n919 , n915 , n918 );
nand ( n920 , n866 , n919 );
nand ( n921 , n914 , n920 );
not ( n922 , n921 );
or ( n923 , n904 , n922 );
not ( n924 , n921 );
nand ( n925 , n924 , n902 );
nand ( n926 , n923 , n925 );
xor ( n927 , n499 , n515 );
not ( n928 , n927 );
and ( n929 , n500 , n501 );
not ( n930 , n500 );
not ( n931 , n501 );
and ( n932 , n930 , n931 );
nor ( n933 , n929 , n932 );
not ( n934 , n933 );
not ( n935 , n500 );
not ( n936 , n499 );
nand ( n937 , n935 , n936 );
nand ( n938 , n500 , n499 );
and ( n939 , n934 , n937 , n938 );
not ( n940 , n939 );
or ( n941 , n928 , n940 );
xor ( n942 , n514 , n499 );
nand ( n943 , n749 , n942 );
nand ( n944 , n941 , n943 );
xnor ( n945 , n926 , n944 );
not ( n946 , n683 );
xor ( n947 , n513 , n503 );
not ( n948 , n947 );
or ( n949 , n946 , n948 );
nand ( n950 , n876 , n504 );
nand ( n951 , n949 , n950 );
not ( n952 , n951 );
nand ( n953 , n867 , n520 );
not ( n954 , n953 );
not ( n955 , n954 );
or ( n956 , n952 , n955 );
not ( n957 , n953 );
not ( n958 , n951 );
not ( n959 , n958 );
or ( n960 , n957 , n959 );
xor ( n961 , n519 , n497 );
not ( n962 , n961 );
buf ( n963 , n832 );
not ( n964 , n963 );
or ( n965 , n962 , n964 );
nand ( n966 , n836 , n886 );
nand ( n967 , n965 , n966 );
nand ( n968 , n960 , n967 );
nand ( n969 , n956 , n968 );
not ( n970 , n969 );
xor ( n971 , n516 , n499 );
not ( n972 , n971 );
xor ( n973 , n500 , n499 );
nand ( n974 , n934 , n973 );
not ( n975 , n974 );
not ( n976 , n975 );
or ( n977 , n972 , n976 );
xor ( n978 , n500 , n501 );
nand ( n979 , n978 , n927 );
nand ( n980 , n977 , n979 );
not ( n981 , n980 );
not ( n982 , n812 );
not ( n983 , n804 );
or ( n984 , n982 , n983 );
or ( n985 , n804 , n812 );
nand ( n986 , n984 , n985 );
nand ( n987 , n981 , n986 );
not ( n988 , n987 );
or ( n989 , n970 , n988 );
not ( n990 , n986 );
nand ( n991 , n990 , n980 );
nand ( n992 , n989 , n991 );
or ( n993 , n945 , n992 );
nand ( n994 , n945 , n992 );
nand ( n995 , n993 , n994 );
not ( n996 , n995 );
and ( n997 , n896 , n996 );
not ( n998 , n896 );
and ( n999 , n998 , n995 );
nor ( n1000 , n997 , n999 );
not ( n1001 , n969 );
not ( n1002 , n1001 );
and ( n1003 , n980 , n986 );
not ( n1004 , n980 );
and ( n1005 , n804 , n811 );
not ( n1006 , n804 );
and ( n1007 , n1006 , n812 );
or ( n1008 , n1005 , n1007 );
and ( n1009 , n1004 , n1008 );
nor ( n1010 , n1003 , n1009 );
not ( n1011 , n1010 );
not ( n1012 , n1011 );
or ( n1013 , n1002 , n1012 );
nand ( n1014 , n1010 , n969 );
nand ( n1015 , n1013 , n1014 );
xor ( n1016 , n515 , n501 );
not ( n1017 , n1016 );
not ( n1018 , n736 );
or ( n1019 , n1017 , n1018 );
nand ( n1020 , n694 , n799 );
nand ( n1021 , n1019 , n1020 );
not ( n1022 , n1021 );
xor ( n1023 , n517 , n499 );
not ( n1024 , n1023 );
not ( n1025 , n975 );
or ( n1026 , n1024 , n1025 );
xor ( n1027 , n500 , n501 );
nand ( n1028 , n1027 , n971 );
nand ( n1029 , n1026 , n1028 );
not ( n1030 , n1029 );
nand ( n1031 , n520 , n498 );
or ( n1032 , n520 , n498 );
nand ( n1033 , n1032 , n499 );
nand ( n1034 , n1031 , n1033 , n497 );
not ( n1035 , n1034 );
xor ( n1036 , n514 , n503 );
not ( n1037 , n1036 );
not ( n1038 , n683 );
or ( n1039 , n1037 , n1038 );
nand ( n1040 , n947 , n504 );
nand ( n1041 , n1039 , n1040 );
nand ( n1042 , n1035 , n1041 );
nand ( n1043 , n1030 , n1042 );
not ( n1044 , n1043 );
or ( n1045 , n1022 , n1044 );
not ( n1046 , n1042 );
nand ( n1047 , n1046 , n1029 );
nand ( n1048 , n1045 , n1047 );
buf ( n1049 , n1048 );
or ( n1050 , n1015 , n1049 );
not ( n1051 , n870 );
not ( n1052 , n882 );
xor ( n1053 , n1052 , n892 );
xnor ( n1054 , n1051 , n1053 );
not ( n1055 , n1054 );
nand ( n1056 , n1050 , n1055 );
nand ( n1057 , n1015 , n1049 );
nand ( n1058 , n1000 , n1056 , n1057 );
not ( n1059 , n1058 );
xor ( n1060 , n520 , n499 );
not ( n1061 , n1060 );
not ( n1062 , n974 );
not ( n1063 , n1062 );
or ( n1064 , n1061 , n1063 );
xor ( n1065 , n519 , n499 );
nand ( n1066 , n978 , n1065 );
nand ( n1067 , n1064 , n1066 );
not ( n1068 , n1067 );
not ( n1069 , n771 );
not ( n1070 , n683 );
or ( n1071 , n1069 , n1070 );
xor ( n1072 , n515 , n503 );
nand ( n1073 , n1072 , n504 );
nand ( n1074 , n1071 , n1073 );
or ( n1075 , n520 , n500 );
nand ( n1076 , n1075 , n501 );
nand ( n1077 , n520 , n500 );
nand ( n1078 , n1076 , n1077 , n499 );
and ( n1079 , n1074 , n1078 );
not ( n1080 , n1074 );
not ( n1081 , n1078 );
and ( n1082 , n1080 , n1081 );
nor ( n1083 , n1079 , n1082 );
not ( n1084 , n1083 );
or ( n1085 , n1068 , n1084 );
or ( n1086 , n1083 , n1067 );
nand ( n1087 , n1085 , n1086 );
xor ( n1088 , n517 , n501 );
and ( n1089 , n1088 , n694 );
not ( n1090 , n760 );
nand ( n1091 , n733 , n734 );
nor ( n1092 , n1090 , n1091 );
nor ( n1093 , n1089 , n1092 );
not ( n1094 , n1093 );
and ( n1095 , n1087 , n1094 );
not ( n1096 , n1087 );
and ( n1097 , n1096 , n1093 );
nor ( n1098 , n1095 , n1097 );
not ( n1099 , n750 );
nand ( n1100 , n1099 , n776 );
buf ( n1101 , n763 );
nand ( n1102 , n1100 , n1101 );
nand ( n1103 , n750 , n775 );
nand ( n1104 , n1102 , n1103 );
nand ( n1105 , n1098 , n1104 );
not ( n1106 , n1105 );
not ( n1107 , n785 );
not ( n1108 , n747 );
or ( n1109 , n1107 , n1108 );
not ( n1110 , n787 );
nand ( n1111 , n1109 , n1110 );
nor ( n1112 , n1106 , n1111 );
not ( n1113 , n1098 );
not ( n1114 , n1101 );
not ( n1115 , n1100 );
or ( n1116 , n1114 , n1115 );
nand ( n1117 , n1116 , n1103 );
not ( n1118 , n1117 );
nand ( n1119 , n1113 , n1118 );
nand ( n1120 , n1074 , n1081 );
not ( n1121 , n1120 );
not ( n1122 , n1121 );
not ( n1123 , n1065 );
not ( n1124 , n1062 );
or ( n1125 , n1123 , n1124 );
xor ( n1126 , n518 , n499 );
nand ( n1127 , n1027 , n1126 );
nand ( n1128 , n1125 , n1127 );
not ( n1129 , n1128 );
not ( n1130 , n1129 );
or ( n1131 , n1122 , n1130 );
nand ( n1132 , n1128 , n1120 );
nand ( n1133 , n1131 , n1132 );
not ( n1134 , n683 );
not ( n1135 , n1072 );
or ( n1136 , n1134 , n1135 );
nand ( n1137 , n1036 , n504 );
nand ( n1138 , n1136 , n1137 );
not ( n1139 , n1138 );
nand ( n1140 , n836 , n520 );
not ( n1141 , n1140 );
not ( n1142 , n1141 );
or ( n1143 , n1139 , n1142 );
not ( n1144 , n1138 );
nand ( n1145 , n1144 , n1140 );
nand ( n1146 , n1143 , n1145 );
not ( n1147 , n1088 );
not ( n1148 , n736 );
or ( n1149 , n1147 , n1148 );
xor ( n1150 , n516 , n501 );
nand ( n1151 , n694 , n1150 );
nand ( n1152 , n1149 , n1151 );
not ( n1153 , n1152 );
and ( n1154 , n1146 , n1153 );
not ( n1155 , n1146 );
and ( n1156 , n1155 , n1152 );
nor ( n1157 , n1154 , n1156 );
not ( n1158 , n1157 );
and ( n1159 , n1133 , n1158 );
not ( n1160 , n1133 );
and ( n1161 , n1160 , n1157 );
nor ( n1162 , n1159 , n1161 );
nand ( n1163 , n1067 , n1094 );
not ( n1164 , n1093 );
not ( n1165 , n1067 );
not ( n1166 , n1165 );
or ( n1167 , n1164 , n1166 );
not ( n1168 , n1083 );
nand ( n1169 , n1167 , n1168 );
nand ( n1170 , n1162 , n1163 , n1169 );
nand ( n1171 , n1119 , n1170 );
nor ( n1172 , n1112 , n1171 );
not ( n1173 , n1172 );
not ( n1174 , n1128 );
not ( n1175 , n1121 );
or ( n1176 , n1174 , n1175 );
nand ( n1177 , n1120 , n1129 );
nand ( n1178 , n1177 , n1157 );
nand ( n1179 , n1176 , n1178 );
not ( n1180 , n1179 );
not ( n1181 , n1140 );
not ( n1182 , n1144 );
or ( n1183 , n1181 , n1182 );
nand ( n1184 , n1183 , n1152 );
nand ( n1185 , n1138 , n1141 );
nand ( n1186 , n1184 , n1185 );
not ( n1187 , n1186 );
not ( n1188 , n1041 );
not ( n1189 , n1034 );
and ( n1190 , n1188 , n1189 );
and ( n1191 , n1041 , n1034 );
nor ( n1192 , n1190 , n1191 );
not ( n1193 , n1192 );
and ( n1194 , n1187 , n1193 );
and ( n1195 , n1186 , n1192 );
nor ( n1196 , n1194 , n1195 );
not ( n1197 , n1126 );
not ( n1198 , n939 );
or ( n1199 , n1197 , n1198 );
nand ( n1200 , n1023 , n749 );
nand ( n1201 , n1199 , n1200 );
not ( n1202 , n1201 );
not ( n1203 , n1150 );
not ( n1204 , n736 );
or ( n1205 , n1203 , n1204 );
nand ( n1206 , n694 , n1016 );
nand ( n1207 , n1205 , n1206 );
not ( n1208 , n1207 );
not ( n1209 , n1208 );
or ( n1210 , n1202 , n1209 );
not ( n1211 , n1201 );
nand ( n1212 , n1207 , n1211 );
nand ( n1213 , n1210 , n1212 );
xor ( n1214 , n520 , n497 );
not ( n1215 , n1214 );
not ( n1216 , n963 );
or ( n1217 , n1215 , n1216 );
nand ( n1218 , n836 , n961 );
nand ( n1219 , n1217 , n1218 );
and ( n1220 , n1213 , n1219 );
not ( n1221 , n1213 );
not ( n1222 , n1219 );
and ( n1223 , n1221 , n1222 );
nor ( n1224 , n1220 , n1223 );
not ( n1225 , n1224 );
and ( n1226 , n1196 , n1225 );
not ( n1227 , n1196 );
and ( n1228 , n1227 , n1224 );
nor ( n1229 , n1226 , n1228 );
not ( n1230 , n1229 );
nand ( n1231 , n1180 , n1230 );
not ( n1232 , n1231 );
or ( n1233 , n1173 , n1232 );
not ( n1234 , n1120 );
nand ( n1235 , n1234 , n1128 );
not ( n1236 , n1235 );
not ( n1237 , n1178 );
or ( n1238 , n1236 , n1237 );
nand ( n1239 , n1238 , n1229 );
not ( n1240 , n1239 );
not ( n1241 , n1162 );
nand ( n1242 , n1163 , n1169 );
nand ( n1243 , n1241 , n1242 );
not ( n1244 , n1243 );
or ( n1245 , n1240 , n1244 );
nand ( n1246 , n1245 , n1231 );
nand ( n1247 , n1233 , n1246 );
not ( n1248 , n1247 );
and ( n1249 , n951 , n953 );
not ( n1250 , n951 );
and ( n1251 , n867 , n520 );
and ( n1252 , n1250 , n1251 );
nor ( n1253 , n1249 , n1252 );
and ( n1254 , n1253 , n967 );
not ( n1255 , n1253 );
not ( n1256 , n967 );
and ( n1257 , n1255 , n1256 );
nor ( n1258 , n1254 , n1257 );
not ( n1259 , n1211 );
not ( n1260 , n1208 );
or ( n1261 , n1259 , n1260 );
nand ( n1262 , n1261 , n1219 );
nand ( n1263 , n1207 , n1201 );
nand ( n1264 , n1258 , n1262 , n1263 );
not ( n1265 , n1264 );
nand ( n1266 , n1047 , n1043 );
xnor ( n1267 , n1266 , n1021 );
not ( n1268 , n1267 );
or ( n1269 , n1265 , n1268 );
not ( n1270 , n1258 );
nand ( n1271 , n1262 , n1263 );
nand ( n1272 , n1270 , n1271 );
nand ( n1273 , n1269 , n1272 );
not ( n1274 , n1273 );
not ( n1275 , n1054 );
not ( n1276 , n1048 );
and ( n1277 , n1275 , n1276 );
and ( n1278 , n1048 , n1054 );
nor ( n1279 , n1277 , n1278 );
xor ( n1280 , n1015 , n1279 );
nand ( n1281 , n1274 , n1280 );
not ( n1282 , n1258 );
not ( n1283 , n1282 );
not ( n1284 , n1271 );
not ( n1285 , n1284 );
or ( n1286 , n1283 , n1285 );
nand ( n1287 , n1271 , n1258 );
nand ( n1288 , n1286 , n1287 );
not ( n1289 , n1267 );
and ( n1290 , n1288 , n1289 );
not ( n1291 , n1288 );
and ( n1292 , n1291 , n1267 );
nor ( n1293 , n1290 , n1292 );
not ( n1294 , n1225 );
not ( n1295 , n1186 );
nand ( n1296 , n1295 , n1192 );
and ( n1297 , n1294 , n1296 );
not ( n1298 , n1186 );
nor ( n1299 , n1298 , n1192 );
nor ( n1300 , n1297 , n1299 );
nand ( n1301 , n1293 , n1300 );
and ( n1302 , n1281 , n1301 );
not ( n1303 , n1302 );
or ( n1304 , n1248 , n1303 );
not ( n1305 , n1280 );
nand ( n1306 , n1305 , n1273 );
not ( n1307 , n1306 );
not ( n1308 , n1293 );
not ( n1309 , n1300 );
nand ( n1310 , n1308 , n1309 );
not ( n1311 , n1310 );
or ( n1312 , n1307 , n1311 );
buf ( n1313 , n1281 );
nand ( n1314 , n1312 , n1313 );
nand ( n1315 , n1304 , n1314 );
not ( n1316 , n1315 );
or ( n1317 , n1059 , n1316 );
nand ( n1318 , n1057 , n1056 );
not ( n1319 , n996 );
buf ( n1320 , n896 );
not ( n1321 , n1320 );
or ( n1322 , n1319 , n1321 );
or ( n1323 , n1320 , n996 );
nand ( n1324 , n1322 , n1323 );
nand ( n1325 , n1318 , n1324 );
nand ( n1326 , n1317 , n1325 );
not ( n1327 , n814 );
not ( n1328 , n1327 );
and ( n1329 , n520 , n1328 );
not ( n1330 , n1329 );
not ( n1331 , n838 );
or ( n1332 , n1330 , n1331 );
nand ( n1333 , n1328 , n520 );
not ( n1334 , n1333 );
not ( n1335 , n838 );
not ( n1336 , n1335 );
or ( n1337 , n1334 , n1336 );
nand ( n1338 , n1337 , n848 );
nand ( n1339 , n1332 , n1338 );
not ( n1340 , n1339 );
or ( n1341 , n921 , n902 );
nand ( n1342 , n1341 , n944 );
nand ( n1343 , n921 , n902 );
nand ( n1344 , n1342 , n1343 );
not ( n1345 , n1344 );
nand ( n1346 , n1340 , n1345 );
not ( n1347 , n1346 );
not ( n1348 , n898 );
not ( n1349 , n683 );
or ( n1350 , n1348 , n1349 );
xor ( n1351 , n503 , n509 );
nand ( n1352 , n504 , n1351 );
nand ( n1353 , n1350 , n1352 );
not ( n1354 , n919 );
and ( n1355 , n497 , n496 );
not ( n1356 , n497 );
not ( n1357 , n496 );
and ( n1358 , n1356 , n1357 );
nor ( n1359 , n1355 , n1358 );
not ( n1360 , n1359 );
nand ( n1361 , n1360 , n857 );
not ( n1362 , n1361 );
not ( n1363 , n1362 );
or ( n1364 , n1354 , n1363 );
xor ( n1365 , n495 , n517 );
nand ( n1366 , n1365 , n1359 );
nand ( n1367 , n1364 , n1366 );
xor ( n1368 , n1353 , n1367 );
not ( n1369 , n516 );
xnor ( n1370 , n1369 , n497 );
not ( n1371 , n1370 );
not ( n1372 , n963 );
or ( n1373 , n1371 , n1372 );
xor ( n1374 , n515 , n497 );
nand ( n1375 , n836 , n1374 );
nand ( n1376 , n1373 , n1375 );
xor ( n1377 , n1368 , n1376 );
not ( n1378 , n1377 );
or ( n1379 , n1347 , n1378 );
nand ( n1380 , n1339 , n1344 );
nand ( n1381 , n1379 , n1380 );
xor ( n1382 , n1353 , n1367 );
and ( n1383 , n1382 , n1376 );
and ( n1384 , n1353 , n1367 );
or ( n1385 , n1383 , n1384 );
not ( n1386 , n1385 );
not ( n1387 , n1091 );
not ( n1388 , n1387 );
not ( n1389 , n846 );
or ( n1390 , n1388 , n1389 );
xor ( n1391 , n511 , n501 );
nand ( n1392 , n694 , n1391 );
nand ( n1393 , n1390 , n1392 );
nand ( n1394 , n520 , n494 );
or ( n1395 , n520 , n494 );
nand ( n1396 , n1395 , n495 );
nand ( n1397 , n1394 , n493 , n1396 );
not ( n1398 , n1397 );
nand ( n1399 , n1393 , n1398 );
not ( n1400 , n1399 );
not ( n1401 , n1400 );
xor ( n1402 , n513 , n499 );
not ( n1403 , n1402 );
not ( n1404 , n1062 );
or ( n1405 , n1403 , n1404 );
not ( n1406 , n512 );
not ( n1407 , n499 );
not ( n1408 , n1407 );
or ( n1409 , n1406 , n1408 );
nand ( n1410 , n874 , n499 );
nand ( n1411 , n1409 , n1410 );
nand ( n1412 , n978 , n1411 );
nand ( n1413 , n1405 , n1412 );
not ( n1414 , n1413 );
not ( n1415 , n1414 );
and ( n1416 , n1401 , n1415 );
and ( n1417 , n1400 , n1414 );
nor ( n1418 , n1416 , n1417 );
not ( n1419 , n1418 );
or ( n1420 , n1386 , n1419 );
or ( n1421 , n1418 , n1385 );
nand ( n1422 , n1420 , n1421 );
not ( n1423 , n1422 );
and ( n1424 , n1381 , n1423 );
not ( n1425 , n1381 );
and ( n1426 , n1425 , n1422 );
nor ( n1427 , n1424 , n1426 );
not ( n1428 , n503 );
nor ( n1429 , n1428 , n504 );
not ( n1430 , n1429 );
not ( n1431 , n1351 );
or ( n1432 , n1430 , n1431 );
xor ( n1433 , n503 , n508 );
nand ( n1434 , n1433 , n504 );
nand ( n1435 , n1432 , n1434 );
not ( n1436 , n1365 );
not ( n1437 , n912 );
or ( n1438 , n1436 , n1437 );
not ( n1439 , n1360 );
xor ( n1440 , n495 , n516 );
nand ( n1441 , n1439 , n1440 );
nand ( n1442 , n1438 , n1441 );
xor ( n1443 , n1435 , n1442 );
xor ( n1444 , n519 , n493 );
not ( n1445 , n1444 );
xor ( n1446 , n494 , n495 );
xor ( n1447 , n493 , n494 );
not ( n1448 , n1447 );
nor ( n1449 , n1446 , n1448 );
not ( n1450 , n1449 );
or ( n1451 , n1445 , n1450 );
xor ( n1452 , n518 , n493 );
nand ( n1453 , n814 , n1452 );
nand ( n1454 , n1451 , n1453 );
xor ( n1455 , n1443 , n1454 );
xor ( n1456 , n492 , n493 );
and ( n1457 , n1456 , n520 );
not ( n1458 , n1391 );
not ( n1459 , n736 );
or ( n1460 , n1458 , n1459 );
xor ( n1461 , n510 , n501 );
nand ( n1462 , n694 , n1461 );
nand ( n1463 , n1460 , n1462 );
xor ( n1464 , n1457 , n1463 );
not ( n1465 , n1374 );
not ( n1466 , n832 );
or ( n1467 , n1465 , n1466 );
xor ( n1468 , n514 , n497 );
nand ( n1469 , n836 , n1468 );
nand ( n1470 , n1467 , n1469 );
xor ( n1471 , n1464 , n1470 );
xor ( n1472 , n1455 , n1471 );
not ( n1473 , n942 );
not ( n1474 , n939 );
or ( n1475 , n1473 , n1474 );
nand ( n1476 , n749 , n1402 );
nand ( n1477 , n1475 , n1476 );
xor ( n1478 , n520 , n493 );
not ( n1479 , n1478 );
not ( n1480 , n1446 );
and ( n1481 , n1480 , n1447 );
not ( n1482 , n1481 );
or ( n1483 , n1479 , n1482 );
nand ( n1484 , n814 , n1444 );
nand ( n1485 , n1483 , n1484 );
or ( n1486 , n1477 , n1485 );
not ( n1487 , n1486 );
and ( n1488 , n1393 , n1397 );
not ( n1489 , n1393 );
and ( n1490 , n1489 , n1398 );
or ( n1491 , n1488 , n1490 );
not ( n1492 , n1491 );
or ( n1493 , n1487 , n1492 );
nand ( n1494 , n1477 , n1485 );
nand ( n1495 , n1493 , n1494 );
not ( n1496 , n1495 );
xor ( n1497 , n1472 , n1496 );
not ( n1498 , n1497 );
and ( n1499 , n1427 , n1498 );
not ( n1500 , n1427 );
and ( n1501 , n1500 , n1497 );
nor ( n1502 , n1499 , n1501 );
xor ( n1503 , n813 , n849 );
and ( n1504 , n1503 , n895 );
and ( n1505 , n813 , n849 );
or ( n1506 , n1504 , n1505 );
not ( n1507 , n1506 );
xor ( n1508 , n1477 , n1485 );
not ( n1509 , n1491 );
xor ( n1510 , n1508 , n1509 );
and ( n1511 , n1339 , n1345 );
not ( n1512 , n1339 );
and ( n1513 , n1512 , n1344 );
nor ( n1514 , n1511 , n1513 );
and ( n1515 , n1514 , n1377 );
not ( n1516 , n1514 );
not ( n1517 , n1377 );
and ( n1518 , n1516 , n1517 );
nor ( n1519 , n1515 , n1518 );
nand ( n1520 , n1510 , n1519 );
not ( n1521 , n1520 );
or ( n1522 , n1507 , n1521 );
not ( n1523 , n1519 );
not ( n1524 , n1510 );
nand ( n1525 , n1523 , n1524 );
nand ( n1526 , n1522 , n1525 );
not ( n1527 , n1526 );
nand ( n1528 , n1502 , n1527 );
not ( n1529 , n992 );
nand ( n1530 , n1529 , n945 );
not ( n1531 , n1530 );
not ( n1532 , n896 );
or ( n1533 , n1531 , n1532 );
not ( n1534 , n945 );
nand ( n1535 , n1534 , n992 );
nand ( n1536 , n1533 , n1535 );
not ( n1537 , n1536 );
and ( n1538 , n1519 , n1524 );
not ( n1539 , n1519 );
and ( n1540 , n1539 , n1510 );
nor ( n1541 , n1538 , n1540 );
xor ( n1542 , n1506 , n1541 );
nand ( n1543 , n1537 , n1542 );
and ( n1544 , n1528 , n1543 );
not ( n1545 , n1498 );
xnor ( n1546 , n1385 , n1418 );
not ( n1547 , n1546 );
or ( n1548 , n1545 , n1547 );
not ( n1549 , n1423 );
not ( n1550 , n1497 );
or ( n1551 , n1549 , n1550 );
nand ( n1552 , n1551 , n1381 );
nand ( n1553 , n1548 , n1552 );
not ( n1554 , n1553 );
not ( n1555 , n1385 );
nand ( n1556 , n1414 , n1399 );
not ( n1557 , n1556 );
or ( n1558 , n1555 , n1557 );
not ( n1559 , n1414 );
nand ( n1560 , n1559 , n1400 );
nand ( n1561 , n1558 , n1560 );
xor ( n1562 , n520 , n491 );
not ( n1563 , n1562 );
xnor ( n1564 , n491 , n492 );
xor ( n1565 , n492 , n493 );
nor ( n1566 , n1564 , n1565 );
not ( n1567 , n1566 );
or ( n1568 , n1563 , n1567 );
xor ( n1569 , n491 , n519 );
nand ( n1570 , n1456 , n1569 );
nand ( n1571 , n1568 , n1570 );
not ( n1572 , n1411 );
not ( n1573 , n975 );
or ( n1574 , n1572 , n1573 );
not ( n1575 , n511 );
not ( n1576 , n499 );
not ( n1577 , n1576 );
or ( n1578 , n1575 , n1577 );
not ( n1579 , n511 );
nand ( n1580 , n1579 , n499 );
nand ( n1581 , n1578 , n1580 );
nand ( n1582 , n1027 , n1581 );
nand ( n1583 , n1574 , n1582 );
xor ( n1584 , n1571 , n1583 );
not ( n1585 , n1452 );
and ( n1586 , n1480 , n1447 );
not ( n1587 , n1586 );
or ( n1588 , n1585 , n1587 );
xor ( n1589 , n517 , n493 );
nand ( n1590 , n814 , n1589 );
nand ( n1591 , n1588 , n1590 );
xor ( n1592 , n1584 , n1591 );
not ( n1593 , n1461 );
not ( n1594 , n1387 );
or ( n1595 , n1593 , n1594 );
and ( n1596 , n509 , n755 );
not ( n1597 , n509 );
and ( n1598 , n1597 , n501 );
or ( n1599 , n1596 , n1598 );
nand ( n1600 , n694 , n1599 );
nand ( n1601 , n1595 , n1600 );
not ( n1602 , n1468 );
not ( n1603 , n888 );
or ( n1604 , n1602 , n1603 );
and ( n1605 , n513 , n497 );
not ( n1606 , n513 );
and ( n1607 , n1606 , n818 );
nor ( n1608 , n1605 , n1607 );
nand ( n1609 , n836 , n1608 );
nand ( n1610 , n1604 , n1609 );
xor ( n1611 , n1601 , n1610 );
not ( n1612 , n1440 );
not ( n1613 , n1362 );
or ( n1614 , n1612 , n1613 );
not ( n1615 , n1360 );
xor ( n1616 , n515 , n495 );
nand ( n1617 , n1615 , n1616 );
nand ( n1618 , n1614 , n1617 );
not ( n1619 , n1618 );
and ( n1620 , n1611 , n1619 );
not ( n1621 , n1611 );
and ( n1622 , n1621 , n1618 );
nor ( n1623 , n1620 , n1622 );
xor ( n1624 , n1592 , n1623 );
xor ( n1625 , n1561 , n1624 );
not ( n1626 , n1625 );
nand ( n1627 , n520 , n492 );
or ( n1628 , n520 , n492 );
nand ( n1629 , n1628 , n493 );
and ( n1630 , n1627 , n1629 , n491 );
not ( n1631 , n1630 );
not ( n1632 , n1429 );
not ( n1633 , n1433 );
or ( n1634 , n1632 , n1633 );
xor ( n1635 , n503 , n507 );
nand ( n1636 , n1635 , n504 );
nand ( n1637 , n1634 , n1636 );
not ( n1638 , n1637 );
or ( n1639 , n1631 , n1638 );
or ( n1640 , n1630 , n1637 );
nand ( n1641 , n1639 , n1640 );
not ( n1642 , n1435 );
not ( n1643 , n1442 );
or ( n1644 , n1642 , n1643 );
not ( n1645 , n1365 );
not ( n1646 , n912 );
or ( n1647 , n1645 , n1646 );
nand ( n1648 , n1647 , n1441 );
or ( n1649 , n1435 , n1648 );
nand ( n1650 , n1649 , n1454 );
nand ( n1651 , n1644 , n1650 );
xor ( n1652 , n1641 , n1651 );
xor ( n1653 , n1457 , n1463 );
and ( n1654 , n1653 , n1470 );
and ( n1655 , n1457 , n1463 );
or ( n1656 , n1654 , n1655 );
xor ( n1657 , n1652 , n1656 );
not ( n1658 , n1657 );
not ( n1659 , n1658 );
not ( n1660 , n1455 );
not ( n1661 , n1660 );
not ( n1662 , n1661 );
not ( n1663 , n1471 );
or ( n1664 , n1662 , n1663 );
not ( n1665 , n1660 );
not ( n1666 , n1471 );
not ( n1667 , n1666 );
or ( n1668 , n1665 , n1667 );
nand ( n1669 , n1668 , n1495 );
nand ( n1670 , n1664 , n1669 );
not ( n1671 , n1670 );
not ( n1672 , n1671 );
or ( n1673 , n1659 , n1672 );
nand ( n1674 , n1657 , n1670 );
nand ( n1675 , n1673 , n1674 );
not ( n1676 , n1675 );
not ( n1677 , n1676 );
or ( n1678 , n1626 , n1677 );
not ( n1679 , n1625 );
nand ( n1680 , n1675 , n1679 );
nand ( n1681 , n1678 , n1680 );
nand ( n1682 , n1554 , n1681 );
not ( n1683 , n1581 );
xor ( n1684 , n500 , n499 );
and ( n1685 , n1684 , n934 );
not ( n1686 , n1685 );
or ( n1687 , n1683 , n1686 );
not ( n1688 , n1027 );
not ( n1689 , n1688 );
and ( n1690 , n510 , n499 );
not ( n1691 , n510 );
not ( n1692 , n499 );
and ( n1693 , n1691 , n1692 );
nor ( n1694 , n1690 , n1693 );
nand ( n1695 , n1689 , n1694 );
nand ( n1696 , n1687 , n1695 );
not ( n1697 , n1608 );
not ( n1698 , n888 );
or ( n1699 , n1697 , n1698 );
xor ( n1700 , n512 , n497 );
nand ( n1701 , n836 , n1700 );
nand ( n1702 , n1699 , n1701 );
xor ( n1703 , n1696 , n1702 );
not ( n1704 , n1616 );
not ( n1705 , n912 );
or ( n1706 , n1704 , n1705 );
xor ( n1707 , n514 , n495 );
nand ( n1708 , n867 , n1707 );
nand ( n1709 , n1706 , n1708 );
xor ( n1710 , n1703 , n1709 );
not ( n1711 , n1569 );
not ( n1712 , n1566 );
or ( n1713 , n1711 , n1712 );
xor ( n1714 , n491 , n518 );
nand ( n1715 , n1456 , n1714 );
nand ( n1716 , n1713 , n1715 );
not ( n1717 , n1716 );
nand ( n1718 , n1637 , n1630 );
xor ( n1719 , n1717 , n1718 );
not ( n1720 , n1480 );
nand ( n1721 , n1589 , n1447 );
not ( n1722 , n1721 );
or ( n1723 , n1720 , n1722 );
xnor ( n1724 , n516 , n493 );
nand ( n1725 , n1724 , n1446 );
nand ( n1726 , n1723 , n1725 );
xor ( n1727 , n1719 , n1726 );
and ( n1728 , n1710 , n1727 );
not ( n1729 , n1710 );
not ( n1730 , n1727 );
and ( n1731 , n1729 , n1730 );
nor ( n1732 , n1728 , n1731 );
not ( n1733 , n1651 );
nand ( n1734 , n1733 , n1641 );
not ( n1735 , n1734 );
not ( n1736 , n1656 );
or ( n1737 , n1735 , n1736 );
not ( n1738 , n1641 );
nand ( n1739 , n1738 , n1651 );
nand ( n1740 , n1737 , n1739 );
xor ( n1741 , n1732 , n1740 );
not ( n1742 , n1583 );
not ( n1743 , n1591 );
or ( n1744 , n1742 , n1743 );
not ( n1745 , n1411 );
not ( n1746 , n975 );
or ( n1747 , n1745 , n1746 );
nand ( n1748 , n749 , n1581 );
nand ( n1749 , n1747 , n1748 );
or ( n1750 , n1591 , n1749 );
nand ( n1751 , n1750 , n1571 );
nand ( n1752 , n1744 , n1751 );
not ( n1753 , n1618 );
not ( n1754 , n1601 );
or ( n1755 , n1753 , n1754 );
or ( n1756 , n1601 , n1618 );
nand ( n1757 , n1756 , n1610 );
nand ( n1758 , n1755 , n1757 );
xor ( n1759 , n1752 , n1758 );
xor ( n1760 , n490 , n491 );
and ( n1761 , n1760 , n520 );
not ( n1762 , n1761 );
not ( n1763 , n1762 );
not ( n1764 , n1635 );
not ( n1765 , n683 );
or ( n1766 , n1764 , n1765 );
and ( n1767 , n503 , n506 );
not ( n1768 , n503 );
not ( n1769 , n506 );
and ( n1770 , n1768 , n1769 );
nor ( n1771 , n1767 , n1770 );
nand ( n1772 , n1771 , n504 );
nand ( n1773 , n1766 , n1772 );
not ( n1774 , n1773 );
or ( n1775 , n1763 , n1774 );
not ( n1776 , n1773 );
nand ( n1777 , n1776 , n1761 );
nand ( n1778 , n1775 , n1777 );
xor ( n1779 , n508 , n501 );
nand ( n1780 , n1779 , n694 );
nand ( n1781 , n736 , n1599 );
nand ( n1782 , n1780 , n1781 );
xor ( n1783 , n1778 , n1782 );
xor ( n1784 , n1759 , n1783 );
or ( n1785 , n1741 , n1784 );
nand ( n1786 , n1741 , n1784 );
nand ( n1787 , n1785 , n1786 );
buf ( n1788 , n1623 );
not ( n1789 , n1592 );
nand ( n1790 , n1788 , n1789 );
not ( n1791 , n1790 );
not ( n1792 , n1561 );
or ( n1793 , n1791 , n1792 );
or ( n1794 , n1788 , n1789 );
nand ( n1795 , n1793 , n1794 );
not ( n1796 , n1795 );
and ( n1797 , n1787 , n1796 );
not ( n1798 , n1787 );
and ( n1799 , n1798 , n1795 );
nor ( n1800 , n1797 , n1799 );
not ( n1801 , n1679 );
not ( n1802 , n1658 );
or ( n1803 , n1801 , n1802 );
not ( n1804 , n1657 );
not ( n1805 , n1625 );
or ( n1806 , n1804 , n1805 );
nand ( n1807 , n1806 , n1670 );
nand ( n1808 , n1803 , n1807 );
not ( n1809 , n1808 );
nand ( n1810 , n1800 , n1809 );
nand ( n1811 , n1326 , n1544 , n1682 , n1810 );
not ( n1812 , n1528 );
nor ( n1813 , n1537 , n1542 );
not ( n1814 , n1813 );
or ( n1815 , n1812 , n1814 );
not ( n1816 , n1502 );
nand ( n1817 , n1816 , n1526 );
nand ( n1818 , n1815 , n1817 );
nand ( n1819 , n1818 , n1682 , n1810 );
not ( n1820 , n1809 );
not ( n1821 , n1800 );
or ( n1822 , n1820 , n1821 );
not ( n1823 , n1553 );
nor ( n1824 , n1681 , n1823 );
nand ( n1825 , n1822 , n1824 );
not ( n1826 , n1800 );
nand ( n1827 , n1826 , n1808 );
nand ( n1828 , n1811 , n1819 , n1825 , n1827 );
xor ( n1829 , n1696 , n1702 );
and ( n1830 , n1829 , n1709 );
and ( n1831 , n1696 , n1702 );
or ( n1832 , n1830 , n1831 );
not ( n1833 , n1700 );
not ( n1834 , n832 );
or ( n1835 , n1833 , n1834 );
xor ( n1836 , n511 , n497 );
nand ( n1837 , n836 , n1836 );
nand ( n1838 , n1835 , n1837 );
not ( n1839 , n1838 );
not ( n1840 , n1779 );
not ( n1841 , n1387 );
or ( n1842 , n1840 , n1841 );
and ( n1843 , n507 , n501 );
not ( n1844 , n507 );
not ( n1845 , n501 );
and ( n1846 , n1844 , n1845 );
nor ( n1847 , n1843 , n1846 );
nand ( n1848 , n694 , n1847 );
nand ( n1849 , n1842 , n1848 );
not ( n1850 , n1849 );
not ( n1851 , n1850 );
or ( n1852 , n1839 , n1851 );
not ( n1853 , n1838 );
nand ( n1854 , n1849 , n1853 );
nand ( n1855 , n1852 , n1854 );
xor ( n1856 , n489 , n490 );
xor ( n1857 , n520 , n489 );
nand ( n1858 , n1856 , n1857 );
buf ( n1859 , n1760 );
or ( n1860 , n1858 , n1859 );
xor ( n1861 , n519 , n489 );
nand ( n1862 , n1859 , n1861 );
nand ( n1863 , n1860 , n1862 );
not ( n1864 , n1863 );
not ( n1865 , n1864 );
and ( n1866 , n1855 , n1865 );
not ( n1867 , n1855 );
and ( n1868 , n1867 , n1864 );
nor ( n1869 , n1866 , n1868 );
xor ( n1870 , n1832 , n1869 );
and ( n1871 , n493 , n1369 );
not ( n1872 , n493 );
and ( n1873 , n1872 , n516 );
nor ( n1874 , n1871 , n1873 );
nor ( n1875 , n1448 , n1874 );
not ( n1876 , n1875 );
not ( n1877 , n1480 );
or ( n1878 , n1876 , n1877 );
xor ( n1879 , n515 , n493 );
nand ( n1880 , n814 , n1879 );
nand ( n1881 , n1878 , n1880 );
not ( n1882 , n1707 );
not ( n1883 , n1362 );
or ( n1884 , n1882 , n1883 );
xor ( n1885 , n513 , n495 );
and ( n1886 , n496 , n497 );
not ( n1887 , n496 );
and ( n1888 , n1887 , n853 );
nor ( n1889 , n1886 , n1888 );
nand ( n1890 , n1885 , n1889 );
nand ( n1891 , n1884 , n1890 );
xor ( n1892 , n1881 , n1891 );
not ( n1893 , n1694 );
not ( n1894 , n1062 );
or ( n1895 , n1893 , n1894 );
and ( n1896 , n509 , n499 );
not ( n1897 , n509 );
and ( n1898 , n1897 , n1692 );
nor ( n1899 , n1896 , n1898 );
nand ( n1900 , n978 , n1899 );
nand ( n1901 , n1895 , n1900 );
xor ( n1902 , n1892 , n1901 );
xor ( n1903 , n1870 , n1902 );
not ( n1904 , n1656 );
not ( n1905 , n1734 );
or ( n1906 , n1904 , n1905 );
nand ( n1907 , n1906 , n1739 );
or ( n1908 , n1730 , n1907 );
buf ( n1909 , n1710 );
nand ( n1910 , n1908 , n1909 );
nand ( n1911 , n1907 , n1730 );
nand ( n1912 , n1910 , n1911 );
not ( n1913 , n1912 );
and ( n1914 , n1903 , n1913 );
not ( n1915 , n1903 );
and ( n1916 , n1915 , n1912 );
nor ( n1917 , n1914 , n1916 );
xor ( n1918 , n1717 , n1718 );
and ( n1919 , n1918 , n1726 );
and ( n1920 , n1717 , n1718 );
or ( n1921 , n1919 , n1920 );
nand ( n1922 , n1776 , n1762 );
not ( n1923 , n1922 );
not ( n1924 , n1782 );
or ( n1925 , n1923 , n1924 );
nand ( n1926 , n1761 , n1773 );
nand ( n1927 , n1925 , n1926 );
not ( n1928 , n1714 );
xnor ( n1929 , n491 , n492 );
nor ( n1930 , n1929 , n1565 );
not ( n1931 , n1930 );
or ( n1932 , n1928 , n1931 );
buf ( n1933 , n1456 );
xor ( n1934 , n517 , n491 );
nand ( n1935 , n1933 , n1934 );
nand ( n1936 , n1932 , n1935 );
not ( n1937 , n1936 );
not ( n1938 , n1771 );
not ( n1939 , n504 );
and ( n1940 , n1939 , n503 );
not ( n1941 , n1940 );
or ( n1942 , n1938 , n1941 );
xor ( n1943 , n503 , n505 );
nand ( n1944 , n1943 , n504 );
nand ( n1945 , n1942 , n1944 );
or ( n1946 , n520 , n490 );
nand ( n1947 , n1946 , n491 );
and ( n1948 , n520 , n490 );
not ( n1949 , n489 );
nor ( n1950 , n1948 , n1949 );
and ( n1951 , n1947 , n1950 );
nor ( n1952 , n1945 , n1951 );
not ( n1953 , n1952 );
nand ( n1954 , n1951 , n1945 );
nand ( n1955 , n1953 , n1954 );
or ( n1956 , n1937 , n1955 );
nand ( n1957 , n1955 , n1937 );
nand ( n1958 , n1956 , n1957 );
xor ( n1959 , n1927 , n1958 );
xor ( n1960 , n1921 , n1959 );
xor ( n1961 , n1752 , n1758 );
and ( n1962 , n1961 , n1783 );
and ( n1963 , n1752 , n1758 );
or ( n1964 , n1962 , n1963 );
xnor ( n1965 , n1960 , n1964 );
and ( n1966 , n1917 , n1965 );
not ( n1967 , n1917 );
not ( n1968 , n1965 );
and ( n1969 , n1967 , n1968 );
nor ( n1970 , n1966 , n1969 );
not ( n1971 , n1784 );
not ( n1972 , n1795 );
or ( n1973 , n1971 , n1972 );
or ( n1974 , n1795 , n1784 );
not ( n1975 , n1741 );
nand ( n1976 , n1974 , n1975 );
nand ( n1977 , n1973 , n1976 );
nand ( n1978 , n1970 , n1977 );
buf ( n1979 , n1978 );
not ( n1980 , n1977 );
not ( n1981 , n1970 );
nand ( n1982 , n1980 , n1981 );
nand ( n1983 , n1979 , n1982 );
xnor ( n1984 , n1828 , n1983 );
nand ( n1985 , n1984 , n793 );
and ( n1986 , n492 , n493 );
not ( n1987 , n492 );
not ( n1988 , n493 );
and ( n1989 , n1987 , n1988 );
nor ( n1990 , n1986 , n1989 );
not ( n1991 , n1990 );
not ( n1992 , n492 );
not ( n1993 , n491 );
not ( n1994 , n1993 );
or ( n1995 , n1992 , n1994 );
not ( n1996 , n492 );
nand ( n1997 , n1996 , n491 );
nand ( n1998 , n1995 , n1997 );
nand ( n1999 , n1991 , n1998 );
not ( n2000 , n1999 );
not ( n2001 , n2000 );
not ( n2002 , n491 );
and ( n2003 , n456 , n464 );
not ( n2004 , n456 );
and ( n2005 , n2004 , n480 );
nor ( n2006 , n2003 , n2005 );
not ( n2007 , n2006 );
or ( n2008 , n2002 , n2007 );
not ( n2009 , n464 );
and ( n2010 , n456 , n2009 );
not ( n2011 , n456 );
not ( n2012 , n480 );
and ( n2013 , n2011 , n2012 );
nor ( n2014 , n2010 , n2013 );
not ( n2015 , n491 );
nand ( n2016 , n2014 , n2015 );
nand ( n2017 , n2008 , n2016 );
not ( n2018 , n2017 );
or ( n2019 , n2001 , n2018 );
not ( n2020 , n2015 );
not ( n2021 , n479 );
not ( n2022 , n456 );
not ( n2023 , n2022 );
or ( n2024 , n2021 , n2023 );
nand ( n2025 , n456 , n463 );
nand ( n2026 , n2024 , n2025 );
not ( n2027 , n2026 );
or ( n2028 , n2020 , n2027 );
and ( n2029 , n456 , n463 );
not ( n2030 , n456 );
and ( n2031 , n2030 , n479 );
nor ( n2032 , n2029 , n2031 );
nand ( n2033 , n2032 , n491 );
nand ( n2034 , n2028 , n2033 );
not ( n2035 , n1990 );
not ( n2036 , n2035 );
nand ( n2037 , n2034 , n2036 );
nand ( n2038 , n2019 , n2037 );
not ( n2039 , n495 );
and ( n2040 , n456 , n460 );
not ( n2041 , n456 );
and ( n2042 , n2041 , n476 );
nor ( n2043 , n2040 , n2042 );
not ( n2044 , n2043 );
or ( n2045 , n2039 , n2044 );
not ( n2046 , n495 );
and ( n2047 , n456 , n460 );
not ( n2048 , n456 );
and ( n2049 , n2048 , n476 );
nor ( n2050 , n2047 , n2049 );
not ( n2051 , n2050 );
nand ( n2052 , n2046 , n2051 );
nand ( n2053 , n2045 , n2052 );
not ( n2054 , n2053 );
not ( n2055 , n495 );
nand ( n2056 , n2055 , n497 , n496 );
not ( n2057 , n497 );
nand ( n2058 , n907 , n2057 , n495 );
nand ( n2059 , n2056 , n2058 );
buf ( n2060 , n2059 );
not ( n2061 , n2060 );
or ( n2062 , n2054 , n2061 );
and ( n2063 , n456 , n459 );
not ( n2064 , n456 );
and ( n2065 , n2064 , n475 );
nor ( n2066 , n2063 , n2065 );
buf ( n2067 , n2066 );
and ( n2068 , n495 , n2067 );
not ( n2069 , n495 );
not ( n2070 , n459 );
and ( n2071 , n456 , n2070 );
not ( n2072 , n456 );
not ( n2073 , n475 );
and ( n2074 , n2072 , n2073 );
nor ( n2075 , n2071 , n2074 );
and ( n2076 , n2069 , n2075 );
or ( n2077 , n2068 , n2076 );
xor ( n2078 , n497 , n496 );
nand ( n2079 , n2077 , n2078 );
nand ( n2080 , n2062 , n2079 );
xor ( n2081 , n2038 , n2080 );
xor ( n2082 , n491 , n490 );
not ( n2083 , n2082 );
not ( n2084 , n2083 );
not ( n2085 , n2084 );
and ( n2086 , n456 , n465 );
not ( n2087 , n456 );
and ( n2088 , n2087 , n481 );
nor ( n2089 , n2086 , n2088 );
not ( n2090 , n2089 );
not ( n2091 , n2090 );
not ( n2092 , n1949 );
or ( n2093 , n2091 , n2092 );
not ( n2094 , n465 );
nand ( n2095 , n2094 , n456 );
not ( n2096 , n2095 );
or ( n2097 , n456 , n481 );
not ( n2098 , n2097 );
or ( n2099 , n2096 , n2098 );
nand ( n2100 , n2099 , n489 );
nand ( n2101 , n2093 , n2100 );
not ( n2102 , n2101 );
or ( n2103 , n2085 , n2102 );
not ( n2104 , n1949 );
and ( n2105 , n456 , n466 );
not ( n2106 , n456 );
and ( n2107 , n2106 , n482 );
nor ( n2108 , n2105 , n2107 );
not ( n2109 , n2108 );
not ( n2110 , n2109 );
or ( n2111 , n2104 , n2110 );
or ( n2112 , n2109 , n1949 );
nand ( n2113 , n2111 , n2112 );
not ( n2114 , n489 );
nor ( n2115 , n490 , n491 );
not ( n2116 , n2115 );
or ( n2117 , n2114 , n2116 );
not ( n2118 , n489 );
nand ( n2119 , n2118 , n491 , n490 );
nand ( n2120 , n2117 , n2119 );
not ( n2121 , n2120 );
not ( n2122 , n2121 );
nand ( n2123 , n2113 , n2122 );
nand ( n2124 , n2103 , n2123 );
and ( n2125 , n2081 , n2124 );
and ( n2126 , n2038 , n2080 );
or ( n2127 , n2125 , n2126 );
xor ( n2128 , n500 , n501 );
not ( n2129 , n499 );
nor ( n2130 , n500 , n501 );
not ( n2131 , n2130 );
or ( n2132 , n2129 , n2131 );
nand ( n2133 , n1576 , n501 , n500 );
nand ( n2134 , n2132 , n2133 );
or ( n2135 , n2128 , n2134 );
nand ( n2136 , n2135 , n499 );
not ( n2137 , n498 );
not ( n2138 , n1407 );
or ( n2139 , n2137 , n2138 );
nand ( n2140 , n825 , n499 );
nand ( n2141 , n2139 , n2140 );
buf ( n2142 , n2141 );
not ( n2143 , n2142 );
and ( n2144 , n456 , n457 );
not ( n2145 , n456 );
and ( n2146 , n2145 , n473 );
nor ( n2147 , n2144 , n2146 );
not ( n2148 , n2147 );
not ( n2149 , n2148 );
and ( n2150 , n497 , n2149 );
not ( n2151 , n497 );
not ( n2152 , n2149 );
and ( n2153 , n2151 , n2152 );
or ( n2154 , n2150 , n2153 );
not ( n2155 , n2154 );
or ( n2156 , n2143 , n2155 );
not ( n2157 , n498 );
not ( n2158 , n499 );
nand ( n2159 , n2157 , n2158 , n497 );
not ( n2160 , n497 );
nand ( n2161 , n2160 , n498 , n499 );
nand ( n2162 , n2159 , n2161 );
buf ( n2163 , n2162 );
buf ( n2164 , n2163 );
and ( n2165 , n456 , n458 );
not ( n2166 , n456 );
and ( n2167 , n2166 , n474 );
nor ( n2168 , n2165 , n2167 );
and ( n2169 , n497 , n2168 );
not ( n2170 , n497 );
and ( n2171 , n456 , n458 );
not ( n2172 , n456 );
and ( n2173 , n2172 , n474 );
nor ( n2174 , n2171 , n2173 );
not ( n2175 , n2174 );
and ( n2176 , n2170 , n2175 );
or ( n2177 , n2169 , n2176 );
nand ( n2178 , n2164 , n2177 );
nand ( n2179 , n2156 , n2178 );
xor ( n2180 , n2136 , n2179 );
and ( n2181 , n917 , n494 );
not ( n2182 , n494 );
and ( n2183 , n2182 , n495 );
nor ( n2184 , n2181 , n2183 );
not ( n2185 , n2184 );
not ( n2186 , n2185 );
and ( n2187 , n456 , n461 );
not ( n2188 , n456 );
and ( n2189 , n2188 , n477 );
nor ( n2190 , n2187 , n2189 );
and ( n2191 , n493 , n2190 );
not ( n2192 , n493 );
not ( n2193 , n2190 );
and ( n2194 , n2192 , n2193 );
or ( n2195 , n2191 , n2194 );
not ( n2196 , n2195 );
or ( n2197 , n2186 , n2196 );
nor ( n2198 , n494 , n495 );
nand ( n2199 , n2198 , n493 );
not ( n2200 , n493 );
nand ( n2201 , n2200 , n495 , n494 );
nand ( n2202 , n2199 , n2201 );
buf ( n2203 , n2202 );
not ( n2204 , n493 );
and ( n2205 , n456 , n462 );
not ( n2206 , n456 );
and ( n2207 , n2206 , n478 );
nor ( n2208 , n2205 , n2207 );
not ( n2209 , n2208 );
or ( n2210 , n2204 , n2209 );
or ( n2211 , n2208 , n493 );
nand ( n2212 , n2210 , n2211 );
nand ( n2213 , n2203 , n2212 );
nand ( n2214 , n2197 , n2213 );
and ( n2215 , n2180 , n2214 );
and ( n2216 , n2136 , n2179 );
or ( n2217 , n2215 , n2216 );
xor ( n2218 , n2127 , n2217 );
xor ( n2219 , n493 , n492 );
not ( n2220 , n2219 );
not ( n2221 , n491 );
not ( n2222 , n2208 );
or ( n2223 , n2221 , n2222 );
not ( n2224 , n462 );
and ( n2225 , n2224 , n456 );
nor ( n2226 , n456 , n478 );
nor ( n2227 , n2225 , n2226 );
nand ( n2228 , n2227 , n2015 );
nand ( n2229 , n2223 , n2228 );
not ( n2230 , n2229 );
or ( n2231 , n2220 , n2230 );
and ( n2232 , n2035 , n1998 );
nand ( n2233 , n2034 , n2232 );
nand ( n2234 , n2231 , n2233 );
not ( n2235 , n2101 );
not ( n2236 , n2122 );
or ( n2237 , n2235 , n2236 );
not ( n2238 , n489 );
not ( n2239 , n2006 );
or ( n2240 , n2238 , n2239 );
nand ( n2241 , n2014 , n1949 );
nand ( n2242 , n2240 , n2241 );
buf ( n2243 , n2082 );
nand ( n2244 , n2242 , n2243 );
nand ( n2245 , n2237 , n2244 );
xor ( n2246 , n2234 , n2245 );
not ( n2247 , n2164 );
not ( n2248 , n2154 );
or ( n2249 , n2247 , n2248 );
buf ( n2250 , n2142 );
nand ( n2251 , n2250 , n497 );
nand ( n2252 , n2249 , n2251 );
xor ( n2253 , n2246 , n2252 );
xor ( n2254 , n2218 , n2253 );
and ( n2255 , n456 , n466 );
not ( n2256 , n456 );
and ( n2257 , n2256 , n482 );
nor ( n2258 , n2255 , n2257 );
not ( n2259 , n2258 );
and ( n2260 , n2259 , n489 );
not ( n2261 , n2203 );
not ( n2262 , n2195 );
or ( n2263 , n2261 , n2262 );
not ( n2264 , n493 );
not ( n2265 , n2264 );
and ( n2266 , n456 , n460 );
not ( n2267 , n456 );
and ( n2268 , n2267 , n476 );
nor ( n2269 , n2266 , n2268 );
not ( n2270 , n2269 );
not ( n2271 , n2270 );
or ( n2272 , n2265 , n2271 );
or ( n2273 , n2270 , n2264 );
nand ( n2274 , n2272 , n2273 );
nand ( n2275 , n2274 , n2185 );
nand ( n2276 , n2263 , n2275 );
xor ( n2277 , n2260 , n2276 );
not ( n2278 , n2060 );
not ( n2279 , n2077 );
or ( n2280 , n2278 , n2279 );
and ( n2281 , n495 , n2168 );
not ( n2282 , n495 );
not ( n2283 , n2168 );
and ( n2284 , n2282 , n2283 );
or ( n2285 , n2281 , n2284 );
nand ( n2286 , n2285 , n2078 );
nand ( n2287 , n2280 , n2286 );
not ( n2288 , n2287 );
xor ( n2289 , n2277 , n2288 );
and ( n2290 , n456 , n467 );
not ( n2291 , n456 );
and ( n2292 , n2291 , n483 );
nor ( n2293 , n2290 , n2292 );
not ( n2294 , n2293 );
and ( n2295 , n2294 , n489 );
buf ( n2296 , n2134 );
not ( n2297 , n473 );
nor ( n2298 , n2297 , n456 );
not ( n2299 , n2298 );
nand ( n2300 , n456 , n457 );
nand ( n2301 , n2299 , n2300 );
or ( n2302 , n2301 , n936 );
nand ( n2303 , n2148 , n936 );
nand ( n2304 , n2302 , n2303 );
and ( n2305 , n2296 , n2304 );
xor ( n2306 , n500 , n501 );
and ( n2307 , n2306 , n499 );
nor ( n2308 , n2305 , n2307 );
not ( n2309 , n2308 );
xor ( n2310 , n2295 , n2309 );
not ( n2311 , n2163 );
and ( n2312 , n456 , n459 );
not ( n2313 , n456 );
and ( n2314 , n2313 , n475 );
or ( n2315 , n2312 , n2314 );
not ( n2316 , n2315 );
not ( n2317 , n2057 );
or ( n2318 , n2316 , n2317 );
nand ( n2319 , n497 , n2066 );
nand ( n2320 , n2318 , n2319 );
not ( n2321 , n2320 );
or ( n2322 , n2311 , n2321 );
nand ( n2323 , n2177 , n2142 );
nand ( n2324 , n2322 , n2323 );
nand ( n2325 , n2182 , n495 );
nand ( n2326 , n917 , n494 );
nand ( n2327 , n2325 , n2326 );
not ( n2328 , n2327 );
not ( n2329 , n2212 );
or ( n2330 , n2328 , n2329 );
not ( n2331 , n2026 );
not ( n2332 , n2264 );
or ( n2333 , n2331 , n2332 );
nand ( n2334 , n2032 , n493 );
nand ( n2335 , n2333 , n2334 );
nand ( n2336 , n2335 , n2202 );
nand ( n2337 , n2330 , n2336 );
xor ( n2338 , n2324 , n2337 );
not ( n2339 , n2219 );
not ( n2340 , n2017 );
or ( n2341 , n2339 , n2340 );
not ( n2342 , n491 );
and ( n2343 , n456 , n465 );
not ( n2344 , n456 );
and ( n2345 , n2344 , n481 );
nor ( n2346 , n2343 , n2345 );
not ( n2347 , n2346 );
or ( n2348 , n2342 , n2347 );
and ( n2349 , n456 , n465 );
not ( n2350 , n456 );
and ( n2351 , n2350 , n481 );
nor ( n2352 , n2349 , n2351 );
not ( n2353 , n2352 );
nand ( n2354 , n2353 , n2015 );
nand ( n2355 , n2348 , n2354 );
nand ( n2356 , n2355 , n2000 );
nand ( n2357 , n2341 , n2356 );
and ( n2358 , n2338 , n2357 );
and ( n2359 , n2324 , n2337 );
or ( n2360 , n2358 , n2359 );
and ( n2361 , n2310 , n2360 );
and ( n2362 , n2295 , n2309 );
or ( n2363 , n2361 , n2362 );
xor ( n2364 , n2289 , n2363 );
not ( n2365 , n2060 );
and ( n2366 , n495 , n2190 );
not ( n2367 , n495 );
not ( n2368 , n461 );
not ( n2369 , n456 );
or ( n2370 , n2368 , n2369 );
not ( n2371 , n456 );
nand ( n2372 , n2371 , n477 );
nand ( n2373 , n2370 , n2372 );
and ( n2374 , n2367 , n2373 );
or ( n2375 , n2366 , n2374 );
not ( n2376 , n2375 );
or ( n2377 , n2365 , n2376 );
nand ( n2378 , n2053 , n2078 );
nand ( n2379 , n2377 , n2378 );
not ( n2380 , n2120 );
not ( n2381 , n1949 );
not ( n2382 , n467 );
and ( n2383 , n456 , n2382 );
not ( n2384 , n456 );
not ( n2385 , n483 );
and ( n2386 , n2384 , n2385 );
nor ( n2387 , n2383 , n2386 );
not ( n2388 , n2387 );
or ( n2389 , n2381 , n2388 );
nand ( n2390 , n2293 , n489 );
nand ( n2391 , n2389 , n2390 );
not ( n2392 , n2391 );
or ( n2393 , n2380 , n2392 );
nand ( n2394 , n2113 , n2082 );
nand ( n2395 , n2393 , n2394 );
xor ( n2396 , n2379 , n2395 );
and ( n2397 , n456 , n468 );
not ( n2398 , n456 );
and ( n2399 , n2398 , n484 );
nor ( n2400 , n2397 , n2399 );
not ( n2401 , n2400 );
and ( n2402 , n489 , n2401 );
and ( n2403 , n2396 , n2402 );
and ( n2404 , n2379 , n2395 );
or ( n2405 , n2403 , n2404 );
xor ( n2406 , n2038 , n2080 );
xor ( n2407 , n2406 , n2124 );
xor ( n2408 , n2405 , n2407 );
xor ( n2409 , n2136 , n2179 );
xor ( n2410 , n2409 , n2214 );
and ( n2411 , n2408 , n2410 );
and ( n2412 , n2405 , n2407 );
or ( n2413 , n2411 , n2412 );
xor ( n2414 , n2364 , n2413 );
xor ( n2415 , n2254 , n2414 );
xor ( n2416 , n2295 , n2309 );
xor ( n2417 , n2416 , n2360 );
not ( n2418 , n502 );
not ( n2419 , n503 );
not ( n2420 , n2419 );
or ( n2421 , n2418 , n2420 );
not ( n2422 , n502 );
nand ( n2423 , n2422 , n503 );
nand ( n2424 , n2421 , n2423 );
not ( n2425 , n2424 );
not ( n2426 , n2425 );
not ( n2427 , n501 );
nand ( n2428 , n2427 , n503 , n502 );
not ( n2429 , n502 );
not ( n2430 , n503 );
nand ( n2431 , n2429 , n2430 , n501 );
and ( n2432 , n2428 , n2431 );
not ( n2433 , n2432 );
or ( n2434 , n2426 , n2433 );
nand ( n2435 , n2434 , n501 );
not ( n2436 , n2128 );
not ( n2437 , n2304 );
or ( n2438 , n2436 , n2437 );
not ( n2439 , n499 );
not ( n2440 , n2168 );
or ( n2441 , n2439 , n2440 );
not ( n2442 , n499 );
nand ( n2443 , n2442 , n2175 );
nand ( n2444 , n2441 , n2443 );
not ( n2445 , n499 );
nor ( n2446 , n500 , n501 );
not ( n2447 , n2446 );
or ( n2448 , n2445 , n2447 );
nand ( n2449 , n2448 , n2133 );
nand ( n2450 , n2444 , n2449 );
nand ( n2451 , n2438 , n2450 );
xor ( n2452 , n2435 , n2451 );
not ( n2453 , n2060 );
not ( n2454 , n495 );
and ( n2455 , n456 , n462 );
not ( n2456 , n456 );
and ( n2457 , n2456 , n478 );
nor ( n2458 , n2455 , n2457 );
not ( n2459 , n2458 );
or ( n2460 , n2454 , n2459 );
or ( n2461 , n2458 , n495 );
nand ( n2462 , n2460 , n2461 );
not ( n2463 , n2462 );
or ( n2464 , n2453 , n2463 );
nand ( n2465 , n2375 , n2078 );
nand ( n2466 , n2464 , n2465 );
and ( n2467 , n2452 , n2466 );
and ( n2468 , n2435 , n2451 );
or ( n2469 , n2467 , n2468 );
xor ( n2470 , n2308 , n2469 );
and ( n2471 , n456 , n469 );
not ( n2472 , n456 );
and ( n2473 , n2472 , n485 );
nor ( n2474 , n2471 , n2473 );
nor ( n2475 , n2474 , n2118 );
not ( n2476 , n2327 );
not ( n2477 , n2335 );
or ( n2478 , n2476 , n2477 );
or ( n2479 , n2012 , n456 );
nand ( n2480 , n456 , n464 );
nand ( n2481 , n2479 , n2480 );
and ( n2482 , n493 , n2481 );
not ( n2483 , n493 );
not ( n2484 , n456 );
and ( n2485 , n2484 , n480 );
not ( n2486 , n2484 );
and ( n2487 , n2486 , n464 );
nor ( n2488 , n2485 , n2487 );
and ( n2489 , n2483 , n2488 );
nor ( n2490 , n2482 , n2489 );
nand ( n2491 , n2202 , n2490 );
nand ( n2492 , n2478 , n2491 );
xor ( n2493 , n2475 , n2492 );
not ( n2494 , n2163 );
not ( n2495 , n497 );
not ( n2496 , n2495 );
not ( n2497 , n2051 );
or ( n2498 , n2496 , n2497 );
or ( n2499 , n2051 , n2495 );
nand ( n2500 , n2498 , n2499 );
not ( n2501 , n2500 );
or ( n2502 , n2494 , n2501 );
nand ( n2503 , n2320 , n2142 );
nand ( n2504 , n2502 , n2503 );
and ( n2505 , n2493 , n2504 );
and ( n2506 , n2475 , n2492 );
or ( n2507 , n2505 , n2506 );
and ( n2508 , n2470 , n2507 );
and ( n2509 , n2308 , n2469 );
or ( n2510 , n2508 , n2509 );
xor ( n2511 , n2417 , n2510 );
xor ( n2512 , n2379 , n2395 );
xor ( n2513 , n2512 , n2402 );
xor ( n2514 , n2324 , n2337 );
xor ( n2515 , n2514 , n2357 );
xor ( n2516 , n2513 , n2515 );
not ( n2517 , n2219 );
not ( n2518 , n2355 );
or ( n2519 , n2517 , n2518 );
and ( n2520 , n493 , n1993 , n492 );
and ( n2521 , n2259 , n2520 );
not ( n2522 , n2259 );
not ( n2523 , n492 );
nand ( n2524 , n2523 , n1988 , n491 );
not ( n2525 , n2524 );
and ( n2526 , n2522 , n2525 );
nor ( n2527 , n2521 , n2526 );
nand ( n2528 , n2519 , n2527 );
not ( n2529 , n2084 );
not ( n2530 , n2391 );
or ( n2531 , n2529 , n2530 );
xor ( n2532 , n489 , n2401 );
nand ( n2533 , n2532 , n2120 );
nand ( n2534 , n2531 , n2533 );
xor ( n2535 , n2528 , n2534 );
nand ( n2536 , n2429 , n2430 , n501 );
nand ( n2537 , n2427 , n503 , n502 );
nand ( n2538 , n2536 , n2537 );
not ( n2539 , n2538 );
not ( n2540 , n501 );
nand ( n2541 , n2148 , n2540 );
nand ( n2542 , n2149 , n501 );
nand ( n2543 , n2541 , n2542 );
not ( n2544 , n2543 );
or ( n2545 , n2539 , n2544 );
and ( n2546 , n502 , n503 );
not ( n2547 , n502 );
not ( n2548 , n503 );
and ( n2549 , n2547 , n2548 );
nor ( n2550 , n2546 , n2549 );
buf ( n2551 , n2550 );
nand ( n2552 , n2551 , n501 );
nand ( n2553 , n2545 , n2552 );
and ( n2554 , n2535 , n2553 );
and ( n2555 , n2528 , n2534 );
or ( n2556 , n2554 , n2555 );
and ( n2557 , n2516 , n2556 );
and ( n2558 , n2513 , n2515 );
or ( n2559 , n2557 , n2558 );
and ( n2560 , n2511 , n2559 );
and ( n2561 , n2417 , n2510 );
or ( n2562 , n2560 , n2561 );
xor ( n2563 , n2415 , n2562 );
xor ( n2564 , n2405 , n2407 );
xor ( n2565 , n2564 , n2410 );
xor ( n2566 , n2417 , n2510 );
xor ( n2567 , n2566 , n2559 );
xor ( n2568 , n2565 , n2567 );
xor ( n2569 , n2308 , n2469 );
xor ( n2570 , n2569 , n2507 );
not ( n2571 , n2327 );
not ( n2572 , n2490 );
or ( n2573 , n2571 , n2572 );
not ( n2574 , n2352 );
not ( n2575 , n493 );
nand ( n2576 , n2575 , n495 , n494 );
not ( n2577 , n2576 );
and ( n2578 , n2574 , n2577 );
not ( n2579 , n2199 );
and ( n2580 , n2579 , n2346 );
nor ( n2581 , n2578 , n2580 );
nand ( n2582 , n2573 , n2581 );
not ( n2583 , n2163 );
not ( n2584 , n828 );
not ( n2585 , n2373 );
or ( n2586 , n2584 , n2585 );
nand ( n2587 , n456 , n461 );
nand ( n2588 , n2371 , n477 );
nand ( n2589 , n2587 , n2588 , n497 );
nand ( n2590 , n2586 , n2589 );
not ( n2591 , n2590 );
or ( n2592 , n2583 , n2591 );
nand ( n2593 , n2500 , n2142 );
nand ( n2594 , n2592 , n2593 );
xor ( n2595 , n2582 , n2594 );
not ( n2596 , n2000 );
not ( n2597 , n2015 );
not ( n2598 , n2294 );
or ( n2599 , n2597 , n2598 );
or ( n2600 , n2294 , n2015 );
nand ( n2601 , n2599 , n2600 );
not ( n2602 , n2601 );
or ( n2603 , n2596 , n2602 );
not ( n2604 , n491 );
not ( n2605 , n2258 );
or ( n2606 , n2604 , n2605 );
nand ( n2607 , n2259 , n2015 );
nand ( n2608 , n2606 , n2607 );
nand ( n2609 , n2608 , n2036 );
nand ( n2610 , n2603 , n2609 );
and ( n2611 , n2595 , n2610 );
and ( n2612 , n2582 , n2594 );
or ( n2613 , n2611 , n2612 );
not ( n2614 , n2306 );
not ( n2615 , n2444 );
or ( n2616 , n2614 , n2615 );
not ( n2617 , n1407 );
and ( n2618 , n456 , n2070 );
not ( n2619 , n456 );
and ( n2620 , n2619 , n2073 );
nor ( n2621 , n2618 , n2620 );
not ( n2622 , n2621 );
or ( n2623 , n2617 , n2622 );
not ( n2624 , n459 );
nand ( n2625 , n2624 , n456 );
not ( n2626 , n2625 );
not ( n2627 , n456 );
nand ( n2628 , n2627 , n2073 );
not ( n2629 , n2628 );
or ( n2630 , n2626 , n2629 );
nand ( n2631 , n2630 , n499 );
nand ( n2632 , n2623 , n2631 );
nand ( n2633 , n2134 , n2632 );
nand ( n2634 , n2616 , n2633 );
not ( n2635 , n470 );
and ( n2636 , n456 , n2635 );
not ( n2637 , n456 );
not ( n2638 , n486 );
and ( n2639 , n2637 , n2638 );
nor ( n2640 , n2636 , n2639 );
and ( n2641 , n2640 , n489 );
xor ( n2642 , n2634 , n2641 );
not ( n2643 , n2078 );
not ( n2644 , n2462 );
or ( n2645 , n2643 , n2644 );
not ( n2646 , n495 );
not ( n2647 , n2032 );
or ( n2648 , n2646 , n2647 );
not ( n2649 , n456 );
not ( n2650 , n463 );
not ( n2651 , n2650 );
or ( n2652 , n2649 , n2651 );
nor ( n2653 , n456 , n479 );
nor ( n2654 , n2653 , n495 );
nand ( n2655 , n2652 , n2654 );
nand ( n2656 , n2648 , n2655 );
nand ( n2657 , n2656 , n2060 );
nand ( n2658 , n2645 , n2657 );
and ( n2659 , n2642 , n2658 );
and ( n2660 , n2634 , n2641 );
or ( n2661 , n2659 , n2660 );
xor ( n2662 , n2613 , n2661 );
xor ( n2663 , n2435 , n2451 );
xor ( n2664 , n2663 , n2466 );
and ( n2665 , n2662 , n2664 );
and ( n2666 , n2613 , n2661 );
or ( n2667 , n2665 , n2666 );
xor ( n2668 , n2570 , n2667 );
xor ( n2669 , n2475 , n2492 );
xor ( n2670 , n2669 , n2504 );
xor ( n2671 , n2528 , n2534 );
xor ( n2672 , n2671 , n2553 );
xor ( n2673 , n2670 , n2672 );
not ( n2674 , n2084 );
not ( n2675 , n2532 );
or ( n2676 , n2674 , n2675 );
and ( n2677 , n456 , n469 );
not ( n2678 , n456 );
and ( n2679 , n2678 , n485 );
nor ( n2680 , n2677 , n2679 );
not ( n2681 , n2680 );
not ( n2682 , n489 );
or ( n2683 , n2681 , n2682 );
and ( n2684 , n456 , n469 );
not ( n2685 , n456 );
and ( n2686 , n2685 , n485 );
nor ( n2687 , n2684 , n2686 );
not ( n2688 , n2687 );
nand ( n2689 , n2688 , n1949 );
nand ( n2690 , n2683 , n2689 );
nand ( n2691 , n2690 , n2122 );
nand ( n2692 , n2676 , n2691 );
not ( n2693 , n2553 );
xor ( n2694 , n2692 , n2693 );
not ( n2695 , n504 );
nand ( n2696 , n2695 , n503 );
not ( n2697 , n2696 );
not ( n2698 , n2697 );
nand ( n2699 , n503 , n504 );
nand ( n2700 , n2698 , n2699 );
not ( n2701 , n2700 );
and ( n2702 , n2694 , n2701 );
and ( n2703 , n2692 , n2693 );
or ( n2704 , n2702 , n2703 );
and ( n2705 , n2673 , n2704 );
and ( n2706 , n2670 , n2672 );
or ( n2707 , n2705 , n2706 );
and ( n2708 , n2668 , n2707 );
and ( n2709 , n2570 , n2667 );
or ( n2710 , n2708 , n2709 );
and ( n2711 , n2568 , n2710 );
and ( n2712 , n2565 , n2567 );
or ( n2713 , n2711 , n2712 );
or ( n2714 , n2563 , n2713 );
nand ( n2715 , n2563 , n2713 );
and ( n2716 , n2714 , n2715 );
xor ( n2717 , n2513 , n2515 );
xor ( n2718 , n2717 , n2556 );
xor ( n2719 , n2570 , n2667 );
xor ( n2720 , n2719 , n2707 );
xor ( n2721 , n2718 , n2720 );
xor ( n2722 , n2613 , n2661 );
xor ( n2723 , n2722 , n2664 );
not ( n2724 , n2142 );
not ( n2725 , n2590 );
or ( n2726 , n2724 , n2725 );
not ( n2727 , n497 );
not ( n2728 , n2208 );
or ( n2729 , n2727 , n2728 );
not ( n2730 , n497 );
and ( n2731 , n456 , n462 );
not ( n2732 , n456 );
and ( n2733 , n2732 , n478 );
or ( n2734 , n2731 , n2733 );
nand ( n2735 , n2730 , n2734 );
nand ( n2736 , n2729 , n2735 );
nand ( n2737 , n2163 , n2736 );
nand ( n2738 , n2726 , n2737 );
not ( n2739 , n2690 );
not ( n2740 , n2243 );
or ( n2741 , n2739 , n2740 );
not ( n2742 , n1949 );
and ( n2743 , n456 , n470 );
not ( n2744 , n456 );
and ( n2745 , n2744 , n486 );
or ( n2746 , n2743 , n2745 );
not ( n2747 , n2746 );
or ( n2748 , n2742 , n2747 );
not ( n2749 , n456 );
nand ( n2750 , n2749 , n486 );
nand ( n2751 , n456 , n470 );
nand ( n2752 , n2750 , n2751 , n489 );
nand ( n2753 , n2748 , n2752 );
nand ( n2754 , n2120 , n2753 );
nand ( n2755 , n2741 , n2754 );
xor ( n2756 , n2738 , n2755 );
and ( n2757 , n456 , n471 );
not ( n2758 , n456 );
and ( n2759 , n2758 , n487 );
nor ( n2760 , n2757 , n2759 );
not ( n2761 , n2760 );
and ( n2762 , n2761 , n489 );
and ( n2763 , n2756 , n2762 );
and ( n2764 , n2738 , n2755 );
or ( n2765 , n2763 , n2764 );
not ( n2766 , n2060 );
and ( n2767 , n495 , n2006 );
not ( n2768 , n495 );
and ( n2769 , n2768 , n2014 );
or ( n2770 , n2767 , n2769 );
not ( n2771 , n2770 );
or ( n2772 , n2766 , n2771 );
nand ( n2773 , n2656 , n2078 );
nand ( n2774 , n2772 , n2773 );
nand ( n2775 , n2431 , n2428 );
not ( n2776 , n2775 );
not ( n2777 , n2540 );
not ( n2778 , n2283 );
or ( n2779 , n2777 , n2778 );
and ( n2780 , n456 , n458 );
not ( n2781 , n456 );
and ( n2782 , n2781 , n474 );
nor ( n2783 , n2780 , n2782 );
nand ( n2784 , n501 , n2783 );
nand ( n2785 , n2779 , n2784 );
not ( n2786 , n2785 );
or ( n2787 , n2776 , n2786 );
nand ( n2788 , n2543 , n2551 );
nand ( n2789 , n2787 , n2788 );
xor ( n2790 , n2774 , n2789 );
not ( n2791 , n499 );
and ( n2792 , n456 , n460 );
not ( n2793 , n456 );
and ( n2794 , n2793 , n476 );
nor ( n2795 , n2792 , n2794 );
not ( n2796 , n2795 );
or ( n2797 , n2791 , n2796 );
not ( n2798 , n476 );
not ( n2799 , n456 );
nand ( n2800 , n2798 , n2799 );
not ( n2801 , n460 );
nand ( n2802 , n2801 , n456 );
nand ( n2803 , n2800 , n2802 , n936 );
nand ( n2804 , n2797 , n2803 );
not ( n2805 , n2804 );
not ( n2806 , n2296 );
or ( n2807 , n2805 , n2806 );
nand ( n2808 , n2632 , n2306 );
nand ( n2809 , n2807 , n2808 );
and ( n2810 , n2790 , n2809 );
and ( n2811 , n2774 , n2789 );
or ( n2812 , n2810 , n2811 );
xor ( n2813 , n2765 , n2812 );
xor ( n2814 , n2582 , n2594 );
xor ( n2815 , n2814 , n2610 );
and ( n2816 , n2813 , n2815 );
and ( n2817 , n2765 , n2812 );
or ( n2818 , n2816 , n2817 );
xor ( n2819 , n2723 , n2818 );
xor ( n2820 , n2634 , n2641 );
xor ( n2821 , n2820 , n2658 );
not ( n2822 , n493 );
not ( n2823 , n2258 );
or ( n2824 , n2822 , n2823 );
not ( n2825 , n482 );
nand ( n2826 , n2627 , n2825 );
not ( n2827 , n466 );
nand ( n2828 , n2827 , n456 );
nand ( n2829 , n2826 , n2828 , n2264 );
nand ( n2830 , n2824 , n2829 );
nand ( n2831 , n2830 , n2202 );
not ( n2832 , n2264 );
not ( n2833 , n2090 );
or ( n2834 , n2832 , n2833 );
or ( n2835 , n2090 , n2264 );
nand ( n2836 , n2834 , n2835 );
nand ( n2837 , n2185 , n2836 );
nand ( n2838 , n2831 , n2837 );
not ( n2839 , n2036 );
not ( n2840 , n2601 );
or ( n2841 , n2839 , n2840 );
and ( n2842 , n456 , n468 );
not ( n2843 , n456 );
and ( n2844 , n2843 , n484 );
nor ( n2845 , n2842 , n2844 );
not ( n2846 , n2845 );
nand ( n2847 , n2846 , n2015 );
and ( n2848 , n456 , n468 );
not ( n2849 , n456 );
and ( n2850 , n2849 , n484 );
nor ( n2851 , n2848 , n2850 );
nand ( n2852 , n2851 , n491 );
nand ( n2853 , n2847 , n2852 );
nand ( n2854 , n2853 , n2000 );
nand ( n2855 , n2841 , n2854 );
xor ( n2856 , n2838 , n2855 );
and ( n2857 , n2856 , n2700 );
and ( n2858 , n2838 , n2855 );
or ( n2859 , n2857 , n2858 );
xor ( n2860 , n2821 , n2859 );
not ( n2861 , n2128 );
not ( n2862 , n2804 );
or ( n2863 , n2861 , n2862 );
and ( n2864 , n2446 , n499 );
and ( n2865 , n456 , n461 );
not ( n2866 , n456 );
and ( n2867 , n2866 , n477 );
or ( n2868 , n2865 , n2867 );
or ( n2869 , n2864 , n2868 );
and ( n2870 , n456 , n461 );
not ( n2871 , n456 );
and ( n2872 , n2871 , n477 );
nor ( n2873 , n2870 , n2872 );
not ( n2874 , n2873 );
not ( n2875 , n499 );
nand ( n2876 , n2875 , n501 , n500 );
nand ( n2877 , n2874 , n2876 );
nand ( n2878 , n2869 , n2877 );
nand ( n2879 , n2863 , n2878 );
not ( n2880 , n493 );
nor ( n2881 , n494 , n495 );
not ( n2882 , n2881 );
or ( n2883 , n2880 , n2882 );
nand ( n2884 , n2883 , n2576 );
not ( n2885 , n2884 );
not ( n2886 , n2264 );
not ( n2887 , n2387 );
or ( n2888 , n2886 , n2887 );
not ( n2889 , n456 );
nand ( n2890 , n2889 , n483 );
nand ( n2891 , n456 , n467 );
nand ( n2892 , n2890 , n2891 , n493 );
nand ( n2893 , n2888 , n2892 );
not ( n2894 , n2893 );
or ( n2895 , n2885 , n2894 );
nand ( n2896 , n2327 , n2830 );
nand ( n2897 , n2895 , n2896 );
xor ( n2898 , n2879 , n2897 );
not ( n2899 , n2219 );
not ( n2900 , n2853 );
or ( n2901 , n2899 , n2900 );
nand ( n2902 , n492 , n493 );
nor ( n2903 , n2902 , n491 );
or ( n2904 , n2474 , n2903 );
not ( n2905 , n491 );
nor ( n2906 , n492 , n493 );
not ( n2907 , n2906 );
or ( n2908 , n2905 , n2907 );
nand ( n2909 , n2908 , n2474 );
nand ( n2910 , n2904 , n2909 );
nand ( n2911 , n2901 , n2910 );
and ( n2912 , n2898 , n2911 );
and ( n2913 , n2879 , n2897 );
or ( n2914 , n2912 , n2913 );
not ( n2915 , n2120 );
not ( n2916 , n489 );
and ( n2917 , n456 , n471 );
not ( n2918 , n456 );
and ( n2919 , n2918 , n487 );
nor ( n2920 , n2917 , n2919 );
not ( n2921 , n2920 );
or ( n2922 , n2916 , n2921 );
or ( n2923 , n2920 , n489 );
nand ( n2924 , n2922 , n2923 );
not ( n2925 , n2924 );
or ( n2926 , n2915 , n2925 );
nand ( n2927 , n2753 , n2082 );
nand ( n2928 , n2926 , n2927 );
not ( n2929 , n2736 );
not ( n2930 , n498 );
not ( n2931 , n1407 );
or ( n2932 , n2930 , n2931 );
nand ( n2933 , n2932 , n2140 );
not ( n2934 , n2933 );
or ( n2935 , n2929 , n2934 );
not ( n2936 , n2057 );
and ( n2937 , n456 , n463 );
not ( n2938 , n456 );
and ( n2939 , n2938 , n479 );
nor ( n2940 , n2937 , n2939 );
not ( n2941 , n2940 );
not ( n2942 , n2941 );
or ( n2943 , n2936 , n2942 );
nand ( n2944 , n2032 , n497 );
nand ( n2945 , n2943 , n2944 );
nand ( n2946 , n2945 , n2163 );
nand ( n2947 , n2935 , n2946 );
xor ( n2948 , n2928 , n2947 );
not ( n2949 , n2060 );
not ( n2950 , n2095 );
not ( n2951 , n456 );
not ( n2952 , n481 );
and ( n2953 , n2951 , n2952 );
nor ( n2954 , n2953 , n495 );
not ( n2955 , n2954 );
or ( n2956 , n2950 , n2955 );
and ( n2957 , n456 , n465 );
not ( n2958 , n456 );
and ( n2959 , n2958 , n481 );
nor ( n2960 , n2957 , n2959 );
nand ( n2961 , n2960 , n495 );
nand ( n2962 , n2956 , n2961 );
not ( n2963 , n2962 );
or ( n2964 , n2949 , n2963 );
nand ( n2965 , n2770 , n2078 );
nand ( n2966 , n2964 , n2965 );
and ( n2967 , n2948 , n2966 );
and ( n2968 , n2928 , n2947 );
or ( n2969 , n2967 , n2968 );
xor ( n2970 , n2914 , n2969 );
and ( n2971 , n456 , n472 );
not ( n2972 , n456 );
and ( n2973 , n2972 , n488 );
or ( n2974 , n2971 , n2973 );
and ( n2975 , n2974 , n489 );
not ( n2976 , n2697 );
not ( n2977 , n2298 );
not ( n2978 , n2977 );
and ( n2979 , n2300 , n503 );
not ( n2980 , n2979 );
or ( n2981 , n2978 , n2980 );
not ( n2982 , n503 );
or ( n2983 , n456 , n473 );
not ( n2984 , n457 );
nand ( n2985 , n2984 , n456 );
nand ( n2986 , n2982 , n2983 , n2985 );
nand ( n2987 , n2981 , n2986 );
not ( n2988 , n2987 );
or ( n2989 , n2976 , n2988 );
nand ( n2990 , n2989 , n2699 );
xor ( n2991 , n2975 , n2990 );
buf ( n2992 , n2550 );
not ( n2993 , n2992 );
not ( n2994 , n2785 );
or ( n2995 , n2993 , n2994 );
and ( n2996 , n456 , n459 );
not ( n2997 , n456 );
and ( n2998 , n2997 , n475 );
nor ( n2999 , n2996 , n2998 );
not ( n3000 , n2999 );
and ( n3001 , n501 , n3000 );
not ( n3002 , n501 );
and ( n3003 , n3002 , n2999 );
nor ( n3004 , n3001 , n3003 );
buf ( n3005 , n3004 );
nand ( n3006 , n3005 , n2775 );
nand ( n3007 , n2995 , n3006 );
and ( n3008 , n2991 , n3007 );
and ( n3009 , n2975 , n2990 );
or ( n3010 , n3008 , n3009 );
and ( n3011 , n2970 , n3010 );
and ( n3012 , n2914 , n2969 );
or ( n3013 , n3011 , n3012 );
and ( n3014 , n2860 , n3013 );
and ( n3015 , n2821 , n2859 );
or ( n3016 , n3014 , n3015 );
and ( n3017 , n2819 , n3016 );
and ( n3018 , n2723 , n2818 );
or ( n3019 , n3017 , n3018 );
xor ( n3020 , n2721 , n3019 );
xor ( n3021 , n2670 , n2672 );
xor ( n3022 , n3021 , n2704 );
xor ( n3023 , n2692 , n2693 );
xor ( n3024 , n3023 , n2701 );
xor ( n3025 , n2765 , n2812 );
xor ( n3026 , n3025 , n2815 );
xor ( n3027 , n3024 , n3026 );
xor ( n3028 , n2738 , n2755 );
xor ( n3029 , n3028 , n2762 );
xor ( n3030 , n2774 , n2789 );
xor ( n3031 , n3030 , n2809 );
xor ( n3032 , n3029 , n3031 );
xor ( n3033 , n2838 , n2855 );
xor ( n3034 , n3033 , n2700 );
and ( n3035 , n3032 , n3034 );
and ( n3036 , n3029 , n3031 );
or ( n3037 , n3035 , n3036 );
and ( n3038 , n3027 , n3037 );
and ( n3039 , n3024 , n3026 );
or ( n3040 , n3038 , n3039 );
xor ( n3041 , n3022 , n3040 );
xor ( n3042 , n2723 , n2818 );
xor ( n3043 , n3042 , n3016 );
and ( n3044 , n3041 , n3043 );
and ( n3045 , n3022 , n3040 );
or ( n3046 , n3044 , n3045 );
nor ( n3047 , n3020 , n3046 );
xor ( n3048 , n2565 , n2567 );
xor ( n3049 , n3048 , n2710 );
xor ( n3050 , n2718 , n2720 );
and ( n3051 , n3050 , n3019 );
and ( n3052 , n2718 , n2720 );
or ( n3053 , n3051 , n3052 );
nor ( n3054 , n3049 , n3053 );
nor ( n3055 , n3047 , n3054 );
xor ( n3056 , n3022 , n3040 );
xor ( n3057 , n3056 , n3043 );
xor ( n3058 , n2821 , n2859 );
xor ( n3059 , n3058 , n3013 );
and ( n3060 , n456 , n472 );
not ( n3061 , n456 );
and ( n3062 , n3061 , n488 );
nor ( n3063 , n3060 , n3062 );
not ( n3064 , n3063 );
not ( n3065 , n2115 );
and ( n3066 , n3064 , n3065 );
nand ( n3067 , n490 , n491 );
nand ( n3068 , n3067 , n489 );
nor ( n3069 , n3066 , n3068 );
not ( n3070 , n504 );
not ( n3071 , n2987 );
or ( n3072 , n3070 , n3071 );
not ( n3073 , n503 );
and ( n3074 , n456 , n458 );
not ( n3075 , n456 );
and ( n3076 , n3075 , n474 );
nor ( n3077 , n3074 , n3076 );
and ( n3078 , n3073 , n3077 );
not ( n3079 , n3073 );
and ( n3080 , n3079 , n2175 );
nor ( n3081 , n3078 , n3080 );
nand ( n3082 , n3081 , n2697 );
nand ( n3083 , n3072 , n3082 );
and ( n3084 , n3069 , n3083 );
not ( n3085 , n2992 );
not ( n3086 , n3004 );
or ( n3087 , n3085 , n3086 );
not ( n3088 , n2043 );
nand ( n3089 , n3088 , n501 );
nand ( n3090 , n2431 , n2428 );
nand ( n3091 , n2269 , n2540 );
nand ( n3092 , n3089 , n3090 , n3091 );
nand ( n3093 , n3087 , n3092 );
not ( n3094 , n2082 );
not ( n3095 , n2924 );
or ( n3096 , n3094 , n3095 );
not ( n3097 , n489 );
and ( n3098 , n456 , n472 );
not ( n3099 , n456 );
and ( n3100 , n3099 , n488 );
nor ( n3101 , n3098 , n3100 );
not ( n3102 , n3101 );
or ( n3103 , n3097 , n3102 );
and ( n3104 , n456 , n472 );
not ( n3105 , n456 );
and ( n3106 , n3105 , n488 );
nor ( n3107 , n3104 , n3106 );
not ( n3108 , n3107 );
nand ( n3109 , n3108 , n1949 );
nand ( n3110 , n3103 , n3109 );
nand ( n3111 , n3110 , n2120 );
nand ( n3112 , n3096 , n3111 );
xor ( n3113 , n3093 , n3112 );
not ( n3114 , n497 );
not ( n3115 , n3114 );
not ( n3116 , n464 );
and ( n3117 , n456 , n3116 );
not ( n3118 , n456 );
not ( n3119 , n480 );
and ( n3120 , n3118 , n3119 );
nor ( n3121 , n3117 , n3120 );
not ( n3122 , n3121 );
or ( n3123 , n3115 , n3122 );
not ( n3124 , n464 );
and ( n3125 , n456 , n3124 );
not ( n3126 , n456 );
and ( n3127 , n3126 , n3119 );
nor ( n3128 , n3125 , n3127 );
or ( n3129 , n3128 , n3114 );
nand ( n3130 , n3123 , n3129 );
not ( n3131 , n3130 );
not ( n3132 , n2163 );
or ( n3133 , n3131 , n3132 );
nand ( n3134 , n2945 , n2142 );
nand ( n3135 , n3133 , n3134 );
and ( n3136 , n3113 , n3135 );
and ( n3137 , n3093 , n3112 );
or ( n3138 , n3136 , n3137 );
xor ( n3139 , n3084 , n3138 );
and ( n3140 , n496 , n497 );
not ( n3141 , n496 );
and ( n3142 , n3141 , n864 );
nor ( n3143 , n3140 , n3142 );
not ( n3144 , n3143 );
not ( n3145 , n2962 );
or ( n3146 , n3144 , n3145 );
not ( n3147 , n495 );
and ( n3148 , n456 , n466 );
not ( n3149 , n456 );
and ( n3150 , n3149 , n482 );
nor ( n3151 , n3148 , n3150 );
not ( n3152 , n3151 );
or ( n3153 , n3147 , n3152 );
not ( n3154 , n2627 );
not ( n3155 , n2825 );
or ( n3156 , n3154 , n3155 );
and ( n3157 , n2827 , n456 );
nor ( n3158 , n3157 , n495 );
nand ( n3159 , n3156 , n3158 );
nand ( n3160 , n3153 , n3159 );
not ( n3161 , n864 );
not ( n3162 , n495 );
nor ( n3163 , n3162 , n496 );
not ( n3164 , n3163 );
or ( n3165 , n3161 , n3164 );
nand ( n3166 , n3165 , n2056 );
nand ( n3167 , n3160 , n3166 );
nand ( n3168 , n3146 , n3167 );
not ( n3169 , n2134 );
and ( n3170 , n499 , n2208 );
not ( n3171 , n499 );
not ( n3172 , n478 );
not ( n3173 , n456 );
not ( n3174 , n3173 );
or ( n3175 , n3172 , n3174 );
nand ( n3176 , n456 , n462 );
nand ( n3177 , n3175 , n3176 );
and ( n3178 , n3171 , n3177 );
or ( n3179 , n3170 , n3178 );
not ( n3180 , n3179 );
or ( n3181 , n3169 , n3180 );
not ( n3182 , n499 );
nand ( n3183 , n3182 , n2373 );
not ( n3184 , n3183 );
nand ( n3185 , n2587 , n2588 , n499 );
not ( n3186 , n3185 );
or ( n3187 , n3184 , n3186 );
nand ( n3188 , n3187 , n2128 );
nand ( n3189 , n3181 , n3188 );
xor ( n3190 , n3168 , n3189 );
not ( n3191 , n2202 );
not ( n3192 , n493 );
nand ( n3193 , n3192 , n2846 );
and ( n3194 , n456 , n468 );
not ( n3195 , n456 );
and ( n3196 , n3195 , n484 );
nor ( n3197 , n3194 , n3196 );
nand ( n3198 , n3197 , n493 );
nand ( n3199 , n3193 , n3198 );
not ( n3200 , n3199 );
or ( n3201 , n3191 , n3200 );
nand ( n3202 , n2893 , n2327 );
nand ( n3203 , n3201 , n3202 );
and ( n3204 , n3190 , n3203 );
and ( n3205 , n3168 , n3189 );
or ( n3206 , n3204 , n3205 );
and ( n3207 , n3139 , n3206 );
and ( n3208 , n3084 , n3138 );
or ( n3209 , n3207 , n3208 );
xor ( n3210 , n2914 , n2969 );
xor ( n3211 , n3210 , n3010 );
xor ( n3212 , n3209 , n3211 );
xor ( n3213 , n2879 , n2897 );
xor ( n3214 , n3213 , n2911 );
xor ( n3215 , n2975 , n2990 );
xor ( n3216 , n3215 , n3007 );
xor ( n3217 , n3214 , n3216 );
xor ( n3218 , n2928 , n2947 );
xor ( n3219 , n3218 , n2966 );
and ( n3220 , n3217 , n3219 );
and ( n3221 , n3214 , n3216 );
or ( n3222 , n3220 , n3221 );
and ( n3223 , n3212 , n3222 );
and ( n3224 , n3209 , n3211 );
or ( n3225 , n3223 , n3224 );
xor ( n3226 , n3059 , n3225 );
xor ( n3227 , n3024 , n3026 );
xor ( n3228 , n3227 , n3037 );
and ( n3229 , n3226 , n3228 );
and ( n3230 , n3059 , n3225 );
or ( n3231 , n3229 , n3230 );
nor ( n3232 , n3057 , n3231 );
not ( n3233 , n3232 );
nand ( n3234 , n3055 , n3233 );
not ( n3235 , n3234 );
xor ( n3236 , n3214 , n3216 );
xor ( n3237 , n3236 , n3219 );
not ( n3238 , n2202 );
nand ( n3239 , n2799 , n485 );
nand ( n3240 , n456 , n469 );
nand ( n3241 , n3239 , n3240 );
xor ( n3242 , n493 , n3241 );
not ( n3243 , n3242 );
or ( n3244 , n3238 , n3243 );
nand ( n3245 , n3199 , n2327 );
nand ( n3246 , n3244 , n3245 );
not ( n3247 , n2219 );
not ( n3248 , n491 );
and ( n3249 , n456 , n470 );
not ( n3250 , n456 );
and ( n3251 , n3250 , n486 );
nor ( n3252 , n3249 , n3251 );
not ( n3253 , n3252 );
or ( n3254 , n3248 , n3253 );
and ( n3255 , n456 , n470 );
not ( n3256 , n456 );
and ( n3257 , n3256 , n486 );
nor ( n3258 , n3255 , n3257 );
not ( n3259 , n3258 );
nand ( n3260 , n3259 , n2015 );
nand ( n3261 , n3254 , n3260 );
not ( n3262 , n3261 );
or ( n3263 , n3247 , n3262 );
not ( n3264 , n491 );
and ( n3265 , n456 , n471 );
not ( n3266 , n456 );
and ( n3267 , n3266 , n487 );
nor ( n3268 , n3265 , n3267 );
not ( n3269 , n3268 );
or ( n3270 , n3264 , n3269 );
nand ( n3271 , n2761 , n2015 );
nand ( n3272 , n3270 , n3271 );
nand ( n3273 , n3272 , n2232 );
nand ( n3274 , n3263 , n3273 );
xor ( n3275 , n3246 , n3274 );
not ( n3276 , n488 );
or ( n3277 , n3276 , n456 );
nand ( n3278 , n456 , n472 );
nand ( n3279 , n3277 , n3278 );
or ( n3280 , n3279 , n492 );
nand ( n3281 , n3280 , n493 );
and ( n3282 , n3279 , n492 );
nor ( n3283 , n3282 , n2015 );
and ( n3284 , n3281 , n3283 );
not ( n3285 , n2697 );
and ( n3286 , n456 , n2801 );
not ( n3287 , n456 );
and ( n3288 , n3287 , n2798 );
nor ( n3289 , n3286 , n3288 );
not ( n3290 , n3289 );
not ( n3291 , n503 );
not ( n3292 , n3291 );
or ( n3293 , n3290 , n3292 );
nand ( n3294 , n2043 , n503 );
nand ( n3295 , n3293 , n3294 );
not ( n3296 , n3295 );
or ( n3297 , n3285 , n3296 );
and ( n3298 , n456 , n459 );
not ( n3299 , n456 );
and ( n3300 , n3299 , n475 );
nor ( n3301 , n3298 , n3300 );
and ( n3302 , n503 , n3301 );
not ( n3303 , n503 );
and ( n3304 , n3303 , n2621 );
or ( n3305 , n3302 , n3304 );
nand ( n3306 , n3305 , n504 );
nand ( n3307 , n3297 , n3306 );
and ( n3308 , n3284 , n3307 );
and ( n3309 , n3275 , n3308 );
and ( n3310 , n3246 , n3274 );
or ( n3311 , n3309 , n3310 );
not ( n3312 , n2219 );
and ( n3313 , n456 , n469 );
not ( n3314 , n456 );
and ( n3315 , n3314 , n485 );
or ( n3316 , n3313 , n3315 );
and ( n3317 , n491 , n3316 );
not ( n3318 , n491 );
and ( n3319 , n3318 , n2474 );
nor ( n3320 , n3317 , n3319 );
not ( n3321 , n3320 );
or ( n3322 , n3312 , n3321 );
nand ( n3323 , n3261 , n2232 );
nand ( n3324 , n3322 , n3323 );
xor ( n3325 , n3069 , n3083 );
xor ( n3326 , n3324 , n3325 );
not ( n3327 , n3107 );
and ( n3328 , n3327 , n2082 );
not ( n3329 , n503 );
nor ( n3330 , n3329 , n504 );
not ( n3331 , n3330 );
not ( n3332 , n3305 );
or ( n3333 , n3331 , n3332 );
nand ( n3334 , n3081 , n504 );
nand ( n3335 , n3333 , n3334 );
xor ( n3336 , n3328 , n3335 );
not ( n3337 , n2424 );
and ( n3338 , n2540 , n2269 );
not ( n3339 , n2540 );
not ( n3340 , n2043 );
and ( n3341 , n3339 , n3340 );
nor ( n3342 , n3338 , n3341 );
not ( n3343 , n3342 );
or ( n3344 , n3337 , n3343 );
not ( n3345 , n501 );
not ( n3346 , n2873 );
or ( n3347 , n3345 , n3346 );
not ( n3348 , n2889 );
not ( n3349 , n477 );
not ( n3350 , n3349 );
or ( n3351 , n3348 , n3350 );
not ( n3352 , n461 );
and ( n3353 , n3352 , n456 );
nor ( n3354 , n3353 , n501 );
nand ( n3355 , n3351 , n3354 );
nand ( n3356 , n3347 , n3355 );
nand ( n3357 , n2775 , n3356 );
nand ( n3358 , n3344 , n3357 );
and ( n3359 , n3336 , n3358 );
and ( n3360 , n3328 , n3335 );
or ( n3361 , n3359 , n3360 );
xor ( n3362 , n3326 , n3361 );
xor ( n3363 , n3311 , n3362 );
not ( n3364 , n3090 );
not ( n3365 , n501 );
and ( n3366 , n456 , n462 );
not ( n3367 , n456 );
and ( n3368 , n3367 , n478 );
nor ( n3369 , n3366 , n3368 );
not ( n3370 , n3369 );
or ( n3371 , n3365 , n3370 );
not ( n3372 , n462 );
and ( n3373 , n456 , n3372 );
not ( n3374 , n456 );
not ( n3375 , n478 );
and ( n3376 , n3374 , n3375 );
nor ( n3377 , n3373 , n3376 );
not ( n3378 , n501 );
nand ( n3379 , n3377 , n3378 );
nand ( n3380 , n3371 , n3379 );
not ( n3381 , n3380 );
or ( n3382 , n3364 , n3381 );
nand ( n3383 , n3356 , n2424 );
nand ( n3384 , n3382 , n3383 );
not ( n3385 , n2163 );
not ( n3386 , n497 );
not ( n3387 , n3151 );
or ( n3388 , n3386 , n3387 );
not ( n3389 , n3151 );
not ( n3390 , n497 );
nand ( n3391 , n3389 , n3390 );
nand ( n3392 , n3388 , n3391 );
not ( n3393 , n3392 );
or ( n3394 , n3385 , n3393 );
not ( n3395 , n3114 );
nand ( n3396 , n3173 , n481 );
nand ( n3397 , n456 , n465 );
nand ( n3398 , n3396 , n3397 );
not ( n3399 , n3398 );
or ( n3400 , n3395 , n3399 );
nand ( n3401 , n2089 , n497 );
nand ( n3402 , n3400 , n3401 );
xor ( n3403 , n498 , n499 );
nand ( n3404 , n3402 , n3403 );
nand ( n3405 , n3394 , n3404 );
xor ( n3406 , n3384 , n3405 );
not ( n3407 , n3143 );
not ( n3408 , n917 );
not ( n3409 , n2387 );
or ( n3410 , n3408 , n3409 );
or ( n3411 , n917 , n2387 );
nand ( n3412 , n3410 , n3411 );
not ( n3413 , n3412 );
or ( n3414 , n3407 , n3413 );
not ( n3415 , n495 );
and ( n3416 , n456 , n468 );
not ( n3417 , n456 );
and ( n3418 , n3417 , n484 );
nor ( n3419 , n3416 , n3418 );
not ( n3420 , n3419 );
or ( n3421 , n3415 , n3420 );
or ( n3422 , n495 , n3197 );
nand ( n3423 , n3421 , n3422 );
nand ( n3424 , n3423 , n2060 );
nand ( n3425 , n3414 , n3424 );
and ( n3426 , n3406 , n3425 );
and ( n3427 , n3384 , n3405 );
or ( n3428 , n3426 , n3427 );
not ( n3429 , n1576 );
not ( n3430 , n3128 );
or ( n3431 , n3429 , n3430 );
or ( n3432 , n2012 , n456 );
or ( n3433 , n2009 , n2371 );
nand ( n3434 , n3432 , n3433 , n499 );
nand ( n3435 , n3431 , n3434 );
not ( n3436 , n3435 );
not ( n3437 , n2134 );
or ( n3438 , n3436 , n3437 );
not ( n3439 , n499 );
not ( n3440 , n2940 );
or ( n3441 , n3439 , n3440 );
or ( n3442 , n2940 , n499 );
nand ( n3443 , n3441 , n3442 );
nand ( n3444 , n3443 , n2128 );
nand ( n3445 , n3438 , n3444 );
not ( n3446 , n2327 );
not ( n3447 , n3242 );
or ( n3448 , n3446 , n3447 );
not ( n3449 , n493 );
not ( n3450 , n3449 );
and ( n3451 , n456 , n2635 );
not ( n3452 , n456 );
and ( n3453 , n3452 , n2638 );
nor ( n3454 , n3451 , n3453 );
not ( n3455 , n3454 );
or ( n3456 , n3450 , n3455 );
or ( n3457 , n3454 , n3449 );
nand ( n3458 , n3456 , n3457 );
nand ( n3459 , n3458 , n2884 );
nand ( n3460 , n3448 , n3459 );
xor ( n3461 , n3445 , n3460 );
not ( n3462 , n2036 );
not ( n3463 , n3272 );
or ( n3464 , n3462 , n3463 );
not ( n3465 , n491 );
not ( n3466 , n3101 );
or ( n3467 , n3465 , n3466 );
or ( n3468 , n3101 , n491 );
nand ( n3469 , n3467 , n3468 );
nand ( n3470 , n2232 , n3469 );
nand ( n3471 , n3464 , n3470 );
and ( n3472 , n3461 , n3471 );
and ( n3473 , n3445 , n3460 );
or ( n3474 , n3472 , n3473 );
xor ( n3475 , n3428 , n3474 );
xor ( n3476 , n3328 , n3335 );
xor ( n3477 , n3476 , n3358 );
and ( n3478 , n3475 , n3477 );
and ( n3479 , n3428 , n3474 );
or ( n3480 , n3478 , n3479 );
and ( n3481 , n3363 , n3480 );
and ( n3482 , n3311 , n3362 );
or ( n3483 , n3481 , n3482 );
xor ( n3484 , n3237 , n3483 );
xor ( n3485 , n3324 , n3325 );
and ( n3486 , n3485 , n3361 );
and ( n3487 , n3324 , n3325 );
or ( n3488 , n3486 , n3487 );
xor ( n3489 , n3084 , n3138 );
xor ( n3490 , n3489 , n3206 );
xor ( n3491 , n3488 , n3490 );
nand ( n3492 , n2163 , n3402 );
nand ( n3493 , n3130 , n3403 );
nand ( n3494 , n3492 , n3493 );
not ( n3495 , n2060 );
not ( n3496 , n3412 );
or ( n3497 , n3495 , n3496 );
and ( n3498 , n496 , n497 );
not ( n3499 , n496 );
and ( n3500 , n3499 , n864 );
nor ( n3501 , n3498 , n3500 );
nand ( n3502 , n3160 , n3501 );
nand ( n3503 , n3497 , n3502 );
xor ( n3504 , n3494 , n3503 );
not ( n3505 , n2449 );
not ( n3506 , n3443 );
or ( n3507 , n3505 , n3506 );
nand ( n3508 , n3179 , n2128 );
nand ( n3509 , n3507 , n3508 );
and ( n3510 , n3504 , n3509 );
and ( n3511 , n3494 , n3503 );
or ( n3512 , n3510 , n3511 );
xor ( n3513 , n3168 , n3189 );
xor ( n3514 , n3513 , n3203 );
xor ( n3515 , n3512 , n3514 );
xor ( n3516 , n3093 , n3112 );
xor ( n3517 , n3516 , n3135 );
and ( n3518 , n3515 , n3517 );
and ( n3519 , n3512 , n3514 );
or ( n3520 , n3518 , n3519 );
xor ( n3521 , n3491 , n3520 );
xor ( n3522 , n3484 , n3521 );
not ( n3523 , n3522 );
xor ( n3524 , n3512 , n3514 );
xor ( n3525 , n3524 , n3517 );
xor ( n3526 , n3494 , n3503 );
xor ( n3527 , n3526 , n3509 );
xor ( n3528 , n3246 , n3274 );
xor ( n3529 , n3528 , n3308 );
xor ( n3530 , n3527 , n3529 );
xor ( n3531 , n3284 , n3307 );
and ( n3532 , n456 , n472 );
not ( n3533 , n456 );
and ( n3534 , n3533 , n488 );
or ( n3535 , n3532 , n3534 );
and ( n3536 , n2219 , n3535 );
not ( n3537 , n501 );
not ( n3538 , n2032 );
or ( n3539 , n3537 , n3538 );
not ( n3540 , n479 );
nand ( n3541 , n3540 , n2627 );
not ( n3542 , n463 );
nand ( n3543 , n3542 , n456 );
nand ( n3544 , n3541 , n3543 , n2540 );
nand ( n3545 , n3539 , n3544 );
not ( n3546 , n3545 );
not ( n3547 , n2538 );
or ( n3548 , n3546 , n3547 );
not ( n3549 , n503 );
not ( n3550 , n2422 );
or ( n3551 , n3549 , n3550 );
nand ( n3552 , n2419 , n502 );
nand ( n3553 , n3551 , n3552 );
nand ( n3554 , n3380 , n3553 );
nand ( n3555 , n3548 , n3554 );
xor ( n3556 , n3536 , n3555 );
not ( n3557 , n2142 );
not ( n3558 , n3392 );
or ( n3559 , n3557 , n3558 );
not ( n3560 , n497 );
and ( n3561 , n456 , n467 );
not ( n3562 , n456 );
and ( n3563 , n3562 , n483 );
nor ( n3564 , n3561 , n3563 );
not ( n3565 , n3564 );
or ( n3566 , n3560 , n3565 );
or ( n3567 , n3564 , n497 );
nand ( n3568 , n3566 , n3567 );
nand ( n3569 , n3568 , n2163 );
nand ( n3570 , n3559 , n3569 );
and ( n3571 , n3556 , n3570 );
and ( n3572 , n3536 , n3555 );
or ( n3573 , n3571 , n3572 );
xor ( n3574 , n3531 , n3573 );
not ( n3575 , n3501 );
not ( n3576 , n3423 );
or ( n3577 , n3575 , n3576 );
not ( n3578 , n485 );
not ( n3579 , n2022 );
or ( n3580 , n3578 , n3579 );
nand ( n3581 , n456 , n469 );
nand ( n3582 , n3580 , n3581 );
not ( n3583 , n495 );
nand ( n3584 , n3582 , n3583 );
and ( n3585 , n456 , n469 );
not ( n3586 , n456 );
and ( n3587 , n3586 , n485 );
nor ( n3588 , n3585 , n3587 );
nand ( n3589 , n3588 , n495 );
nand ( n3590 , n3584 , n3589 );
nand ( n3591 , n3166 , n3590 );
nand ( n3592 , n3577 , n3591 );
not ( n3593 , n3330 );
not ( n3594 , n2548 );
not ( n3595 , n2373 );
or ( n3596 , n3594 , n3595 );
nand ( n3597 , n2190 , n503 );
nand ( n3598 , n3596 , n3597 );
not ( n3599 , n3598 );
or ( n3600 , n3593 , n3599 );
nand ( n3601 , n3295 , n504 );
nand ( n3602 , n3600 , n3601 );
xor ( n3603 , n3592 , n3602 );
not ( n3604 , n2185 );
not ( n3605 , n3458 );
or ( n3606 , n3604 , n3605 );
and ( n3607 , n493 , n3268 );
not ( n3608 , n493 );
and ( n3609 , n3608 , n2761 );
or ( n3610 , n3607 , n3609 );
nand ( n3611 , n3610 , n2884 );
nand ( n3612 , n3606 , n3611 );
and ( n3613 , n3603 , n3612 );
and ( n3614 , n3592 , n3602 );
or ( n3615 , n3613 , n3614 );
and ( n3616 , n3574 , n3615 );
and ( n3617 , n3531 , n3573 );
or ( n3618 , n3616 , n3617 );
and ( n3619 , n3530 , n3618 );
and ( n3620 , n3527 , n3529 );
or ( n3621 , n3619 , n3620 );
xor ( n3622 , n3525 , n3621 );
xor ( n3623 , n3311 , n3362 );
xor ( n3624 , n3623 , n3480 );
and ( n3625 , n3622 , n3624 );
and ( n3626 , n3525 , n3621 );
or ( n3627 , n3625 , n3626 );
not ( n3628 , n3627 );
nand ( n3629 , n3523 , n3628 );
buf ( n3630 , n3629 );
xor ( n3631 , n3059 , n3225 );
xor ( n3632 , n3631 , n3228 );
not ( n3633 , n3632 );
xor ( n3634 , n3029 , n3031 );
xor ( n3635 , n3634 , n3034 );
xor ( n3636 , n3488 , n3490 );
and ( n3637 , n3636 , n3520 );
and ( n3638 , n3488 , n3490 );
or ( n3639 , n3637 , n3638 );
xor ( n3640 , n3635 , n3639 );
xor ( n3641 , n3209 , n3211 );
xor ( n3642 , n3641 , n3222 );
and ( n3643 , n3640 , n3642 );
and ( n3644 , n3635 , n3639 );
or ( n3645 , n3643 , n3644 );
not ( n3646 , n3645 );
nand ( n3647 , n3633 , n3646 );
xor ( n3648 , n3635 , n3639 );
xor ( n3649 , n3648 , n3642 );
not ( n3650 , n3649 );
xor ( n3651 , n3237 , n3483 );
and ( n3652 , n3651 , n3521 );
and ( n3653 , n3237 , n3483 );
or ( n3654 , n3652 , n3653 );
not ( n3655 , n3654 );
nand ( n3656 , n3650 , n3655 );
and ( n3657 , n3630 , n3647 , n3656 );
xor ( n3658 , n3428 , n3474 );
xor ( n3659 , n3658 , n3477 );
xor ( n3660 , n3527 , n3529 );
xor ( n3661 , n3660 , n3618 );
xor ( n3662 , n3659 , n3661 );
xor ( n3663 , n3445 , n3460 );
xor ( n3664 , n3663 , n3471 );
xor ( n3665 , n3384 , n3405 );
xor ( n3666 , n3665 , n3425 );
xor ( n3667 , n3664 , n3666 );
not ( n3668 , n499 );
not ( n3669 , n2960 );
or ( n3670 , n3668 , n3669 );
nand ( n3671 , n3398 , n2158 );
nand ( n3672 , n3670 , n3671 );
not ( n3673 , n3672 );
not ( n3674 , n2296 );
or ( n3675 , n3673 , n3674 );
nand ( n3676 , n3435 , n2306 );
nand ( n3677 , n3675 , n3676 );
nand ( n3678 , n2182 , n917 );
nand ( n3679 , n3678 , n3327 );
nand ( n3680 , n494 , n495 );
and ( n3681 , n3679 , n3680 , n493 );
not ( n3682 , n3553 );
not ( n3683 , n3545 );
or ( n3684 , n3682 , n3683 );
not ( n3685 , n3121 );
not ( n3686 , n2540 );
or ( n3687 , n3685 , n3686 );
nand ( n3688 , n2006 , n501 );
nand ( n3689 , n3687 , n3688 );
nand ( n3690 , n2538 , n3689 );
nand ( n3691 , n3684 , n3690 );
and ( n3692 , n3681 , n3691 );
xor ( n3693 , n3677 , n3692 );
not ( n3694 , n3403 );
not ( n3695 , n3568 );
or ( n3696 , n3694 , n3695 );
not ( n3697 , n2495 );
not ( n3698 , n3419 );
not ( n3699 , n3698 );
or ( n3700 , n3697 , n3699 );
nand ( n3701 , n2851 , n497 );
nand ( n3702 , n3700 , n3701 );
nand ( n3703 , n2163 , n3702 );
nand ( n3704 , n3696 , n3703 );
not ( n3705 , n2060 );
not ( n3706 , n495 );
not ( n3707 , n3252 );
or ( n3708 , n3706 , n3707 );
not ( n3709 , n495 );
and ( n3710 , n456 , n470 );
not ( n3711 , n456 );
and ( n3712 , n3711 , n486 );
or ( n3713 , n3710 , n3712 );
nand ( n3714 , n3709 , n3713 );
nand ( n3715 , n3708 , n3714 );
not ( n3716 , n3715 );
or ( n3717 , n3705 , n3716 );
nand ( n3718 , n3590 , n3143 );
nand ( n3719 , n3717 , n3718 );
xor ( n3720 , n3704 , n3719 );
not ( n3721 , n504 );
not ( n3722 , n3598 );
or ( n3723 , n3721 , n3722 );
not ( n3724 , n3176 );
nand ( n3725 , n3724 , n3291 );
nand ( n3726 , n3369 , n503 );
nand ( n3727 , n478 , n3291 , n2889 );
nand ( n3728 , n3725 , n3726 , n3727 );
nand ( n3729 , n3728 , n2697 );
nand ( n3730 , n3723 , n3729 );
and ( n3731 , n3720 , n3730 );
and ( n3732 , n3704 , n3719 );
or ( n3733 , n3731 , n3732 );
and ( n3734 , n3693 , n3733 );
and ( n3735 , n3677 , n3692 );
or ( n3736 , n3734 , n3735 );
and ( n3737 , n3667 , n3736 );
and ( n3738 , n3664 , n3666 );
or ( n3739 , n3737 , n3738 );
xor ( n3740 , n3662 , n3739 );
not ( n3741 , n3740 );
xor ( n3742 , n3531 , n3573 );
xor ( n3743 , n3742 , n3615 );
xor ( n3744 , n3592 , n3602 );
xor ( n3745 , n3744 , n3612 );
xor ( n3746 , n3536 , n3555 );
xor ( n3747 , n3746 , n3570 );
xor ( n3748 , n3745 , n3747 );
not ( n3749 , n2327 );
not ( n3750 , n3610 );
or ( n3751 , n3749 , n3750 );
and ( n3752 , n493 , n3101 );
not ( n3753 , n493 );
and ( n3754 , n3753 , n3535 );
or ( n3755 , n3752 , n3754 );
nand ( n3756 , n3755 , n2884 );
nand ( n3757 , n3751 , n3756 );
not ( n3758 , n2296 );
not ( n3759 , n1407 );
not ( n3760 , n2259 );
or ( n3761 , n3759 , n3760 );
nand ( n3762 , n2108 , n499 );
nand ( n3763 , n3761 , n3762 );
not ( n3764 , n3763 );
or ( n3765 , n3758 , n3764 );
nand ( n3766 , n3672 , n2306 );
nand ( n3767 , n3765 , n3766 );
xor ( n3768 , n3757 , n3767 );
xor ( n3769 , n3681 , n3691 );
and ( n3770 , n3768 , n3769 );
and ( n3771 , n3757 , n3767 );
or ( n3772 , n3770 , n3771 );
and ( n3773 , n3748 , n3772 );
and ( n3774 , n3745 , n3747 );
or ( n3775 , n3773 , n3774 );
xor ( n3776 , n3743 , n3775 );
xor ( n3777 , n3664 , n3666 );
xor ( n3778 , n3777 , n3736 );
and ( n3779 , n3776 , n3778 );
and ( n3780 , n3743 , n3775 );
or ( n3781 , n3779 , n3780 );
not ( n3782 , n3781 );
nor ( n3783 , n3741 , n3782 );
not ( n3784 , n3783 );
xor ( n3785 , n3525 , n3621 );
xor ( n3786 , n3785 , n3624 );
not ( n3787 , n3786 );
xor ( n3788 , n3659 , n3661 );
and ( n3789 , n3788 , n3739 );
and ( n3790 , n3659 , n3661 );
or ( n3791 , n3789 , n3790 );
not ( n3792 , n3791 );
nand ( n3793 , n3787 , n3792 );
not ( n3794 , n3793 );
or ( n3795 , n3784 , n3794 );
not ( n3796 , n3627 );
not ( n3797 , n3522 );
or ( n3798 , n3796 , n3797 );
nand ( n3799 , n3786 , n3791 );
nand ( n3800 , n3798 , n3799 );
not ( n3801 , n3800 );
nand ( n3802 , n3795 , n3801 );
not ( n3803 , n3802 );
not ( n3804 , n3143 );
not ( n3805 , n3715 );
or ( n3806 , n3804 , n3805 );
nor ( n3807 , n456 , n487 );
not ( n3808 , n3807 );
not ( n3809 , n471 );
nand ( n3810 , n3809 , n456 );
nand ( n3811 , n3808 , n3810 , n3583 );
not ( n3812 , n917 );
nand ( n3813 , n3812 , n3268 );
nand ( n3814 , n3811 , n3813 );
nand ( n3815 , n3814 , n3166 );
nand ( n3816 , n3806 , n3815 );
not ( n3817 , n504 );
not ( n3818 , n3728 );
or ( n3819 , n3817 , n3818 );
xor ( n3820 , n503 , n2941 );
nand ( n3821 , n3820 , n3330 );
nand ( n3822 , n3819 , n3821 );
xor ( n3823 , n3816 , n3822 );
not ( n3824 , n2449 );
not ( n3825 , n499 );
not ( n3826 , n2293 );
or ( n3827 , n3825 , n3826 );
and ( n3828 , n456 , n467 );
not ( n3829 , n456 );
and ( n3830 , n3829 , n483 );
nor ( n3831 , n3828 , n3830 );
not ( n3832 , n3831 );
nand ( n3833 , n1407 , n3832 );
nand ( n3834 , n3827 , n3833 );
not ( n3835 , n3834 );
or ( n3836 , n3824 , n3835 );
nand ( n3837 , n3763 , n2128 );
nand ( n3838 , n3836 , n3837 );
xor ( n3839 , n3823 , n3838 );
not ( n3840 , n2306 );
not ( n3841 , n3834 );
or ( n3842 , n3840 , n3841 );
not ( n3843 , n499 );
not ( n3844 , n2400 );
or ( n3845 , n3843 , n3844 );
or ( n3846 , n499 , n3197 );
nand ( n3847 , n3845 , n3846 );
nand ( n3848 , n3847 , n2134 );
nand ( n3849 , n3842 , n3848 );
or ( n3850 , n496 , n497 );
and ( n3851 , n3850 , n3279 );
nand ( n3852 , n496 , n497 );
nand ( n3853 , n3852 , n495 );
nor ( n3854 , n3851 , n3853 );
not ( n3855 , n2538 );
not ( n3856 , n501 );
not ( n3857 , n2258 );
or ( n3858 , n3856 , n3857 );
not ( n3859 , n456 );
not ( n3860 , n482 );
and ( n3861 , n3859 , n3860 );
nor ( n3862 , n3861 , n501 );
nand ( n3863 , n2827 , n456 );
nand ( n3864 , n3862 , n3863 );
nand ( n3865 , n3858 , n3864 );
not ( n3866 , n3865 );
or ( n3867 , n3855 , n3866 );
not ( n3868 , n501 );
not ( n3869 , n2960 );
or ( n3870 , n3868 , n3869 );
not ( n3871 , n3397 );
not ( n3872 , n3396 );
or ( n3873 , n3871 , n3872 );
nand ( n3874 , n3873 , n2540 );
nand ( n3875 , n3870 , n3874 );
nand ( n3876 , n3875 , n2551 );
nand ( n3877 , n3867 , n3876 );
xor ( n3878 , n3854 , n3877 );
xor ( n3879 , n3849 , n3878 );
and ( n3880 , n3327 , n3501 );
not ( n3881 , n504 );
nand ( n3882 , n2006 , n503 );
nand ( n3883 , n3073 , n456 , n464 );
not ( n3884 , n503 );
nand ( n3885 , n3884 , n2484 , n480 );
nand ( n3886 , n3882 , n3883 , n3885 );
not ( n3887 , n3886 );
or ( n3888 , n3881 , n3887 );
not ( n3889 , n503 );
not ( n3890 , n2960 );
or ( n3891 , n3889 , n3890 );
and ( n3892 , n456 , n465 );
not ( n3893 , n456 );
and ( n3894 , n3893 , n481 );
or ( n3895 , n3892 , n3894 );
nand ( n3896 , n3895 , n3884 );
nand ( n3897 , n3891 , n3896 );
nand ( n3898 , n3897 , n3330 );
nand ( n3899 , n3888 , n3898 );
xor ( n3900 , n3880 , n3899 );
not ( n3901 , n2142 );
not ( n3902 , n2627 );
not ( n3903 , n486 );
or ( n3904 , n3902 , n3903 );
nand ( n3905 , n456 , n470 );
nand ( n3906 , n3904 , n3905 );
and ( n3907 , n497 , n3906 );
not ( n3908 , n497 );
and ( n3909 , n456 , n2635 );
not ( n3910 , n456 );
and ( n3911 , n3910 , n2638 );
nor ( n3912 , n3909 , n3911 );
not ( n3913 , n3912 );
and ( n3914 , n3908 , n3913 );
nor ( n3915 , n3907 , n3914 );
not ( n3916 , n3915 );
or ( n3917 , n3901 , n3916 );
not ( n3918 , n497 );
not ( n3919 , n3268 );
or ( n3920 , n3918 , n3919 );
and ( n3921 , n456 , n3809 );
not ( n3922 , n456 );
not ( n3923 , n487 );
and ( n3924 , n3922 , n3923 );
nor ( n3925 , n3921 , n3924 );
nand ( n3926 , n3925 , n3390 );
nand ( n3927 , n3920 , n3926 );
nand ( n3928 , n3927 , n2163 );
nand ( n3929 , n3917 , n3928 );
and ( n3930 , n3900 , n3929 );
and ( n3931 , n3880 , n3899 );
or ( n3932 , n3930 , n3931 );
and ( n3933 , n3879 , n3932 );
and ( n3934 , n3849 , n3878 );
or ( n3935 , n3933 , n3934 );
xor ( n3936 , n3839 , n3935 );
and ( n3937 , n3854 , n3877 );
not ( n3938 , n3403 );
and ( n3939 , n3588 , n497 );
not ( n3940 , n3588 );
and ( n3941 , n3940 , n2057 );
or ( n3942 , n3939 , n3941 );
not ( n3943 , n3942 );
or ( n3944 , n3938 , n3943 );
nand ( n3945 , n2163 , n3915 );
nand ( n3946 , n3944 , n3945 );
not ( n3947 , n2060 );
not ( n3948 , n495 );
not ( n3949 , n3948 );
not ( n3950 , n3108 );
or ( n3951 , n3949 , n3950 );
or ( n3952 , n3948 , n3327 );
nand ( n3953 , n3951 , n3952 );
not ( n3954 , n3953 );
or ( n3955 , n3947 , n3954 );
nand ( n3956 , n3143 , n3814 );
nand ( n3957 , n3955 , n3956 );
xor ( n3958 , n3946 , n3957 );
not ( n3959 , n2697 );
not ( n3960 , n3886 );
or ( n3961 , n3959 , n3960 );
nand ( n3962 , n3820 , n504 );
nand ( n3963 , n3961 , n3962 );
and ( n3964 , n3958 , n3963 );
and ( n3965 , n3946 , n3957 );
or ( n3966 , n3964 , n3965 );
xor ( n3967 , n3937 , n3966 );
not ( n3968 , n488 );
nor ( n3969 , n3968 , n456 );
not ( n3970 , n3969 );
and ( n3971 , n472 , n456 );
not ( n3972 , n3971 );
and ( n3973 , n3970 , n3972 );
nand ( n3974 , n917 , n494 );
and ( n3975 , n3974 , n2325 );
nor ( n3976 , n3973 , n3975 );
not ( n3977 , n2992 );
not ( n3978 , n3689 );
or ( n3979 , n3977 , n3978 );
nand ( n3980 , n3875 , n3090 );
nand ( n3981 , n3979 , n3980 );
xor ( n3982 , n3976 , n3981 );
not ( n3983 , n2163 );
not ( n3984 , n3942 );
or ( n3985 , n3983 , n3984 );
nand ( n3986 , n3702 , n2142 );
nand ( n3987 , n3985 , n3986 );
xor ( n3988 , n3982 , n3987 );
xor ( n3989 , n3967 , n3988 );
xor ( n3990 , n3936 , n3989 );
not ( n3991 , n3990 );
xor ( n3992 , n3946 , n3957 );
xor ( n3993 , n3992 , n3963 );
not ( n3994 , n2538 );
and ( n3995 , n3831 , n3378 );
not ( n3996 , n3831 );
and ( n3997 , n3996 , n501 );
nor ( n3998 , n3995 , n3997 );
not ( n3999 , n3998 );
or ( n4000 , n3994 , n3999 );
nand ( n4001 , n3865 , n2551 );
nand ( n4002 , n4000 , n4001 );
not ( n4003 , n2449 );
nand ( n4004 , n499 , n2680 );
or ( n4005 , n456 , n485 );
not ( n4006 , n469 );
nand ( n4007 , n4006 , n456 );
nand ( n4008 , n4005 , n4007 , n1692 );
nand ( n4009 , n4004 , n4008 );
not ( n4010 , n4009 );
or ( n4011 , n4003 , n4010 );
nand ( n4012 , n3847 , n2306 );
nand ( n4013 , n4011 , n4012 );
xor ( n4014 , n4002 , n4013 );
nor ( n4015 , n498 , n499 );
not ( n4016 , n4015 );
and ( n4017 , n4016 , n3535 );
not ( n4018 , n498 );
not ( n4019 , n499 );
or ( n4020 , n4018 , n4019 );
nand ( n4021 , n4020 , n497 );
nor ( n4022 , n4017 , n4021 );
not ( n4023 , n504 );
not ( n4024 , n3897 );
or ( n4025 , n4023 , n4024 );
and ( n4026 , n3389 , n503 );
not ( n4027 , n3389 );
not ( n4028 , n503 );
and ( n4029 , n4027 , n4028 );
nor ( n4030 , n4026 , n4029 );
nand ( n4031 , n4030 , n2697 );
nand ( n4032 , n4025 , n4031 );
and ( n4033 , n4022 , n4032 );
and ( n4034 , n4014 , n4033 );
and ( n4035 , n4002 , n4013 );
or ( n4036 , n4034 , n4035 );
xor ( n4037 , n3993 , n4036 );
xor ( n4038 , n3849 , n3878 );
xor ( n4039 , n4038 , n3932 );
and ( n4040 , n4037 , n4039 );
and ( n4041 , n3993 , n4036 );
or ( n4042 , n4040 , n4041 );
not ( n4043 , n4042 );
nand ( n4044 , n3991 , n4043 );
not ( n4045 , n4044 );
xor ( n4046 , n3993 , n4036 );
xor ( n4047 , n4046 , n4039 );
nand ( n4048 , n4015 , n497 );
not ( n4049 , n4048 );
not ( n4050 , n3101 );
or ( n4051 , n4049 , n4050 );
not ( n4052 , n498 );
nor ( n4053 , n4052 , n1692 , n497 );
or ( n4054 , n3101 , n4053 );
nand ( n4055 , n4051 , n4054 );
and ( n4056 , n498 , n1407 );
not ( n4057 , n498 );
and ( n4058 , n4057 , n499 );
or ( n4059 , n4056 , n4058 );
nand ( n4060 , n4059 , n3927 );
nand ( n4061 , n4055 , n4060 );
not ( n4062 , n2538 );
not ( n4063 , n501 );
not ( n4064 , n3197 );
or ( n4065 , n4063 , n4064 );
nand ( n4066 , n2846 , n2540 );
nand ( n4067 , n4065 , n4066 );
not ( n4068 , n4067 );
or ( n4069 , n4062 , n4068 );
nand ( n4070 , n3998 , n3553 );
nand ( n4071 , n4069 , n4070 );
xor ( n4072 , n4061 , n4071 );
not ( n4073 , n2134 );
not ( n4074 , n499 );
and ( n4075 , n456 , n470 );
not ( n4076 , n456 );
and ( n4077 , n4076 , n486 );
nor ( n4078 , n4075 , n4077 );
not ( n4079 , n4078 );
or ( n4080 , n4074 , n4079 );
or ( n4081 , n4078 , n499 );
nand ( n4082 , n4080 , n4081 );
not ( n4083 , n4082 );
or ( n4084 , n4073 , n4083 );
nand ( n4085 , n4009 , n2306 );
nand ( n4086 , n4084 , n4085 );
and ( n4087 , n4072 , n4086 );
and ( n4088 , n4061 , n4071 );
or ( n4089 , n4087 , n4088 );
xor ( n4090 , n3880 , n3899 );
xor ( n4091 , n4090 , n3929 );
xor ( n4092 , n4089 , n4091 );
xor ( n4093 , n4002 , n4013 );
xor ( n4094 , n4093 , n4033 );
and ( n4095 , n4092 , n4094 );
and ( n4096 , n4089 , n4091 );
or ( n4097 , n4095 , n4096 );
nor ( n4098 , n4047 , n4097 );
xor ( n4099 , n4089 , n4091 );
xor ( n4100 , n4099 , n4094 );
xor ( n4101 , n4022 , n4032 );
and ( n4102 , n3327 , n3403 );
not ( n4103 , n504 );
not ( n4104 , n4030 );
or ( n4105 , n4103 , n4104 );
and ( n4106 , n456 , n467 );
not ( n4107 , n456 );
and ( n4108 , n4107 , n483 );
nor ( n4109 , n4106 , n4108 );
and ( n4110 , n4109 , n2548 );
not ( n4111 , n4109 );
and ( n4112 , n4111 , n503 );
nor ( n4113 , n4110 , n4112 );
nand ( n4114 , n4113 , n3330 );
nand ( n4115 , n4105 , n4114 );
xor ( n4116 , n4102 , n4115 );
not ( n4117 , n2538 );
not ( n4118 , n501 );
not ( n4119 , n2687 );
or ( n4120 , n4118 , n4119 );
not ( n4121 , n3581 );
not ( n4122 , n3239 );
or ( n4123 , n4121 , n4122 );
nand ( n4124 , n4123 , n2540 );
nand ( n4125 , n4120 , n4124 );
not ( n4126 , n4125 );
or ( n4127 , n4117 , n4126 );
nand ( n4128 , n4067 , n2551 );
nand ( n4129 , n4127 , n4128 );
and ( n4130 , n4116 , n4129 );
and ( n4131 , n4102 , n4115 );
or ( n4132 , n4130 , n4131 );
xor ( n4133 , n4101 , n4132 );
xor ( n4134 , n4061 , n4071 );
xor ( n4135 , n4134 , n4086 );
and ( n4136 , n4133 , n4135 );
and ( n4137 , n4101 , n4132 );
or ( n4138 , n4136 , n4137 );
nor ( n4139 , n4100 , n4138 );
nor ( n4140 , n4098 , n4139 );
not ( n4141 , n4140 );
xor ( n4142 , n4101 , n4132 );
xor ( n4143 , n4142 , n4135 );
not ( n4144 , n2296 );
xor ( n4145 , n499 , n2761 );
not ( n4146 , n4145 );
or ( n4147 , n4144 , n4146 );
nand ( n4148 , n4082 , n2306 );
nand ( n4149 , n4147 , n4148 );
not ( n4150 , n2130 );
nand ( n4151 , n4150 , n2974 );
nand ( n4152 , n500 , n501 );
and ( n4153 , n4151 , n4152 , n499 );
not ( n4154 , n3330 );
and ( n4155 , n503 , n2400 );
not ( n4156 , n503 );
and ( n4157 , n4156 , n2846 );
or ( n4158 , n4155 , n4157 );
not ( n4159 , n4158 );
or ( n4160 , n4154 , n4159 );
nand ( n4161 , n4113 , n504 );
nand ( n4162 , n4160 , n4161 );
and ( n4163 , n4153 , n4162 );
xor ( n4164 , n4149 , n4163 );
xor ( n4165 , n4102 , n4115 );
xor ( n4166 , n4165 , n4129 );
and ( n4167 , n4164 , n4166 );
and ( n4168 , n4149 , n4163 );
or ( n4169 , n4167 , n4168 );
nor ( n4170 , n4143 , n4169 );
xor ( n4171 , n4149 , n4163 );
xor ( n4172 , n4171 , n4166 );
not ( n4173 , n2538 );
not ( n4174 , n501 );
not ( n4175 , n3252 );
or ( n4176 , n4174 , n4175 );
nand ( n4177 , n3259 , n2540 );
nand ( n4178 , n4176 , n4177 );
not ( n4179 , n4178 );
or ( n4180 , n4173 , n4179 );
nand ( n4181 , n4125 , n3553 );
nand ( n4182 , n4180 , n4181 );
not ( n4183 , n499 );
not ( n4184 , n3063 );
or ( n4185 , n4183 , n4184 );
not ( n4186 , n499 );
nand ( n4187 , n4186 , n2974 );
nand ( n4188 , n4185 , n4187 );
not ( n4189 , n4188 );
not ( n4190 , n2449 );
or ( n4191 , n4189 , n4190 );
nand ( n4192 , n4145 , n2306 );
nand ( n4193 , n4191 , n4192 );
xor ( n4194 , n4182 , n4193 );
xor ( n4195 , n4153 , n4162 );
and ( n4196 , n4194 , n4195 );
and ( n4197 , n4182 , n4193 );
or ( n4198 , n4196 , n4197 );
nor ( n4199 , n4172 , n4198 );
nor ( n4200 , n4170 , n4199 );
and ( n4201 , n3252 , n503 );
and ( n4202 , n4201 , n1939 );
not ( n4203 , n2687 );
not ( n4204 , n2699 );
not ( n4205 , n4204 );
or ( n4206 , n4203 , n4205 );
not ( n4207 , n504 );
nor ( n4208 , n4207 , n503 );
nand ( n4209 , n3241 , n4208 );
nand ( n4210 , n4206 , n4209 );
nor ( n4211 , n4202 , n4210 );
not ( n4212 , n4211 );
not ( n4213 , n502 );
nand ( n4214 , n4213 , n3063 );
and ( n4215 , n4214 , n503 );
not ( n4216 , n502 );
not ( n4217 , n3108 );
or ( n4218 , n4216 , n4217 );
nand ( n4219 , n4218 , n501 );
nor ( n4220 , n4215 , n4219 );
not ( n4221 , n4220 );
and ( n4222 , n4212 , n4221 );
and ( n4223 , n4220 , n4211 );
nor ( n4224 , n4222 , n4223 );
not ( n4225 , n501 );
not ( n4226 , n2920 );
or ( n4227 , n4225 , n4226 );
nand ( n4228 , n2761 , n2540 );
nand ( n4229 , n4227 , n4228 );
not ( n4230 , n4229 );
not ( n4231 , n4230 );
not ( n4232 , n2425 );
and ( n4233 , n4231 , n4232 );
not ( n4234 , n501 );
not ( n4235 , n3101 );
or ( n4236 , n4234 , n4235 );
nand ( n4237 , n3327 , n2540 );
nand ( n4238 , n4236 , n4237 );
and ( n4239 , n4238 , n2775 );
nor ( n4240 , n4233 , n4239 );
nand ( n4241 , n4224 , n4240 );
not ( n4242 , n4241 );
nor ( n4243 , n2974 , n2699 );
not ( n4244 , n4243 );
buf ( n4245 , n3268 );
not ( n4246 , n4245 );
or ( n4247 , n4244 , n4246 );
nand ( n4248 , n3063 , n2697 );
nand ( n4249 , n4247 , n4248 );
and ( n4250 , n3279 , n3553 );
nor ( n4251 , n4249 , n4250 );
not ( n4252 , n2548 );
not ( n4253 , n2640 );
or ( n4254 , n4252 , n4253 );
not ( n4255 , n4201 );
nand ( n4256 , n4254 , n4255 );
and ( n4257 , n4256 , n504 );
not ( n4258 , n4245 );
nor ( n4259 , n4258 , n2696 );
nor ( n4260 , n4257 , n4259 );
or ( n4261 , n4251 , n4260 );
nand ( n4262 , n4261 , C1 );
not ( n4263 , n4262 );
or ( n4264 , n4242 , n4263 );
not ( n4265 , n4224 );
not ( n4266 , n4240 );
nand ( n4267 , n4265 , n4266 );
nand ( n4268 , n4264 , n4267 );
not ( n4269 , n4268 );
and ( n4270 , n2128 , n3535 );
not ( n4271 , n2992 );
not ( n4272 , n4178 );
or ( n4273 , n4271 , n4272 );
nand ( n4274 , n4229 , n2538 );
nand ( n4275 , n4273 , n4274 );
xor ( n4276 , n4270 , n4275 );
not ( n4277 , n2697 );
not ( n4278 , n503 );
not ( n4279 , n2687 );
or ( n4280 , n4278 , n4279 );
not ( n4281 , n503 );
nand ( n4282 , n4281 , n3241 );
nand ( n4283 , n4280 , n4282 );
not ( n4284 , n4283 );
or ( n4285 , n4277 , n4284 );
nand ( n4286 , n504 , n4158 );
nand ( n4287 , n4285 , n4286 );
xor ( n4288 , n4276 , n4287 );
not ( n4289 , n4288 );
and ( n4290 , n3252 , n503 , n1939 );
or ( n4291 , n4290 , n4210 );
nand ( n4292 , n4291 , n4220 );
nand ( n4293 , n4289 , n4292 );
not ( n4294 , n4293 );
or ( n4295 , n4269 , n4294 );
buf ( n4296 , n4288 );
not ( n4297 , n4292 );
nand ( n4298 , n4296 , n4297 );
nand ( n4299 , n4295 , n4298 );
xor ( n4300 , n4182 , n4193 );
xor ( n4301 , n4300 , n4195 );
not ( n4302 , n4301 );
xor ( n4303 , n4270 , n4275 );
and ( n4304 , n4303 , n4287 );
and ( n4305 , n4270 , n4275 );
or ( n4306 , n4304 , n4305 );
not ( n4307 , n4306 );
nand ( n4308 , n4302 , n4307 );
nand ( n4309 , n4299 , n4308 );
buf ( n4310 , n4301 );
nand ( n4311 , n4310 , n4306 );
nand ( n4312 , n4172 , n4198 );
nand ( n4313 , n4309 , n4311 , n4312 );
nand ( n4314 , n4200 , n4313 );
and ( n4315 , n4100 , n4138 );
and ( n4316 , n4143 , n4169 );
nor ( n4317 , n4315 , n4316 );
nand ( n4318 , n4314 , n4317 );
not ( n4319 , n4318 );
or ( n4320 , n4141 , n4319 );
buf ( n4321 , n4047 );
nand ( n4322 , n4321 , n4097 );
nand ( n4323 , n4320 , n4322 );
not ( n4324 , n4323 );
or ( n4325 , n4045 , n4324 );
buf ( n4326 , n3990 );
nand ( n4327 , n4326 , n4042 );
nand ( n4328 , n4325 , n4327 );
xor ( n4329 , n3757 , n3767 );
xor ( n4330 , n4329 , n3769 );
xor ( n4331 , n3976 , n3981 );
and ( n4332 , n4331 , n3987 );
and ( n4333 , n3976 , n3981 );
or ( n4334 , n4332 , n4333 );
xor ( n4335 , n3816 , n3822 );
and ( n4336 , n4335 , n3838 );
and ( n4337 , n3816 , n3822 );
or ( n4338 , n4336 , n4337 );
xor ( n4339 , n4334 , n4338 );
xor ( n4340 , n3704 , n3719 );
xor ( n4341 , n4340 , n3730 );
xor ( n4342 , n4339 , n4341 );
xor ( n4343 , n4330 , n4342 );
xor ( n4344 , n3937 , n3966 );
and ( n4345 , n4344 , n3988 );
and ( n4346 , n3937 , n3966 );
or ( n4347 , n4345 , n4346 );
xor ( n4348 , n4343 , n4347 );
not ( n4349 , n4348 );
xor ( n4350 , n3839 , n3935 );
and ( n4351 , n4350 , n3989 );
and ( n4352 , n3839 , n3935 );
or ( n4353 , n4351 , n4352 );
not ( n4354 , n4353 );
and ( n4355 , n4349 , n4354 );
xor ( n4356 , n3677 , n3692 );
xor ( n4357 , n4356 , n3733 );
xor ( n4358 , n4334 , n4338 );
and ( n4359 , n4358 , n4341 );
and ( n4360 , n4334 , n4338 );
or ( n4361 , n4359 , n4360 );
xor ( n4362 , n4357 , n4361 );
xor ( n4363 , n3745 , n3747 );
xor ( n4364 , n4363 , n3772 );
xor ( n4365 , n4362 , n4364 );
xor ( n4366 , n4330 , n4342 );
and ( n4367 , n4366 , n4347 );
and ( n4368 , n4330 , n4342 );
or ( n4369 , n4367 , n4368 );
nor ( n4370 , n4365 , n4369 );
nor ( n4371 , n4355 , n4370 );
xor ( n4372 , n3743 , n3775 );
xor ( n4373 , n4372 , n3778 );
not ( n4374 , n4373 );
xor ( n4375 , n4357 , n4361 );
and ( n4376 , n4375 , n4364 );
and ( n4377 , n4357 , n4361 );
or ( n4378 , n4376 , n4377 );
not ( n4379 , n4378 );
nand ( n4380 , n4374 , n4379 );
nand ( n4381 , n4328 , n4371 , n4380 );
nand ( n4382 , n4373 , n4378 );
not ( n4383 , n4382 );
nand ( n4384 , n4348 , n4353 );
not ( n4385 , n4384 );
nand ( n4386 , n4369 , n4365 );
not ( n4387 , n4386 );
or ( n4388 , n4385 , n4387 );
not ( n4389 , n4365 );
not ( n4390 , n4369 );
nand ( n4391 , n4389 , n4390 );
nand ( n4392 , n4388 , n4391 );
not ( n4393 , n4392 );
or ( n4394 , n4383 , n4393 );
not ( n4395 , n4373 );
nand ( n4396 , n4395 , n4379 );
nand ( n4397 , n4394 , n4396 );
nand ( n4398 , n4381 , n4397 );
not ( n4399 , n3786 );
nand ( n4400 , n4399 , n3792 );
nand ( n4401 , n3741 , n3782 );
nand ( n4402 , n4398 , n4400 , n4401 );
nand ( n4403 , n3803 , n4402 );
nand ( n4404 , n3235 , n3657 , n4403 );
not ( n4405 , n3053 );
not ( n4406 , n3049 );
and ( n4407 , n4405 , n4406 );
nand ( n4408 , n3020 , n3046 );
or ( n4409 , n4407 , n4408 );
not ( n4410 , n4405 );
not ( n4411 , n4406 );
nand ( n4412 , n4410 , n4411 );
nand ( n4413 , n4409 , n4412 );
not ( n4414 , n4413 );
not ( n4415 , n3020 );
not ( n4416 , n3046 );
and ( n4417 , n4415 , n4416 );
nor ( n4418 , n4417 , n3054 );
and ( n4419 , n3057 , n3231 );
nand ( n4420 , n4418 , n4419 );
nor ( n4421 , n3057 , n3231 );
not ( n4422 , n4421 );
nor ( n4423 , n3645 , n3632 );
nand ( n4424 , n3649 , n3654 );
or ( n4425 , n4423 , n4424 );
nand ( n4426 , n3632 , n3645 );
nand ( n4427 , n4425 , n4426 );
nand ( n4428 , n4422 , n3055 , n4427 );
nand ( n4429 , n4404 , n4414 , n4420 , n4428 );
xor ( n4430 , n2716 , n4429 );
nand ( n4431 , n4430 , n455 );
buf ( n4432 , n4100 );
nor ( n4433 , n4432 , n4138 );
not ( n4434 , n4433 );
buf ( n4435 , n4318 );
nand ( n4436 , n4434 , n4435 );
or ( n4437 , n4321 , n4097 );
nand ( n4438 , n4437 , n4322 );
xor ( n4439 , n4436 , n4438 );
nand ( n4440 , n4439 , n455 );
not ( n4441 , n454 );
and ( n4442 , n539 , n540 );
and ( n4443 , n540 , n541 );
not ( n4444 , n540 );
not ( n4445 , n541 );
and ( n4446 , n4444 , n4445 );
nor ( n4447 , n4443 , n4446 );
nor ( n4448 , n539 , n540 );
nor ( n4449 , n4442 , n4447 , n4448 );
buf ( n4450 , n4449 );
not ( n4451 , n4450 );
not ( n4452 , n539 );
buf ( n4453 , n4401 );
not ( n4454 , n4453 );
nand ( n4455 , n4381 , n4397 );
buf ( n4456 , n4455 );
not ( n4457 , n4456 );
or ( n4458 , n4454 , n4457 );
nand ( n4459 , n3740 , n3781 );
nand ( n4460 , n4458 , n4459 );
not ( n4461 , n4400 );
nand ( n4462 , n3786 , n3791 );
not ( n4463 , n4462 );
nor ( n4464 , n4461 , n4463 );
not ( n4465 , n455 );
nor ( n4466 , n4464 , n4465 );
and ( n4467 , n4460 , n4466 );
not ( n4468 , n4460 );
and ( n4469 , n455 , n4400 , n4462 );
and ( n4470 , n4468 , n4469 );
nor ( n4471 , n4467 , n4470 );
nand ( n4472 , n4471 , n1985 );
buf ( n4473 , n4472 );
not ( n4474 , n4473 );
not ( n4475 , n4474 );
or ( n4476 , n4452 , n4475 );
not ( n4477 , n539 );
nand ( n4478 , n4473 , n4477 );
nand ( n4479 , n4476 , n4478 );
not ( n4480 , n4479 );
or ( n4481 , n4451 , n4480 );
nand ( n4482 , n4462 , n4459 );
not ( n4483 , n4482 );
not ( n4484 , n4400 );
or ( n4485 , n4483 , n4484 );
nand ( n4486 , n4485 , n4402 );
nand ( n4487 , n3627 , n3522 );
buf ( n4488 , n4487 );
nor ( n4489 , n3522 , n3627 );
not ( n4490 , n4489 );
and ( n4491 , n4488 , n4490 );
and ( n4492 , n4486 , n4491 );
not ( n4493 , n455 );
nor ( n4494 , n4492 , n4493 );
not ( n4495 , n4494 );
not ( n4496 , n4486 );
nand ( n4497 , n3630 , n4488 );
nand ( n4498 , n4496 , n4497 );
not ( n4499 , n4498 );
or ( n4500 , n4495 , n4499 );
not ( n4501 , n1982 );
not ( n4502 , n1828 );
or ( n4503 , n4501 , n4502 );
nand ( n4504 , n4503 , n1979 );
not ( n4505 , n1936 );
nand ( n4506 , n4505 , n1955 );
not ( n4507 , n4506 );
not ( n4508 , n1927 );
or ( n4509 , n4507 , n4508 );
not ( n4510 , n1955 );
nand ( n4511 , n4510 , n1936 );
nand ( n4512 , n4509 , n4511 );
not ( n4513 , n1954 );
not ( n4514 , n1863 );
not ( n4515 , n1849 );
or ( n4516 , n4514 , n4515 );
or ( n4517 , n1849 , n1863 );
nand ( n4518 , n4517 , n1838 );
nand ( n4519 , n4516 , n4518 );
xor ( n4520 , n4513 , n4519 );
xor ( n4521 , n1881 , n1891 );
and ( n4522 , n4521 , n1901 );
and ( n4523 , n1881 , n1891 );
or ( n4524 , n4522 , n4523 );
xor ( n4525 , n4520 , n4524 );
xor ( n4526 , n4512 , n4525 );
or ( n4527 , n1902 , n1869 );
nand ( n4528 , n4527 , n1832 );
nand ( n4529 , n1902 , n1869 );
nand ( n4530 , n4528 , n4529 );
xor ( n4531 , n4526 , n4530 );
not ( n4532 , n4531 );
not ( n4533 , n1921 );
not ( n4534 , n4533 );
not ( n4535 , n1959 );
not ( n4536 , n4535 );
or ( n4537 , n4534 , n4536 );
not ( n4538 , n1921 );
not ( n4539 , n1959 );
or ( n4540 , n4538 , n4539 );
nand ( n4541 , n4540 , n1964 );
nand ( n4542 , n4537 , n4541 );
not ( n4543 , n4542 );
not ( n4544 , n4543 );
not ( n4545 , n1879 );
not ( n4546 , n1586 );
or ( n4547 , n4545 , n4546 );
xor ( n4548 , n514 , n493 );
nand ( n4549 , n814 , n4548 );
nand ( n4550 , n4547 , n4549 );
not ( n4551 , n1899 );
not ( n4552 , n975 );
or ( n4553 , n4551 , n4552 );
and ( n4554 , n508 , n499 );
not ( n4555 , n508 );
not ( n4556 , n499 );
and ( n4557 , n4555 , n4556 );
nor ( n4558 , n4554 , n4557 );
nand ( n4559 , n749 , n4558 );
nand ( n4560 , n4553 , n4559 );
xor ( n4561 , n4550 , n4560 );
not ( n4562 , n1934 );
nor ( n4563 , n1929 , n1565 );
not ( n4564 , n4563 );
or ( n4565 , n4562 , n4564 );
xor ( n4566 , n516 , n491 );
nand ( n4567 , n1933 , n4566 );
nand ( n4568 , n4565 , n4567 );
xor ( n4569 , n4561 , n4568 );
not ( n4570 , n1847 );
not ( n4571 , n736 );
or ( n4572 , n4570 , n4571 );
xor ( n4573 , n506 , n501 );
nand ( n4574 , n4573 , n694 );
nand ( n4575 , n4572 , n4574 );
nand ( n4576 , n520 , n489 );
not ( n4577 , n683 );
not ( n4578 , n1943 );
or ( n4579 , n4577 , n4578 );
nand ( n4580 , n4579 , n699 );
xnor ( n4581 , n4576 , n4580 );
xor ( n4582 , n4575 , n4581 );
not ( n4583 , n4582 );
and ( n4584 , n4569 , n4583 );
not ( n4585 , n4569 );
and ( n4586 , n4585 , n4582 );
nor ( n4587 , n4584 , n4586 );
not ( n4588 , n1861 );
not ( n4589 , n1856 );
nor ( n4590 , n4589 , n1760 );
not ( n4591 , n4590 );
or ( n4592 , n4588 , n4591 );
xor ( n4593 , n518 , n489 );
nand ( n4594 , n1859 , n4593 );
nand ( n4595 , n4592 , n4594 );
not ( n4596 , n1885 );
not ( n4597 , n859 );
or ( n4598 , n4596 , n4597 );
xor ( n4599 , n512 , n495 );
nand ( n4600 , n867 , n4599 );
nand ( n4601 , n4598 , n4600 );
xor ( n4602 , n4595 , n4601 );
not ( n4603 , n1836 );
not ( n4604 , n963 );
or ( n4605 , n4603 , n4604 );
xor ( n4606 , n510 , n497 );
nand ( n4607 , n836 , n4606 );
nand ( n4608 , n4605 , n4607 );
xor ( n4609 , n4602 , n4608 );
buf ( n4610 , n4609 );
and ( n4611 , n4587 , n4610 );
not ( n4612 , n4587 );
not ( n4613 , n4610 );
and ( n4614 , n4612 , n4613 );
nor ( n4615 , n4611 , n4614 );
not ( n4616 , n4615 );
not ( n4617 , n4616 );
or ( n4618 , n4544 , n4617 );
nand ( n4619 , n4542 , n4615 );
nand ( n4620 , n4618 , n4619 );
not ( n4621 , n4620 );
not ( n4622 , n4621 );
or ( n4623 , n4532 , n4622 );
not ( n4624 , n4531 );
nand ( n4625 , n4620 , n4624 );
nand ( n4626 , n4623 , n4625 );
not ( n4627 , n4626 );
not ( n4628 , n1903 );
not ( n4629 , n1968 );
or ( n4630 , n4628 , n4629 );
not ( n4631 , n1965 );
not ( n4632 , n1903 );
not ( n4633 , n4632 );
or ( n4634 , n4631 , n4633 );
nand ( n4635 , n4634 , n1912 );
nand ( n4636 , n4630 , n4635 );
not ( n4637 , n4636 );
not ( n4638 , n4637 );
and ( n4639 , n4627 , n4638 );
not ( n4640 , n4627 );
and ( n4641 , n4640 , n4637 );
nor ( n4642 , n4639 , n4641 );
not ( n4643 , n4642 );
and ( n4644 , n4504 , n4643 );
not ( n4645 , n4504 );
and ( n4646 , n4645 , n4642 );
nor ( n4647 , n4644 , n4646 );
nand ( n4648 , n4647 , n793 );
nand ( n4649 , n4500 , n4648 );
not ( n4650 , n4649 );
not ( n4651 , n4650 );
not ( n4652 , n4651 );
not ( n4653 , n4477 );
and ( n4654 , n4652 , n4653 );
buf ( n4655 , n4649 );
and ( n4656 , n4655 , n4477 );
nor ( n4657 , n4654 , n4656 );
not ( n4658 , n4657 );
buf ( n4659 , n4447 );
buf ( n4660 , n4659 );
nand ( n4661 , n4658 , n4660 );
nand ( n4662 , n4481 , n4661 );
xnor ( n4663 , n543 , n544 );
not ( n4664 , n544 );
or ( n4665 , n4664 , n545 );
not ( n4666 , n545 );
or ( n4667 , n4666 , n544 );
nand ( n4668 , n4665 , n4667 );
buf ( n4669 , n4668 );
nor ( n4670 , n4663 , n4669 );
buf ( n4671 , n4670 );
not ( n4672 , n4671 );
not ( n4673 , n543 );
xor ( n4674 , n507 , n499 );
not ( n4675 , n4674 );
not ( n4676 , n975 );
or ( n4677 , n4675 , n4676 );
and ( n4678 , n506 , n499 );
not ( n4679 , n506 );
and ( n4680 , n4679 , n2158 );
nor ( n4681 , n4678 , n4680 );
nand ( n4682 , n1027 , n4681 );
nand ( n4683 , n4677 , n4682 );
nand ( n4684 , n518 , n489 );
not ( n4685 , n4684 );
and ( n4686 , n4683 , n4685 );
not ( n4687 , n4683 );
and ( n4688 , n4687 , n4684 );
nor ( n4689 , n4686 , n4688 );
xor ( n4690 , n511 , n495 );
not ( n4691 , n4690 );
not ( n4692 , n1361 );
not ( n4693 , n4692 );
or ( n4694 , n4691 , n4693 );
xor ( n4695 , n510 , n495 );
nand ( n4696 , n867 , n4695 );
nand ( n4697 , n4694 , n4696 );
xor ( n4698 , n4689 , n4697 );
xor ( n4699 , n505 , n501 );
not ( n4700 , n4699 );
not ( n4701 , n736 );
or ( n4702 , n4700 , n4701 );
nand ( n4703 , n694 , n501 );
nand ( n4704 , n4702 , n4703 );
xor ( n4705 , n517 , n489 );
not ( n4706 , n4705 );
not ( n4707 , n4590 );
or ( n4708 , n4706 , n4707 );
xor ( n4709 , n516 , n489 );
nand ( n4710 , n1859 , n4709 );
nand ( n4711 , n4708 , n4710 );
and ( n4712 , n4704 , n4711 );
not ( n4713 , n4704 );
not ( n4714 , n4711 );
and ( n4715 , n4713 , n4714 );
or ( n4716 , n4712 , n4715 );
not ( n4717 , n4606 );
not ( n4718 , n963 );
or ( n4719 , n4717 , n4718 );
xor ( n4720 , n509 , n497 );
nand ( n4721 , n836 , n4720 );
nand ( n4722 , n4719 , n4721 );
not ( n4723 , n4722 );
and ( n4724 , n4716 , n4723 );
not ( n4725 , n4716 );
and ( n4726 , n4725 , n4722 );
nor ( n4727 , n4724 , n4726 );
not ( n4728 , n4727 );
xor ( n4729 , n4698 , n4728 );
not ( n4730 , n4580 );
nand ( n4731 , n4730 , n4576 );
not ( n4732 , n4731 );
not ( n4733 , n4575 );
or ( n4734 , n4732 , n4733 );
not ( n4735 , n4576 );
nand ( n4736 , n4735 , n4580 );
nand ( n4737 , n4734 , n4736 );
xor ( n4738 , n4550 , n4560 );
and ( n4739 , n4738 , n4568 );
and ( n4740 , n4550 , n4560 );
or ( n4741 , n4739 , n4740 );
xor ( n4742 , n4737 , n4741 );
xor ( n4743 , n4595 , n4601 );
and ( n4744 , n4743 , n4608 );
and ( n4745 , n4595 , n4601 );
or ( n4746 , n4744 , n4745 );
and ( n4747 , n4742 , n4746 );
and ( n4748 , n4737 , n4741 );
or ( n4749 , n4747 , n4748 );
xnor ( n4750 , n4729 , n4749 );
not ( n4751 , n4722 );
not ( n4752 , n1586 );
not ( n4753 , n4548 );
or ( n4754 , n4752 , n4753 );
xor ( n4755 , n513 , n493 );
nand ( n4756 , n814 , n4755 );
nand ( n4757 , n4754 , n4756 );
not ( n4758 , n4757 );
not ( n4759 , n4566 );
not ( n4760 , n1930 );
or ( n4761 , n4759 , n4760 );
and ( n4762 , n515 , n1993 );
not ( n4763 , n515 );
and ( n4764 , n4763 , n491 );
or ( n4765 , n4762 , n4764 );
nand ( n4766 , n1933 , n4765 );
nand ( n4767 , n4761 , n4766 );
not ( n4768 , n4767 );
not ( n4769 , n4768 );
or ( n4770 , n4758 , n4769 );
or ( n4771 , n4768 , n4757 );
nand ( n4772 , n4770 , n4771 );
not ( n4773 , n4772 );
or ( n4774 , n4751 , n4773 );
or ( n4775 , n4772 , n4722 );
nand ( n4776 , n4774 , n4775 );
not ( n4777 , n4776 );
xor ( n4778 , n4737 , n4741 );
xor ( n4779 , n4778 , n4746 );
not ( n4780 , n4779 );
or ( n4781 , n4777 , n4780 );
or ( n4782 , n4776 , n4779 );
not ( n4783 , n4582 );
not ( n4784 , n4569 );
or ( n4785 , n4783 , n4784 );
or ( n4786 , n4582 , n4569 );
nand ( n4787 , n4786 , n4609 );
nand ( n4788 , n4785 , n4787 );
nand ( n4789 , n4782 , n4788 );
nand ( n4790 , n4781 , n4789 );
not ( n4791 , n4790 );
xor ( n4792 , n4750 , n4791 );
not ( n4793 , n4767 );
not ( n4794 , n4757 );
or ( n4795 , n4793 , n4794 );
not ( n4796 , n4768 );
not ( n4797 , n4757 );
not ( n4798 , n4797 );
or ( n4799 , n4796 , n4798 );
nand ( n4800 , n4799 , n4723 );
nand ( n4801 , n4795 , n4800 );
not ( n4802 , n4801 );
not ( n4803 , n1933 );
xor ( n4804 , n514 , n491 );
not ( n4805 , n4804 );
or ( n4806 , n4803 , n4805 );
xnor ( n4807 , n491 , n492 );
not ( n4808 , n4807 );
not ( n4809 , n1565 );
nand ( n4810 , n4808 , n4765 , n4809 );
nand ( n4811 , n4806 , n4810 );
not ( n4812 , n4811 );
not ( n4813 , n4755 );
not ( n4814 , n1481 );
or ( n4815 , n4813 , n4814 );
xor ( n4816 , n512 , n493 );
nand ( n4817 , n814 , n4816 );
nand ( n4818 , n4815 , n4817 );
not ( n4819 , n4818 );
and ( n4820 , n4812 , n4819 );
not ( n4821 , n4812 );
and ( n4822 , n4821 , n4818 );
nor ( n4823 , n4820 , n4822 );
not ( n4824 , n4720 );
not ( n4825 , n963 );
or ( n4826 , n4824 , n4825 );
xor ( n4827 , n508 , n497 );
nand ( n4828 , n836 , n4827 );
nand ( n4829 , n4826 , n4828 );
xor ( n4830 , n4823 , n4829 );
not ( n4831 , n4830 );
or ( n4832 , n4802 , n4831 );
not ( n4833 , n4830 );
not ( n4834 , n4801 );
nand ( n4835 , n4833 , n4834 );
nand ( n4836 , n4832 , n4835 );
nand ( n4837 , n519 , n489 );
not ( n4838 , n4837 );
not ( n4839 , n503 );
not ( n4840 , n683 );
or ( n4841 , n4839 , n4840 );
nand ( n4842 , n4841 , n699 );
not ( n4843 , n4842 );
or ( n4844 , n4838 , n4843 );
not ( n4845 , n4593 );
not ( n4846 , n4590 );
or ( n4847 , n4845 , n4846 );
nand ( n4848 , n1859 , n4705 );
nand ( n4849 , n4847 , n4848 );
nand ( n4850 , n4844 , n4849 );
not ( n4851 , n4842 );
not ( n4852 , n4837 );
nand ( n4853 , n4851 , n4852 );
nand ( n4854 , n4850 , n4853 );
not ( n4855 , n4854 );
not ( n4856 , n4599 );
not ( n4857 , n859 );
or ( n4858 , n4856 , n4857 );
nand ( n4859 , n867 , n4690 );
nand ( n4860 , n4858 , n4859 );
not ( n4861 , n4860 );
not ( n4862 , n4674 );
not ( n4863 , n749 );
or ( n4864 , n4862 , n4863 );
nand ( n4865 , n934 , n938 , n4558 , n937 );
nand ( n4866 , n4864 , n4865 );
not ( n4867 , n4866 );
or ( n4868 , n4861 , n4867 );
not ( n4869 , n4860 );
not ( n4870 , n4869 );
not ( n4871 , n4866 );
not ( n4872 , n4871 );
or ( n4873 , n4870 , n4872 );
not ( n4874 , n4573 );
not ( n4875 , n736 );
or ( n4876 , n4874 , n4875 );
nand ( n4877 , n694 , n4699 );
nand ( n4878 , n4876 , n4877 );
nand ( n4879 , n4873 , n4878 );
nand ( n4880 , n4868 , n4879 );
not ( n4881 , n4880 );
not ( n4882 , n4881 );
or ( n4883 , n4855 , n4882 );
not ( n4884 , n4854 );
nand ( n4885 , n4884 , n4880 );
nand ( n4886 , n4883 , n4885 );
and ( n4887 , n4836 , n4886 );
not ( n4888 , n4836 );
not ( n4889 , n4886 );
and ( n4890 , n4888 , n4889 );
nor ( n4891 , n4887 , n4890 );
xor ( n4892 , n4852 , n4842 );
xnor ( n4893 , n4892 , n4849 );
not ( n4894 , n4871 );
not ( n4895 , n4869 );
nand ( n4896 , n4894 , n4895 , n4878 );
not ( n4897 , n4878 );
nand ( n4898 , n4895 , n4897 , n4871 );
not ( n4899 , n4871 );
not ( n4900 , n4860 );
nand ( n4901 , n4899 , n4900 , n4897 );
nand ( n4902 , n4900 , n4871 , n4878 );
nand ( n4903 , n4896 , n4898 , n4901 , n4902 );
or ( n4904 , n4893 , n4903 );
not ( n4905 , n4904 );
xor ( n4906 , n4513 , n4519 );
and ( n4907 , n4906 , n4524 );
and ( n4908 , n4513 , n4519 );
or ( n4909 , n4907 , n4908 );
not ( n4910 , n4909 );
or ( n4911 , n4905 , n4910 );
nand ( n4912 , n4893 , n4903 );
nand ( n4913 , n4911 , n4912 );
and ( n4914 , n4891 , n4913 );
not ( n4915 , n4891 );
not ( n4916 , n4913 );
and ( n4917 , n4915 , n4916 );
nor ( n4918 , n4914 , n4917 );
xor ( n4919 , n4792 , n4918 );
or ( n4920 , n4893 , n4903 );
nand ( n4921 , n4920 , n4912 );
not ( n4922 , n4921 );
not ( n4923 , n4909 );
and ( n4924 , n4922 , n4923 );
and ( n4925 , n4909 , n4921 );
nor ( n4926 , n4924 , n4925 );
not ( n4927 , n4926 );
not ( n4928 , n4927 );
xor ( n4929 , n4776 , n4788 );
xnor ( n4930 , n4929 , n4779 );
not ( n4931 , n4930 );
not ( n4932 , n4931 );
or ( n4933 , n4928 , n4932 );
not ( n4934 , n4926 );
not ( n4935 , n4930 );
or ( n4936 , n4934 , n4935 );
xor ( n4937 , n4512 , n4525 );
and ( n4938 , n4937 , n4530 );
and ( n4939 , n4512 , n4525 );
or ( n4940 , n4938 , n4939 );
buf ( n4941 , n4940 );
nand ( n4942 , n4936 , n4941 );
nand ( n4943 , n4933 , n4942 );
not ( n4944 , n4943 );
nand ( n4945 , n4919 , n4944 );
not ( n4946 , n4945 );
not ( n4947 , n4926 );
not ( n4948 , n4940 );
or ( n4949 , n4947 , n4948 );
not ( n4950 , n4940 );
nand ( n4951 , n4950 , n4927 );
nand ( n4952 , n4949 , n4951 );
or ( n4953 , n4931 , n4952 );
nand ( n4954 , n4952 , n4931 );
nand ( n4955 , n4953 , n4954 );
not ( n4956 , n4624 );
buf ( n4957 , n4615 );
not ( n4958 , n4957 );
and ( n4959 , n4956 , n4958 );
nand ( n4960 , n4624 , n4957 );
buf ( n4961 , n4542 );
and ( n4962 , n4960 , n4961 );
nor ( n4963 , n4959 , n4962 );
nand ( n4964 , n4955 , n4963 );
not ( n4965 , n4964 );
not ( n4966 , n1980 );
not ( n4967 , n1981 );
or ( n4968 , n4966 , n4967 );
or ( n4969 , n4620 , n4624 );
nand ( n4970 , n4969 , n4625 );
not ( n4971 , n4970 );
not ( n4972 , n4636 );
nand ( n4973 , n4971 , n4972 );
nand ( n4974 , n4968 , n4973 );
nor ( n4975 , n4965 , n4974 );
not ( n4976 , n4975 );
not ( n4977 , n1828 );
or ( n4978 , n4976 , n4977 );
or ( n4979 , n4955 , n4963 );
nand ( n4980 , n4627 , n4972 );
not ( n4981 , n4636 );
not ( n4982 , n4970 );
or ( n4983 , n4981 , n4982 );
nand ( n4984 , n4983 , n1978 );
nand ( n4985 , n4964 , n4980 , n4984 );
nand ( n4986 , n4979 , n4985 );
not ( n4987 , n4986 );
nand ( n4988 , n4978 , n4987 );
not ( n4989 , n4988 );
or ( n4990 , n4946 , n4989 );
not ( n4991 , n4919 );
nand ( n4992 , n4991 , n4943 );
nand ( n4993 , n4990 , n4992 );
not ( n4994 , n455 );
not ( n4995 , n4994 );
not ( n4996 , n4711 );
nand ( n4997 , n4996 , n4704 );
not ( n4998 , n4997 );
not ( n4999 , n4722 );
or ( n5000 , n4998 , n4999 );
not ( n5001 , n4704 );
nand ( n5002 , n5001 , n4711 );
nand ( n5003 , n5000 , n5002 );
not ( n5004 , n4816 );
not ( n5005 , n1586 );
or ( n5006 , n5004 , n5005 );
and ( n5007 , n493 , n1579 );
not ( n5008 , n493 );
and ( n5009 , n5008 , n511 );
or ( n5010 , n5007 , n5009 );
nand ( n5011 , n814 , n5010 );
nand ( n5012 , n5006 , n5011 );
nand ( n5013 , n517 , n489 );
xor ( n5014 , n5012 , n5013 );
not ( n5015 , n836 );
xor ( n5016 , n497 , n507 );
not ( n5017 , n5016 );
or ( n5018 , n5015 , n5017 );
nand ( n5019 , n4827 , n963 );
nand ( n5020 , n5018 , n5019 );
xnor ( n5021 , n5014 , n5020 );
xor ( n5022 , n5003 , n5021 );
not ( n5023 , n4804 );
not ( n5024 , n1930 );
or ( n5025 , n5023 , n5024 );
xor ( n5026 , n491 , n513 );
nand ( n5027 , n1933 , n5026 );
nand ( n5028 , n5025 , n5027 );
not ( n5029 , n4709 );
not ( n5030 , n4590 );
or ( n5031 , n5029 , n5030 );
xor ( n5032 , n515 , n489 );
nand ( n5033 , n1859 , n5032 );
nand ( n5034 , n5031 , n5033 );
xnor ( n5035 , n5028 , n5034 );
and ( n5036 , n5035 , n5001 );
not ( n5037 , n5035 );
and ( n5038 , n5037 , n4704 );
nor ( n5039 , n5036 , n5038 );
xor ( n5040 , n5022 , n5039 );
xnor ( n5041 , n4886 , n4830 );
nand ( n5042 , n5041 , n4834 );
not ( n5043 , n5042 );
not ( n5044 , n4913 );
or ( n5045 , n5043 , n5044 );
not ( n5046 , n5041 );
nand ( n5047 , n5046 , n4801 );
nand ( n5048 , n5045 , n5047 );
xor ( n5049 , n5040 , n5048 );
not ( n5050 , n4884 );
not ( n5051 , n4881 );
or ( n5052 , n5050 , n5051 );
nand ( n5053 , n5052 , n4830 );
nand ( n5054 , n4880 , n4854 );
nand ( n5055 , n5053 , n5054 );
not ( n5056 , n4829 );
nand ( n5057 , n4819 , n4812 );
not ( n5058 , n5057 );
or ( n5059 , n5056 , n5058 );
nand ( n5060 , n4811 , n4818 );
nand ( n5061 , n5059 , n5060 );
or ( n5062 , n4683 , n4685 );
nand ( n5063 , n5062 , n4697 );
nand ( n5064 , n4683 , n4685 );
nand ( n5065 , n5063 , n5064 );
not ( n5066 , n5065 );
and ( n5067 , n5061 , n5066 );
not ( n5068 , n5061 );
and ( n5069 , n5068 , n5065 );
or ( n5070 , n5067 , n5069 );
not ( n5071 , n1027 );
and ( n5072 , n499 , n505 );
not ( n5073 , n499 );
not ( n5074 , n505 );
and ( n5075 , n5073 , n5074 );
nor ( n5076 , n5072 , n5075 );
not ( n5077 , n5076 );
or ( n5078 , n5071 , n5077 );
nand ( n5079 , n4681 , n973 , n1688 );
nand ( n5080 , n5078 , n5079 );
not ( n5081 , n5080 );
not ( n5082 , n734 );
nand ( n5083 , n5082 , n801 , n802 );
nand ( n5084 , n5083 , n501 );
and ( n5085 , n5081 , n5084 );
not ( n5086 , n5081 );
not ( n5087 , n5084 );
and ( n5088 , n5086 , n5087 );
nor ( n5089 , n5085 , n5088 );
not ( n5090 , n4695 );
not ( n5091 , n859 );
or ( n5092 , n5090 , n5091 );
xor ( n5093 , n509 , n495 );
nand ( n5094 , n867 , n5093 );
nand ( n5095 , n5092 , n5094 );
xor ( n5096 , n5089 , n5095 );
not ( n5097 , n5096 );
and ( n5098 , n5070 , n5097 );
not ( n5099 , n5070 );
and ( n5100 , n5099 , n5096 );
nor ( n5101 , n5098 , n5100 );
xor ( n5102 , n5055 , n5101 );
not ( n5103 , n4698 );
nand ( n5104 , n4727 , n5103 );
not ( n5105 , n5104 );
not ( n5106 , n4749 );
or ( n5107 , n5105 , n5106 );
not ( n5108 , n5103 );
nand ( n5109 , n5108 , n4728 );
nand ( n5110 , n5107 , n5109 );
xor ( n5111 , n5102 , n5110 );
xnor ( n5112 , n5049 , n5111 );
not ( n5113 , n5112 );
xor ( n5114 , n4750 , n4791 );
and ( n5115 , n5114 , n4918 );
and ( n5116 , n4750 , n4791 );
or ( n5117 , n5115 , n5116 );
not ( n5118 , n5117 );
xnor ( n5119 , n5113 , n5118 );
nor ( n5120 , n4995 , n5119 );
and ( n5121 , n4993 , n5120 );
not ( n5122 , n4993 );
and ( n5123 , n5119 , n4493 );
and ( n5124 , n5122 , n5123 );
nor ( n5125 , n5121 , n5124 );
not ( n5126 , n4403 );
not ( n5127 , n3657 );
or ( n5128 , n5126 , n5127 );
not ( n5129 , n4427 );
nand ( n5130 , n5128 , n5129 );
not ( n5131 , n4419 );
and ( n5132 , n3233 , n5131 , n455 );
and ( n5133 , n5130 , n5132 );
not ( n5134 , n5130 );
not ( n5135 , n4419 );
nand ( n5136 , n5135 , n3233 );
not ( n5137 , n5136 );
nor ( n5138 , n5137 , n4493 );
and ( n5139 , n5134 , n5138 );
nor ( n5140 , n5133 , n5139 );
nand ( n5141 , n5125 , n5140 );
not ( n5142 , n5141 );
or ( n5143 , n4673 , n5142 );
nand ( n5144 , n5125 , n5140 );
not ( n5145 , n5144 );
not ( n5146 , n543 );
nand ( n5147 , n5145 , n5146 );
nand ( n5148 , n5143 , n5147 );
not ( n5149 , n5148 );
or ( n5150 , n4672 , n5149 );
not ( n5151 , n543 );
nand ( n5152 , n5112 , n5117 );
nand ( n5153 , n5152 , n4945 );
not ( n5154 , n5153 );
not ( n5155 , n5154 );
and ( n5156 , n1828 , n4975 );
not ( n5157 , n5156 );
or ( n5158 , n5155 , n5157 );
buf ( n5159 , n4986 );
and ( n5160 , n5159 , n5154 );
not ( n5161 , n5118 );
not ( n5162 , n5113 );
or ( n5163 , n5161 , n5162 );
not ( n5164 , n5117 );
not ( n5165 , n5112 );
or ( n5166 , n5164 , n5165 );
nor ( n5167 , n4919 , n4944 );
nand ( n5168 , n5166 , n5167 );
nand ( n5169 , n5163 , n5168 );
nor ( n5170 , n5160 , n5169 );
nand ( n5171 , n5158 , n5170 );
not ( n5172 , n5171 );
xor ( n5173 , n5003 , n5021 );
and ( n5174 , n5173 , n5039 );
and ( n5175 , n5003 , n5021 );
or ( n5176 , n5174 , n5175 );
not ( n5177 , n5076 );
not ( n5178 , n1062 );
or ( n5179 , n5177 , n5178 );
nand ( n5180 , n978 , n499 );
nand ( n5181 , n5179 , n5180 );
not ( n5182 , n5181 );
not ( n5183 , n5087 );
not ( n5184 , n5081 );
or ( n5185 , n5183 , n5184 );
nand ( n5186 , n5185 , n5095 );
nand ( n5187 , n5084 , n5080 );
nand ( n5188 , n5186 , n5187 );
xor ( n5189 , n5182 , n5188 );
not ( n5190 , n5012 );
nand ( n5191 , n5190 , n5013 );
not ( n5192 , n5191 );
not ( n5193 , n5020 );
or ( n5194 , n5192 , n5193 );
not ( n5195 , n5013 );
nand ( n5196 , n5012 , n5195 );
nand ( n5197 , n5194 , n5196 );
xor ( n5198 , n5189 , n5197 );
not ( n5199 , n5065 );
not ( n5200 , n5097 );
or ( n5201 , n5199 , n5200 );
not ( n5202 , n5096 );
not ( n5203 , n5066 );
or ( n5204 , n5202 , n5203 );
nand ( n5205 , n5204 , n5061 );
nand ( n5206 , n5201 , n5205 );
xor ( n5207 , n5198 , n5206 );
and ( n5208 , n516 , n489 );
not ( n5209 , n5032 );
not ( n5210 , n1856 );
nor ( n5211 , n5210 , n1760 );
not ( n5212 , n5211 );
or ( n5213 , n5209 , n5212 );
xor ( n5214 , n514 , n489 );
nand ( n5215 , n1760 , n5214 );
nand ( n5216 , n5213 , n5215 );
xor ( n5217 , n5208 , n5216 );
not ( n5218 , n5093 );
not ( n5219 , n4692 );
or ( n5220 , n5218 , n5219 );
xor ( n5221 , n508 , n495 );
nand ( n5222 , n867 , n5221 );
nand ( n5223 , n5220 , n5222 );
xor ( n5224 , n5217 , n5223 );
not ( n5225 , n5026 );
not ( n5226 , n1930 );
or ( n5227 , n5225 , n5226 );
xor ( n5228 , n512 , n491 );
nand ( n5229 , n1933 , n5228 );
nand ( n5230 , n5227 , n5229 );
buf ( n5231 , n5230 );
not ( n5232 , n5016 );
not ( n5233 , n832 );
or ( n5234 , n5232 , n5233 );
and ( n5235 , n506 , n497 );
not ( n5236 , n506 );
and ( n5237 , n5236 , n2057 );
nor ( n5238 , n5235 , n5237 );
nand ( n5239 , n836 , n5238 );
nand ( n5240 , n5234 , n5239 );
not ( n5241 , n5240 );
not ( n5242 , n5010 );
not ( n5243 , n1449 );
or ( n5244 , n5242 , n5243 );
not ( n5245 , n1327 );
xor ( n5246 , n510 , n493 );
nand ( n5247 , n5245 , n5246 );
nand ( n5248 , n5244 , n5247 );
not ( n5249 , n5248 );
or ( n5250 , n5241 , n5249 );
or ( n5251 , n5248 , n5240 );
nand ( n5252 , n5250 , n5251 );
and ( n5253 , n5231 , n5252 );
not ( n5254 , n5231 );
not ( n5255 , n5248 );
not ( n5256 , n5240 );
not ( n5257 , n5256 );
or ( n5258 , n5255 , n5257 );
not ( n5259 , n5010 );
not ( n5260 , n1449 );
or ( n5261 , n5259 , n5260 );
nand ( n5262 , n5261 , n5247 );
not ( n5263 , n5240 );
or ( n5264 , n5262 , n5263 );
nand ( n5265 , n5258 , n5264 );
and ( n5266 , n5254 , n5265 );
nor ( n5267 , n5253 , n5266 );
xor ( n5268 , n5224 , n5267 );
not ( n5269 , n5028 );
not ( n5270 , n5034 );
or ( n5271 , n5269 , n5270 );
or ( n5272 , n5034 , n5028 );
nand ( n5273 , n5272 , n4704 );
nand ( n5274 , n5271 , n5273 );
xnor ( n5275 , n5268 , n5274 );
xor ( n5276 , n5207 , n5275 );
xor ( n5277 , n5176 , n5276 );
xor ( n5278 , n5055 , n5101 );
and ( n5279 , n5278 , n5110 );
and ( n5280 , n5055 , n5101 );
or ( n5281 , n5279 , n5280 );
xor ( n5282 , n5277 , n5281 );
not ( n5283 , n5040 );
not ( n5284 , n5111 );
or ( n5285 , n5283 , n5284 );
or ( n5286 , n5111 , n5040 );
not ( n5287 , n5042 );
not ( n5288 , n4913 );
or ( n5289 , n5287 , n5288 );
nand ( n5290 , n5289 , n5047 );
nand ( n5291 , n5286 , n5290 );
nand ( n5292 , n5285 , n5291 );
nand ( n5293 , n5282 , n5292 );
not ( n5294 , n5282 );
not ( n5295 , n5292 );
nand ( n5296 , n5294 , n5295 );
nand ( n5297 , n5293 , n5296 );
not ( n5298 , n5297 );
nand ( n5299 , n5172 , n5298 );
nand ( n5300 , n5171 , n5297 );
not ( n5301 , n455 );
nand ( n5302 , n5299 , n5300 , n5301 );
not ( n5303 , n3649 );
nand ( n5304 , n5303 , n3655 );
nand ( n5305 , n5304 , n3629 );
not ( n5306 , n5305 );
and ( n5307 , n3233 , n5306 , n3647 );
nand ( n5308 , n5307 , n4403 );
and ( n5309 , n4427 , n3233 );
nor ( n5310 , n5309 , n4419 );
nand ( n5311 , n5308 , n5310 );
not ( n5312 , n5311 );
nand ( n5313 , n3046 , n3020 );
or ( n5314 , n3020 , n3046 );
nand ( n5315 , n5313 , n5314 );
and ( n5316 , n5315 , n455 );
nand ( n5317 , n5312 , n5316 );
not ( n5318 , n5315 );
nand ( n5319 , n5318 , n5311 , n455 );
nand ( n5320 , n5302 , n5317 , n5319 );
not ( n5321 , n5320 );
not ( n5322 , n5321 );
not ( n5323 , n5322 );
or ( n5324 , n5151 , n5323 );
nand ( n5325 , n5302 , n5317 , n5319 );
not ( n5326 , n5325 );
nand ( n5327 , n5326 , n5146 );
nand ( n5328 , n5324 , n5327 );
buf ( n5329 , n4669 );
buf ( n5330 , n5329 );
nand ( n5331 , n5328 , n5330 );
nand ( n5332 , n5150 , n5331 );
xor ( n5333 , n4662 , n5332 );
xor ( n5334 , n546 , n547 );
not ( n5335 , n5334 );
and ( n5336 , n545 , n546 );
nor ( n5337 , n545 , n546 );
nor ( n5338 , n5336 , n5337 );
and ( n5339 , n5335 , n5338 );
not ( n5340 , n5339 );
not ( n5341 , n5340 );
not ( n5342 , n5341 );
not ( n5343 , n545 );
not ( n5344 , n455 );
not ( n5345 , n5313 );
not ( n5346 , n5314 );
not ( n5347 , n5346 );
or ( n5348 , n5345 , n5347 );
not ( n5349 , n4407 );
nand ( n5350 , n4410 , n4411 );
nand ( n5351 , n5349 , n5350 );
nand ( n5352 , n5348 , n5351 );
not ( n5353 , n5352 );
not ( n5354 , n5353 );
nand ( n5355 , n5310 , n5308 , n5313 );
not ( n5356 , n5355 );
or ( n5357 , n5354 , n5356 );
not ( n5358 , n5314 );
not ( n5359 , n5311 );
or ( n5360 , n5358 , n5359 );
not ( n5361 , n5313 );
nor ( n5362 , n5361 , n5351 );
nand ( n5363 , n5360 , n5362 );
nand ( n5364 , n5357 , n5363 );
not ( n5365 , n5364 );
or ( n5366 , n5344 , n5365 );
not ( n5367 , n5296 );
not ( n5368 , n5154 );
not ( n5369 , n5156 );
or ( n5370 , n5368 , n5369 );
nand ( n5371 , n5370 , n5170 );
not ( n5372 , n5371 );
or ( n5373 , n5367 , n5372 );
nand ( n5374 , n5373 , n5293 );
xor ( n5375 , n5176 , n5276 );
and ( n5376 , n5375 , n5281 );
and ( n5377 , n5176 , n5276 );
or ( n5378 , n5376 , n5377 );
xor ( n5379 , n5208 , n5216 );
and ( n5380 , n5379 , n5223 );
and ( n5381 , n5208 , n5216 );
or ( n5382 , n5380 , n5381 );
not ( n5383 , n5382 );
not ( n5384 , n5214 );
not ( n5385 , n4590 );
or ( n5386 , n5384 , n5385 );
xor ( n5387 , n513 , n489 );
nand ( n5388 , n1859 , n5387 );
nand ( n5389 , n5386 , n5388 );
not ( n5390 , n5221 );
not ( n5391 , n4692 );
or ( n5392 , n5390 , n5391 );
xor ( n5393 , n507 , n495 );
nand ( n5394 , n867 , n5393 );
nand ( n5395 , n5392 , n5394 );
xor ( n5396 , n5389 , n5395 );
not ( n5397 , n5228 );
not ( n5398 , n1930 );
or ( n5399 , n5397 , n5398 );
xor ( n5400 , n511 , n491 );
nand ( n5401 , n1933 , n5400 );
nand ( n5402 , n5399 , n5401 );
xor ( n5403 , n5396 , n5402 );
xor ( n5404 , n5383 , n5403 );
or ( n5405 , n978 , n1062 );
nand ( n5406 , n5405 , n499 );
not ( n5407 , n5246 );
not ( n5408 , n1481 );
or ( n5409 , n5407 , n5408 );
xor ( n5410 , n509 , n493 );
nand ( n5411 , n1328 , n5410 );
nand ( n5412 , n5409 , n5411 );
xor ( n5413 , n5406 , n5412 );
not ( n5414 , n5238 );
not ( n5415 , n963 );
or ( n5416 , n5414 , n5415 );
xor ( n5417 , n497 , n505 );
nand ( n5418 , n836 , n5417 );
nand ( n5419 , n5416 , n5418 );
xor ( n5420 , n5413 , n5419 );
xnor ( n5421 , n5404 , n5420 );
not ( n5422 , n5248 );
not ( n5423 , n5230 );
or ( n5424 , n5422 , n5423 );
or ( n5425 , n5230 , n5248 );
nand ( n5426 , n5425 , n5240 );
nand ( n5427 , n5424 , n5426 );
nand ( n5428 , n515 , n489 );
and ( n5429 , n5428 , n5182 );
not ( n5430 , n5428 );
and ( n5431 , n5430 , n5181 );
nor ( n5432 , n5429 , n5431 );
xor ( n5433 , n5427 , n5432 );
xor ( n5434 , n5182 , n5188 );
and ( n5435 , n5434 , n5197 );
and ( n5436 , n5182 , n5188 );
or ( n5437 , n5435 , n5436 );
xor ( n5438 , n5433 , n5437 );
not ( n5439 , n5224 );
not ( n5440 , n5439 );
not ( n5441 , n5274 );
not ( n5442 , n5441 );
or ( n5443 , n5440 , n5442 );
not ( n5444 , n5267 );
nand ( n5445 , n5443 , n5444 );
not ( n5446 , n5439 );
nand ( n5447 , n5446 , n5274 );
nand ( n5448 , n5445 , n5447 );
xor ( n5449 , n5438 , n5448 );
xor ( n5450 , n5421 , n5449 );
xor ( n5451 , n5198 , n5206 );
and ( n5452 , n5451 , n5275 );
and ( n5453 , n5198 , n5206 );
or ( n5454 , n5452 , n5453 );
xor ( n5455 , n5450 , n5454 );
or ( n5456 , n5378 , n5455 );
nand ( n5457 , n5378 , n5455 );
nand ( n5458 , n5456 , n5457 );
not ( n5459 , n5458 );
and ( n5460 , n5374 , n5459 );
not ( n5461 , n5374 );
and ( n5462 , n5461 , n5458 );
nor ( n5463 , n5460 , n5462 );
nand ( n5464 , n5463 , n793 );
nand ( n5465 , n5366 , n5464 );
buf ( n5466 , n5465 );
not ( n5467 , n5466 );
not ( n5468 , n5467 );
or ( n5469 , n5343 , n5468 );
not ( n5470 , n545 );
nand ( n5471 , n5470 , n5466 );
nand ( n5472 , n5469 , n5471 );
not ( n5473 , n5472 );
or ( n5474 , n5342 , n5473 );
not ( n5475 , n545 );
not ( n5476 , n793 );
xor ( n5477 , n5389 , n5395 );
and ( n5478 , n5477 , n5402 );
and ( n5479 , n5389 , n5395 );
or ( n5480 , n5478 , n5479 );
not ( n5481 , n5387 );
not ( n5482 , n5211 );
or ( n5483 , n5481 , n5482 );
xor ( n5484 , n512 , n489 );
nand ( n5485 , n1760 , n5484 );
nand ( n5486 , n5483 , n5485 );
not ( n5487 , n5400 );
nor ( n5488 , n4807 , n1565 );
not ( n5489 , n5488 );
or ( n5490 , n5487 , n5489 );
xor ( n5491 , n510 , n491 );
nand ( n5492 , n1456 , n5491 );
nand ( n5493 , n5490 , n5492 );
xor ( n5494 , n5486 , n5493 );
not ( n5495 , n832 );
not ( n5496 , n5495 );
and ( n5497 , n5496 , n5417 );
and ( n5498 , n836 , n497 );
nor ( n5499 , n5497 , n5498 );
xnor ( n5500 , n5494 , n5499 );
xor ( n5501 , n5480 , n5500 );
xor ( n5502 , n5406 , n5412 );
and ( n5503 , n5502 , n5419 );
and ( n5504 , n5406 , n5412 );
or ( n5505 , n5503 , n5504 );
xor ( n5506 , n5501 , n5505 );
xor ( n5507 , n5433 , n5437 );
and ( n5508 , n5507 , n5448 );
and ( n5509 , n5433 , n5437 );
or ( n5510 , n5508 , n5509 );
xor ( n5511 , n5506 , n5510 );
not ( n5512 , n5382 );
not ( n5513 , n5403 );
or ( n5514 , n5512 , n5513 );
not ( n5515 , n5383 );
not ( n5516 , n5403 );
not ( n5517 , n5516 );
or ( n5518 , n5515 , n5517 );
nand ( n5519 , n5518 , n5420 );
nand ( n5520 , n5514 , n5519 );
nand ( n5521 , n514 , n489 );
not ( n5522 , n5393 );
not ( n5523 , n859 );
or ( n5524 , n5522 , n5523 );
xor ( n5525 , n506 , n495 );
nand ( n5526 , n867 , n5525 );
nand ( n5527 , n5524 , n5526 );
xor ( n5528 , n5521 , n5527 );
xor ( n5529 , n508 , n493 );
and ( n5530 , n5529 , n1328 );
not ( n5531 , n5410 );
not ( n5532 , n1481 );
nor ( n5533 , n5531 , n5532 );
nor ( n5534 , n5530 , n5533 );
xor ( n5535 , n5528 , n5534 );
not ( n5536 , n5535 );
nand ( n5537 , n5182 , n5428 );
not ( n5538 , n5537 );
not ( n5539 , n5427 );
or ( n5540 , n5538 , n5539 );
or ( n5541 , n5182 , n5428 );
nand ( n5542 , n5540 , n5541 );
not ( n5543 , n5542 );
not ( n5544 , n5543 );
or ( n5545 , n5536 , n5544 );
not ( n5546 , n5535 );
nand ( n5547 , n5546 , n5542 );
nand ( n5548 , n5545 , n5547 );
not ( n5549 , n5548 );
and ( n5550 , n5520 , n5549 );
not ( n5551 , n5520 );
and ( n5552 , n5551 , n5548 );
nor ( n5553 , n5550 , n5552 );
xor ( n5554 , n5511 , n5553 );
not ( n5555 , n5554 );
xor ( n5556 , n5421 , n5449 );
and ( n5557 , n5556 , n5454 );
and ( n5558 , n5421 , n5449 );
or ( n5559 , n5557 , n5558 );
not ( n5560 , n5559 );
nand ( n5561 , n5555 , n5560 );
and ( n5562 , n5559 , n5554 );
not ( n5563 , n5562 );
nand ( n5564 , n5561 , n5563 );
not ( n5565 , n4975 );
not ( n5566 , n1828 );
or ( n5567 , n5565 , n5566 );
nand ( n5568 , n5567 , n4987 );
not ( n5569 , n5568 );
and ( n5570 , n5152 , n5456 , n5296 , n4945 );
not ( n5571 , n5570 );
or ( n5572 , n5569 , n5571 );
not ( n5573 , n5292 );
not ( n5574 , n5282 );
and ( n5575 , n5573 , n5574 );
nor ( n5576 , n5378 , n5455 );
nor ( n5577 , n5575 , n5576 );
and ( n5578 , n5169 , n5577 );
or ( n5579 , n5293 , n5576 );
nand ( n5580 , n5579 , n5457 );
buf ( n5581 , n5580 );
nor ( n5582 , n5578 , n5581 );
nand ( n5583 , n5572 , n5582 );
xnor ( n5584 , n5564 , n5583 );
not ( n5585 , n5584 );
or ( n5586 , n5476 , n5585 );
nand ( n5587 , n5586 , n4431 );
buf ( n5588 , n5587 );
not ( n5589 , n5588 );
not ( n5590 , n5589 );
or ( n5591 , n5475 , n5590 );
nand ( n5592 , n5588 , n4666 );
nand ( n5593 , n5591 , n5592 );
buf ( n5594 , n5334 );
buf ( n5595 , n5594 );
nand ( n5596 , n5593 , n5595 );
nand ( n5597 , n5474 , n5596 );
xor ( n5598 , n5333 , n5597 );
not ( n5599 , n538 );
not ( n5600 , n5599 );
not ( n5601 , n539 );
and ( n5602 , n5600 , n5601 );
nor ( n5603 , n4477 , n538 );
nor ( n5604 , n5602 , n5603 );
not ( n5605 , n537 );
and ( n5606 , n5599 , n5605 );
and ( n5607 , n537 , n538 );
nor ( n5608 , n5606 , n5607 );
and ( n5609 , n5604 , n5608 );
not ( n5610 , n5609 );
not ( n5611 , n537 );
not ( n5612 , n793 );
not ( n5613 , n1813 );
nand ( n5614 , n5613 , n1543 );
not ( n5615 , n1058 );
not ( n5616 , n1315 );
or ( n5617 , n5615 , n5616 );
nand ( n5618 , n5617 , n1325 );
not ( n5619 , n5618 );
not ( n5620 , n5619 );
and ( n5621 , n5614 , n5620 );
not ( n5622 , n5614 );
and ( n5623 , n5622 , n5619 );
nor ( n5624 , n5621 , n5623 );
not ( n5625 , n5624 );
or ( n5626 , n5612 , n5625 );
buf ( n5627 , n4328 );
not ( n5628 , n5627 );
buf ( n5629 , n4348 );
not ( n5630 , n5629 );
not ( n5631 , n4353 );
nand ( n5632 , n5630 , n5631 );
nand ( n5633 , n5629 , n4353 );
nand ( n5634 , n5632 , n5633 );
or ( n5635 , n5634 , n793 );
not ( n5636 , n5635 );
or ( n5637 , n5628 , n5636 );
not ( n5638 , n455 );
not ( n5639 , n5634 );
or ( n5640 , n5638 , n5639 );
not ( n5641 , n5627 );
nand ( n5642 , n5640 , n5641 );
nand ( n5643 , n5637 , n5642 );
nand ( n5644 , n5626 , n5643 );
not ( n5645 , n5644 );
or ( n5646 , n5611 , n5645 );
not ( n5647 , n5644 );
nand ( n5648 , n5647 , n5605 );
nand ( n5649 , n5646 , n5648 );
not ( n5650 , n5649 );
or ( n5651 , n5610 , n5650 );
not ( n5652 , n537 );
not ( n5653 , n455 );
not ( n5654 , n4389 );
not ( n5655 , n5654 );
not ( n5656 , n4390 );
not ( n5657 , n5656 );
or ( n5658 , n5655 , n5657 );
buf ( n5659 , n4391 );
nand ( n5660 , n5658 , n5659 );
not ( n5661 , n5660 );
not ( n5662 , n5661 );
not ( n5663 , n5632 );
not ( n5664 , n4328 );
or ( n5665 , n5663 , n5664 );
nand ( n5666 , n5665 , n5633 );
not ( n5667 , n5666 );
not ( n5668 , n5667 );
or ( n5669 , n5662 , n5668 );
not ( n5670 , n4370 );
not ( n5671 , n5670 );
nand ( n5672 , n5654 , n5656 );
not ( n5673 , n5672 );
or ( n5674 , n5671 , n5673 );
nand ( n5675 , n5674 , n5666 );
nand ( n5676 , n5669 , n5675 );
not ( n5677 , n5676 );
or ( n5678 , n5653 , n5677 );
not ( n5679 , n5618 );
not ( n5680 , n1543 );
or ( n5681 , n5679 , n5680 );
nand ( n5682 , n5681 , n5613 );
nand ( n5683 , n1817 , n1528 );
not ( n5684 , n5683 );
and ( n5685 , n5682 , n5684 );
not ( n5686 , n5682 );
buf ( n5687 , n5683 );
and ( n5688 , n5686 , n5687 );
nor ( n5689 , n5685 , n5688 );
nand ( n5690 , n5689 , n793 );
nand ( n5691 , n5678 , n5690 );
not ( n5692 , n5691 );
not ( n5693 , n5692 );
or ( n5694 , n5652 , n5693 );
or ( n5695 , n537 , n5692 );
nand ( n5696 , n5694 , n5695 );
not ( n5697 , n5604 );
nand ( n5698 , n5696 , n5697 );
nand ( n5699 , n5651 , n5698 );
not ( n5700 , n3990 );
nand ( n5701 , n5700 , n4043 );
nand ( n5702 , n4327 , n5701 );
not ( n5703 , n5702 );
buf ( n5704 , n4323 );
not ( n5705 , n455 );
nor ( n5706 , n5704 , n5705 );
not ( n5707 , n5706 );
or ( n5708 , n5703 , n5707 );
nand ( n5709 , n4327 , n5701 , n455 );
not ( n5710 , n5704 );
or ( n5711 , n5709 , n5710 );
nand ( n5712 , n5708 , n5711 );
not ( n5713 , n1315 );
and ( n5714 , n1324 , n1318 );
not ( n5715 , n1324 );
not ( n5716 , n1318 );
and ( n5717 , n5715 , n5716 );
nor ( n5718 , n5714 , n5717 );
not ( n5719 , n5718 );
and ( n5720 , n5713 , n5719 );
not ( n5721 , n5713 );
and ( n5722 , n5721 , n5718 );
nor ( n5723 , n5720 , n5722 );
nor ( n5724 , n5723 , n455 );
nor ( n5725 , n5712 , n5724 );
not ( n5726 , n5725 );
not ( n5727 , n5726 );
and ( n5728 , n5727 , n537 );
and ( n5729 , n5699 , n5728 );
not ( n5730 , n541 );
not ( n5731 , n4655 );
not ( n5732 , n5731 );
or ( n5733 , n5730 , n5732 );
not ( n5734 , n541 );
nand ( n5735 , n4651 , n5734 );
nand ( n5736 , n5733 , n5735 );
not ( n5737 , n5736 );
and ( n5738 , n542 , n543 );
not ( n5739 , n542 );
and ( n5740 , n5739 , n5146 );
nor ( n5741 , n5738 , n5740 );
not ( n5742 , n5741 );
and ( n5743 , n541 , n542 );
nor ( n5744 , n541 , n542 );
nor ( n5745 , n5743 , n5744 );
and ( n5746 , n5742 , n5745 );
buf ( n5747 , n5746 );
not ( n5748 , n5747 );
or ( n5749 , n5737 , n5748 );
and ( n5750 , n4627 , n4972 );
and ( n5751 , n1980 , n1981 );
nor ( n5752 , n5750 , n5751 );
not ( n5753 , n5752 );
not ( n5754 , n1828 );
or ( n5755 , n5753 , n5754 );
nand ( n5756 , n4980 , n4984 );
nand ( n5757 , n5755 , n5756 );
not ( n5758 , n5757 );
nand ( n5759 , n4979 , n4964 );
and ( n5760 , n5759 , n4465 );
nand ( n5761 , n5758 , n5760 );
nand ( n5762 , n4398 , n3629 , n4400 , n4401 );
nand ( n5763 , n3802 , n3629 );
nand ( n5764 , n5762 , n5763 );
not ( n5765 , n5764 );
nand ( n5766 , n3656 , n4424 );
and ( n5767 , n5766 , n455 );
nand ( n5768 , n5765 , n5767 );
nor ( n5769 , n5759 , n455 );
nand ( n5770 , n5757 , n5769 );
not ( n5771 , n5763 );
not ( n5772 , n5762 );
or ( n5773 , n5771 , n5772 );
and ( n5774 , n3656 , n4424 , n455 );
nand ( n5775 , n5773 , n5774 );
nand ( n5776 , n5761 , n5768 , n5770 , n5775 );
not ( n5777 , n5776 );
not ( n5778 , n5777 );
nand ( n5779 , n5778 , n541 );
not ( n5780 , n5779 );
nand ( n5781 , n5777 , n4445 );
not ( n5782 , n5781 );
or ( n5783 , n5780 , n5782 );
buf ( n5784 , n5741 );
buf ( n5785 , n5784 );
buf ( n5786 , n5785 );
nand ( n5787 , n5783 , n5786 );
nand ( n5788 , n5749 , n5787 );
xor ( n5789 , n5729 , n5788 );
not ( n5790 , n5697 );
not ( n5791 , n455 );
not ( n5792 , n5791 );
buf ( n5793 , n1682 );
or ( n5794 , n1823 , n1681 );
nand ( n5795 , n5793 , n5794 );
not ( n5796 , n1544 );
not ( n5797 , n5618 );
or ( n5798 , n5796 , n5797 );
not ( n5799 , n1818 );
nand ( n5800 , n5798 , n5799 );
and ( n5801 , n5795 , n5800 );
not ( n5802 , n5795 );
not ( n5803 , n5800 );
and ( n5804 , n5802 , n5803 );
nor ( n5805 , n5801 , n5804 );
not ( n5806 , n5805 );
or ( n5807 , n5792 , n5806 );
not ( n5808 , n5659 );
not ( n5809 , n5666 );
or ( n5810 , n5808 , n5809 );
nand ( n5811 , n5654 , n4369 );
buf ( n5812 , n5811 );
nand ( n5813 , n5810 , n5812 );
nand ( n5814 , n4396 , n4382 );
not ( n5815 , n5814 );
and ( n5816 , n5815 , n455 );
and ( n5817 , n5813 , n5816 );
and ( n5818 , n5811 , n5814 , n455 );
nand ( n5819 , n5659 , n5666 );
and ( n5820 , n5818 , n5819 );
nor ( n5821 , n5817 , n5820 );
nand ( n5822 , n5807 , n5821 );
not ( n5823 , n5822 );
not ( n5824 , n5823 );
not ( n5825 , n5824 );
not ( n5826 , n537 );
nand ( n5827 , n5825 , n5826 );
nand ( n5828 , n5824 , n537 );
nand ( n5829 , n5827 , n5828 );
not ( n5830 , n5829 );
or ( n5831 , n5790 , n5830 );
nand ( n5832 , n5609 , n5696 );
nand ( n5833 , n5831 , n5832 );
not ( n5834 , n455 );
nand ( n5835 , n5834 , n5624 );
nand ( n5836 , n5835 , n5643 );
not ( n5837 , n5836 );
nand ( n5838 , n5837 , n537 );
xnor ( n5839 , n5833 , n5838 );
and ( n5840 , n5789 , n5839 );
and ( n5841 , n5729 , n5788 );
or ( n5842 , n5840 , n5841 );
not ( n5843 , n541 );
not ( n5844 , n5791 );
nand ( n5845 , n4992 , n4945 );
xor ( n5846 , n5568 , n5845 );
not ( n5847 , n5846 );
or ( n5848 , n5844 , n5847 );
not ( n5849 , n4455 );
nor ( n5850 , n3740 , n3781 );
nor ( n5851 , n4489 , n5850 );
nand ( n5852 , n4400 , n5304 , n5851 );
nor ( n5853 , n5849 , n5852 );
not ( n5854 , n5853 );
not ( n5855 , n5854 );
not ( n5856 , n3793 );
nor ( n5857 , n5856 , n4459 );
nor ( n5858 , n5857 , n4463 );
or ( n5859 , n5858 , n5305 );
not ( n5860 , n4487 );
nand ( n5861 , n3654 , n3649 );
not ( n5862 , n5861 );
or ( n5863 , n5860 , n5862 );
nand ( n5864 , n5863 , n3656 );
nand ( n5865 , n5859 , n5864 );
not ( n5866 , n5865 );
not ( n5867 , n5866 );
or ( n5868 , n5855 , n5867 );
nand ( n5869 , n3632 , n3645 );
nand ( n5870 , n3647 , n5869 );
not ( n5871 , n5870 );
not ( n5872 , n5871 );
nand ( n5873 , n5868 , n5872 );
nand ( n5874 , n5871 , n5854 , n5866 );
nand ( n5875 , n5873 , n5874 , n455 );
nand ( n5876 , n5848 , n5875 );
not ( n5877 , n5876 );
or ( n5878 , n5843 , n5877 );
not ( n5879 , n5568 );
nand ( n5880 , n5879 , n5845 , n5301 );
not ( n5881 , n5854 );
not ( n5882 , n5866 );
or ( n5883 , n5881 , n5882 );
not ( n5884 , n455 );
nor ( n5885 , n5884 , n5870 );
nand ( n5886 , n5883 , n5885 );
nand ( n5887 , n5866 , n5854 , n5870 , n455 );
nor ( n5888 , n5845 , n455 );
nand ( n5889 , n5888 , n5568 );
nand ( n5890 , n5880 , n5886 , n5887 , n5889 );
not ( n5891 , n5890 );
nand ( n5892 , n5891 , n5734 );
nand ( n5893 , n5878 , n5892 );
nand ( n5894 , n5893 , n5785 );
not ( n5895 , n5781 );
nand ( n5896 , n5778 , n541 );
not ( n5897 , n5896 );
or ( n5898 , n5895 , n5897 );
nand ( n5899 , n5898 , n5747 );
nand ( n5900 , n5894 , n5899 );
not ( n5901 , n5696 );
not ( n5902 , n5901 );
not ( n5903 , n5609 );
not ( n5904 , n5903 );
and ( n5905 , n5902 , n5904 );
and ( n5906 , n5829 , n5697 );
nor ( n5907 , n5905 , n5906 );
nor ( n5908 , n5907 , n5838 );
xor ( n5909 , n5900 , n5908 );
not ( n5910 , n455 );
not ( n5911 , n5676 );
or ( n5912 , n5910 , n5911 );
nand ( n5913 , n5912 , n5690 );
buf ( n5914 , n5913 );
and ( n5915 , n5914 , n537 );
not ( n5916 , n5697 );
not ( n5917 , n537 );
not ( n5918 , n455 );
nand ( n5919 , n4401 , n4459 );
not ( n5920 , n5919 );
and ( n5921 , n4456 , n5920 );
not ( n5922 , n4456 );
and ( n5923 , n5922 , n5919 );
nor ( n5924 , n5921 , n5923 );
not ( n5925 , n5924 );
or ( n5926 , n5918 , n5925 );
not ( n5927 , n5793 );
not ( n5928 , n5800 );
or ( n5929 , n5927 , n5928 );
buf ( n5930 , n5794 );
nand ( n5931 , n5929 , n5930 );
and ( n5932 , n1808 , n1800 );
not ( n5933 , n1808 );
and ( n5934 , n5933 , n1826 );
nor ( n5935 , n5932 , n5934 );
not ( n5936 , n5935 );
and ( n5937 , n5931 , n5936 );
not ( n5938 , n5931 );
and ( n5939 , n5938 , n5935 );
nor ( n5940 , n5937 , n5939 );
nand ( n5941 , n5940 , n793 );
nand ( n5942 , n5926 , n5941 );
buf ( n5943 , n5942 );
not ( n5944 , n5943 );
not ( n5945 , n5944 );
or ( n5946 , n5917 , n5945 );
nand ( n5947 , n5943 , n5605 );
nand ( n5948 , n5946 , n5947 );
not ( n5949 , n5948 );
or ( n5950 , n5916 , n5949 );
nand ( n5951 , n5609 , n5829 );
nand ( n5952 , n5950 , n5951 );
xor ( n5953 , n5915 , n5952 );
xor ( n5954 , n5909 , n5953 );
xor ( n5955 , n5842 , n5954 );
not ( n5956 , n4660 );
not ( n5957 , n4479 );
or ( n5958 , n5956 , n5957 );
not ( n5959 , n5943 );
not ( n5960 , n5959 );
not ( n5961 , n4450 );
nor ( n5962 , n5961 , n539 );
and ( n5963 , n5960 , n5962 );
nand ( n5964 , n4450 , n539 );
not ( n5965 , n5964 );
and ( n5966 , n5959 , n5965 );
nor ( n5967 , n5963 , n5966 );
nand ( n5968 , n5958 , n5967 );
not ( n5969 , n5943 );
not ( n5970 , n4660 );
nor ( n5971 , n5970 , n4477 );
nand ( n5972 , n5969 , n5971 );
not ( n5973 , n455 );
not ( n5974 , n5924 );
or ( n5975 , n5973 , n5974 );
nand ( n5976 , n5975 , n5941 );
nor ( n5977 , n5970 , n539 );
nand ( n5978 , n5976 , n5977 );
and ( n5979 , n5823 , n539 );
not ( n5980 , n5823 );
and ( n5981 , n5980 , n4477 );
nor ( n5982 , n5979 , n5981 );
nand ( n5983 , n5982 , n4450 );
nand ( n5984 , n5972 , n5978 , n5983 );
not ( n5985 , n537 );
not ( n5986 , n5726 );
or ( n5987 , n5985 , n5986 );
nand ( n5988 , n5605 , n5725 );
nand ( n5989 , n5987 , n5988 );
not ( n5990 , n5989 );
not ( n5991 , n5990 );
not ( n5992 , n5903 );
and ( n5993 , n5991 , n5992 );
and ( n5994 , n5649 , n5697 );
nor ( n5995 , n5993 , n5994 );
not ( n5996 , n793 );
not ( n5997 , n1301 );
buf ( n5998 , n1247 );
not ( n5999 , n5998 );
or ( n6000 , n5997 , n5999 );
nand ( n6001 , n1308 , n1309 );
nand ( n6002 , n6000 , n6001 );
nand ( n6003 , n1306 , n1313 );
not ( n6004 , n6003 );
and ( n6005 , n6002 , n6004 );
not ( n6006 , n6002 );
and ( n6007 , n6006 , n6003 );
nor ( n6008 , n6005 , n6007 );
not ( n6009 , n6008 );
or ( n6010 , n5996 , n6009 );
nand ( n6011 , n6010 , n4440 );
buf ( n6012 , n6011 );
not ( n6013 , n6012 );
not ( n6014 , n6013 );
nand ( n6015 , n6014 , n537 );
nor ( n6016 , n5995 , n6015 );
xor ( n6017 , n5984 , n6016 );
and ( n6018 , n5609 , n5649 );
and ( n6019 , n5696 , n5697 );
nor ( n6020 , n6018 , n6019 );
and ( n6021 , n5728 , n6020 );
not ( n6022 , n5728 );
and ( n6023 , n6022 , n5699 );
or ( n6024 , n6021 , n6023 );
and ( n6025 , n6017 , n6024 );
and ( n6026 , n5984 , n6016 );
or ( n6027 , n6025 , n6026 );
xor ( n6028 , n5968 , n6027 );
not ( n6029 , n5330 );
not ( n6030 , n5148 );
or ( n6031 , n6029 , n6030 );
not ( n6032 , n5146 );
not ( n6033 , n5891 );
not ( n6034 , n6033 );
not ( n6035 , n6034 );
or ( n6036 , n6032 , n6035 );
nand ( n6037 , n6033 , n543 );
nand ( n6038 , n6036 , n6037 );
nand ( n6039 , n6038 , n4671 );
nand ( n6040 , n6031 , n6039 );
and ( n6041 , n6028 , n6040 );
and ( n6042 , n5968 , n6027 );
or ( n6043 , n6041 , n6042 );
xor ( n6044 , n5955 , n6043 );
xor ( n6045 , n5598 , n6044 );
not ( n6046 , n5595 );
not ( n6047 , n5472 );
or ( n6048 , n6046 , n6047 );
xor ( n6049 , n545 , n5321 );
nand ( n6050 , n6049 , n5341 );
nand ( n6051 , n6048 , n6050 );
xor ( n6052 , n5729 , n5788 );
xor ( n6053 , n6052 , n5839 );
xor ( n6054 , n6051 , n6053 );
not ( n6055 , n4671 );
buf ( n6056 , n5776 );
and ( n6057 , n5146 , n6056 );
not ( n6058 , n5146 );
not ( n6059 , n6056 );
and ( n6060 , n6058 , n6059 );
nor ( n6061 , n6057 , n6060 );
not ( n6062 , n6061 );
or ( n6063 , n6055 , n6062 );
nand ( n6064 , n6038 , n5330 );
nand ( n6065 , n6063 , n6064 );
not ( n6066 , n5747 );
and ( n6067 , n4473 , n5734 );
not ( n6068 , n4473 );
and ( n6069 , n6068 , n541 );
or ( n6070 , n6067 , n6069 );
not ( n6071 , n6070 );
or ( n6072 , n6066 , n6071 );
nand ( n6073 , n5736 , n5786 );
nand ( n6074 , n6072 , n6073 );
xor ( n6075 , n6065 , n6074 );
not ( n6076 , n5339 );
not ( n6077 , n545 );
not ( n6078 , n5141 );
or ( n6079 , n6077 , n6078 );
nand ( n6080 , n5145 , n4666 );
nand ( n6081 , n6079 , n6080 );
not ( n6082 , n6081 );
or ( n6083 , n6076 , n6082 );
nand ( n6084 , n6049 , n5595 );
nand ( n6085 , n6083 , n6084 );
and ( n6086 , n6075 , n6085 );
and ( n6087 , n6065 , n6074 );
or ( n6088 , n6086 , n6087 );
and ( n6089 , n6054 , n6088 );
and ( n6090 , n6051 , n6053 );
or ( n6091 , n6089 , n6090 );
xor ( n6092 , n6045 , n6091 );
xor ( n6093 , n6051 , n6053 );
xor ( n6094 , n6093 , n6088 );
xor ( n6095 , n550 , n551 );
not ( n6096 , n6095 );
not ( n6097 , n2713 );
not ( n6098 , n2563 );
and ( n6099 , n6097 , n6098 );
xor ( n6100 , n2254 , n2414 );
and ( n6101 , n6100 , n2562 );
and ( n6102 , n2254 , n2414 );
or ( n6103 , n6101 , n6102 );
xor ( n6104 , n2127 , n2217 );
and ( n6105 , n6104 , n2253 );
and ( n6106 , n2127 , n2217 );
or ( n6107 , n6105 , n6106 );
or ( n6108 , n2142 , n2164 );
nand ( n6109 , n6108 , n497 );
not ( n6110 , n2078 );
and ( n6111 , n495 , n2149 );
not ( n6112 , n495 );
and ( n6113 , n6112 , n2152 );
or ( n6114 , n6111 , n6113 );
not ( n6115 , n6114 );
or ( n6116 , n6110 , n6115 );
nand ( n6117 , n2285 , n2060 );
nand ( n6118 , n6116 , n6117 );
xor ( n6119 , n6109 , n6118 );
not ( n6120 , n2000 );
not ( n6121 , n2229 );
or ( n6122 , n6120 , n6121 );
not ( n6123 , n491 );
not ( n6124 , n2190 );
or ( n6125 , n6123 , n6124 );
nand ( n6126 , n2193 , n2015 );
nand ( n6127 , n6125 , n6126 );
nand ( n6128 , n6127 , n2036 );
nand ( n6129 , n6122 , n6128 );
xor ( n6130 , n6119 , n6129 );
xor ( n6131 , n2260 , n2276 );
and ( n6132 , n6131 , n2288 );
and ( n6133 , n2260 , n2276 );
or ( n6134 , n6132 , n6133 );
xor ( n6135 , n6130 , n6134 );
xor ( n6136 , n2234 , n2245 );
and ( n6137 , n6136 , n2252 );
and ( n6138 , n2234 , n2245 );
or ( n6139 , n6137 , n6138 );
xor ( n6140 , n2287 , n6139 );
not ( n6141 , n2120 );
not ( n6142 , n2242 );
or ( n6143 , n6141 , n6142 );
xor ( n6144 , n489 , n2026 );
nand ( n6145 , n6144 , n2243 );
nand ( n6146 , n6143 , n6145 );
not ( n6147 , n2274 );
not ( n6148 , n2202 );
or ( n6149 , n6147 , n6148 );
not ( n6150 , n3301 );
not ( n6151 , n6150 );
nand ( n6152 , n2185 , n2264 );
not ( n6153 , n6152 );
or ( n6154 , n6151 , n6153 );
not ( n6155 , n493 );
not ( n6156 , n2185 );
or ( n6157 , n6155 , n6156 );
nand ( n6158 , n6157 , n2067 );
nand ( n6159 , n6154 , n6158 );
nand ( n6160 , n6149 , n6159 );
xor ( n6161 , n6146 , n6160 );
and ( n6162 , n2090 , n489 );
xor ( n6163 , n6161 , n6162 );
xor ( n6164 , n6140 , n6163 );
xor ( n6165 , n6135 , n6164 );
xor ( n6166 , n6107 , n6165 );
xor ( n6167 , n2289 , n2363 );
and ( n6168 , n6167 , n2413 );
and ( n6169 , n2289 , n2363 );
or ( n6170 , n6168 , n6169 );
xor ( n6171 , n6166 , n6170 );
nor ( n6172 , n6103 , n6171 );
nor ( n6173 , n6099 , n6172 );
buf ( n6174 , n6173 );
xor ( n6175 , n2287 , n6139 );
and ( n6176 , n6175 , n6163 );
and ( n6177 , n2287 , n6139 );
or ( n6178 , n6176 , n6177 );
xor ( n6179 , n6109 , n6118 );
and ( n6180 , n6179 , n6129 );
and ( n6181 , n6109 , n6118 );
or ( n6182 , n6180 , n6181 );
not ( n6183 , n2084 );
not ( n6184 , n489 );
not ( n6185 , n2208 );
or ( n6186 , n6184 , n6185 );
nand ( n6187 , n2227 , n1949 );
nand ( n6188 , n6186 , n6187 );
not ( n6189 , n6188 );
or ( n6190 , n6183 , n6189 );
nand ( n6191 , n6144 , n2122 );
nand ( n6192 , n6190 , n6191 );
and ( n6193 , n2481 , n489 );
xor ( n6194 , n6192 , n6193 );
not ( n6195 , n2060 );
not ( n6196 , n6114 );
or ( n6197 , n6195 , n6196 );
nand ( n6198 , n2078 , n495 );
nand ( n6199 , n6197 , n6198 );
xor ( n6200 , n6194 , n6199 );
xor ( n6201 , n6182 , n6200 );
not ( n6202 , n2000 );
not ( n6203 , n6127 );
or ( n6204 , n6202 , n6203 );
not ( n6205 , n491 );
not ( n6206 , n2270 );
not ( n6207 , n6206 );
or ( n6208 , n6205 , n6207 );
nand ( n6209 , n2270 , n2015 );
nand ( n6210 , n6208 , n6209 );
nand ( n6211 , n6210 , n2036 );
nand ( n6212 , n6204 , n6211 );
and ( n6213 , n2264 , n3301 );
not ( n6214 , n2264 );
and ( n6215 , n6214 , n6150 );
nor ( n6216 , n6213 , n6215 );
not ( n6217 , n6216 );
not ( n6218 , n2203 );
or ( n6219 , n6217 , n6218 );
and ( n6220 , n456 , n458 );
not ( n6221 , n456 );
and ( n6222 , n6221 , n474 );
nor ( n6223 , n6220 , n6222 );
and ( n6224 , n493 , n6223 );
not ( n6225 , n493 );
and ( n6226 , n6225 , n2283 );
or ( n6227 , n6224 , n6226 );
nand ( n6228 , n6227 , n2185 );
nand ( n6229 , n6219 , n6228 );
not ( n6230 , n6229 );
xor ( n6231 , n6212 , n6230 );
xor ( n6232 , n6146 , n6160 );
and ( n6233 , n6232 , n6162 );
and ( n6234 , n6146 , n6160 );
or ( n6235 , n6233 , n6234 );
xor ( n6236 , n6231 , n6235 );
xor ( n6237 , n6201 , n6236 );
xor ( n6238 , n6178 , n6237 );
xor ( n6239 , n6130 , n6134 );
and ( n6240 , n6239 , n6164 );
and ( n6241 , n6130 , n6134 );
or ( n6242 , n6240 , n6241 );
xor ( n6243 , n6238 , n6242 );
xor ( n6244 , n6107 , n6165 );
and ( n6245 , n6244 , n6170 );
and ( n6246 , n6107 , n6165 );
or ( n6247 , n6245 , n6246 );
nor ( n6248 , n6243 , n6247 );
not ( n6249 , n6248 );
and ( n6250 , n6174 , n6249 );
not ( n6251 , n6250 );
not ( n6252 , n4429 );
or ( n6253 , n6251 , n6252 );
not ( n6254 , n6103 );
not ( n6255 , n6171 );
or ( n6256 , n6254 , n6255 );
nor ( n6257 , n6171 , n6103 );
nand ( n6258 , n2563 , n2713 );
or ( n6259 , n6257 , n6258 );
nand ( n6260 , n6256 , n6259 );
buf ( n6261 , n6260 );
not ( n6262 , n6247 );
not ( n6263 , n6243 );
nand ( n6264 , n6262 , n6263 );
and ( n6265 , n6261 , n6264 );
nand ( n6266 , n6247 , n6243 );
not ( n6267 , n6266 );
nor ( n6268 , n6265 , n6267 );
nand ( n6269 , n6253 , n6268 );
xor ( n6270 , n6212 , n6230 );
and ( n6271 , n6270 , n6235 );
and ( n6272 , n6212 , n6230 );
or ( n6273 , n6271 , n6272 );
xor ( n6274 , n6192 , n6193 );
and ( n6275 , n6274 , n6199 );
and ( n6276 , n6192 , n6193 );
or ( n6277 , n6275 , n6276 );
or ( n6278 , n2078 , n2060 );
nand ( n6279 , n6278 , n495 );
not ( n6280 , n2185 );
and ( n6281 , n493 , n2149 );
not ( n6282 , n493 );
and ( n6283 , n6282 , n2152 );
or ( n6284 , n6281 , n6283 );
not ( n6285 , n6284 );
or ( n6286 , n6280 , n6285 );
nand ( n6287 , n6227 , n2203 );
nand ( n6288 , n6286 , n6287 );
xor ( n6289 , n6279 , n6288 );
not ( n6290 , n2084 );
xor ( n6291 , n489 , n2193 );
not ( n6292 , n6291 );
or ( n6293 , n6290 , n6292 );
nand ( n6294 , n6188 , n2122 );
nand ( n6295 , n6293 , n6294 );
xor ( n6296 , n6289 , n6295 );
xor ( n6297 , n6277 , n6296 );
and ( n6298 , n489 , n2026 );
not ( n6299 , n2036 );
not ( n6300 , n491 );
not ( n6301 , n2067 );
or ( n6302 , n6300 , n6301 );
not ( n6303 , n2075 );
not ( n6304 , n6303 );
nand ( n6305 , n6304 , n2015 );
nand ( n6306 , n6302 , n6305 );
not ( n6307 , n6306 );
or ( n6308 , n6299 , n6307 );
nand ( n6309 , n6210 , n2000 );
nand ( n6310 , n6308 , n6309 );
xor ( n6311 , n6298 , n6310 );
xor ( n6312 , n6311 , n6229 );
xor ( n6313 , n6297 , n6312 );
xor ( n6314 , n6273 , n6313 );
xor ( n6315 , n6182 , n6200 );
and ( n6316 , n6315 , n6236 );
and ( n6317 , n6182 , n6200 );
or ( n6318 , n6316 , n6317 );
xor ( n6319 , n6314 , n6318 );
not ( n6320 , n6319 );
xor ( n6321 , n6178 , n6237 );
and ( n6322 , n6321 , n6242 );
and ( n6323 , n6178 , n6237 );
or ( n6324 , n6322 , n6323 );
not ( n6325 , n6324 );
nand ( n6326 , n6320 , n6325 );
not ( n6327 , n6325 );
nand ( n6328 , n6327 , n6319 );
nand ( n6329 , n6326 , n6328 );
not ( n6330 , n6329 );
and ( n6331 , n6330 , n455 );
and ( n6332 , n6269 , n6331 );
not ( n6333 , n6269 );
and ( n6334 , n6329 , n455 );
and ( n6335 , n6333 , n6334 );
nor ( n6336 , n6332 , n6335 );
not ( n6337 , n5560 );
not ( n6338 , n5555 );
or ( n6339 , n6337 , n6338 );
xor ( n6340 , n5506 , n5510 );
and ( n6341 , n6340 , n5553 );
and ( n6342 , n5506 , n5510 );
or ( n6343 , n6341 , n6342 );
not ( n6344 , n6343 );
xor ( n6345 , n5480 , n5500 );
and ( n6346 , n6345 , n5505 );
and ( n6347 , n5480 , n5500 );
or ( n6348 , n6346 , n6347 );
not ( n6349 , n6348 );
not ( n6350 , n6349 );
xor ( n6351 , n5521 , n5527 );
and ( n6352 , n6351 , n5534 );
and ( n6353 , n5521 , n5527 );
or ( n6354 , n6352 , n6353 );
not ( n6355 , n6354 );
not ( n6356 , n6355 );
not ( n6357 , n5525 );
not ( n6358 , n859 );
or ( n6359 , n6357 , n6358 );
xor ( n6360 , n505 , n495 );
nand ( n6361 , n867 , n6360 );
nand ( n6362 , n6359 , n6361 );
not ( n6363 , n836 );
not ( n6364 , n6363 );
not ( n6365 , n5495 );
or ( n6366 , n6364 , n6365 );
nand ( n6367 , n6366 , n497 );
xor ( n6368 , n6362 , n6367 );
not ( n6369 , n5491 );
not ( n6370 , n1930 );
or ( n6371 , n6369 , n6370 );
xor ( n6372 , n509 , n491 );
nand ( n6373 , n1933 , n6372 );
nand ( n6374 , n6371 , n6373 );
not ( n6375 , n6374 );
and ( n6376 , n6368 , n6375 );
not ( n6377 , n6368 );
and ( n6378 , n6377 , n6374 );
nor ( n6379 , n6376 , n6378 );
not ( n6380 , n6379 );
not ( n6381 , n6380 );
or ( n6382 , n6356 , n6381 );
nand ( n6383 , n6379 , n6354 );
nand ( n6384 , n6382 , n6383 );
not ( n6385 , n5527 );
not ( n6386 , n6385 );
not ( n6387 , n5493 );
not ( n6388 , n5486 );
or ( n6389 , n6387 , n6388 );
nor ( n6390 , n5493 , n5486 );
or ( n6391 , n5499 , n6390 );
nand ( n6392 , n6389 , n6391 );
not ( n6393 , n6392 );
not ( n6394 , n6393 );
or ( n6395 , n6386 , n6394 );
not ( n6396 , n6385 );
nand ( n6397 , n6396 , n6392 );
nand ( n6398 , n6395 , n6397 );
nand ( n6399 , n513 , n489 );
xor ( n6400 , n489 , n511 );
nand ( n6401 , n1859 , n6400 );
nand ( n6402 , n5211 , n5484 );
and ( n6403 , n6401 , n6402 );
xor ( n6404 , n6399 , n6403 );
not ( n6405 , n5532 );
xnor ( n6406 , n508 , n493 );
not ( n6407 , n6406 );
and ( n6408 , n6405 , n6407 );
xor ( n6409 , n493 , n507 );
and ( n6410 , n814 , n6409 );
nor ( n6411 , n6408 , n6410 );
xor ( n6412 , n6404 , n6411 );
not ( n6413 , n6412 );
not ( n6414 , n6413 );
and ( n6415 , n6398 , n6414 );
not ( n6416 , n6398 );
and ( n6417 , n6416 , n6413 );
nor ( n6418 , n6415 , n6417 );
and ( n6419 , n6384 , n6418 );
not ( n6420 , n6384 );
not ( n6421 , n6418 );
and ( n6422 , n6420 , n6421 );
nor ( n6423 , n6419 , n6422 );
not ( n6424 , n6423 );
or ( n6425 , n6350 , n6424 );
or ( n6426 , n6423 , n6349 );
nand ( n6427 , n6425 , n6426 );
not ( n6428 , n5542 );
nand ( n6429 , n6428 , n5535 );
not ( n6430 , n6429 );
not ( n6431 , n5520 );
or ( n6432 , n6430 , n6431 );
nand ( n6433 , n6432 , n5547 );
xor ( n6434 , n6427 , n6433 );
nand ( n6435 , n6344 , n6434 );
nand ( n6436 , n6339 , n6435 );
buf ( n6437 , n6436 );
nand ( n6438 , n6423 , n6349 );
not ( n6439 , n6438 );
not ( n6440 , n6433 );
or ( n6441 , n6439 , n6440 );
or ( n6442 , n6349 , n6423 );
nand ( n6443 , n6441 , n6442 );
not ( n6444 , n6385 );
not ( n6445 , n6412 );
or ( n6446 , n6444 , n6445 );
nand ( n6447 , n6446 , n6392 );
nand ( n6448 , n6413 , n5527 );
nand ( n6449 , n6447 , n6448 );
not ( n6450 , n6449 );
nand ( n6451 , n512 , n489 );
not ( n6452 , n6451 );
not ( n6453 , n6400 );
not ( n6454 , n4590 );
or ( n6455 , n6453 , n6454 );
xor ( n6456 , n489 , n510 );
nand ( n6457 , n1859 , n6456 );
nand ( n6458 , n6455 , n6457 );
not ( n6459 , n6458 );
xor ( n6460 , n6452 , n6459 );
not ( n6461 , n6360 );
not ( n6462 , n4692 );
or ( n6463 , n6461 , n6462 );
nand ( n6464 , n867 , n495 );
nand ( n6465 , n6463 , n6464 );
xor ( n6466 , n6460 , n6465 );
not ( n6467 , n6374 );
not ( n6468 , n6362 );
or ( n6469 , n6467 , n6468 );
not ( n6470 , n6375 );
not ( n6471 , n6362 );
not ( n6472 , n6471 );
or ( n6473 , n6470 , n6472 );
nand ( n6474 , n6473 , n6367 );
nand ( n6475 , n6469 , n6474 );
not ( n6476 , n6475 );
xor ( n6477 , n6466 , n6476 );
not ( n6478 , n6409 );
not ( n6479 , n1481 );
or ( n6480 , n6478 , n6479 );
xor ( n6481 , n506 , n493 );
nand ( n6482 , n814 , n6481 );
nand ( n6483 , n6480 , n6482 );
not ( n6484 , n6372 );
not ( n6485 , n1930 );
or ( n6486 , n6484 , n6485 );
xor ( n6487 , n508 , n491 );
nand ( n6488 , n1933 , n6487 );
nand ( n6489 , n6486 , n6488 );
xor ( n6490 , n6483 , n6489 );
xor ( n6491 , n6399 , n6403 );
and ( n6492 , n6491 , n6411 );
and ( n6493 , n6399 , n6403 );
or ( n6494 , n6492 , n6493 );
not ( n6495 , n6494 );
and ( n6496 , n6490 , n6495 );
not ( n6497 , n6490 );
and ( n6498 , n6497 , n6494 );
nor ( n6499 , n6496 , n6498 );
xor ( n6500 , n6477 , n6499 );
xor ( n6501 , n6450 , n6500 );
not ( n6502 , n6383 );
not ( n6503 , n6418 );
or ( n6504 , n6502 , n6503 );
or ( n6505 , n6379 , n6354 );
nand ( n6506 , n6504 , n6505 );
xnor ( n6507 , n6501 , n6506 );
not ( n6508 , n6507 );
nor ( n6509 , n6443 , n6508 );
nor ( n6510 , n6437 , n6509 );
and ( n6511 , n6510 , n5296 , n5456 );
not ( n6512 , n6511 );
not ( n6513 , n5371 );
or ( n6514 , n6512 , n6513 );
nor ( n6515 , n6436 , n6509 );
not ( n6516 , n6515 );
not ( n6517 , n5580 );
or ( n6518 , n6516 , n6517 );
not ( n6519 , n6435 );
not ( n6520 , n5562 );
or ( n6521 , n6519 , n6520 );
not ( n6522 , n6434 );
nand ( n6523 , n6522 , n6343 );
nand ( n6524 , n6521 , n6523 );
not ( n6525 , n6443 );
buf ( n6526 , n6507 );
nand ( n6527 , n6525 , n6526 );
and ( n6528 , n6524 , n6527 );
nand ( n6529 , n6443 , n6508 );
not ( n6530 , n6529 );
nor ( n6531 , n6528 , n6530 );
nand ( n6532 , n6518 , n6531 );
not ( n6533 , n6532 );
nand ( n6534 , n6514 , n6533 );
and ( n6535 , n489 , n511 );
xor ( n6536 , n6535 , n6483 );
xor ( n6537 , n507 , n491 );
nand ( n6538 , n1933 , n6537 );
nand ( n6539 , n6487 , n1930 );
nand ( n6540 , n6538 , n6539 );
xor ( n6541 , n6536 , n6540 );
not ( n6542 , n6541 );
not ( n6543 , n6542 );
not ( n6544 , n6451 );
not ( n6545 , n6459 );
or ( n6546 , n6544 , n6545 );
nand ( n6547 , n6546 , n6465 );
nand ( n6548 , n6452 , n6458 );
nand ( n6549 , n6547 , n6548 );
not ( n6550 , n6549 );
or ( n6551 , n6543 , n6550 );
not ( n6552 , n6549 );
nand ( n6553 , n6541 , n6552 );
nand ( n6554 , n6551 , n6553 );
not ( n6555 , n6481 );
not ( n6556 , n1586 );
or ( n6557 , n6555 , n6556 );
xor ( n6558 , n505 , n493 );
nand ( n6559 , n1328 , n6558 );
nand ( n6560 , n6557 , n6559 );
not ( n6561 , n6456 );
buf ( n6562 , n4590 );
not ( n6563 , n6562 );
or ( n6564 , n6561 , n6563 );
xor ( n6565 , n489 , n509 );
nand ( n6566 , n1859 , n6565 );
nand ( n6567 , n6564 , n6566 );
not ( n6568 , n6567 );
xor ( n6569 , n6560 , n6568 );
or ( n6570 , n4692 , n867 );
nand ( n6571 , n6570 , n495 );
xnor ( n6572 , n6569 , n6571 );
xor ( n6573 , n6554 , n6572 );
not ( n6574 , n6573 );
not ( n6575 , n6489 );
nand ( n6576 , n6575 , n6483 );
not ( n6577 , n6576 );
not ( n6578 , n6495 );
or ( n6579 , n6577 , n6578 );
not ( n6580 , n6483 );
nand ( n6581 , n6580 , n6489 );
nand ( n6582 , n6579 , n6581 );
not ( n6583 , n6582 );
not ( n6584 , n6583 );
and ( n6585 , n6574 , n6584 );
and ( n6586 , n6573 , n6583 );
nor ( n6587 , n6585 , n6586 );
not ( n6588 , n6499 );
not ( n6589 , n6466 );
or ( n6590 , n6588 , n6589 );
nand ( n6591 , n6590 , n6475 );
not ( n6592 , n6499 );
nand ( n6593 , n6592 , n6589 );
nand ( n6594 , n6591 , n6593 );
xor ( n6595 , n6587 , n6594 );
not ( n6596 , n6450 );
not ( n6597 , n6500 );
or ( n6598 , n6596 , n6597 );
nand ( n6599 , n6598 , n6506 );
not ( n6600 , n6500 );
nand ( n6601 , n6600 , n6449 );
and ( n6602 , n6599 , n6601 );
nor ( n6603 , n6595 , n6602 );
not ( n6604 , n6603 );
not ( n6605 , n6602 );
not ( n6606 , n6605 );
nand ( n6607 , n6606 , n6595 );
nand ( n6608 , n6604 , n6607 );
not ( n6609 , n6608 );
and ( n6610 , n6609 , n4994 );
and ( n6611 , n6534 , n6610 );
not ( n6612 , n6534 );
not ( n6613 , n6608 );
nor ( n6614 , n6613 , n455 );
and ( n6615 , n6612 , n6614 );
nor ( n6616 , n6611 , n6615 );
nand ( n6617 , n6336 , n6616 );
not ( n6618 , n6617 );
xor ( n6619 , n549 , n6618 );
not ( n6620 , n6619 );
or ( n6621 , n6096 , n6620 );
not ( n6622 , n549 );
not ( n6623 , n6174 );
not ( n6624 , n3656 );
nor ( n6625 , n6624 , n4423 );
nand ( n6626 , n5764 , n6625 , n4418 , n3233 );
nand ( n6627 , n6626 , n4428 , n4420 );
not ( n6628 , n6627 );
or ( n6629 , n6623 , n6628 );
not ( n6630 , n4414 );
and ( n6631 , n6630 , n6174 );
nor ( n6632 , n6631 , n6261 );
nand ( n6633 , n6629 , n6632 );
not ( n6634 , n6633 );
nand ( n6635 , n6266 , n6264 );
nand ( n6636 , n6634 , n6635 );
not ( n6637 , n6636 );
not ( n6638 , n6635 );
and ( n6639 , n6633 , n6638 );
nor ( n6640 , n6639 , n5705 );
not ( n6641 , n6640 );
or ( n6642 , n6637 , n6641 );
not ( n6643 , n6436 );
not ( n6644 , n6643 );
not ( n6645 , n5583 );
or ( n6646 , n6644 , n6645 );
not ( n6647 , n6524 );
nand ( n6648 , n6646 , n6647 );
nand ( n6649 , n6527 , n6529 );
not ( n6650 , n6649 );
and ( n6651 , n6648 , n6650 );
not ( n6652 , n6648 );
and ( n6653 , n6652 , n6649 );
nor ( n6654 , n6651 , n6653 );
nand ( n6655 , n6654 , n793 );
nand ( n6656 , n6642 , n6655 );
not ( n6657 , n6656 );
not ( n6658 , n6657 );
or ( n6659 , n6622 , n6658 );
not ( n6660 , n549 );
nand ( n6661 , n6660 , n6656 );
nand ( n6662 , n6659 , n6661 );
and ( n6663 , n549 , n550 );
nor ( n6664 , n549 , n550 );
nor ( n6665 , n6663 , n6095 , n6664 );
not ( n6666 , n6665 );
not ( n6667 , n6666 );
nand ( n6668 , n6662 , n6667 );
nand ( n6669 , n6621 , n6668 );
not ( n6670 , n552 );
not ( n6671 , n5154 );
not ( n6672 , n4988 );
or ( n6673 , n6671 , n6672 );
not ( n6674 , n5169 );
nand ( n6675 , n6673 , n6674 );
nor ( n6676 , n6436 , n6509 );
nand ( n6677 , n5577 , n6607 , n6676 );
not ( n6678 , n6677 );
and ( n6679 , n6675 , n6678 );
not ( n6680 , n6607 );
not ( n6681 , n6532 );
or ( n6682 , n6680 , n6681 );
buf ( n6683 , n6604 );
nand ( n6684 , n6682 , n6683 );
or ( n6685 , n6679 , n6684 );
not ( n6686 , n6582 );
not ( n6687 , n6573 );
or ( n6688 , n6686 , n6687 );
not ( n6689 , n6583 );
not ( n6690 , n6573 );
not ( n6691 , n6690 );
or ( n6692 , n6689 , n6691 );
nand ( n6693 , n6692 , n6594 );
nand ( n6694 , n6688 , n6693 );
xor ( n6695 , n6535 , n6483 );
and ( n6696 , n6695 , n6540 );
and ( n6697 , n6535 , n6483 );
or ( n6698 , n6696 , n6697 );
not ( n6699 , n6698 );
not ( n6700 , n6541 );
not ( n6701 , n6549 );
or ( n6702 , n6700 , n6701 );
not ( n6703 , n6552 );
not ( n6704 , n6542 );
or ( n6705 , n6703 , n6704 );
nand ( n6706 , n6705 , n6572 );
nand ( n6707 , n6702 , n6706 );
xor ( n6708 , n6699 , n6707 );
not ( n6709 , n6558 );
not ( n6710 , n1481 );
or ( n6711 , n6709 , n6710 );
nand ( n6712 , n1328 , n493 );
nand ( n6713 , n6711 , n6712 );
not ( n6714 , n6713 );
and ( n6715 , n489 , n510 );
not ( n6716 , n6565 );
not ( n6717 , n6562 );
or ( n6718 , n6716 , n6717 );
xnor ( n6719 , n489 , n508 );
not ( n6720 , n6719 );
nand ( n6721 , n6720 , n1859 );
nand ( n6722 , n6718 , n6721 );
xor ( n6723 , n6715 , n6722 );
not ( n6724 , n6537 );
not ( n6725 , n4563 );
or ( n6726 , n6724 , n6725 );
xnor ( n6727 , n491 , n506 );
not ( n6728 , n6727 );
nand ( n6729 , n6728 , n1933 );
nand ( n6730 , n6726 , n6729 );
xor ( n6731 , n6723 , n6730 );
xor ( n6732 , n6714 , n6731 );
not ( n6733 , n6568 );
not ( n6734 , n6571 );
not ( n6735 , n6734 );
or ( n6736 , n6733 , n6735 );
nand ( n6737 , n6736 , n6560 );
nand ( n6738 , n6571 , n6567 );
nand ( n6739 , n6737 , n6738 );
xor ( n6740 , n6732 , n6739 );
not ( n6741 , n6740 );
not ( n6742 , n6741 );
xnor ( n6743 , n6708 , n6742 );
nor ( n6744 , n6694 , n6743 );
not ( n6745 , n6744 );
nand ( n6746 , n6685 , n6745 );
nand ( n6747 , n6743 , n6694 );
buf ( n6748 , n6747 );
not ( n6749 , n6742 );
not ( n6750 , n6698 );
or ( n6751 , n6749 , n6750 );
not ( n6752 , n6741 );
not ( n6753 , n6699 );
or ( n6754 , n6752 , n6753 );
nand ( n6755 , n6754 , n6707 );
nand ( n6756 , n6751 , n6755 );
and ( n6757 , n489 , n509 );
not ( n6758 , n4563 );
or ( n6759 , n6758 , n6727 );
not ( n6760 , n1933 );
and ( n6761 , n491 , n5074 );
not ( n6762 , n491 );
and ( n6763 , n6762 , n505 );
nor ( n6764 , n6761 , n6763 );
or ( n6765 , n6760 , n6764 );
nand ( n6766 , n6759 , n6765 );
xor ( n6767 , n6757 , n6766 );
not ( n6768 , n1327 );
not ( n6769 , n5532 );
or ( n6770 , n6768 , n6769 );
nand ( n6771 , n6770 , n493 );
xor ( n6772 , n6767 , n6771 );
not ( n6773 , n6562 );
or ( n6774 , n6773 , n6719 );
not ( n6775 , n1859 );
xnor ( n6776 , n507 , n489 );
or ( n6777 , n6775 , n6776 );
nand ( n6778 , n6774 , n6777 );
and ( n6779 , n6778 , n6713 );
not ( n6780 , n6778 );
and ( n6781 , n6780 , n6714 );
nor ( n6782 , n6779 , n6781 );
xor ( n6783 , n6715 , n6722 );
and ( n6784 , n6783 , n6730 );
and ( n6785 , n6715 , n6722 );
or ( n6786 , n6784 , n6785 );
and ( n6787 , n6782 , n6786 );
not ( n6788 , n6782 );
not ( n6789 , n6786 );
and ( n6790 , n6788 , n6789 );
or ( n6791 , n6787 , n6790 );
xor ( n6792 , n6772 , n6791 );
xor ( n6793 , n6714 , n6731 );
and ( n6794 , n6793 , n6739 );
and ( n6795 , n6714 , n6731 );
or ( n6796 , n6794 , n6795 );
xnor ( n6797 , n6792 , n6796 );
nor ( n6798 , n6756 , n6797 );
not ( n6799 , n6798 );
nand ( n6800 , n6756 , n6797 );
and ( n6801 , n6748 , n6799 , n6800 , n793 );
and ( n6802 , n6746 , n6801 );
and ( n6803 , n6748 , n6746 );
not ( n6804 , n6799 );
not ( n6805 , n6800 );
or ( n6806 , n6804 , n6805 );
nand ( n6807 , n6806 , n793 );
nor ( n6808 , n6803 , n6807 );
nor ( n6809 , n6802 , n6808 );
nor ( n6810 , n6324 , n6319 );
nor ( n6811 , n6248 , n6810 );
nand ( n6812 , n6173 , n6811 );
xor ( n6813 , n6273 , n6313 );
and ( n6814 , n6813 , n6318 );
and ( n6815 , n6273 , n6313 );
or ( n6816 , n6814 , n6815 );
xor ( n6817 , n6298 , n6310 );
and ( n6818 , n6817 , n6229 );
and ( n6819 , n6298 , n6310 );
or ( n6820 , n6818 , n6819 );
and ( n6821 , n6284 , n2203 );
and ( n6822 , n2185 , n493 );
nor ( n6823 , n6821 , n6822 );
xor ( n6824 , n6279 , n6288 );
and ( n6825 , n6824 , n6295 );
and ( n6826 , n6279 , n6288 );
or ( n6827 , n6825 , n6826 );
xor ( n6828 , n6823 , n6827 );
and ( n6829 , n2227 , n489 );
not ( n6830 , n2036 );
not ( n6831 , n491 );
not ( n6832 , n2168 );
or ( n6833 , n6831 , n6832 );
nand ( n6834 , n2283 , n2015 );
nand ( n6835 , n6833 , n6834 );
not ( n6836 , n6835 );
or ( n6837 , n6830 , n6836 );
nand ( n6838 , n6306 , n2000 );
nand ( n6839 , n6837 , n6838 );
xor ( n6840 , n6829 , n6839 );
not ( n6841 , n2122 );
not ( n6842 , n6291 );
or ( n6843 , n6841 , n6842 );
xor ( n6844 , n489 , n2270 );
nand ( n6845 , n6844 , n2084 );
nand ( n6846 , n6843 , n6845 );
xor ( n6847 , n6840 , n6846 );
xor ( n6848 , n6828 , n6847 );
xor ( n6849 , n6820 , n6848 );
xor ( n6850 , n6277 , n6296 );
and ( n6851 , n6850 , n6312 );
and ( n6852 , n6277 , n6296 );
or ( n6853 , n6851 , n6852 );
xor ( n6854 , n6849 , n6853 );
nor ( n6855 , n6816 , n6854 );
nor ( n6856 , n6812 , n6855 );
not ( n6857 , n6856 );
not ( n6858 , n4429 );
or ( n6859 , n6857 , n6858 );
not ( n6860 , n6855 );
not ( n6861 , n6811 );
not ( n6862 , n6260 );
or ( n6863 , n6861 , n6862 );
or ( n6864 , n6266 , n6810 );
nand ( n6865 , n6324 , n6319 );
nand ( n6866 , n6864 , n6865 );
not ( n6867 , n6866 );
nand ( n6868 , n6863 , n6867 );
and ( n6869 , n6860 , n6868 );
nand ( n6870 , n6854 , n6816 );
not ( n6871 , n6870 );
nor ( n6872 , n6869 , n6871 );
nand ( n6873 , n6859 , n6872 );
or ( n6874 , n2185 , n2203 );
nand ( n6875 , n6874 , n493 );
not ( n6876 , n2000 );
not ( n6877 , n6835 );
or ( n6878 , n6876 , n6877 );
not ( n6879 , n491 );
not ( n6880 , n2149 );
or ( n6881 , n6879 , n6880 );
nand ( n6882 , n2152 , n2015 );
nand ( n6883 , n6881 , n6882 );
nand ( n6884 , n6883 , n2036 );
nand ( n6885 , n6878 , n6884 );
xor ( n6886 , n6875 , n6885 );
and ( n6887 , n489 , n2193 );
xor ( n6888 , n6886 , n6887 );
not ( n6889 , n2084 );
xor ( n6890 , n489 , n6304 );
not ( n6891 , n6890 );
or ( n6892 , n6889 , n6891 );
nand ( n6893 , n6844 , n2122 );
nand ( n6894 , n6892 , n6893 );
not ( n6895 , n6823 );
xor ( n6896 , n6894 , n6895 );
xor ( n6897 , n6829 , n6839 );
and ( n6898 , n6897 , n6846 );
and ( n6899 , n6829 , n6839 );
or ( n6900 , n6898 , n6899 );
xor ( n6901 , n6896 , n6900 );
xor ( n6902 , n6888 , n6901 );
xor ( n6903 , n6823 , n6827 );
and ( n6904 , n6903 , n6847 );
and ( n6905 , n6823 , n6827 );
or ( n6906 , n6904 , n6905 );
xor ( n6907 , n6902 , n6906 );
xor ( n6908 , n6820 , n6848 );
and ( n6909 , n6908 , n6853 );
and ( n6910 , n6820 , n6848 );
or ( n6911 , n6909 , n6910 );
nor ( n6912 , n6907 , n6911 );
not ( n6913 , n6912 );
nand ( n6914 , n6907 , n6911 );
nand ( n6915 , n6913 , n6914 );
and ( n6916 , n6915 , n455 );
and ( n6917 , n6873 , n6916 );
not ( n6918 , n6873 );
not ( n6919 , n455 );
nor ( n6920 , n6919 , n6915 );
and ( n6921 , n6918 , n6920 );
nor ( n6922 , n6917 , n6921 );
nand ( n6923 , n6809 , n6922 );
not ( n6924 , n551 );
and ( n6925 , n6923 , n6924 );
not ( n6926 , n6923 );
and ( n6927 , n6926 , n551 );
or ( n6928 , n6925 , n6927 );
not ( n6929 , n6928 );
or ( n6930 , n6670 , n6929 );
not ( n6931 , n551 );
not ( n6932 , n793 );
not ( n6933 , n6674 );
nand ( n6934 , n6678 , n6933 );
not ( n6935 , n6677 );
buf ( n6936 , n4988 );
nand ( n6937 , n6935 , n6936 , n5154 );
not ( n6938 , n6595 );
not ( n6939 , n6602 );
and ( n6940 , n6938 , n6939 );
and ( n6941 , n6532 , n6607 );
nor ( n6942 , n6940 , n6941 );
nand ( n6943 , n6934 , n6937 , n6942 );
nand ( n6944 , n6745 , n6747 );
not ( n6945 , n6944 );
and ( n6946 , n6943 , n6945 );
not ( n6947 , n6943 );
and ( n6948 , n6947 , n6944 );
nor ( n6949 , n6946 , n6948 );
not ( n6950 , n6949 );
or ( n6951 , n6932 , n6950 );
not ( n6952 , n6812 );
not ( n6953 , n6952 );
not ( n6954 , n4429 );
or ( n6955 , n6953 , n6954 );
not ( n6956 , n6868 );
nand ( n6957 , n6955 , n6956 );
nand ( n6958 , n6860 , n6870 );
and ( n6959 , n455 , n6958 );
and ( n6960 , n6957 , n6959 );
not ( n6961 , n6957 );
not ( n6962 , n455 );
nor ( n6963 , n6962 , n6958 );
and ( n6964 , n6961 , n6963 );
nor ( n6965 , n6960 , n6964 );
nand ( n6966 , n6951 , n6965 );
buf ( n6967 , n6966 );
not ( n6968 , n6967 );
not ( n6969 , n6968 );
or ( n6970 , n6931 , n6969 );
nand ( n6971 , n6967 , n6924 );
nand ( n6972 , n6970 , n6971 );
not ( n6973 , n552 );
and ( n6974 , n6973 , n551 );
nand ( n6975 , n6972 , n6974 );
nand ( n6976 , n6930 , n6975 );
xor ( n6977 , n6669 , n6976 );
not ( n6978 , n549 );
not ( n6979 , n548 );
or ( n6980 , n6978 , n6979 );
or ( n6981 , n548 , n549 );
nand ( n6982 , n6980 , n6981 );
not ( n6983 , n6982 );
not ( n6984 , n6983 );
not ( n6985 , n6626 );
nand ( n6986 , n4428 , n4420 );
nor ( n6987 , n6985 , n6986 );
not ( n6988 , n2714 );
or ( n6989 , n6987 , n6988 );
not ( n6990 , n2715 );
nor ( n6991 , n4414 , n6988 );
nor ( n6992 , n6990 , n6991 );
nand ( n6993 , n6989 , n6992 );
not ( n6994 , n6172 );
nand ( n6995 , n6103 , n6171 );
nand ( n6996 , n6994 , n6995 );
nand ( n6997 , n6996 , n455 );
nor ( n6998 , n6993 , n6997 );
not ( n6999 , n6998 );
not ( n7000 , n5561 );
not ( n7001 , n5583 );
or ( n7002 , n7000 , n7001 );
nand ( n7003 , n7002 , n5563 );
not ( n7004 , n7003 );
nand ( n7005 , n6435 , n6523 );
not ( n7006 , n7005 );
nor ( n7007 , n7006 , n455 );
nand ( n7008 , n7004 , n7007 );
nor ( n7009 , n7005 , n455 );
nand ( n7010 , n7003 , n7009 );
not ( n7011 , n455 );
nor ( n7012 , n7011 , n6996 );
nand ( n7013 , n7012 , n6993 );
nand ( n7014 , n6999 , n7008 , n7010 , n7013 );
not ( n7015 , n7014 );
not ( n7016 , n7015 );
and ( n7017 , n547 , n7016 );
not ( n7018 , n547 );
not ( n7019 , n7015 );
not ( n7020 , n7019 );
and ( n7021 , n7018 , n7020 );
or ( n7022 , n7017 , n7021 );
not ( n7023 , n7022 );
or ( n7024 , n6984 , n7023 );
xor ( n7025 , n548 , n547 );
and ( n7026 , n7025 , n6982 );
and ( n7027 , n5588 , n547 );
not ( n7028 , n5588 );
not ( n7029 , n547 );
and ( n7030 , n7028 , n7029 );
nor ( n7031 , n7027 , n7030 );
nand ( n7032 , n7026 , n7031 );
nand ( n7033 , n7024 , n7032 );
xor ( n7034 , n6977 , n7033 );
xor ( n7035 , n6094 , n7034 );
not ( n7036 , n6972 );
not ( n7037 , n552 );
or ( n7038 , n7036 , n7037 );
not ( n7039 , n6618 );
buf ( n7040 , n6974 );
nand ( n7041 , n7039 , n7040 );
nand ( n7042 , n7038 , n7041 );
not ( n7043 , n5595 );
not ( n7044 , n6081 );
or ( n7045 , n7043 , n7044 );
not ( n7046 , n545 );
not ( n7047 , n5891 );
not ( n7048 , n7047 );
or ( n7049 , n7046 , n7048 );
nand ( n7050 , n5891 , n4666 );
nand ( n7051 , n7049 , n7050 );
nand ( n7052 , n7051 , n5339 );
nand ( n7053 , n7045 , n7052 );
not ( n7054 , n5697 );
not ( n7055 , n5989 );
or ( n7056 , n7054 , n7055 );
not ( n7057 , n537 );
or ( n7058 , n7057 , n6012 );
nand ( n7059 , n6012 , n5605 );
nand ( n7060 , n7058 , n7059 );
nand ( n7061 , n7060 , n5609 );
nand ( n7062 , n7056 , n7061 );
not ( n7063 , n7062 );
not ( n7064 , n793 );
nand ( n7065 , n6001 , n1301 );
xor ( n7066 , n7065 , n5998 );
not ( n7067 , n7066 );
or ( n7068 , n7064 , n7067 );
and ( n7069 , n4432 , n4138 );
nor ( n7070 , n7069 , n4433 );
not ( n7071 , n7070 );
buf ( n7072 , n4314 );
nand ( n7073 , n4143 , n4169 );
buf ( n7074 , n7073 );
nand ( n7075 , n7072 , n7074 );
or ( n7076 , n7071 , n7075 );
not ( n7077 , n7070 );
nand ( n7078 , n7077 , n7075 );
nand ( n7079 , n7076 , n7078 , n455 );
nand ( n7080 , n7068 , n7079 );
buf ( n7081 , n7080 );
not ( n7082 , n7081 );
nand ( n7083 , n7082 , n537 );
nor ( n7084 , n7063 , n7083 );
not ( n7085 , n4659 );
not ( n7086 , n5982 );
or ( n7087 , n7085 , n7086 );
not ( n7088 , n5913 );
and ( n7089 , n539 , n7088 );
not ( n7090 , n539 );
and ( n7091 , n7090 , n5913 );
nor ( n7092 , n7089 , n7091 );
not ( n7093 , n7092 );
nand ( n7094 , n7093 , n4450 );
nand ( n7095 , n7087 , n7094 );
xor ( n7096 , n7084 , n7095 );
xor ( n7097 , n5995 , n6015 );
xor ( n7098 , n7096 , n7097 );
xor ( n7099 , n7053 , n7098 );
not ( n7100 , n6983 );
and ( n7101 , n5466 , n547 );
not ( n7102 , n5466 );
and ( n7103 , n7102 , n7029 );
nor ( n7104 , n7101 , n7103 );
not ( n7105 , n7104 );
or ( n7106 , n7100 , n7105 );
and ( n7107 , n547 , n5325 );
not ( n7108 , n547 );
buf ( n7109 , n5321 );
and ( n7110 , n7108 , n7109 );
nor ( n7111 , n7107 , n7110 );
not ( n7112 , n7111 );
nand ( n7113 , n7112 , n7026 );
nand ( n7114 , n7106 , n7113 );
and ( n7115 , n7099 , n7114 );
and ( n7116 , n7053 , n7098 );
or ( n7117 , n7115 , n7116 );
xor ( n7118 , n7042 , n7117 );
xor ( n7119 , n7084 , n7095 );
and ( n7120 , n7119 , n7097 );
and ( n7121 , n7084 , n7095 );
or ( n7122 , n7120 , n7121 );
not ( n7123 , n6983 );
not ( n7124 , n7031 );
or ( n7125 , n7123 , n7124 );
not ( n7126 , n7026 );
not ( n7127 , n7126 );
nand ( n7128 , n7104 , n7127 );
nand ( n7129 , n7125 , n7128 );
xor ( n7130 , n7122 , n7129 );
not ( n7131 , n7083 );
not ( n7132 , n7062 );
not ( n7133 , n7132 );
or ( n7134 , n7131 , n7133 );
not ( n7135 , n7083 );
nand ( n7136 , n7135 , n7062 );
nand ( n7137 , n7134 , n7136 );
not ( n7138 , n7092 );
not ( n7139 , n5970 );
and ( n7140 , n7138 , n7139 );
not ( n7141 , n539 );
not ( n7142 , n5644 );
or ( n7143 , n7141 , n7142 );
not ( n7144 , n793 );
not ( n7145 , n5624 );
or ( n7146 , n7144 , n7145 );
nand ( n7147 , n7146 , n5643 );
not ( n7148 , n7147 );
nand ( n7149 , n7148 , n4477 );
nand ( n7150 , n7143 , n7149 );
and ( n7151 , n7150 , n4450 );
nor ( n7152 , n7140 , n7151 );
nor ( n7153 , n7137 , n7152 );
not ( n7154 , n5330 );
not ( n7155 , n6061 );
or ( n7156 , n7154 , n7155 );
not ( n7157 , n5146 );
not ( n7158 , n4655 );
or ( n7159 , n7157 , n7158 );
nand ( n7160 , n4650 , n543 );
nand ( n7161 , n7159 , n7160 );
nand ( n7162 , n7161 , n4671 );
nand ( n7163 , n7156 , n7162 );
xor ( n7164 , n7153 , n7163 );
not ( n7165 , n5786 );
not ( n7166 , n6070 );
or ( n7167 , n7165 , n7166 );
and ( n7168 , n5734 , n5969 );
not ( n7169 , n5734 );
and ( n7170 , n7169 , n5943 );
nor ( n7171 , n7168 , n7170 );
nand ( n7172 , n7171 , n5747 );
nand ( n7173 , n7167 , n7172 );
and ( n7174 , n7164 , n7173 );
and ( n7175 , n7153 , n7163 );
or ( n7176 , n7174 , n7175 );
xor ( n7177 , n7130 , n7176 );
and ( n7178 , n7118 , n7177 );
and ( n7179 , n7042 , n7117 );
or ( n7180 , n7178 , n7179 );
and ( n7181 , n7035 , n7180 );
and ( n7182 , n6094 , n7034 );
or ( n7183 , n7181 , n7182 );
xor ( n7184 , n6092 , n7183 );
xor ( n7185 , n6669 , n6976 );
and ( n7186 , n7185 , n7033 );
and ( n7187 , n6669 , n6976 );
or ( n7188 , n7186 , n7187 );
not ( n7189 , n6095 );
not ( n7190 , n549 );
nor ( n7191 , n7189 , n7190 );
not ( n7192 , n7191 );
not ( n7193 , n7192 );
not ( n7194 , n6967 );
not ( n7195 , n7194 );
or ( n7196 , n7193 , n7195 );
nor ( n7197 , n7189 , n549 );
or ( n7198 , n7194 , n7197 );
nand ( n7199 , n7196 , n7198 );
nand ( n7200 , n6619 , n6667 );
nand ( n7201 , n7199 , n7200 );
not ( n7202 , n6974 );
not ( n7203 , n6928 );
or ( n7204 , n7202 , n7203 );
not ( n7205 , n6924 );
not ( n7206 , n6816 );
not ( n7207 , n6854 );
and ( n7208 , n7206 , n7207 );
nor ( n7209 , n7208 , n6912 );
not ( n7210 , n7209 );
nor ( n7211 , n7210 , n6812 );
not ( n7212 , n7211 );
not ( n7213 , n4429 );
or ( n7214 , n7212 , n7213 );
and ( n7215 , n6868 , n7209 );
nor ( n7216 , n6911 , n6907 );
or ( n7217 , n7216 , n6870 );
nand ( n7218 , n7217 , n6914 );
nor ( n7219 , n7215 , n7218 );
nand ( n7220 , n7214 , n7219 );
not ( n7221 , n7220 );
xor ( n7222 , n6888 , n6901 );
and ( n7223 , n7222 , n6906 );
and ( n7224 , n6888 , n6901 );
or ( n7225 , n7223 , n7224 );
xor ( n7226 , n6875 , n6885 );
and ( n7227 , n7226 , n6887 );
and ( n7228 , n6875 , n6885 );
or ( n7229 , n7227 , n7228 );
not ( n7230 , n2122 );
not ( n7231 , n6890 );
or ( n7232 , n7230 , n7231 );
not ( n7233 , n489 );
not ( n7234 , n2168 );
or ( n7235 , n7233 , n7234 );
nand ( n7236 , n2283 , n1949 );
nand ( n7237 , n7235 , n7236 );
nand ( n7238 , n7237 , n2084 );
nand ( n7239 , n7232 , n7238 );
and ( n7240 , n489 , n2270 );
xor ( n7241 , n7239 , n7240 );
not ( n7242 , n6883 );
not ( n7243 , n7242 );
not ( n7244 , n1999 );
and ( n7245 , n7243 , n7244 );
and ( n7246 , n2036 , n491 );
nor ( n7247 , n7245 , n7246 );
xor ( n7248 , n7241 , n7247 );
xor ( n7249 , n7229 , n7248 );
xor ( n7250 , n6894 , n6895 );
and ( n7251 , n7250 , n6900 );
and ( n7252 , n6894 , n6895 );
or ( n7253 , n7251 , n7252 );
xor ( n7254 , n7249 , n7253 );
or ( n7255 , n7225 , n7254 );
nand ( n7256 , n7225 , n7254 );
nand ( n7257 , n7255 , n7256 );
and ( n7258 , n7257 , n455 );
nand ( n7259 , n7221 , n7258 );
nor ( n7260 , n6744 , n6798 );
not ( n7261 , n7260 );
not ( n7262 , n6943 );
or ( n7263 , n7261 , n7262 );
or ( n7264 , n6747 , n6798 );
nand ( n7265 , n7264 , n6800 );
not ( n7266 , n7265 );
nand ( n7267 , n7263 , n7266 );
not ( n7268 , n7267 );
not ( n7269 , n6778 );
nand ( n7270 , n7269 , n6714 );
not ( n7271 , n7270 );
not ( n7272 , n6786 );
or ( n7273 , n7271 , n7272 );
nand ( n7274 , n6713 , n6778 );
nand ( n7275 , n7273 , n7274 );
and ( n7276 , n508 , n489 );
xor ( n7277 , n489 , n506 );
not ( n7278 , n7277 );
not ( n7279 , n1859 );
or ( n7280 , n7278 , n7279 );
not ( n7281 , n6776 );
nand ( n7282 , n7281 , n6562 );
nand ( n7283 , n7280 , n7282 );
xor ( n7284 , n7276 , n7283 );
not ( n7285 , n6758 );
not ( n7286 , n6764 );
and ( n7287 , n7285 , n7286 );
and ( n7288 , n1933 , n491 );
nor ( n7289 , n7287 , n7288 );
xor ( n7290 , n7284 , n7289 );
xor ( n7291 , n6757 , n6766 );
and ( n7292 , n7291 , n6771 );
and ( n7293 , n6757 , n6766 );
or ( n7294 , n7292 , n7293 );
and ( n7295 , n7290 , n7294 );
not ( n7296 , n7290 );
not ( n7297 , n7294 );
and ( n7298 , n7296 , n7297 );
nor ( n7299 , n7295 , n7298 );
xor ( n7300 , n7275 , n7299 );
not ( n7301 , n7300 );
not ( n7302 , n6796 );
not ( n7303 , n7302 );
not ( n7304 , n6772 );
not ( n7305 , n7304 );
and ( n7306 , n7303 , n7305 );
nand ( n7307 , n7302 , n7304 );
not ( n7308 , n6791 );
and ( n7309 , n7307 , n7308 );
nor ( n7310 , n7306 , n7309 );
nand ( n7311 , n7301 , n7310 );
not ( n7312 , n7300 );
nor ( n7313 , n7312 , n7310 );
not ( n7314 , n7313 );
nand ( n7315 , n7311 , n7314 );
not ( n7316 , n7315 );
nor ( n7317 , n7316 , n455 );
nand ( n7318 , n7268 , n7317 );
not ( n7319 , n7257 );
and ( n7320 , n7319 , n455 );
nand ( n7321 , n7220 , n7320 );
not ( n7322 , n4994 );
nor ( n7323 , n7322 , n7315 );
nand ( n7324 , n7323 , n7267 );
nand ( n7325 , n7259 , n7318 , n7321 , n7324 );
not ( n7326 , n7325 );
not ( n7327 , n7326 );
or ( n7328 , n7205 , n7327 );
or ( n7329 , n7326 , n6924 );
nand ( n7330 , n7328 , n7329 );
nand ( n7331 , n7330 , n552 );
nand ( n7332 , n7204 , n7331 );
xor ( n7333 , n7201 , n7332 );
not ( n7334 , n7127 );
not ( n7335 , n7022 );
or ( n7336 , n7334 , n7335 );
not ( n7337 , n6640 );
not ( n7338 , n6636 );
or ( n7339 , n7337 , n7338 );
nand ( n7340 , n7339 , n6655 );
not ( n7341 , n7340 );
and ( n7342 , n547 , n7341 );
not ( n7343 , n547 );
and ( n7344 , n7343 , n6656 );
or ( n7345 , n7342 , n7344 );
nand ( n7346 , n7345 , n6983 );
nand ( n7347 , n7336 , n7346 );
xor ( n7348 , n7333 , n7347 );
xor ( n7349 , n7188 , n7348 );
xor ( n7350 , n5968 , n6027 );
xor ( n7351 , n7350 , n6040 );
xor ( n7352 , n7122 , n7129 );
and ( n7353 , n7352 , n7176 );
and ( n7354 , n7122 , n7129 );
or ( n7355 , n7353 , n7354 );
xor ( n7356 , n7351 , n7355 );
xor ( n7357 , n5984 , n6016 );
xor ( n7358 , n7357 , n6024 );
xor ( n7359 , n6065 , n6074 );
xor ( n7360 , n7359 , n6085 );
xor ( n7361 , n7358 , n7360 );
not ( n7362 , n6667 );
and ( n7363 , n549 , n7015 );
not ( n7364 , n549 );
and ( n7365 , n7364 , n7019 );
nor ( n7366 , n7363 , n7365 );
not ( n7367 , n7366 );
or ( n7368 , n7362 , n7367 );
nand ( n7369 , n6662 , n6095 );
nand ( n7370 , n7368 , n7369 );
and ( n7371 , n7361 , n7370 );
and ( n7372 , n7358 , n7360 );
or ( n7373 , n7371 , n7372 );
and ( n7374 , n7356 , n7373 );
and ( n7375 , n7351 , n7355 );
or ( n7376 , n7374 , n7375 );
xor ( n7377 , n7349 , n7376 );
xor ( n7378 , n7184 , n7377 );
not ( n7379 , n7378 );
xor ( n7380 , n7351 , n7355 );
xor ( n7381 , n7380 , n7373 );
not ( n7382 , n5785 );
not ( n7383 , n7171 );
or ( n7384 , n7382 , n7383 );
not ( n7385 , n5822 );
not ( n7386 , n7385 );
not ( n7387 , n5734 );
or ( n7388 , n7386 , n7387 );
nand ( n7389 , n5824 , n541 );
nand ( n7390 , n7388 , n7389 );
nand ( n7391 , n7390 , n5747 );
nand ( n7392 , n7384 , n7391 );
not ( n7393 , n5330 );
not ( n7394 , n7161 );
or ( n7395 , n7393 , n7394 );
nand ( n7396 , n4670 , n543 );
not ( n7397 , n7396 );
not ( n7398 , n4473 );
and ( n7399 , n7397 , n7398 );
buf ( n7400 , n4473 );
not ( n7401 , n4670 );
nor ( n7402 , n7401 , n543 );
and ( n7403 , n7400 , n7402 );
nor ( n7404 , n7399 , n7403 );
nand ( n7405 , n7395 , n7404 );
xor ( n7406 , n7392 , n7405 );
not ( n7407 , n5609 );
not ( n7408 , n5605 );
not ( n7409 , n7081 );
not ( n7410 , n7409 );
or ( n7411 , n7408 , n7410 );
nand ( n7412 , n537 , n7081 );
nand ( n7413 , n7411 , n7412 );
not ( n7414 , n7413 );
or ( n7415 , n7407 , n7414 );
nand ( n7416 , n7060 , n5697 );
nand ( n7417 , n7415 , n7416 );
not ( n7418 , n1172 );
nand ( n7419 , n7418 , n1243 );
not ( n7420 , n455 );
nand ( n7421 , n7419 , n1231 , n1239 , n7420 );
nand ( n7422 , n4172 , n4198 );
not ( n7423 , n7422 );
not ( n7424 , n4199 );
not ( n7425 , n4306 );
not ( n7426 , n4310 );
or ( n7427 , n7425 , n7426 );
nand ( n7428 , n7427 , n4309 );
nand ( n7429 , n7424 , n7428 );
not ( n7430 , n7429 );
or ( n7431 , n7423 , n7430 );
nor ( n7432 , n7420 , n4170 );
and ( n7433 , n7073 , n7432 );
nand ( n7434 , n7431 , n7433 );
not ( n7435 , n4170 );
nand ( n7436 , n7435 , n7073 );
nand ( n7437 , n7436 , n7422 , n455 , n7429 );
not ( n7438 , n7419 );
nand ( n7439 , n1231 , n1239 );
nand ( n7440 , n7438 , n7439 , n7420 );
nand ( n7441 , n7421 , n7434 , n7437 , n7440 );
not ( n7442 , n7441 );
not ( n7443 , n7442 );
not ( n7444 , n7443 );
and ( n7445 , n7444 , n537 );
xor ( n7446 , n7417 , n7445 );
not ( n7447 , n4659 );
not ( n7448 , n7150 );
or ( n7449 , n7447 , n7448 );
not ( n7450 , n539 );
not ( n7451 , n5726 );
or ( n7452 , n7450 , n7451 );
nand ( n7453 , n5727 , n4477 );
nand ( n7454 , n7452 , n7453 );
nand ( n7455 , n7454 , n4450 );
nand ( n7456 , n7449 , n7455 );
and ( n7457 , n7446 , n7456 );
and ( n7458 , n7417 , n7445 );
or ( n7459 , n7457 , n7458 );
and ( n7460 , n7406 , n7459 );
and ( n7461 , n7392 , n7405 );
or ( n7462 , n7460 , n7461 );
xor ( n7463 , n7153 , n7163 );
xor ( n7464 , n7463 , n7173 );
xor ( n7465 , n7462 , n7464 );
not ( n7466 , n6095 );
not ( n7467 , n7366 );
or ( n7468 , n7466 , n7467 );
not ( n7469 , n5588 );
not ( n7470 , n7469 );
nor ( n7471 , n6666 , n549 );
and ( n7472 , n7470 , n7471 );
nor ( n7473 , n6666 , n7190 );
and ( n7474 , n7469 , n7473 );
nor ( n7475 , n7472 , n7474 );
nand ( n7476 , n7468 , n7475 );
and ( n7477 , n7465 , n7476 );
and ( n7478 , n7462 , n7464 );
or ( n7479 , n7477 , n7478 );
xor ( n7480 , n7358 , n7360 );
xor ( n7481 , n7480 , n7370 );
xor ( n7482 , n7479 , n7481 );
not ( n7483 , n551 );
not ( n7484 , n7340 );
not ( n7485 , n7484 );
or ( n7486 , n7483 , n7485 );
nand ( n7487 , n6656 , n6924 );
nand ( n7488 , n7486 , n7487 );
nand ( n7489 , n7488 , n6974 );
not ( n7490 , n6618 );
nor ( n7491 , n6924 , n6973 );
nand ( n7492 , n7490 , n7491 );
not ( n7493 , n7490 );
nor ( n7494 , n6973 , n551 );
nand ( n7495 , n7493 , n7494 );
nand ( n7496 , n7489 , n7492 , n7495 );
not ( n7497 , n5339 );
not ( n7498 , n545 );
not ( n7499 , n6059 );
not ( n7500 , n7499 );
or ( n7501 , n7498 , n7500 );
not ( n7502 , n6056 );
nand ( n7503 , n7502 , n4666 );
nand ( n7504 , n7501 , n7503 );
not ( n7505 , n7504 );
or ( n7506 , n7497 , n7505 );
nand ( n7507 , n5595 , n7051 );
nand ( n7508 , n7506 , n7507 );
xor ( n7509 , n7137 , n7152 );
xor ( n7510 , n7508 , n7509 );
and ( n7511 , n547 , n5141 );
not ( n7512 , n547 );
and ( n7513 , n7512 , n5145 );
or ( n7514 , n7511 , n7513 );
not ( n7515 , n7514 );
or ( n7516 , n7515 , n7126 );
or ( n7517 , n7111 , n6982 );
nand ( n7518 , n7516 , n7517 );
and ( n7519 , n7510 , n7518 );
and ( n7520 , n7508 , n7509 );
or ( n7521 , n7519 , n7520 );
xor ( n7522 , n7496 , n7521 );
xor ( n7523 , n7053 , n7098 );
xor ( n7524 , n7523 , n7114 );
and ( n7525 , n7522 , n7524 );
and ( n7526 , n7496 , n7521 );
or ( n7527 , n7525 , n7526 );
and ( n7528 , n7482 , n7527 );
and ( n7529 , n7479 , n7481 );
or ( n7530 , n7528 , n7529 );
xor ( n7531 , n7381 , n7530 );
xor ( n7532 , n6094 , n7034 );
xor ( n7533 , n7532 , n7180 );
and ( n7534 , n7531 , n7533 );
and ( n7535 , n7381 , n7530 );
or ( n7536 , n7534 , n7535 );
not ( n7537 , n7536 );
and ( n7538 , n7379 , n7537 );
xor ( n7539 , n7381 , n7530 );
xor ( n7540 , n7539 , n7533 );
not ( n7541 , n7540 );
xor ( n7542 , n7042 , n7117 );
xor ( n7543 , n7542 , n7177 );
not ( n7544 , n5466 );
nand ( n7545 , n7544 , n7473 );
nand ( n7546 , n5589 , n7191 );
nand ( n7547 , n5588 , n7197 );
nand ( n7548 , n5466 , n7471 );
nand ( n7549 , n7545 , n7546 , n7547 , n7548 );
not ( n7550 , n5697 );
not ( n7551 , n7413 );
or ( n7552 , n7550 , n7551 );
not ( n7553 , n537 );
not ( n7554 , n7441 );
or ( n7555 , n7553 , n7554 );
nand ( n7556 , n7442 , n5605 );
nand ( n7557 , n7555 , n7556 );
nand ( n7558 , n7557 , n5609 );
nand ( n7559 , n7552 , n7558 );
buf ( n7560 , n7428 );
nand ( n7561 , n7424 , n7422 );
not ( n7562 , n7561 );
and ( n7563 , n7560 , n7562 );
not ( n7564 , n7560 );
and ( n7565 , n7564 , n7561 );
nor ( n7566 , n7563 , n7565 );
and ( n7567 , n455 , n7566 );
not ( n7568 , n455 );
not ( n7569 , n1119 );
buf ( n7570 , n1111 );
not ( n7571 , n7570 );
or ( n7572 , n7569 , n7571 );
nand ( n7573 , n7572 , n1105 );
nand ( n7574 , n1170 , n1243 );
or ( n7575 , n7573 , n7574 );
nand ( n7576 , n7573 , n7574 );
nand ( n7577 , n7575 , n7576 );
and ( n7578 , n7568 , n7577 );
nor ( n7579 , n7567 , n7578 );
not ( n7580 , n7579 );
and ( n7581 , n7580 , n537 );
xor ( n7582 , n7559 , n7581 );
not ( n7583 , n4660 );
not ( n7584 , n7454 );
or ( n7585 , n7583 , n7584 );
not ( n7586 , n539 );
not ( n7587 , n6012 );
not ( n7588 , n7587 );
or ( n7589 , n7586 , n7588 );
nand ( n7590 , n6012 , n4477 );
nand ( n7591 , n7589 , n7590 );
nand ( n7592 , n7591 , n4450 );
nand ( n7593 , n7585 , n7592 );
and ( n7594 , n7582 , n7593 );
and ( n7595 , n7559 , n7581 );
or ( n7596 , n7594 , n7595 );
not ( n7597 , n541 );
not ( n7598 , n7088 );
or ( n7599 , n7597 , n7598 );
nand ( n7600 , n5734 , n5691 );
nand ( n7601 , n7599 , n7600 );
not ( n7602 , n7601 );
not ( n7603 , n5747 );
or ( n7604 , n7602 , n7603 );
not ( n7605 , n7390 );
not ( n7606 , n5786 );
or ( n7607 , n7605 , n7606 );
nand ( n7608 , n7604 , n7607 );
xor ( n7609 , n7596 , n7608 );
nand ( n7610 , n4669 , n543 );
or ( n7611 , n7610 , n7400 );
not ( n7612 , n4474 );
not ( n7613 , n4669 );
nor ( n7614 , n7613 , n543 );
nand ( n7615 , n7612 , n7614 );
not ( n7616 , n543 );
not ( n7617 , n5943 );
not ( n7618 , n7617 );
or ( n7619 , n7616 , n7618 );
nand ( n7620 , n5943 , n5146 );
nand ( n7621 , n7619 , n7620 );
nand ( n7622 , n7621 , n4671 );
nand ( n7623 , n7611 , n7615 , n7622 );
and ( n7624 , n7609 , n7623 );
and ( n7625 , n7596 , n7608 );
or ( n7626 , n7624 , n7625 );
xor ( n7627 , n7549 , n7626 );
xor ( n7628 , n7417 , n7445 );
xor ( n7629 , n7628 , n7456 );
not ( n7630 , n5595 );
not ( n7631 , n7504 );
or ( n7632 , n7630 , n7631 );
not ( n7633 , n545 );
not ( n7634 , n5731 );
or ( n7635 , n7633 , n7634 );
nand ( n7636 , n4655 , n4666 );
nand ( n7637 , n7635 , n7636 );
nand ( n7638 , n7637 , n5339 );
nand ( n7639 , n7632 , n7638 );
xor ( n7640 , n7629 , n7639 );
not ( n7641 , n7601 );
not ( n7642 , n5784 );
or ( n7643 , n7641 , n7642 );
not ( n7644 , n541 );
not ( n7645 , n7147 );
or ( n7646 , n7644 , n7645 );
nand ( n7647 , n5734 , n5835 , n5643 );
nand ( n7648 , n7646 , n7647 );
nand ( n7649 , n7648 , n5747 );
nand ( n7650 , n7643 , n7649 );
not ( n7651 , n5697 );
not ( n7652 , n7557 );
or ( n7653 , n7651 , n7652 );
and ( n7654 , n7580 , n537 );
not ( n7655 , n7580 );
and ( n7656 , n7655 , n7057 );
nor ( n7657 , n7654 , n7656 );
nand ( n7658 , n7657 , n5609 );
nand ( n7659 , n7653 , n7658 );
not ( n7660 , n455 );
not ( n7661 , n4306 );
not ( n7662 , n4310 );
or ( n7663 , n7661 , n7662 );
nand ( n7664 , n7663 , n4308 );
not ( n7665 , n4268 );
not ( n7666 , n4293 );
or ( n7667 , n7665 , n7666 );
nand ( n7668 , n7667 , n4298 );
not ( n7669 , n7668 );
and ( n7670 , n7664 , n7669 );
not ( n7671 , n7664 );
and ( n7672 , n7671 , n7668 );
nor ( n7673 , n7670 , n7672 );
not ( n7674 , n7673 );
or ( n7675 , n7660 , n7674 );
not ( n7676 , n1087 );
not ( n7677 , n7676 );
not ( n7678 , n1117 );
not ( n7679 , n1093 );
and ( n7680 , n7678 , n7679 );
and ( n7681 , n1117 , n1093 );
nor ( n7682 , n7680 , n7681 );
not ( n7683 , n7682 );
not ( n7684 , n7683 );
or ( n7685 , n7677 , n7684 );
not ( n7686 , n7676 );
nand ( n7687 , n7686 , n7682 );
nand ( n7688 , n7685 , n7687 );
and ( n7689 , n7688 , n7570 );
not ( n7690 , n7688 );
not ( n7691 , n7570 );
and ( n7692 , n7690 , n7691 );
nor ( n7693 , n7689 , n7692 );
nand ( n7694 , n7693 , n793 );
nand ( n7695 , n7675 , n7694 );
buf ( n7696 , n7695 );
buf ( n7697 , n7696 );
and ( n7698 , n7697 , n537 );
xor ( n7699 , n7659 , n7698 );
not ( n7700 , n4660 );
not ( n7701 , n7591 );
or ( n7702 , n7700 , n7701 );
or ( n7703 , n539 , n7081 );
nand ( n7704 , n7081 , n539 );
nand ( n7705 , n7703 , n7704 );
nand ( n7706 , n7705 , n4450 );
nand ( n7707 , n7702 , n7706 );
and ( n7708 , n7699 , n7707 );
and ( n7709 , n7659 , n7698 );
or ( n7710 , n7708 , n7709 );
xor ( n7711 , n7650 , n7710 );
not ( n7712 , n4671 );
not ( n7713 , n543 );
not ( n7714 , n7385 );
not ( n7715 , n7714 );
or ( n7716 , n7713 , n7715 );
nand ( n7717 , n7385 , n5146 );
nand ( n7718 , n7716 , n7717 );
not ( n7719 , n7718 );
or ( n7720 , n7712 , n7719 );
nand ( n7721 , n7621 , n5330 );
nand ( n7722 , n7720 , n7721 );
and ( n7723 , n7711 , n7722 );
and ( n7724 , n7650 , n7710 );
or ( n7725 , n7723 , n7724 );
and ( n7726 , n7640 , n7725 );
and ( n7727 , n7629 , n7639 );
or ( n7728 , n7726 , n7727 );
and ( n7729 , n7627 , n7728 );
and ( n7730 , n7549 , n7626 );
or ( n7731 , n7729 , n7730 );
xor ( n7732 , n7462 , n7464 );
xor ( n7733 , n7732 , n7476 );
xor ( n7734 , n7731 , n7733 );
xor ( n7735 , n7392 , n7405 );
xor ( n7736 , n7735 , n7459 );
not ( n7737 , n6974 );
and ( n7738 , n7016 , n551 );
not ( n7739 , n7016 );
and ( n7740 , n7739 , n6924 );
or ( n7741 , n7738 , n7740 );
not ( n7742 , n7741 );
or ( n7743 , n7737 , n7742 );
nand ( n7744 , n7488 , n552 );
nand ( n7745 , n7743 , n7744 );
xor ( n7746 , n7736 , n7745 );
xor ( n7747 , n7508 , n7509 );
xor ( n7748 , n7747 , n7518 );
and ( n7749 , n7746 , n7748 );
and ( n7750 , n7736 , n7745 );
or ( n7751 , n7749 , n7750 );
and ( n7752 , n7734 , n7751 );
and ( n7753 , n7731 , n7733 );
or ( n7754 , n7752 , n7753 );
xor ( n7755 , n7543 , n7754 );
xor ( n7756 , n7479 , n7481 );
xor ( n7757 , n7756 , n7527 );
and ( n7758 , n7755 , n7757 );
and ( n7759 , n7543 , n7754 );
or ( n7760 , n7758 , n7759 );
not ( n7761 , n7760 );
and ( n7762 , n7541 , n7761 );
nor ( n7763 , n7538 , n7762 );
not ( n7764 , n7763 );
xor ( n7765 , n7736 , n7745 );
xor ( n7766 , n7765 , n7748 );
not ( n7767 , n552 );
not ( n7768 , n7741 );
or ( n7769 , n7767 , n7768 );
not ( n7770 , n551 );
not ( n7771 , n7469 );
or ( n7772 , n7770 , n7771 );
nand ( n7773 , n5588 , n6924 );
nand ( n7774 , n7772 , n7773 );
nand ( n7775 , n7774 , n6974 );
nand ( n7776 , n7769 , n7775 );
not ( n7777 , n6983 );
not ( n7778 , n7514 );
or ( n7779 , n7777 , n7778 );
not ( n7780 , n6033 );
buf ( n7781 , n7780 );
nor ( n7782 , n7126 , n547 );
and ( n7783 , n7781 , n7782 );
not ( n7784 , n7780 );
not ( n7785 , n547 );
nor ( n7786 , n7785 , n7126 );
and ( n7787 , n7784 , n7786 );
nor ( n7788 , n7783 , n7787 );
nand ( n7789 , n7779 , n7788 );
xor ( n7790 , n7559 , n7581 );
xor ( n7791 , n7790 , n7593 );
nand ( n7792 , n7499 , n7786 );
not ( n7793 , n6033 );
nor ( n7794 , n6982 , n547 );
nand ( n7795 , n7793 , n7794 );
nand ( n7796 , n6059 , n7782 );
nand ( n7797 , n6983 , n547 );
not ( n7798 , n7797 );
nand ( n7799 , n7798 , n7047 );
nand ( n7800 , n7792 , n7795 , n7796 , n7799 );
xor ( n7801 , n7791 , n7800 );
and ( n7802 , n4473 , n4666 );
not ( n7803 , n4473 );
and ( n7804 , n7803 , n545 );
or ( n7805 , n7802 , n7804 );
not ( n7806 , n7805 );
or ( n7807 , n7806 , n5340 );
not ( n7808 , n7637 );
not ( n7809 , n5595 );
or ( n7810 , n7808 , n7809 );
nand ( n7811 , n7807 , n7810 );
and ( n7812 , n7801 , n7811 );
and ( n7813 , n7791 , n7800 );
or ( n7814 , n7812 , n7813 );
xor ( n7815 , n7789 , n7814 );
xor ( n7816 , n7596 , n7608 );
xor ( n7817 , n7816 , n7623 );
xor ( n7818 , n7815 , n7817 );
xor ( n7819 , n7776 , n7818 );
not ( n7820 , n6974 );
not ( n7821 , n551 );
not ( n7822 , n5467 );
or ( n7823 , n7821 , n7822 );
nand ( n7824 , n6924 , n5466 );
nand ( n7825 , n7823 , n7824 );
not ( n7826 , n7825 );
or ( n7827 , n7820 , n7826 );
nand ( n7828 , n7774 , n552 );
nand ( n7829 , n7827 , n7828 );
not ( n7830 , n5330 );
not ( n7831 , n7718 );
or ( n7832 , n7830 , n7831 );
not ( n7833 , n543 );
not ( n7834 , n7088 );
or ( n7835 , n7833 , n7834 );
nand ( n7836 , n5146 , n5691 );
nand ( n7837 , n7835 , n7836 );
nand ( n7838 , n7837 , n4671 );
nand ( n7839 , n7832 , n7838 );
not ( n7840 , n742 );
nand ( n7841 , n7840 , n746 );
not ( n7842 , n709 );
and ( n7843 , n7841 , n7842 );
not ( n7844 , n7841 );
and ( n7845 , n7844 , n709 );
nor ( n7846 , n7843 , n7845 );
nand ( n7847 , n7846 , n793 );
nand ( n7848 , n4267 , n4241 );
not ( n7849 , n7848 );
nor ( n7850 , n4262 , n5791 );
and ( n7851 , n7849 , n7850 );
and ( n7852 , n4262 , n455 );
and ( n7853 , n7852 , n7848 );
nor ( n7854 , n7851 , n7853 );
nand ( n7855 , n7847 , n7854 );
buf ( n7856 , n7855 );
and ( n7857 , n537 , n7856 );
not ( n7858 , n5697 );
not ( n7859 , n537 );
not ( n7860 , n7696 );
not ( n7861 , n7860 );
or ( n7862 , n7859 , n7861 );
nand ( n7863 , n7696 , n5605 );
nand ( n7864 , n7862 , n7863 );
not ( n7865 , n7864 );
or ( n7866 , n7858 , n7865 );
not ( n7867 , n4297 );
not ( n7868 , n4296 );
or ( n7869 , n7867 , n7868 );
nand ( n7870 , n7869 , n4293 );
not ( n7871 , n7870 );
buf ( n7872 , n4268 );
nand ( n7873 , n7871 , n7872 );
not ( n7874 , n7872 );
nand ( n7875 , n7870 , n7874 );
nand ( n7876 , n7873 , n7875 , n455 );
nand ( n7877 , n7876 , n794 );
buf ( n7878 , n7877 );
xor ( n7879 , n537 , n7878 );
nand ( n7880 , n7879 , n5609 );
nand ( n7881 , n7866 , n7880 );
xor ( n7882 , n7857 , n7881 );
not ( n7883 , n5697 );
not ( n7884 , n7879 );
or ( n7885 , n7883 , n7884 );
xor ( n7886 , n537 , n7856 );
nand ( n7887 , n7886 , n5609 );
nand ( n7888 , n7885 , n7887 );
not ( n7889 , n7888 );
not ( n7890 , n5599 );
not ( n7891 , n7856 );
not ( n7892 , n7891 );
or ( n7893 , n7890 , n7892 );
nand ( n7894 , n7893 , n539 );
not ( n7895 , n7856 );
not ( n7896 , n7895 );
and ( n7897 , n7896 , n538 );
nor ( n7898 , n7897 , n5605 );
nand ( n7899 , n7894 , n7898 );
nor ( n7900 , n7889 , n7899 );
and ( n7901 , n7882 , n7900 );
and ( n7902 , n7857 , n7881 );
or ( n7903 , n7901 , n7902 );
not ( n7904 , n5746 );
not ( n7905 , n541 );
not ( n7906 , n7587 );
or ( n7907 , n7905 , n7906 );
nand ( n7908 , n6012 , n5734 );
nand ( n7909 , n7907 , n7908 );
not ( n7910 , n7909 );
or ( n7911 , n7904 , n7910 );
not ( n7912 , n541 );
not ( n7913 , n5726 );
or ( n7914 , n7912 , n7913 );
not ( n7915 , n5712 );
nor ( n7916 , n5723 , n455 );
not ( n7917 , n7916 );
nand ( n7918 , n7915 , n7917 , n5734 );
nand ( n7919 , n7914 , n7918 );
nand ( n7920 , n7919 , n5741 );
nand ( n7921 , n7911 , n7920 );
xor ( n7922 , n7903 , n7921 );
and ( n7923 , n537 , n7878 );
not ( n7924 , n5697 );
not ( n7925 , n7657 );
or ( n7926 , n7924 , n7925 );
nand ( n7927 , n7864 , n5609 );
nand ( n7928 , n7926 , n7927 );
xor ( n7929 , n7923 , n7928 );
not ( n7930 , n4660 );
not ( n7931 , n7705 );
or ( n7932 , n7930 , n7931 );
not ( n7933 , n539 );
not ( n7934 , n7441 );
or ( n7935 , n7933 , n7934 );
nand ( n7936 , n7442 , n4477 );
nand ( n7937 , n7935 , n7936 );
nand ( n7938 , n7937 , n4450 );
nand ( n7939 , n7932 , n7938 );
xor ( n7940 , n7929 , n7939 );
and ( n7941 , n7922 , n7940 );
and ( n7942 , n7903 , n7921 );
or ( n7943 , n7941 , n7942 );
xor ( n7944 , n7839 , n7943 );
not ( n7945 , n6983 );
not ( n7946 , n6056 );
and ( n7947 , n547 , n7946 );
not ( n7948 , n547 );
buf ( n7949 , n6056 );
and ( n7950 , n7948 , n7949 );
nor ( n7951 , n7947 , n7950 );
not ( n7952 , n7951 );
or ( n7953 , n7945 , n7952 );
not ( n7954 , n547 );
not ( n7955 , n5731 );
or ( n7956 , n7954 , n7955 );
not ( n7957 , n547 );
not ( n7958 , n4650 );
nand ( n7959 , n7957 , n7958 );
nand ( n7960 , n7956 , n7959 );
nand ( n7961 , n7960 , n7127 );
nand ( n7962 , n7953 , n7961 );
and ( n7963 , n7944 , n7962 );
and ( n7964 , n7839 , n7943 );
or ( n7965 , n7963 , n7964 );
xor ( n7966 , n7829 , n7965 );
not ( n7967 , n5595 );
not ( n7968 , n7805 );
or ( n7969 , n7967 , n7968 );
and ( n7970 , n5976 , n4666 );
not ( n7971 , n5976 );
and ( n7972 , n7971 , n545 );
or ( n7973 , n7970 , n7972 );
nand ( n7974 , n7973 , n5339 );
nand ( n7975 , n7969 , n7974 );
xor ( n7976 , n7923 , n7928 );
and ( n7977 , n7976 , n7939 );
and ( n7978 , n7923 , n7928 );
or ( n7979 , n7977 , n7978 );
not ( n7980 , n5785 );
not ( n7981 , n7648 );
or ( n7982 , n7980 , n7981 );
nand ( n7983 , n5747 , n7919 );
nand ( n7984 , n7982 , n7983 );
xor ( n7985 , n7979 , n7984 );
xor ( n7986 , n7659 , n7698 );
xor ( n7987 , n7986 , n7707 );
xor ( n7988 , n7985 , n7987 );
xor ( n7989 , n7975 , n7988 );
not ( n7990 , n4670 );
not ( n7991 , n543 );
not ( n7992 , n5836 );
or ( n7993 , n7991 , n7992 );
nand ( n7994 , n5837 , n5146 );
nand ( n7995 , n7993 , n7994 );
not ( n7996 , n7995 );
or ( n7997 , n7990 , n7996 );
nand ( n7998 , n7837 , n5329 );
nand ( n7999 , n7997 , n7998 );
not ( n8000 , n5595 );
not ( n8001 , n7973 );
or ( n8002 , n8000 , n8001 );
not ( n8003 , n545 );
not ( n8004 , n7714 );
or ( n8005 , n8003 , n8004 );
nand ( n8006 , n7385 , n4666 );
nand ( n8007 , n8005 , n8006 );
nand ( n8008 , n8007 , n5339 );
nand ( n8009 , n8002 , n8008 );
xor ( n8010 , n7999 , n8009 );
not ( n8011 , n4660 );
not ( n8012 , n7937 );
or ( n8013 , n8011 , n8012 );
and ( n8014 , n4465 , n7577 );
not ( n8015 , n4465 );
and ( n8016 , n8015 , n7566 );
nor ( n8017 , n8014 , n8016 );
and ( n8018 , n8017 , n539 );
not ( n8019 , n8017 );
and ( n8020 , n8019 , n4477 );
or ( n8021 , n8018 , n8020 );
nand ( n8022 , n8021 , n4450 );
nand ( n8023 , n8013 , n8022 );
xor ( n8024 , n7857 , n7881 );
xor ( n8025 , n8024 , n7900 );
xor ( n8026 , n8023 , n8025 );
not ( n8027 , n5741 );
not ( n8028 , n7909 );
or ( n8029 , n8027 , n8028 );
not ( n8030 , n541 );
not ( n8031 , n7081 );
or ( n8032 , n8030 , n8031 );
nand ( n8033 , n7409 , n5734 );
nand ( n8034 , n8032 , n8033 );
nand ( n8035 , n8034 , n5747 );
nand ( n8036 , n8029 , n8035 );
and ( n8037 , n8026 , n8036 );
and ( n8038 , n8023 , n8025 );
or ( n8039 , n8037 , n8038 );
and ( n8040 , n8010 , n8039 );
and ( n8041 , n7999 , n8009 );
or ( n8042 , n8040 , n8041 );
and ( n8043 , n7989 , n8042 );
and ( n8044 , n7975 , n7988 );
or ( n8045 , n8043 , n8044 );
and ( n8046 , n7966 , n8045 );
and ( n8047 , n7829 , n7965 );
or ( n8048 , n8046 , n8047 );
and ( n8049 , n7819 , n8048 );
and ( n8050 , n7776 , n7818 );
or ( n8051 , n8049 , n8050 );
xor ( n8052 , n7766 , n8051 );
xor ( n8053 , n7789 , n7814 );
and ( n8054 , n8053 , n7817 );
and ( n8055 , n7789 , n7814 );
or ( n8056 , n8054 , n8055 );
xor ( n8057 , n7549 , n7626 );
xor ( n8058 , n8057 , n7728 );
xor ( n8059 , n8056 , n8058 );
not ( n8060 , n6095 );
and ( n8061 , n549 , n5466 );
not ( n8062 , n549 );
and ( n8063 , n8062 , n7544 );
nor ( n8064 , n8061 , n8063 );
not ( n8065 , n8064 );
or ( n8066 , n8060 , n8065 );
not ( n8067 , n549 );
not ( n8068 , n7109 );
not ( n8069 , n8068 );
or ( n8070 , n8067 , n8069 );
not ( n8071 , n549 );
nand ( n8072 , n8071 , n7109 );
nand ( n8073 , n8070 , n8072 );
nand ( n8074 , n8073 , n6667 );
nand ( n8075 , n8066 , n8074 );
xor ( n8076 , n7629 , n7639 );
xor ( n8077 , n8076 , n7725 );
xor ( n8078 , n8075 , n8077 );
xor ( n8079 , n7979 , n7984 );
and ( n8080 , n8079 , n7987 );
and ( n8081 , n7979 , n7984 );
or ( n8082 , n8080 , n8081 );
xor ( n8083 , n7650 , n7710 );
xor ( n8084 , n8083 , n7722 );
xor ( n8085 , n8082 , n8084 );
not ( n8086 , n6667 );
not ( n8087 , n5145 );
and ( n8088 , n549 , n8087 );
not ( n8089 , n549 );
not ( n8090 , n5141 );
and ( n8091 , n8089 , n8090 );
or ( n8092 , n8088 , n8091 );
not ( n8093 , n8092 );
or ( n8094 , n8086 , n8093 );
nand ( n8095 , n8073 , n6095 );
nand ( n8096 , n8094 , n8095 );
and ( n8097 , n8085 , n8096 );
and ( n8098 , n8082 , n8084 );
or ( n8099 , n8097 , n8098 );
and ( n8100 , n8078 , n8099 );
and ( n8101 , n8075 , n8077 );
or ( n8102 , n8100 , n8101 );
xor ( n8103 , n8059 , n8102 );
xor ( n8104 , n8052 , n8103 );
xor ( n8105 , n8075 , n8077 );
xor ( n8106 , n8105 , n8099 );
xor ( n8107 , n7791 , n7800 );
xor ( n8108 , n8107 , n7811 );
not ( n8109 , n6095 );
not ( n8110 , n8092 );
or ( n8111 , n8109 , n8110 );
and ( n8112 , n549 , n7047 );
not ( n8113 , n549 );
and ( n8114 , n8113 , n7793 );
or ( n8115 , n8112 , n8114 );
nand ( n8116 , n8115 , n6667 );
nand ( n8117 , n8111 , n8116 );
xor ( n8118 , n7903 , n7921 );
xor ( n8119 , n8118 , n7940 );
not ( n8120 , n7026 );
xor ( n8121 , n4473 , n547 );
not ( n8122 , n8121 );
or ( n8123 , n8120 , n8122 );
nand ( n8124 , n7960 , n6983 );
nand ( n8125 , n8123 , n8124 );
xor ( n8126 , n8119 , n8125 );
not ( n8127 , n6667 );
not ( n8128 , n549 );
not ( n8129 , n7499 );
or ( n8130 , n8128 , n8129 );
not ( n8131 , n549 );
nand ( n8132 , n8131 , n7946 );
nand ( n8133 , n8130 , n8132 );
not ( n8134 , n8133 );
or ( n8135 , n8127 , n8134 );
nand ( n8136 , n8115 , n6095 );
nand ( n8137 , n8135 , n8136 );
and ( n8138 , n8126 , n8137 );
and ( n8139 , n8119 , n8125 );
or ( n8140 , n8138 , n8139 );
xor ( n8141 , n8117 , n8140 );
not ( n8142 , n551 );
not ( n8143 , n8068 );
or ( n8144 , n8142 , n8143 );
nand ( n8145 , n7109 , n6924 );
nand ( n8146 , n8144 , n8145 );
not ( n8147 , n8146 );
not ( n8148 , n6974 );
or ( n8149 , n8147 , n8148 );
not ( n8150 , n7825 );
or ( n8151 , n8150 , n6973 );
nand ( n8152 , n8149 , n8151 );
and ( n8153 , n8141 , n8152 );
and ( n8154 , n8117 , n8140 );
or ( n8155 , n8153 , n8154 );
xor ( n8156 , n8108 , n8155 );
xor ( n8157 , n8082 , n8084 );
xor ( n8158 , n8157 , n8096 );
and ( n8159 , n8156 , n8158 );
and ( n8160 , n8108 , n8155 );
or ( n8161 , n8159 , n8160 );
xor ( n8162 , n8106 , n8161 );
xor ( n8163 , n7776 , n7818 );
xor ( n8164 , n8163 , n8048 );
and ( n8165 , n8162 , n8164 );
and ( n8166 , n8106 , n8161 );
or ( n8167 , n8165 , n8166 );
nor ( n8168 , n8104 , n8167 );
xor ( n8169 , n8106 , n8161 );
xor ( n8170 , n8169 , n8164 );
xor ( n8171 , n7829 , n7965 );
xor ( n8172 , n8171 , n8045 );
xor ( n8173 , n7839 , n7943 );
xor ( n8174 , n8173 , n7962 );
xor ( n8175 , n7975 , n7988 );
xor ( n8176 , n8175 , n8042 );
xor ( n8177 , n8174 , n8176 );
xnor ( n8178 , n7888 , n7899 );
not ( n8179 , n4660 );
not ( n8180 , n8021 );
or ( n8181 , n8179 , n8180 );
not ( n8182 , n539 );
not ( n8183 , n7860 );
or ( n8184 , n8182 , n8183 );
nand ( n8185 , n7696 , n4477 );
nand ( n8186 , n8184 , n8185 );
nand ( n8187 , n4450 , n8186 );
nand ( n8188 , n8181 , n8187 );
xor ( n8189 , n8178 , n8188 );
buf ( n8190 , n7856 );
and ( n8191 , n8190 , n5697 );
not ( n8192 , n4659 );
not ( n8193 , n8186 );
or ( n8194 , n8192 , n8193 );
not ( n8195 , n539 );
not ( n8196 , n7878 );
not ( n8197 , n8196 );
or ( n8198 , n8195 , n8197 );
nand ( n8199 , n7878 , n4477 );
nand ( n8200 , n8198 , n8199 );
nand ( n8201 , n8200 , n4450 );
nand ( n8202 , n8194 , n8201 );
xor ( n8203 , n8191 , n8202 );
not ( n8204 , n540 );
nand ( n8205 , n8204 , n7891 );
and ( n8206 , n8205 , n541 );
not ( n8207 , n540 );
not ( n8208 , n7856 );
or ( n8209 , n8207 , n8208 );
nand ( n8210 , n8209 , n539 );
nor ( n8211 , n8206 , n8210 );
not ( n8212 , n4660 );
not ( n8213 , n8200 );
or ( n8214 , n8212 , n8213 );
and ( n8215 , n7896 , n5962 );
nor ( n8216 , n7855 , n5964 );
nor ( n8217 , n8215 , n8216 );
nand ( n8218 , n8214 , n8217 );
and ( n8219 , n8211 , n8218 );
and ( n8220 , n8203 , n8219 );
and ( n8221 , n8191 , n8202 );
or ( n8222 , n8220 , n8221 );
and ( n8223 , n8189 , n8222 );
and ( n8224 , n8178 , n8188 );
or ( n8225 , n8223 , n8224 );
not ( n8226 , n4669 );
not ( n8227 , n7995 );
or ( n8228 , n8226 , n8227 );
not ( n8229 , n543 );
nor ( n8230 , n7916 , n5712 );
not ( n8231 , n8230 );
not ( n8232 , n8231 );
or ( n8233 , n8229 , n8232 );
nand ( n8234 , n8230 , n5146 );
nand ( n8235 , n8233 , n8234 );
nand ( n8236 , n8235 , n4670 );
nand ( n8237 , n8228 , n8236 );
xor ( n8238 , n8225 , n8237 );
not ( n8239 , n5595 );
not ( n8240 , n8007 );
or ( n8241 , n8239 , n8240 );
not ( n8242 , n545 );
not ( n8243 , n7088 );
or ( n8244 , n8242 , n8243 );
nand ( n8245 , n5914 , n4666 );
nand ( n8246 , n8244 , n8245 );
nand ( n8247 , n8246 , n5339 );
nand ( n8248 , n8241 , n8247 );
and ( n8249 , n8238 , n8248 );
and ( n8250 , n8225 , n8237 );
or ( n8251 , n8249 , n8250 );
not ( n8252 , n6974 );
not ( n8253 , n551 );
not ( n8254 , n8087 );
or ( n8255 , n8253 , n8254 );
nand ( n8256 , n8090 , n6924 );
nand ( n8257 , n8255 , n8256 );
not ( n8258 , n8257 );
or ( n8259 , n8252 , n8258 );
nand ( n8260 , n8146 , n552 );
nand ( n8261 , n8259 , n8260 );
xor ( n8262 , n8251 , n8261 );
xor ( n8263 , n7999 , n8009 );
xor ( n8264 , n8263 , n8039 );
and ( n8265 , n8262 , n8264 );
and ( n8266 , n8251 , n8261 );
or ( n8267 , n8265 , n8266 );
and ( n8268 , n8177 , n8267 );
and ( n8269 , n8174 , n8176 );
or ( n8270 , n8268 , n8269 );
xor ( n8271 , n8172 , n8270 );
xor ( n8272 , n8108 , n8155 );
xor ( n8273 , n8272 , n8158 );
and ( n8274 , n8271 , n8273 );
and ( n8275 , n8172 , n8270 );
or ( n8276 , n8274 , n8275 );
nand ( n8277 , n8170 , n8276 );
or ( n8278 , n8168 , n8277 );
nand ( n8279 , n8104 , n8167 );
nand ( n8280 , n8278 , n8279 );
not ( n8281 , n8280 );
xor ( n8282 , n7543 , n7754 );
xor ( n8283 , n8282 , n7757 );
xor ( n8284 , n7496 , n7521 );
xor ( n8285 , n8284 , n7524 );
xor ( n8286 , n8056 , n8058 );
and ( n8287 , n8286 , n8102 );
and ( n8288 , n8056 , n8058 );
or ( n8289 , n8287 , n8288 );
xor ( n8290 , n8285 , n8289 );
xor ( n8291 , n7731 , n7733 );
xor ( n8292 , n8291 , n7751 );
and ( n8293 , n8290 , n8292 );
and ( n8294 , n8285 , n8289 );
or ( n8295 , n8293 , n8294 );
nor ( n8296 , n8283 , n8295 );
xor ( n8297 , n8285 , n8289 );
xor ( n8298 , n8297 , n8292 );
xor ( n8299 , n7766 , n8051 );
and ( n8300 , n8299 , n8103 );
and ( n8301 , n7766 , n8051 );
or ( n8302 , n8300 , n8301 );
nor ( n8303 , n8298 , n8302 );
nor ( n8304 , n8296 , n8303 );
not ( n8305 , n8304 );
or ( n8306 , n8281 , n8305 );
not ( n8307 , n8296 );
nand ( n8308 , n8298 , n8302 );
not ( n8309 , n8308 );
and ( n8310 , n8307 , n8309 );
not ( n8311 , n8283 );
not ( n8312 , n8295 );
nor ( n8313 , n8311 , n8312 );
nor ( n8314 , n8310 , n8313 );
nand ( n8315 , n8306 , n8314 );
not ( n8316 , n8315 );
or ( n8317 , n7764 , n8316 );
nor ( n8318 , n7378 , n7536 );
not ( n8319 , n8318 );
nand ( n8320 , n7540 , n7760 );
not ( n8321 , n8320 );
and ( n8322 , n8319 , n8321 );
and ( n8323 , n7378 , n7536 );
nor ( n8324 , n8322 , n8323 );
nand ( n8325 , n8317 , n8324 );
not ( n8326 , n8283 );
nand ( n8327 , n8326 , n8312 );
not ( n8328 , n8298 );
not ( n8329 , n8302 );
nand ( n8330 , n8328 , n8329 );
nand ( n8331 , n8327 , n8330 );
not ( n8332 , n8331 );
not ( n8333 , n8104 );
not ( n8334 , n8167 );
nand ( n8335 , n8333 , n8334 );
not ( n8336 , n8170 );
not ( n8337 , n8276 );
nand ( n8338 , n8336 , n8337 );
nand ( n8339 , n8335 , n8338 );
not ( n8340 , n8339 );
not ( n8341 , n552 );
not ( n8342 , n551 );
not ( n8343 , n7949 );
or ( n8344 , n8342 , n8343 );
nand ( n8345 , n7946 , n6924 );
nand ( n8346 , n8344 , n8345 );
not ( n8347 , n8346 );
or ( n8348 , n8341 , n8347 );
buf ( n8349 , n4651 );
nand ( n8350 , n8349 , n6924 );
nand ( n8351 , n551 , n5731 );
nand ( n8352 , n8350 , n8351 );
nand ( n8353 , n8352 , n6974 );
nand ( n8354 , n8348 , n8353 );
not ( n8355 , n7026 );
and ( n8356 , n547 , n7147 );
not ( n8357 , n547 );
and ( n8358 , n8357 , n5837 );
or ( n8359 , n8356 , n8358 );
not ( n8360 , n8359 );
or ( n8361 , n8355 , n8360 );
and ( n8362 , n5914 , n7029 );
not ( n8363 , n5914 );
and ( n8364 , n8363 , n547 );
or ( n8365 , n8362 , n8364 );
nand ( n8366 , n8365 , n6983 );
nand ( n8367 , n8361 , n8366 );
not ( n8368 , n543 );
not ( n8369 , n7443 );
or ( n8370 , n8368 , n8369 );
nand ( n8371 , n7442 , n5146 );
nand ( n8372 , n8370 , n8371 );
nand ( n8373 , n8372 , n4669 );
not ( n8374 , n543 );
not ( n8375 , n8017 );
or ( n8376 , n8374 , n8375 );
not ( n8377 , n8017 );
nand ( n8378 , n8377 , n5146 );
nand ( n8379 , n8376 , n8378 );
nand ( n8380 , n8379 , n4670 );
nand ( n8381 , n8373 , n8380 );
and ( n8382 , n8190 , n4659 );
not ( n8383 , n5741 );
not ( n8384 , n5734 );
not ( n8385 , n7696 );
or ( n8386 , n8384 , n8385 );
or ( n8387 , n7696 , n4445 );
nand ( n8388 , n8386 , n8387 );
not ( n8389 , n8388 );
or ( n8390 , n8383 , n8389 );
not ( n8391 , n541 );
not ( n8392 , n8196 );
or ( n8393 , n8391 , n8392 );
nand ( n8394 , n7878 , n5734 );
nand ( n8395 , n8393 , n8394 );
nand ( n8396 , n8395 , n5746 );
nand ( n8397 , n8390 , n8396 );
xor ( n8398 , n8382 , n8397 );
not ( n8399 , n5741 );
not ( n8400 , n8395 );
or ( n8401 , n8399 , n8400 );
not ( n8402 , n7856 );
not ( n8403 , n4445 );
or ( n8404 , n8402 , n8403 );
or ( n8405 , n7856 , n4445 );
nand ( n8406 , n8404 , n8405 );
nand ( n8407 , n8406 , n5746 );
nand ( n8408 , n8401 , n8407 );
not ( n8409 , n8408 );
not ( n8410 , n542 );
not ( n8411 , n8410 );
not ( n8412 , n7891 );
or ( n8413 , n8411 , n8412 );
nand ( n8414 , n8413 , n543 );
and ( n8415 , n7896 , n542 );
nor ( n8416 , n8415 , n5734 );
nand ( n8417 , n8414 , n8416 );
nor ( n8418 , n8409 , n8417 );
xor ( n8419 , n8398 , n8418 );
xor ( n8420 , n8381 , n8419 );
not ( n8421 , n5595 );
not ( n8422 , n545 );
not ( n8423 , n6012 );
not ( n8424 , n8423 );
or ( n8425 , n8422 , n8424 );
nand ( n8426 , n6012 , n4666 );
nand ( n8427 , n8425 , n8426 );
not ( n8428 , n8427 );
or ( n8429 , n8421 , n8428 );
not ( n8430 , n545 );
not ( n8431 , n7081 );
or ( n8432 , n8430 , n8431 );
nand ( n8433 , n7409 , n4666 );
nand ( n8434 , n8432 , n8433 );
nand ( n8435 , n8434 , n5339 );
nand ( n8436 , n8429 , n8435 );
and ( n8437 , n8420 , n8436 );
and ( n8438 , n8381 , n8419 );
or ( n8439 , n8437 , n8438 );
xor ( n8440 , n8367 , n8439 );
not ( n8441 , n6095 );
and ( n8442 , n549 , n5959 );
not ( n8443 , n549 );
not ( n8444 , n7617 );
and ( n8445 , n8443 , n8444 );
or ( n8446 , n8442 , n8445 );
not ( n8447 , n8446 );
or ( n8448 , n8441 , n8447 );
not ( n8449 , n549 );
not ( n8450 , n7714 );
or ( n8451 , n8449 , n8450 );
not ( n8452 , n549 );
not ( n8453 , n7714 );
nand ( n8454 , n8452 , n8453 );
nand ( n8455 , n8451 , n8454 );
nand ( n8456 , n8455 , n6667 );
nand ( n8457 , n8448 , n8456 );
and ( n8458 , n8440 , n8457 );
and ( n8459 , n8367 , n8439 );
or ( n8460 , n8458 , n8459 );
xor ( n8461 , n8354 , n8460 );
xor ( n8462 , n8211 , n8218 );
xor ( n8463 , n7580 , n541 );
not ( n8464 , n8463 );
not ( n8465 , n5741 );
or ( n8466 , n8464 , n8465 );
nand ( n8467 , n8388 , n5746 );
nand ( n8468 , n8466 , n8467 );
xor ( n8469 , n8462 , n8468 );
xor ( n8470 , n8382 , n8397 );
and ( n8471 , n8470 , n8418 );
and ( n8472 , n8382 , n8397 );
or ( n8473 , n8471 , n8472 );
and ( n8474 , n8469 , n8473 );
and ( n8475 , n8462 , n8468 );
or ( n8476 , n8474 , n8475 );
not ( n8477 , n5595 );
not ( n8478 , n545 );
not ( n8479 , n5836 );
or ( n8480 , n8478 , n8479 );
nand ( n8481 , n5837 , n4666 );
nand ( n8482 , n8480 , n8481 );
not ( n8483 , n8482 );
or ( n8484 , n8477 , n8483 );
not ( n8485 , n545 );
not ( n8486 , n8231 );
or ( n8487 , n8485 , n8486 );
nand ( n8488 , n8230 , n4666 );
nand ( n8489 , n8487 , n8488 );
nand ( n8490 , n8489 , n5339 );
nand ( n8491 , n8484 , n8490 );
xor ( n8492 , n8476 , n8491 );
not ( n8493 , n5784 );
not ( n8494 , n541 );
not ( n8495 , n7443 );
or ( n8496 , n8494 , n8495 );
nand ( n8497 , n7442 , n5734 );
nand ( n8498 , n8496 , n8497 );
not ( n8499 , n8498 );
or ( n8500 , n8493 , n8499 );
nand ( n8501 , n8463 , n5747 );
nand ( n8502 , n8500 , n8501 );
xor ( n8503 , n8191 , n8202 );
xor ( n8504 , n8503 , n8219 );
xor ( n8505 , n8502 , n8504 );
not ( n8506 , n543 );
not ( n8507 , n7081 );
or ( n8508 , n8506 , n8507 );
nand ( n8509 , n7409 , n5146 );
nand ( n8510 , n8508 , n8509 );
nand ( n8511 , n8510 , n4670 );
not ( n8512 , n543 );
not ( n8513 , n8423 );
or ( n8514 , n8512 , n8513 );
nand ( n8515 , n6012 , n5146 );
nand ( n8516 , n8514 , n8515 );
nand ( n8517 , n8516 , n4669 );
nand ( n8518 , n8511 , n8517 );
xor ( n8519 , n8505 , n8518 );
xor ( n8520 , n8492 , n8519 );
and ( n8521 , n8461 , n8520 );
and ( n8522 , n8354 , n8460 );
or ( n8523 , n8521 , n8522 );
not ( n8524 , n5741 );
not ( n8525 , n8034 );
or ( n8526 , n8524 , n8525 );
nand ( n8527 , n8498 , n5746 );
nand ( n8528 , n8526 , n8527 );
not ( n8529 , n4670 );
not ( n8530 , n8516 );
or ( n8531 , n8529 , n8530 );
nand ( n8532 , n8235 , n4669 );
nand ( n8533 , n8531 , n8532 );
xor ( n8534 , n8528 , n8533 );
xor ( n8535 , n8178 , n8188 );
xor ( n8536 , n8535 , n8222 );
xor ( n8537 , n8534 , n8536 );
not ( n8538 , n6667 );
not ( n8539 , n549 );
not ( n8540 , n4474 );
or ( n8541 , n8539 , n8540 );
not ( n8542 , n549 );
nand ( n8543 , n8542 , n7612 );
nand ( n8544 , n8541 , n8543 );
not ( n8545 , n8544 );
or ( n8546 , n8538 , n8545 );
and ( n8547 , n549 , n5731 );
not ( n8548 , n549 );
and ( n8549 , n8548 , n4651 );
or ( n8550 , n8547 , n8549 );
nand ( n8551 , n8550 , n6095 );
nand ( n8552 , n8546 , n8551 );
xor ( n8553 , n8537 , n8552 );
not ( n8554 , n552 );
not ( n8555 , n6924 );
not ( n8556 , n7781 );
or ( n8557 , n8555 , n8556 );
nand ( n8558 , n7784 , n551 );
nand ( n8559 , n8557 , n8558 );
not ( n8560 , n8559 );
or ( n8561 , n8554 , n8560 );
nand ( n8562 , n8346 , n6974 );
nand ( n8563 , n8561 , n8562 );
xor ( n8564 , n8553 , n8563 );
xor ( n8565 , n8523 , n8564 );
xor ( n8566 , n8476 , n8491 );
and ( n8567 , n8566 , n8519 );
and ( n8568 , n8476 , n8491 );
or ( n8569 , n8567 , n8568 );
not ( n8570 , n5339 );
not ( n8571 , n8482 );
or ( n8572 , n8570 , n8571 );
nand ( n8573 , n8246 , n5595 );
nand ( n8574 , n8572 , n8573 );
not ( n8575 , n7026 );
not ( n8576 , n547 );
not ( n8577 , n8576 );
not ( n8578 , n8453 );
or ( n8579 , n8577 , n8578 );
nand ( n8580 , n7714 , n547 );
nand ( n8581 , n8579 , n8580 );
not ( n8582 , n8581 );
or ( n8583 , n8575 , n8582 );
and ( n8584 , n547 , n5944 );
not ( n8585 , n547 );
and ( n8586 , n8585 , n5976 );
or ( n8587 , n8584 , n8586 );
nand ( n8588 , n8587 , n6983 );
nand ( n8589 , n8583 , n8588 );
xor ( n8590 , n8574 , n8589 );
xor ( n8591 , n8502 , n8504 );
and ( n8592 , n8591 , n8518 );
and ( n8593 , n8502 , n8504 );
or ( n8594 , n8592 , n8593 );
xor ( n8595 , n8590 , n8594 );
xor ( n8596 , n8569 , n8595 );
not ( n8597 , n6983 );
not ( n8598 , n8581 );
or ( n8599 , n8597 , n8598 );
nand ( n8600 , n8365 , n7127 );
nand ( n8601 , n8599 , n8600 );
not ( n8602 , n5329 );
not ( n8603 , n8510 );
or ( n8604 , n8602 , n8603 );
nand ( n8605 , n8372 , n4670 );
nand ( n8606 , n8604 , n8605 );
not ( n8607 , n5339 );
not ( n8608 , n8427 );
or ( n8609 , n8607 , n8608 );
nand ( n8610 , n8489 , n5595 );
nand ( n8611 , n8609 , n8610 );
xor ( n8612 , n8606 , n8611 );
xor ( n8613 , n8462 , n8468 );
xor ( n8614 , n8613 , n8473 );
and ( n8615 , n8612 , n8614 );
and ( n8616 , n8606 , n8611 );
or ( n8617 , n8615 , n8616 );
xor ( n8618 , n8601 , n8617 );
not ( n8619 , n6095 );
not ( n8620 , n8544 );
or ( n8621 , n8619 , n8620 );
nand ( n8622 , n6667 , n8446 );
nand ( n8623 , n8621 , n8622 );
and ( n8624 , n8618 , n8623 );
and ( n8625 , n8601 , n8617 );
or ( n8626 , n8624 , n8625 );
xor ( n8627 , n8596 , n8626 );
and ( n8628 , n8565 , n8627 );
and ( n8629 , n8523 , n8564 );
or ( n8630 , n8628 , n8629 );
not ( n8631 , n6095 );
not ( n8632 , n8133 );
or ( n8633 , n8631 , n8632 );
nand ( n8634 , n8550 , n6667 );
nand ( n8635 , n8633 , n8634 );
xor ( n8636 , n8225 , n8237 );
xor ( n8637 , n8636 , n8248 );
xor ( n8638 , n8635 , n8637 );
xor ( n8639 , n8574 , n8589 );
and ( n8640 , n8639 , n8594 );
and ( n8641 , n8574 , n8589 );
or ( n8642 , n8640 , n8641 );
xor ( n8643 , n8638 , n8642 );
xor ( n8644 , n8569 , n8595 );
and ( n8645 , n8644 , n8626 );
and ( n8646 , n8569 , n8595 );
or ( n8647 , n8645 , n8646 );
xor ( n8648 , n8643 , n8647 );
not ( n8649 , n552 );
not ( n8650 , n8257 );
or ( n8651 , n8649 , n8650 );
nand ( n8652 , n8559 , n6974 );
nand ( n8653 , n8651 , n8652 );
xor ( n8654 , n8023 , n8025 );
xor ( n8655 , n8654 , n8036 );
xor ( n8656 , n8528 , n8533 );
and ( n8657 , n8656 , n8536 );
and ( n8658 , n8528 , n8533 );
or ( n8659 , n8657 , n8658 );
xor ( n8660 , n8655 , n8659 );
not ( n8661 , n6983 );
not ( n8662 , n8121 );
or ( n8663 , n8661 , n8662 );
nand ( n8664 , n8587 , n7127 );
nand ( n8665 , n8663 , n8664 );
xor ( n8666 , n8660 , n8665 );
xor ( n8667 , n8653 , n8666 );
xor ( n8668 , n8537 , n8552 );
and ( n8669 , n8668 , n8563 );
and ( n8670 , n8537 , n8552 );
or ( n8671 , n8669 , n8670 );
xor ( n8672 , n8667 , n8671 );
xor ( n8673 , n8648 , n8672 );
nor ( n8674 , n8630 , n8673 );
xor ( n8675 , n8523 , n8564 );
xor ( n8676 , n8675 , n8627 );
xor ( n8677 , n8601 , n8617 );
xor ( n8678 , n8677 , n8623 );
xor ( n8679 , n8606 , n8611 );
xor ( n8680 , n8679 , n8614 );
not ( n8681 , n6974 );
not ( n8682 , n551 );
not ( n8683 , n4474 );
or ( n8684 , n8682 , n8683 );
nand ( n8685 , n7612 , n6924 );
nand ( n8686 , n8684 , n8685 );
not ( n8687 , n8686 );
or ( n8688 , n8681 , n8687 );
not ( n8689 , n8351 );
not ( n8690 , n8350 );
or ( n8691 , n8689 , n8690 );
nand ( n8692 , n8691 , n552 );
nand ( n8693 , n8688 , n8692 );
xor ( n8694 , n8680 , n8693 );
xnor ( n8695 , n8408 , n8417 );
not ( n8696 , n4669 );
not ( n8697 , n8379 );
or ( n8698 , n8696 , n8697 );
not ( n8699 , n543 );
not ( n8700 , n7860 );
or ( n8701 , n8699 , n8700 );
nand ( n8702 , n7696 , n5146 );
nand ( n8703 , n8701 , n8702 );
nand ( n8704 , n8703 , n4670 );
nand ( n8705 , n8698 , n8704 );
xor ( n8706 , n8695 , n8705 );
and ( n8707 , n8190 , n5741 );
not ( n8708 , n4669 );
not ( n8709 , n8703 );
or ( n8710 , n8708 , n8709 );
not ( n8711 , n543 );
not ( n8712 , n8196 );
or ( n8713 , n8711 , n8712 );
nand ( n8714 , n7878 , n5146 );
nand ( n8715 , n8713 , n8714 );
nand ( n8716 , n8715 , n4670 );
nand ( n8717 , n8710 , n8716 );
xor ( n8718 , n8707 , n8717 );
not ( n8719 , n4664 );
not ( n8720 , n7891 );
or ( n8721 , n8719 , n8720 );
nand ( n8722 , n8721 , n545 );
and ( n8723 , n7896 , n544 );
nor ( n8724 , n8723 , n5146 );
and ( n8725 , n8722 , n8724 );
not ( n8726 , n4669 );
not ( n8727 , n8715 );
or ( n8728 , n8726 , n8727 );
not ( n8729 , n7891 );
not ( n8730 , n7402 );
not ( n8731 , n8730 );
and ( n8732 , n8729 , n8731 );
nor ( n8733 , n7896 , n7396 );
nor ( n8734 , n8732 , n8733 );
nand ( n8735 , n8728 , n8734 );
and ( n8736 , n8725 , n8735 );
and ( n8737 , n8718 , n8736 );
and ( n8738 , n8707 , n8717 );
or ( n8739 , n8737 , n8738 );
and ( n8740 , n8706 , n8739 );
and ( n8741 , n8695 , n8705 );
or ( n8742 , n8740 , n8741 );
not ( n8743 , n6983 );
not ( n8744 , n8359 );
or ( n8745 , n8743 , n8744 );
and ( n8746 , n547 , n5726 );
not ( n8747 , n547 );
and ( n8748 , n8747 , n8230 );
or ( n8749 , n8746 , n8748 );
nand ( n8750 , n8749 , n7127 );
nand ( n8751 , n8745 , n8750 );
xor ( n8752 , n8742 , n8751 );
xor ( n8753 , n8381 , n8419 );
xor ( n8754 , n8753 , n8436 );
and ( n8755 , n8752 , n8754 );
and ( n8756 , n8742 , n8751 );
or ( n8757 , n8755 , n8756 );
and ( n8758 , n8694 , n8757 );
and ( n8759 , n8680 , n8693 );
or ( n8760 , n8758 , n8759 );
xor ( n8761 , n8678 , n8760 );
xor ( n8762 , n8354 , n8460 );
xor ( n8763 , n8762 , n8520 );
and ( n8764 , n8761 , n8763 );
and ( n8765 , n8678 , n8760 );
or ( n8766 , n8764 , n8765 );
nor ( n8767 , n8676 , n8766 );
nor ( n8768 , n8674 , n8767 );
not ( n8769 , n8768 );
xor ( n8770 , n8678 , n8760 );
xor ( n8771 , n8770 , n8763 );
not ( n8772 , n8771 );
xor ( n8773 , n8367 , n8439 );
xor ( n8774 , n8773 , n8457 );
not ( n8775 , n6095 );
not ( n8776 , n8455 );
or ( n8777 , n8775 , n8776 );
not ( n8778 , n549 );
not ( n8779 , n7088 );
or ( n8780 , n8778 , n8779 );
nand ( n8781 , n5914 , n7190 );
nand ( n8782 , n8780 , n8781 );
nand ( n8783 , n8782 , n6667 );
nand ( n8784 , n8777 , n8783 );
not ( n8785 , n5595 );
not ( n8786 , n8434 );
or ( n8787 , n8785 , n8786 );
not ( n8788 , n545 );
not ( n8789 , n7443 );
or ( n8790 , n8788 , n8789 );
nand ( n8791 , n4666 , n7444 );
nand ( n8792 , n8790 , n8791 );
nand ( n8793 , n5339 , n8792 );
nand ( n8794 , n8787 , n8793 );
not ( n8795 , n6983 );
not ( n8796 , n8749 );
or ( n8797 , n8795 , n8796 );
not ( n8798 , n6012 );
not ( n8799 , n8576 );
or ( n8800 , n8798 , n8799 );
or ( n8801 , n8576 , n6012 );
nand ( n8802 , n8800 , n8801 );
nand ( n8803 , n8802 , n7026 );
nand ( n8804 , n8797 , n8803 );
xor ( n8805 , n8794 , n8804 );
xor ( n8806 , n8695 , n8705 );
xor ( n8807 , n8806 , n8739 );
and ( n8808 , n8805 , n8807 );
and ( n8809 , n8794 , n8804 );
or ( n8810 , n8808 , n8809 );
xor ( n8811 , n8784 , n8810 );
not ( n8812 , n552 );
not ( n8813 , n8686 );
or ( n8814 , n8812 , n8813 );
not ( n8815 , n551 );
not ( n8816 , n5944 );
or ( n8817 , n8815 , n8816 );
nand ( n8818 , n5943 , n6924 );
nand ( n8819 , n8817 , n8818 );
nand ( n8820 , n8819 , n6974 );
nand ( n8821 , n8814 , n8820 );
and ( n8822 , n8811 , n8821 );
and ( n8823 , n8784 , n8810 );
or ( n8824 , n8822 , n8823 );
xor ( n8825 , n8774 , n8824 );
xor ( n8826 , n8680 , n8693 );
xor ( n8827 , n8826 , n8757 );
and ( n8828 , n8825 , n8827 );
and ( n8829 , n8774 , n8824 );
or ( n8830 , n8828 , n8829 );
not ( n8831 , n8830 );
nand ( n8832 , n8772 , n8831 );
not ( n8833 , n8832 );
xor ( n8834 , n8774 , n8824 );
xor ( n8835 , n8834 , n8827 );
not ( n8836 , n8835 );
not ( n8837 , n6095 );
not ( n8838 , n8782 );
or ( n8839 , n8837 , n8838 );
not ( n8840 , n5644 );
not ( n8841 , n549 );
or ( n8842 , n8840 , n8841 );
or ( n8843 , n7147 , n549 );
nand ( n8844 , n8842 , n8843 );
nand ( n8845 , n8844 , n6667 );
nand ( n8846 , n8839 , n8845 );
not ( n8847 , n552 );
not ( n8848 , n8819 );
or ( n8849 , n8847 , n8848 );
and ( n8850 , n7714 , n7040 );
nor ( n8851 , C0 , n8850 );
nand ( n8852 , n8849 , n8851 );
xor ( n8853 , n8846 , n8852 );
not ( n8854 , n5595 );
not ( n8855 , n8792 );
or ( n8856 , n8854 , n8855 );
not ( n8857 , n545 );
not ( n8858 , n8017 );
or ( n8859 , n8857 , n8858 );
nand ( n8860 , n8377 , n4666 );
nand ( n8861 , n8859 , n8860 );
nand ( n8862 , n8861 , n5339 );
nand ( n8863 , n8856 , n8862 );
xor ( n8864 , n8707 , n8717 );
xor ( n8865 , n8864 , n8736 );
xor ( n8866 , n8863 , n8865 );
not ( n8867 , n6983 );
not ( n8868 , n8802 );
or ( n8869 , n8867 , n8868 );
and ( n8870 , n547 , n7081 );
not ( n8871 , n547 );
and ( n8872 , n8871 , n7409 );
or ( n8873 , n8870 , n8872 );
nand ( n8874 , n8873 , n7026 );
nand ( n8875 , n8869 , n8874 );
and ( n8876 , n8866 , n8875 );
and ( n8877 , n8863 , n8865 );
or ( n8878 , n8876 , n8877 );
and ( n8879 , n8853 , n8878 );
and ( n8880 , n8846 , n8852 );
or ( n8881 , n8879 , n8880 );
xor ( n8882 , n8742 , n8751 );
xor ( n8883 , n8882 , n8754 );
xor ( n8884 , n8881 , n8883 );
xor ( n8885 , n8784 , n8810 );
xor ( n8886 , n8885 , n8821 );
and ( n8887 , n8884 , n8886 );
and ( n8888 , n8881 , n8883 );
or ( n8889 , n8887 , n8888 );
not ( n8890 , n8889 );
and ( n8891 , n8836 , n8890 );
xor ( n8892 , n8881 , n8883 );
xor ( n8893 , n8892 , n8886 );
xor ( n8894 , n8794 , n8804 );
xor ( n8895 , n8894 , n8807 );
xor ( n8896 , n8725 , n8735 );
not ( n8897 , n5594 );
not ( n8898 , n8861 );
or ( n8899 , n8897 , n8898 );
not ( n8900 , n545 );
not ( n8901 , n7860 );
or ( n8902 , n8900 , n8901 );
nand ( n8903 , n7696 , n4666 );
nand ( n8904 , n8902 , n8903 );
nand ( n8905 , n8904 , n5339 );
nand ( n8906 , n8899 , n8905 );
xor ( n8907 , n8896 , n8906 );
not ( n8908 , n6983 );
not ( n8909 , n8873 );
or ( n8910 , n8908 , n8909 );
not ( n8911 , n547 );
not ( n8912 , n7443 );
or ( n8913 , n8911 , n8912 );
not ( n8914 , n547 );
nand ( n8915 , n8914 , n7442 );
nand ( n8916 , n8913 , n8915 );
nand ( n8917 , n8916 , n7127 );
nand ( n8918 , n8910 , n8917 );
and ( n8919 , n8907 , n8918 );
and ( n8920 , n8896 , n8906 );
or ( n8921 , n8919 , n8920 );
not ( n8922 , n6095 );
not ( n8923 , n8844 );
or ( n8924 , n8922 , n8923 );
and ( n8925 , n549 , n8230 );
not ( n8926 , n549 );
and ( n8927 , n8926 , n5726 );
nor ( n8928 , n8925 , n8927 );
nand ( n8929 , n8928 , n6667 );
nand ( n8930 , n8924 , n8929 );
xor ( n8931 , n8921 , n8930 );
nand ( n8932 , n8453 , n7494 );
nand ( n8933 , n7714 , n7491 );
and ( n8934 , n6924 , n7088 );
not ( n8935 , n6924 );
and ( n8936 , n8935 , n5914 );
nor ( n8937 , n8934 , n8936 );
nand ( n8938 , n8937 , n6974 );
nand ( n8939 , n8932 , n8933 , n8938 );
and ( n8940 , n8931 , n8939 );
and ( n8941 , n8921 , n8930 );
or ( n8942 , n8940 , n8941 );
xor ( n8943 , n8895 , n8942 );
xor ( n8944 , n8846 , n8852 );
xor ( n8945 , n8944 , n8878 );
and ( n8946 , n8943 , n8945 );
and ( n8947 , n8895 , n8942 );
or ( n8948 , n8946 , n8947 );
nor ( n8949 , n8893 , n8948 );
nor ( n8950 , n8891 , n8949 );
not ( n8951 , n8950 );
xor ( n8952 , n8895 , n8942 );
xor ( n8953 , n8952 , n8945 );
not ( n8954 , n8953 );
xor ( n8955 , n8863 , n8865 );
xor ( n8956 , n8955 , n8875 );
and ( n8957 , n8190 , n4669 );
not ( n8958 , n5594 );
not ( n8959 , n8904 );
or ( n8960 , n8958 , n8959 );
not ( n8961 , n545 );
not ( n8962 , n8196 );
or ( n8963 , n8961 , n8962 );
nand ( n8964 , n7878 , n4666 );
nand ( n8965 , n8963 , n8964 );
nand ( n8966 , n5339 , n8965 );
nand ( n8967 , n8960 , n8966 );
xor ( n8968 , n8957 , n8967 );
and ( n8969 , n7896 , n546 );
nor ( n8970 , n8969 , n4666 );
not ( n8971 , n546 );
not ( n8972 , n8971 );
not ( n8973 , n7891 );
or ( n8974 , n8972 , n8973 );
nand ( n8975 , n8974 , n547 );
and ( n8976 , n8970 , n8975 );
not ( n8977 , n5594 );
not ( n8978 , n8965 );
or ( n8979 , n8977 , n8978 );
and ( n8980 , n545 , n7856 );
not ( n8981 , n545 );
and ( n8982 , n8981 , n7891 );
nor ( n8983 , n8980 , n8982 );
nand ( n8984 , n8983 , n5339 );
nand ( n8985 , n8979 , n8984 );
and ( n8986 , n8976 , n8985 );
and ( n8987 , n8968 , n8986 );
and ( n8988 , n8957 , n8967 );
or ( n8989 , n8987 , n8988 );
not ( n8990 , n6012 );
and ( n8991 , n549 , n8990 );
not ( n8992 , n549 );
and ( n8993 , n8992 , n6012 );
or ( n8994 , n8991 , n8993 );
not ( n8995 , n8994 );
not ( n8996 , n6667 );
or ( n8997 , n8995 , n8996 );
nand ( n8998 , n8928 , n6095 );
nand ( n8999 , n8997 , n8998 );
xor ( n9000 , n8989 , n8999 );
xor ( n9001 , n8896 , n8906 );
xor ( n9002 , n9001 , n8918 );
and ( n9003 , n9000 , n9002 );
and ( n9004 , n8989 , n8999 );
or ( n9005 , n9003 , n9004 );
xor ( n9006 , n8956 , n9005 );
xor ( n9007 , n8921 , n8930 );
xor ( n9008 , n9007 , n8939 );
and ( n9009 , n9006 , n9008 );
and ( n9010 , n8956 , n9005 );
or ( n9011 , n9009 , n9010 );
not ( n9012 , n9011 );
nand ( n9013 , n8954 , n9012 );
not ( n9014 , n9013 );
xor ( n9015 , n8956 , n9005 );
xor ( n9016 , n9015 , n9008 );
not ( n9017 , n8937 );
not ( n9018 , n552 );
or ( n9019 , n9017 , n9018 );
not ( n9020 , n7040 );
or ( n9021 , n5837 , n9020 );
nand ( n9022 , n9019 , n9021 );
not ( n9023 , n6983 );
not ( n9024 , n8916 );
or ( n9025 , n9023 , n9024 );
and ( n9026 , n547 , n8017 );
not ( n9027 , n547 );
and ( n9028 , n9027 , n7580 );
or ( n9029 , n9026 , n9028 );
nand ( n9030 , n9029 , n7127 );
nand ( n9031 , n9025 , n9030 );
xor ( n9032 , n8957 , n8967 );
xor ( n9033 , n9032 , n8986 );
xor ( n9034 , n9031 , n9033 );
not ( n9035 , n6095 );
not ( n9036 , n8994 );
or ( n9037 , n9035 , n9036 );
and ( n9038 , n549 , n7081 );
not ( n9039 , n549 );
and ( n9040 , n9039 , n7082 );
or ( n9041 , n9038 , n9040 );
nand ( n9042 , n9041 , n6667 );
nand ( n9043 , n9037 , n9042 );
and ( n9044 , n9034 , n9043 );
and ( n9045 , n9031 , n9033 );
or ( n9046 , n9044 , n9045 );
xor ( n9047 , n9022 , n9046 );
xor ( n9048 , n8989 , n8999 );
xor ( n9049 , n9048 , n9002 );
and ( n9050 , n9047 , n9049 );
and ( n9051 , n9022 , n9046 );
or ( n9052 , n9050 , n9051 );
nor ( n9053 , n9016 , n9052 );
xor ( n9054 , n9022 , n9046 );
xor ( n9055 , n9054 , n9049 );
not ( n9056 , n9055 );
xor ( n9057 , n8976 , n8985 );
not ( n9058 , n6983 );
not ( n9059 , n9029 );
or ( n9060 , n9058 , n9059 );
xor ( n9061 , n547 , n7696 );
nand ( n9062 , n9061 , n7026 );
nand ( n9063 , n9060 , n9062 );
xor ( n9064 , n9057 , n9063 );
and ( n9065 , n8190 , n5594 );
not ( n9066 , n6983 );
not ( n9067 , n9061 );
or ( n9068 , n9066 , n9067 );
xor ( n9069 , n7878 , n547 );
nand ( n9070 , n9069 , n7026 );
nand ( n9071 , n9068 , n9070 );
xor ( n9072 , n9065 , n9071 );
and ( n9073 , n9069 , n6983 );
not ( n9074 , n7786 );
not ( n9075 , n7891 );
or ( n9076 , n9074 , n9075 );
nand ( n9077 , n7856 , n7782 );
nand ( n9078 , n9076 , n9077 );
nor ( n9079 , n9073 , n9078 );
and ( n9080 , n7856 , n548 );
nor ( n9081 , n9080 , n8576 );
not ( n9082 , n548 );
not ( n9083 , n9082 );
not ( n9084 , n7891 );
or ( n9085 , n9083 , n9084 );
nand ( n9086 , n9085 , n549 );
nand ( n9087 , n9081 , n9086 );
nor ( n9088 , n9079 , n9087 );
and ( n9089 , n9072 , n9088 );
and ( n9090 , n9065 , n9071 );
or ( n9091 , n9089 , n9090 );
and ( n9092 , n9064 , n9091 );
and ( n9093 , n9057 , n9063 );
or ( n9094 , n9092 , n9093 );
not ( n9095 , n552 );
and ( n9096 , n551 , n5837 );
not ( n9097 , n551 );
and ( n9098 , n9097 , n5836 );
nor ( n9099 , n9096 , n9098 );
not ( n9100 , n9099 );
or ( n9101 , n9095 , n9100 );
not ( n9102 , n551 );
not ( n9103 , n5726 );
or ( n9104 , n9102 , n9103 );
nand ( n9105 , n8230 , n6924 );
nand ( n9106 , n9104 , n9105 );
nand ( n9107 , n9106 , n6974 );
nand ( n9108 , n9101 , n9107 );
xor ( n9109 , n9094 , n9108 );
xor ( n9110 , n9031 , n9033 );
xor ( n9111 , n9110 , n9043 );
and ( n9112 , n9109 , n9111 );
and ( n9113 , n9094 , n9108 );
or ( n9114 , n9112 , n9113 );
not ( n9115 , n9114 );
nand ( n9116 , n9056 , n9115 );
xor ( n9117 , n9094 , n9108 );
xor ( n9118 , n9117 , n9111 );
not ( n9119 , n6095 );
not ( n9120 , n9041 );
or ( n9121 , n9119 , n9120 );
and ( n9122 , n549 , n7443 );
not ( n9123 , n549 );
and ( n9124 , n9123 , n7442 );
or ( n9125 , n9122 , n9124 );
nand ( n9126 , n9125 , n6667 );
nand ( n9127 , n9121 , n9126 );
not ( n9128 , n6974 );
not ( n9129 , n6013 );
or ( n9130 , n9128 , n9129 );
nand ( n9131 , n9106 , n552 );
nand ( n9132 , n9130 , n9131 );
xor ( n9133 , n9127 , n9132 );
xor ( n9134 , n9057 , n9063 );
xor ( n9135 , n9134 , n9091 );
and ( n9136 , n9133 , n9135 );
and ( n9137 , n9127 , n9132 );
or ( n9138 , n9136 , n9137 );
nor ( n9139 , n9118 , n9138 );
not ( n9140 , n6095 );
not ( n9141 , n9125 );
or ( n9142 , n9140 , n9141 );
and ( n9143 , n549 , n8017 );
not ( n9144 , n549 );
and ( n9145 , n9144 , n7580 );
or ( n9146 , n9143 , n9145 );
nand ( n9147 , n9146 , n6667 );
nand ( n9148 , n9142 , n9147 );
xor ( n9149 , n9065 , n9071 );
xor ( n9150 , n9149 , n9088 );
xor ( n9151 , n9148 , n9150 );
not ( n9152 , n7494 );
not ( n9153 , n9152 );
nand ( n9154 , n9153 , n6012 );
nand ( n9155 , n7081 , n6974 );
nand ( n9156 , n8990 , n7491 );
nand ( n9157 , n9154 , n9155 , n9156 );
and ( n9158 , n9151 , n9157 );
and ( n9159 , n9148 , n9150 );
or ( n9160 , n9158 , n9159 );
not ( n9161 , n9160 );
xor ( n9162 , n9127 , n9132 );
xor ( n9163 , n9162 , n9135 );
not ( n9164 , n9163 );
nand ( n9165 , n9161 , n9164 );
nor ( n9166 , n7895 , n6982 );
not ( n9167 , n6095 );
and ( n9168 , n549 , n7860 );
not ( n9169 , n549 );
and ( n9170 , n9169 , n7696 );
or ( n9171 , n9168 , n9170 );
not ( n9172 , n9171 );
or ( n9173 , n9167 , n9172 );
not ( n9174 , n549 );
not ( n9175 , n8196 );
or ( n9176 , n9174 , n9175 );
not ( n9177 , n549 );
nand ( n9178 , n9177 , n7878 );
nand ( n9179 , n9176 , n9178 );
nand ( n9180 , n9179 , n6667 );
nand ( n9181 , n9173 , n9180 );
xor ( n9182 , n9166 , n9181 );
and ( n9183 , n7896 , n550 );
nor ( n9184 , n9183 , n7190 );
not ( n9185 , n550 );
not ( n9186 , n9185 );
not ( n9187 , n7891 );
or ( n9188 , n9186 , n9187 );
nand ( n9189 , n9188 , n551 );
and ( n9190 , n9184 , n9189 );
not ( n9191 , n6095 );
not ( n9192 , n9179 );
or ( n9193 , n9191 , n9192 );
and ( n9194 , n7896 , n7471 );
and ( n9195 , n7891 , n7473 );
nor ( n9196 , n9194 , n9195 );
nand ( n9197 , n9193 , n9196 );
and ( n9198 , n9190 , n9197 );
xor ( n9199 , n9182 , n9198 );
not ( n9200 , n552 );
and ( n9201 , n7441 , n551 );
not ( n9202 , n7441 );
and ( n9203 , n9202 , n6924 );
or ( n9204 , n9201 , n9203 );
not ( n9205 , n9204 );
or ( n9206 , n9200 , n9205 );
and ( n9207 , n7580 , n6924 );
not ( n9208 , n7580 );
and ( n9209 , n9208 , n551 );
or ( n9210 , n9207 , n9209 );
nand ( n9211 , n9210 , n6974 );
nand ( n9212 , n9206 , n9211 );
or ( n9213 , n9199 , n9212 );
xor ( n9214 , n9190 , n9197 );
not ( n9215 , n9214 );
not ( n9216 , n7697 );
not ( n9217 , n6974 );
not ( n9218 , n9217 );
and ( n9219 , n9216 , n9218 );
and ( n9220 , n9210 , n552 );
nor ( n9221 , n9219 , n9220 );
nand ( n9222 , n9215 , n9221 );
not ( n9223 , n9222 );
and ( n9224 , n8190 , n6095 );
not ( n9225 , n551 );
not ( n9226 , n8196 );
or ( n9227 , n9225 , n9226 );
nand ( n9228 , n7878 , n6924 );
nand ( n9229 , n9227 , n9228 );
and ( n9230 , n552 , n9229 );
and ( n9231 , n7891 , n7040 );
nor ( n9232 , n9230 , n9231 );
nand ( n9233 , n7855 , n552 );
nand ( n9234 , n551 , n9233 );
nor ( n9235 , n9232 , n9234 );
xor ( n9236 , n9224 , n9235 );
not ( n9237 , n7697 );
nand ( n9238 , n9237 , n7491 );
nand ( n9239 , n9229 , n6974 );
nand ( n9240 , n7697 , n7494 );
nand ( n9241 , n9238 , n9239 , n9240 );
and ( n9242 , n9236 , n9241 );
or ( n9243 , n9242 , C0 );
not ( n9244 , n9243 );
or ( n9245 , n9223 , n9244 );
not ( n9246 , n9221 );
nand ( n9247 , n9246 , n9214 );
nand ( n9248 , n9245 , n9247 );
and ( n9249 , n9213 , n9248 );
and ( n9250 , n9199 , n9212 );
nor ( n9251 , n9249 , n9250 );
xor ( n9252 , n9079 , n9087 );
not ( n9253 , n6095 );
not ( n9254 , n9146 );
or ( n9255 , n9253 , n9254 );
nand ( n9256 , n9171 , n6667 );
nand ( n9257 , n9255 , n9256 );
xor ( n9258 , n9252 , n9257 );
nand ( n9259 , n7494 , n7409 );
nand ( n9260 , n7081 , n7491 );
nand ( n9261 , n9204 , n6974 );
nand ( n9262 , n9259 , n9260 , n9261 );
xor ( n9263 , n9258 , n9262 );
xor ( n9264 , n9166 , n9181 );
and ( n9265 , n9264 , n9198 );
and ( n9266 , n9166 , n9181 );
or ( n9267 , n9265 , n9266 );
nor ( n9268 , n9263 , n9267 );
or ( n9269 , n9251 , n9268 );
nand ( n9270 , n9263 , n9267 );
nand ( n9271 , n9269 , n9270 );
not ( n9272 , n9271 );
xor ( n9273 , n9148 , n9150 );
xor ( n9274 , n9273 , n9157 );
not ( n9275 , n9274 );
xor ( n9276 , n9252 , n9257 );
and ( n9277 , n9276 , n9262 );
and ( n9278 , n9252 , n9257 );
or ( n9279 , n9277 , n9278 );
not ( n9280 , n9279 );
nand ( n9281 , n9275 , n9280 );
not ( n9282 , n9281 );
or ( n9283 , n9272 , n9282 );
nand ( n9284 , n9274 , n9279 );
nand ( n9285 , n9283 , n9284 );
and ( n9286 , n9165 , n9285 );
nand ( n9287 , n9163 , n9160 );
not ( n9288 , n9287 );
nor ( n9289 , n9286 , n9288 );
or ( n9290 , n9139 , n9289 );
nand ( n9291 , n9118 , n9138 );
nand ( n9292 , n9290 , n9291 );
and ( n9293 , n9116 , n9292 );
nand ( n9294 , n9055 , n9114 );
not ( n9295 , n9294 );
nor ( n9296 , n9293 , n9295 );
or ( n9297 , n9053 , n9296 );
nand ( n9298 , n9016 , n9052 );
nand ( n9299 , n9297 , n9298 );
not ( n9300 , n9299 );
or ( n9301 , n9014 , n9300 );
nand ( n9302 , n8953 , n9011 );
nand ( n9303 , n9301 , n9302 );
not ( n9304 , n9303 );
or ( n9305 , n8951 , n9304 );
not ( n9306 , n8835 );
not ( n9307 , n8889 );
nand ( n9308 , n9306 , n9307 );
and ( n9309 , n8893 , n8948 );
and ( n9310 , n9308 , n9309 );
not ( n9311 , n8835 );
nor ( n9312 , n9311 , n9307 );
nor ( n9313 , n9310 , n9312 );
nand ( n9314 , n9305 , n9313 );
not ( n9315 , n9314 );
or ( n9316 , n8833 , n9315 );
buf ( n9317 , n8771 );
nand ( n9318 , n9317 , n8830 );
nand ( n9319 , n9316 , n9318 );
not ( n9320 , n9319 );
or ( n9321 , n8769 , n9320 );
nand ( n9322 , n8676 , n8766 );
not ( n9323 , n9322 );
nor ( n9324 , n8673 , n8630 );
not ( n9325 , n9324 );
and ( n9326 , n9323 , n9325 );
nand ( n9327 , n8673 , n8630 );
not ( n9328 , n9327 );
nor ( n9329 , n9326 , n9328 );
nand ( n9330 , n9321 , n9329 );
not ( n9331 , n9330 );
xor ( n9332 , n8653 , n8666 );
and ( n9333 , n9332 , n8671 );
and ( n9334 , n8653 , n8666 );
or ( n9335 , n9333 , n9334 );
xor ( n9336 , n8251 , n8261 );
xor ( n9337 , n9336 , n8264 );
xor ( n9338 , n9335 , n9337 );
xor ( n9339 , n8655 , n8659 );
and ( n9340 , n9339 , n8665 );
and ( n9341 , n8655 , n8659 );
or ( n9342 , n9340 , n9341 );
xor ( n9343 , n8119 , n8125 );
xor ( n9344 , n9343 , n8137 );
xor ( n9345 , n9342 , n9344 );
xor ( n9346 , n8635 , n8637 );
and ( n9347 , n9346 , n8642 );
and ( n9348 , n8635 , n8637 );
or ( n9349 , n9347 , n9348 );
xor ( n9350 , n9345 , n9349 );
and ( n9351 , n9338 , n9350 );
and ( n9352 , n9335 , n9337 );
or ( n9353 , n9351 , n9352 );
not ( n9354 , n9353 );
not ( n9355 , n9354 );
xor ( n9356 , n9342 , n9344 );
and ( n9357 , n9356 , n9349 );
and ( n9358 , n9342 , n9344 );
or ( n9359 , n9357 , n9358 );
xor ( n9360 , n8117 , n8140 );
xor ( n9361 , n9360 , n8152 );
xor ( n9362 , n9359 , n9361 );
xor ( n9363 , n8174 , n8176 );
xor ( n9364 , n9363 , n8267 );
xor ( n9365 , n9362 , n9364 );
not ( n9366 , n9365 );
not ( n9367 , n9366 );
or ( n9368 , n9355 , n9367 );
xor ( n9369 , n9335 , n9337 );
xor ( n9370 , n9369 , n9350 );
xor ( n9371 , n8643 , n8647 );
and ( n9372 , n9371 , n8672 );
and ( n9373 , n8643 , n8647 );
or ( n9374 , n9372 , n9373 );
or ( n9375 , n9370 , n9374 );
nand ( n9376 , n9368 , n9375 );
xor ( n9377 , n8172 , n8270 );
xor ( n9378 , n9377 , n8273 );
xor ( n9379 , n9359 , n9361 );
and ( n9380 , n9379 , n9364 );
and ( n9381 , n9359 , n9361 );
or ( n9382 , n9380 , n9381 );
nor ( n9383 , n9378 , n9382 );
nor ( n9384 , n9376 , n9383 );
not ( n9385 , n9384 );
or ( n9386 , n9331 , n9385 );
not ( n9387 , n9378 );
not ( n9388 , n9382 );
nand ( n9389 , n9387 , n9388 );
nor ( n9390 , n9353 , n9365 );
nand ( n9391 , n9370 , n9374 );
or ( n9392 , n9390 , n9391 );
nand ( n9393 , n9365 , n9353 );
nand ( n9394 , n9392 , n9393 );
and ( n9395 , n9389 , n9394 );
nand ( n9396 , n9378 , n9382 );
not ( n9397 , n9396 );
nor ( n9398 , n9395 , n9397 );
nand ( n9399 , n9386 , n9398 );
and ( n9400 , n7763 , n8332 , n8340 , n9399 );
nor ( n9401 , n8325 , n9400 );
not ( n9402 , n545 );
not ( n9403 , n6998 );
nand ( n9404 , n9403 , n7008 , n7010 , n7013 );
not ( n9405 , n9404 );
or ( n9406 , n9402 , n9405 );
nand ( n9407 , n7015 , n4666 );
nand ( n9408 , n9406 , n9407 );
nand ( n9409 , n9408 , n5595 );
nand ( n9410 , n5593 , n5341 );
nand ( n9411 , n9409 , n9410 );
not ( n9412 , n552 );
and ( n9413 , n7260 , n7311 );
not ( n9414 , n9413 );
not ( n9415 , n6943 );
or ( n9416 , n9414 , n9415 );
not ( n9417 , n7311 );
not ( n9418 , n7265 );
or ( n9419 , n9417 , n9418 );
nand ( n9420 , n9419 , n7314 );
not ( n9421 , n9420 );
nand ( n9422 , n9416 , n9421 );
not ( n9423 , n9422 );
xor ( n9424 , n7276 , n7283 );
and ( n9425 , n9424 , n7289 );
and ( n9426 , n7276 , n7283 );
or ( n9427 , n9425 , n9426 );
and ( n9428 , n507 , n489 );
not ( n9429 , n7277 );
not ( n9430 , n6562 );
or ( n9431 , n9429 , n9430 );
xnor ( n9432 , n489 , n505 );
not ( n9433 , n9432 );
nand ( n9434 , n9433 , n1859 );
nand ( n9435 , n9431 , n9434 );
xor ( n9436 , n9428 , n9435 );
not ( n9437 , n6760 );
not ( n9438 , n6758 );
or ( n9439 , n9437 , n9438 );
nand ( n9440 , n9439 , n491 );
xor ( n9441 , n9436 , n9440 );
xor ( n9442 , n9427 , n9441 );
not ( n9443 , n7289 );
xor ( n9444 , n9442 , n9443 );
not ( n9445 , n9444 );
not ( n9446 , n7290 );
nand ( n9447 , n9446 , n7297 );
and ( n9448 , n7275 , n9447 );
and ( n9449 , n7294 , n7290 );
nor ( n9450 , n9448 , n9449 );
nand ( n9451 , n9445 , n9450 );
or ( n9452 , n9445 , n9450 );
nand ( n9453 , n9451 , n9452 );
nor ( n9454 , n9453 , n455 );
nand ( n9455 , n9423 , n9454 );
nand ( n9456 , n7209 , n7255 );
nor ( n9457 , n6812 , n9456 );
not ( n9458 , n9457 );
not ( n9459 , n6627 );
or ( n9460 , n9458 , n9459 );
not ( n9461 , n6173 );
not ( n9462 , n4413 );
or ( n9463 , n9461 , n9462 );
nor ( n9464 , n6260 , n6866 );
nand ( n9465 , n9463 , n9464 );
nand ( n9466 , n6264 , n6326 );
and ( n9467 , n6867 , n9466 );
nor ( n9468 , n9467 , n9456 );
and ( n9469 , n9465 , n9468 );
not ( n9470 , n7255 );
not ( n9471 , n7218 );
or ( n9472 , n9470 , n9471 );
nand ( n9473 , n9472 , n7256 );
nor ( n9474 , n9469 , n9473 );
nand ( n9475 , n9460 , n9474 );
not ( n9476 , n9475 );
xor ( n9477 , n7229 , n7248 );
and ( n9478 , n9477 , n7253 );
and ( n9479 , n7229 , n7248 );
or ( n9480 , n9478 , n9479 );
not ( n9481 , n9480 );
not ( n9482 , n7247 );
not ( n9483 , n2035 );
not ( n9484 , n1999 );
or ( n9485 , n9483 , n9484 );
nand ( n9486 , n9485 , n491 );
not ( n9487 , n2122 );
not ( n9488 , n7237 );
or ( n9489 , n9487 , n9488 );
xor ( n9490 , n489 , n2152 );
nand ( n9491 , n9490 , n2084 );
nand ( n9492 , n9489 , n9491 );
xor ( n9493 , n9486 , n9492 );
and ( n9494 , n489 , n6304 );
xor ( n9495 , n9493 , n9494 );
xor ( n9496 , n9482 , n9495 );
xor ( n9497 , n7239 , n7240 );
and ( n9498 , n9497 , n7247 );
and ( n9499 , n7239 , n7240 );
or ( n9500 , n9498 , n9499 );
xor ( n9501 , n9496 , n9500 );
not ( n9502 , n9501 );
xnor ( n9503 , n9481 , n9502 );
nor ( n9504 , n9503 , n5791 );
nand ( n9505 , n9476 , n9504 );
not ( n9506 , n9453 );
nor ( n9507 , n9506 , n455 );
nand ( n9508 , n9507 , n9422 );
nand ( n9509 , n9475 , n9503 , n455 );
nand ( n9510 , n9455 , n9505 , n9508 , n9509 );
and ( n9511 , n9510 , n6924 );
not ( n9512 , n9510 );
and ( n9513 , n9512 , n551 );
or ( n9514 , n9511 , n9513 );
not ( n9515 , n9514 );
or ( n9516 , n9412 , n9515 );
nand ( n9517 , n7259 , n7318 , n7321 , n7324 );
nand ( n9518 , n9517 , n7040 );
nand ( n9519 , n9516 , n9518 );
xor ( n9520 , n9411 , n9519 );
and ( n9521 , n6967 , n7471 );
not ( n9522 , n6967 );
and ( n9523 , n9522 , n7473 );
nor ( n9524 , n9521 , n9523 );
xor ( n9525 , n549 , n6923 );
nand ( n9526 , n9525 , n6095 );
nand ( n9527 , n9524 , n9526 );
and ( n9528 , n9520 , n9527 );
and ( n9529 , n9411 , n9519 );
or ( n9530 , n9528 , n9529 );
not ( n9531 , n541 );
not ( n9532 , n5322 );
or ( n9533 , n9531 , n9532 );
nand ( n9534 , n7109 , n5734 );
nand ( n9535 , n9533 , n9534 );
not ( n9536 , n9535 );
not ( n9537 , n5786 );
or ( n9538 , n9536 , n9537 );
not ( n9539 , n5145 );
not ( n9540 , n5734 );
or ( n9541 , n9539 , n9540 );
nand ( n9542 , n541 , n5141 );
nand ( n9543 , n9541 , n9542 );
nand ( n9544 , n9543 , n5747 );
nand ( n9545 , n9538 , n9544 );
not ( n9546 , n4671 );
not ( n9547 , n543 );
not ( n9548 , n7544 );
or ( n9549 , n9547 , n9548 );
nand ( n9550 , n5146 , n5466 );
nand ( n9551 , n9549 , n9550 );
not ( n9552 , n9551 );
or ( n9553 , n9546 , n9552 );
not ( n9554 , n543 );
not ( n9555 , n5589 );
or ( n9556 , n9554 , n9555 );
nand ( n9557 , n5588 , n5146 );
nand ( n9558 , n9556 , n9557 );
nand ( n9559 , n9558 , n5330 );
nand ( n9560 , n9553 , n9559 );
xor ( n9561 , n9545 , n9560 );
not ( n9562 , n545 );
not ( n9563 , n6657 );
or ( n9564 , n9562 , n9563 );
nand ( n9565 , n6656 , n4666 );
nand ( n9566 , n9564 , n9565 );
nand ( n9567 , n9566 , n5595 );
nand ( n9568 , n9408 , n5341 );
nand ( n9569 , n9567 , n9568 );
xor ( n9570 , n9561 , n9569 );
xor ( n9571 , n9530 , n9570 );
not ( n9572 , n6983 );
and ( n9573 , n547 , n7039 );
not ( n9574 , n547 );
and ( n9575 , n9574 , n7493 );
or ( n9576 , n9573 , n9575 );
not ( n9577 , n9576 );
or ( n9578 , n9572 , n9577 );
nand ( n9579 , n7345 , n7127 );
nand ( n9580 , n9578 , n9579 );
not ( n9581 , n5697 );
not ( n9582 , n537 );
not ( n9583 , n4474 );
or ( n9584 , n9582 , n9583 );
nand ( n9585 , n4473 , n5605 );
nand ( n9586 , n9584 , n9585 );
not ( n9587 , n9586 );
or ( n9588 , n9581 , n9587 );
nand ( n9589 , n5609 , n5948 );
nand ( n9590 , n9588 , n9589 );
and ( n9591 , n5915 , n5952 );
xor ( n9592 , n9590 , n9591 );
not ( n9593 , n539 );
not ( n9594 , n6056 );
or ( n9595 , n9593 , n9594 );
nand ( n9596 , n5777 , n4477 );
nand ( n9597 , n9595 , n9596 );
and ( n9598 , n9597 , n4659 );
not ( n9599 , n4450 );
nor ( n9600 , n9599 , n4657 );
nor ( n9601 , n9598 , n9600 );
nand ( n9602 , n8453 , n537 );
and ( n9603 , n9601 , n9602 );
not ( n9604 , n9601 );
not ( n9605 , n9602 );
and ( n9606 , n9604 , n9605 );
nor ( n9607 , n9603 , n9606 );
xor ( n9608 , n9592 , n9607 );
xor ( n9609 , n9580 , n9608 );
xor ( n9610 , n4662 , n5332 );
and ( n9611 , n9610 , n5597 );
and ( n9612 , n4662 , n5332 );
or ( n9613 , n9611 , n9612 );
and ( n9614 , n9609 , n9613 );
and ( n9615 , n9580 , n9608 );
or ( n9616 , n9614 , n9615 );
xor ( n9617 , n9571 , n9616 );
and ( n9618 , n7311 , n9451 );
and ( n9619 , n7260 , n9618 );
not ( n9620 , n9619 );
not ( n9621 , n6943 );
or ( n9622 , n9620 , n9621 );
and ( n9623 , n9420 , n9451 );
not ( n9624 , n9452 );
nor ( n9625 , n9623 , n9624 );
nand ( n9626 , n9622 , n9625 );
xor ( n9627 , n9427 , n9441 );
not ( n9628 , n7289 );
and ( n9629 , n9627 , n9628 );
and ( n9630 , n9427 , n9441 );
or ( n9631 , n9629 , n9630 );
or ( n9632 , n6773 , n9432 );
or ( n9633 , n6775 , n2118 );
nand ( n9634 , n9632 , n9633 );
nand ( n9635 , n506 , n489 );
xor ( n9636 , n9634 , n9635 );
xor ( n9637 , n9428 , n9435 );
and ( n9638 , n9637 , n9440 );
and ( n9639 , n9428 , n9435 );
or ( n9640 , n9638 , n9639 );
xor ( n9641 , n9636 , n9640 );
or ( n9642 , n9631 , n9641 );
nand ( n9643 , n9631 , n9641 );
nand ( n9644 , n9642 , n9643 );
and ( n9645 , n9626 , n9644 );
nor ( n9646 , n9645 , n455 );
not ( n9647 , n9646 );
not ( n9648 , n9626 );
not ( n9649 , n9644 );
nand ( n9650 , n9648 , n9649 );
not ( n9651 , n9650 );
or ( n9652 , n9647 , n9651 );
nor ( n9653 , n9502 , n9481 );
nor ( n9654 , n9475 , n9653 );
xor ( n9655 , n9482 , n9495 );
and ( n9656 , n9655 , n9500 );
and ( n9657 , n9482 , n9495 );
or ( n9658 , n9656 , n9657 );
not ( n9659 , n9658 );
not ( n9660 , n2122 );
not ( n9661 , n9490 );
or ( n9662 , n9660 , n9661 );
or ( n9663 , n2083 , n1949 );
nand ( n9664 , n9662 , n9663 );
nand ( n9665 , n2283 , n489 );
xor ( n9666 , n9664 , n9665 );
xor ( n9667 , n9486 , n9492 );
and ( n9668 , n9667 , n9494 );
and ( n9669 , n9486 , n9492 );
or ( n9670 , n9668 , n9669 );
xor ( n9671 , n9666 , n9670 );
not ( n9672 , n9671 );
or ( n9673 , n9659 , n9672 );
not ( n9674 , n9673 );
nand ( n9675 , n9659 , n9672 );
not ( n9676 , n9675 );
or ( n9677 , n9674 , n9676 );
nand ( n9678 , n9677 , n455 );
nand ( n9679 , n9654 , n9678 );
nand ( n9680 , n9675 , n9673 , n455 );
nand ( n9681 , n9481 , n9502 );
nand ( n9682 , n9475 , n9680 , n9681 );
nor ( n9683 , n9653 , n9681 );
nand ( n9684 , n9678 , n9683 );
nand ( n9685 , n9680 , n9653 );
nand ( n9686 , n9679 , n9682 , n9684 , n9685 );
nand ( n9687 , n9652 , n9686 );
not ( n9688 , n9687 );
not ( n9689 , n9688 );
nand ( n9690 , n9689 , n7491 );
nand ( n9691 , n9688 , n7494 );
not ( n9692 , n9510 );
nand ( n9693 , n9692 , n7040 );
nand ( n9694 , n9690 , n9691 , n9693 );
not ( n9695 , n6095 );
not ( n9696 , n549 );
not ( n9697 , n9696 );
not ( n9698 , n7326 );
or ( n9699 , n9697 , n9698 );
not ( n9700 , n7325 );
or ( n9701 , n9696 , n9700 );
nand ( n9702 , n9699 , n9701 );
not ( n9703 , n9702 );
or ( n9704 , n9695 , n9703 );
nand ( n9705 , n9525 , n6667 );
nand ( n9706 , n9704 , n9705 );
xor ( n9707 , n9694 , n9706 );
xor ( n9708 , n9590 , n9591 );
and ( n9709 , n9708 , n9607 );
and ( n9710 , n9590 , n9591 );
or ( n9711 , n9709 , n9710 );
xor ( n9712 , n9707 , n9711 );
not ( n9713 , n7127 );
not ( n9714 , n9576 );
or ( n9715 , n9713 , n9714 );
xor ( n9716 , n547 , n6967 );
nand ( n9717 , n9716 , n6983 );
nand ( n9718 , n9715 , n9717 );
not ( n9719 , n5786 );
not ( n9720 , n9543 );
or ( n9721 , n9719 , n9720 );
buf ( n9722 , n5893 );
nand ( n9723 , n5747 , n9722 );
nand ( n9724 , n9721 , n9723 );
xor ( n9725 , n5900 , n5908 );
and ( n9726 , n9725 , n5953 );
and ( n9727 , n5900 , n5908 );
or ( n9728 , n9726 , n9727 );
xor ( n9729 , n9724 , n9728 );
buf ( n9730 , n5330 );
not ( n9731 , n9730 );
not ( n9732 , n9551 );
or ( n9733 , n9731 , n9732 );
nand ( n9734 , n5328 , n4671 );
nand ( n9735 , n9733 , n9734 );
and ( n9736 , n9729 , n9735 );
and ( n9737 , n9724 , n9728 );
or ( n9738 , n9736 , n9737 );
xor ( n9739 , n9718 , n9738 );
not ( n9740 , n5609 );
not ( n9741 , n9586 );
or ( n9742 , n9740 , n9741 );
not ( n9743 , n4651 );
not ( n9744 , n5605 );
and ( n9745 , n9743 , n9744 );
and ( n9746 , n7958 , n5605 );
nor ( n9747 , n9745 , n9746 );
not ( n9748 , n9747 );
nand ( n9749 , n9748 , n5697 );
nand ( n9750 , n9742 , n9749 );
nor ( n9751 , n9601 , n9602 );
xor ( n9752 , n9750 , n9751 );
and ( n9753 , n8444 , n537 );
not ( n9754 , n9753 );
not ( n9755 , n9754 );
not ( n9756 , n4659 );
not ( n9757 , n539 );
not ( n9758 , n6033 );
or ( n9759 , n9757 , n9758 );
nand ( n9760 , n5891 , n4477 );
nand ( n9761 , n9759 , n9760 );
not ( n9762 , n9761 );
or ( n9763 , n9756 , n9762 );
nand ( n9764 , n9597 , n4450 );
nand ( n9765 , n9763 , n9764 );
not ( n9766 , n9765 );
or ( n9767 , n9755 , n9766 );
buf ( n9768 , n9754 );
or ( n9769 , n9768 , n9765 );
nand ( n9770 , n9767 , n9769 );
xor ( n9771 , n9752 , n9770 );
xor ( n9772 , n9739 , n9771 );
xor ( n9773 , n9712 , n9772 );
xor ( n9774 , n9724 , n9728 );
xor ( n9775 , n9774 , n9735 );
xor ( n9776 , n5842 , n5954 );
and ( n9777 , n9776 , n6043 );
and ( n9778 , n5842 , n5954 );
or ( n9779 , n9777 , n9778 );
xor ( n9780 , n9775 , n9779 );
xor ( n9781 , n7201 , n7332 );
and ( n9782 , n9781 , n7347 );
and ( n9783 , n7201 , n7332 );
or ( n9784 , n9782 , n9783 );
and ( n9785 , n9780 , n9784 );
and ( n9786 , n9775 , n9779 );
or ( n9787 , n9785 , n9786 );
xor ( n9788 , n9773 , n9787 );
xor ( n9789 , n9617 , n9788 );
xor ( n9790 , n9580 , n9608 );
xor ( n9791 , n9790 , n9613 );
xor ( n9792 , n9411 , n9519 );
xor ( n9793 , n9792 , n9527 );
xor ( n9794 , n9791 , n9793 );
xor ( n9795 , n5598 , n6044 );
and ( n9796 , n9795 , n6091 );
and ( n9797 , n5598 , n6044 );
or ( n9798 , n9796 , n9797 );
and ( n9799 , n9794 , n9798 );
and ( n9800 , n9791 , n9793 );
or ( n9801 , n9799 , n9800 );
xor ( n9802 , n9789 , n9801 );
xor ( n9803 , n9775 , n9779 );
xor ( n9804 , n9803 , n9784 );
xor ( n9805 , n9791 , n9793 );
xor ( n9806 , n9805 , n9798 );
xor ( n9807 , n9804 , n9806 );
xor ( n9808 , n7188 , n7348 );
and ( n9809 , n9808 , n7376 );
and ( n9810 , n7188 , n7348 );
or ( n9811 , n9809 , n9810 );
and ( n9812 , n9807 , n9811 );
and ( n9813 , n9804 , n9806 );
or ( n9814 , n9812 , n9813 );
nor ( n9815 , n9802 , n9814 );
not ( n9816 , n9815 );
xor ( n9817 , n9545 , n9560 );
and ( n9818 , n9817 , n9569 );
and ( n9819 , n9545 , n9560 );
or ( n9820 , n9818 , n9819 );
not ( n9821 , n5786 );
not ( n9822 , n541 );
not ( n9823 , n5467 );
or ( n9824 , n9822 , n9823 );
nand ( n9825 , n5466 , n5734 );
nand ( n9826 , n9824 , n9825 );
not ( n9827 , n9826 );
or ( n9828 , n9821 , n9827 );
nand ( n9829 , n9535 , n5747 );
nand ( n9830 , n9828 , n9829 );
not ( n9831 , n5595 );
not ( n9832 , n545 );
not ( n9833 , n7490 );
or ( n9834 , n9832 , n9833 );
nand ( n9835 , n6618 , n4666 );
nand ( n9836 , n9834 , n9835 );
not ( n9837 , n9836 );
or ( n9838 , n9831 , n9837 );
nand ( n9839 , n9566 , n5341 );
nand ( n9840 , n9838 , n9839 );
xor ( n9841 , n9830 , n9840 );
not ( n9842 , n6095 );
and ( n9843 , n549 , n9692 );
not ( n9844 , n549 );
and ( n9845 , n9844 , n9510 );
or ( n9846 , n9843 , n9845 );
not ( n9847 , n9846 );
or ( n9848 , n9842 , n9847 );
nand ( n9849 , n9702 , n6667 );
nand ( n9850 , n9848 , n9849 );
xor ( n9851 , n9841 , n9850 );
xor ( n9852 , n9820 , n9851 );
nand ( n9853 , n7020 , n7614 );
nand ( n9854 , n9558 , n4671 );
not ( n9855 , n7610 );
nand ( n9856 , n9855 , n7019 );
nand ( n9857 , n9853 , n9854 , n9856 );
xor ( n9858 , n9750 , n9751 );
and ( n9859 , n9858 , n9770 );
and ( n9860 , n9750 , n9751 );
or ( n9861 , n9859 , n9860 );
xor ( n9862 , n9857 , n9861 );
not ( n9863 , n7127 );
not ( n9864 , n9716 );
or ( n9865 , n9863 , n9864 );
nand ( n9866 , n6922 , n6809 );
not ( n9867 , n9866 );
and ( n9868 , n547 , n9867 );
not ( n9869 , n547 );
and ( n9870 , n9869 , n6923 );
or ( n9871 , n9868 , n9870 );
nand ( n9872 , n9871 , n6983 );
nand ( n9873 , n9865 , n9872 );
xor ( n9874 , n9862 , n9873 );
xor ( n9875 , n9852 , n9874 );
xor ( n9876 , n9712 , n9772 );
and ( n9877 , n9876 , n9787 );
and ( n9878 , n9712 , n9772 );
or ( n9879 , n9877 , n9878 );
xor ( n9880 , n9875 , n9879 );
xor ( n9881 , n9718 , n9738 );
and ( n9882 , n9881 , n9771 );
and ( n9883 , n9718 , n9738 );
or ( n9884 , n9882 , n9883 );
not ( n9885 , n7040 );
not ( n9886 , n9689 );
not ( n9887 , n9886 );
not ( n9888 , n9887 );
or ( n9889 , n9885 , n9888 );
not ( n9890 , n551 );
not ( n9891 , n455 );
not ( n9892 , n9475 );
not ( n9893 , n9675 );
not ( n9894 , n9653 );
or ( n9895 , n9893 , n9894 );
nand ( n9896 , n9895 , n9673 );
or ( n9897 , n2122 , n2084 );
nand ( n9898 , n9897 , n489 );
and ( n9899 , n489 , n2152 );
xor ( n9900 , n9898 , n9899 );
not ( n9901 , n9665 );
xor ( n9902 , n9900 , n9901 );
not ( n9903 , n9902 );
xor ( n9904 , n9664 , n9665 );
and ( n9905 , n9904 , n9670 );
and ( n9906 , n9664 , n9665 );
or ( n9907 , n9905 , n9906 );
not ( n9908 , n9907 );
or ( n9909 , n9903 , n9908 );
or ( n9910 , n9907 , n9902 );
nand ( n9911 , n9909 , n9910 );
nor ( n9912 , n9896 , n9911 );
nand ( n9913 , n9892 , n9912 );
nand ( n9914 , n9681 , n9675 );
not ( n9915 , n9911 );
nor ( n9916 , n9914 , n9915 );
nand ( n9917 , n9916 , n9475 );
not ( n9918 , n9911 );
not ( n9919 , n9896 );
nand ( n9920 , n9918 , n9919 , n9914 );
not ( n9921 , n9915 );
nand ( n9922 , n9921 , n9896 );
nand ( n9923 , n9913 , n9917 , n9920 , n9922 );
not ( n9924 , n9923 );
or ( n9925 , n9891 , n9924 );
xor ( n9926 , n9634 , n9635 );
and ( n9927 , n9926 , n9640 );
and ( n9928 , n9634 , n9635 );
or ( n9929 , n9927 , n9928 );
not ( n9930 , n9929 );
not ( n9931 , n9635 );
nand ( n9932 , n505 , n489 );
not ( n9933 , n9932 );
or ( n9934 , n6562 , n1859 );
nand ( n9935 , n9934 , n489 );
not ( n9936 , n9935 );
or ( n9937 , n9933 , n9936 );
or ( n9938 , n9935 , n9932 );
nand ( n9939 , n9937 , n9938 );
not ( n9940 , n9939 );
or ( n9941 , n9931 , n9940 );
or ( n9942 , n9939 , n9635 );
nand ( n9943 , n9941 , n9942 );
not ( n9944 , n9943 );
and ( n9945 , n9930 , n9944 );
and ( n9946 , n9929 , n9943 );
nor ( n9947 , n9945 , n9946 );
not ( n9948 , n9947 );
not ( n9949 , n9948 );
not ( n9950 , n6934 );
not ( n9951 , n6937 );
or ( n9952 , n9950 , n9951 );
and ( n9953 , n9618 , n9642 );
and ( n9954 , n9953 , n7260 );
nand ( n9955 , n9952 , n9954 );
not ( n9956 , n7260 );
not ( n9957 , n6684 );
or ( n9958 , n9956 , n9957 );
nand ( n9959 , n9958 , n7266 );
nand ( n9960 , n9959 , n9953 );
not ( n9961 , n9451 );
not ( n9962 , n7313 );
or ( n9963 , n9961 , n9962 );
nand ( n9964 , n9963 , n9452 );
and ( n9965 , n9964 , n9642 );
not ( n9966 , n9643 );
nor ( n9967 , n9965 , n9966 );
nand ( n9968 , n9955 , n9960 , n9967 );
not ( n9969 , n9968 );
or ( n9970 , n9949 , n9969 );
not ( n9971 , n9967 );
nor ( n9972 , n9971 , n9948 );
nand ( n9973 , n9955 , n9960 , n9972 );
nand ( n9974 , n9970 , n9973 );
nand ( n9975 , n9974 , n793 );
nand ( n9976 , n9925 , n9975 );
not ( n9977 , n9976 );
not ( n9978 , n9977 );
or ( n9979 , n9890 , n9978 );
or ( n9980 , n551 , n9977 );
nand ( n9981 , n9979 , n9980 );
nand ( n9982 , n9981 , n552 );
nand ( n9983 , n9889 , n9982 );
buf ( n9984 , n4450 );
nand ( n9985 , n9761 , n9984 );
nand ( n9986 , n5141 , n5971 );
nand ( n9987 , n5145 , n5977 );
nand ( n9988 , n9985 , n9986 , n9987 );
not ( n9989 , n4450 );
not ( n9990 , n9597 );
or ( n9991 , n9989 , n9990 );
nand ( n9992 , n9761 , n4659 );
nand ( n9993 , n9991 , n9992 );
nand ( n9994 , n9993 , n9753 );
not ( n9995 , n9994 );
xor ( n9996 , n9988 , n9995 );
and ( n9997 , n7400 , n537 );
not ( n9998 , n9997 );
not ( n9999 , n9998 );
or ( n10000 , n9747 , n5903 );
not ( n10001 , n537 );
not ( n10002 , n6056 );
or ( n10003 , n10001 , n10002 );
nand ( n10004 , n6059 , n5605 );
nand ( n10005 , n10003 , n10004 );
nand ( n10006 , n10005 , n5697 );
nand ( n10007 , n10000 , n10006 );
not ( n10008 , n10007 );
or ( n10009 , n9999 , n10008 );
nand ( n10010 , n10006 , n9997 , n10000 );
nand ( n10011 , n10009 , n10010 );
xor ( n10012 , n9996 , n10011 );
xor ( n10013 , n9983 , n10012 );
xor ( n10014 , n9694 , n9706 );
and ( n10015 , n10014 , n9711 );
and ( n10016 , n9694 , n9706 );
or ( n10017 , n10015 , n10016 );
xor ( n10018 , n10013 , n10017 );
xor ( n10019 , n9884 , n10018 );
xor ( n10020 , n9530 , n9570 );
and ( n10021 , n10020 , n9616 );
and ( n10022 , n9530 , n9570 );
or ( n10023 , n10021 , n10022 );
xor ( n10024 , n10019 , n10023 );
xor ( n10025 , n9880 , n10024 );
xor ( n10026 , n9617 , n9788 );
and ( n10027 , n10026 , n9801 );
and ( n10028 , n9617 , n9788 );
or ( n10029 , n10027 , n10028 );
nor ( n10030 , n10025 , n10029 );
not ( n10031 , n10030 );
xor ( n10032 , n9804 , n9806 );
xor ( n10033 , n10032 , n9811 );
not ( n10034 , n10033 );
xor ( n10035 , n6092 , n7183 );
and ( n10036 , n10035 , n7377 );
and ( n10037 , n6092 , n7183 );
or ( n10038 , n10036 , n10037 );
not ( n10039 , n10038 );
nand ( n10040 , n10034 , n10039 );
nand ( n10041 , n9816 , n10031 , n10040 );
or ( n10042 , n9401 , n10041 );
nor ( n10043 , n10030 , n9815 );
nand ( n10044 , n10033 , n10038 );
nand ( n10045 , n9802 , n9814 );
nand ( n10046 , n10044 , n10045 );
and ( n10047 , n10043 , n10046 );
nand ( n10048 , n10025 , n10029 );
not ( n10049 , n10048 );
nor ( n10050 , n10047 , n10049 );
nand ( n10051 , n10042 , n10050 );
buf ( n10052 , n10051 );
buf ( n10053 , n10052 );
xor ( n10054 , n9830 , n9840 );
and ( n10055 , n10054 , n9850 );
and ( n10056 , n9830 , n9840 );
or ( n10057 , n10055 , n10056 );
not ( n10058 , n5786 );
not ( n10059 , n541 );
not ( n10060 , n5588 );
not ( n10061 , n10060 );
or ( n10062 , n10059 , n10061 );
nand ( n10063 , n5588 , n5734 );
nand ( n10064 , n10062 , n10063 );
not ( n10065 , n10064 );
or ( n10066 , n10058 , n10065 );
buf ( n10067 , n5747 );
nand ( n10068 , n9826 , n10067 );
nand ( n10069 , n10066 , n10068 );
not ( n10070 , n5341 );
not ( n10071 , n9836 );
or ( n10072 , n10070 , n10071 );
not ( n10073 , n545 );
not ( n10074 , n6967 );
not ( n10075 , n10074 );
or ( n10076 , n10073 , n10075 );
nand ( n10077 , n6967 , n4666 );
nand ( n10078 , n10076 , n10077 );
nand ( n10079 , n10078 , n5595 );
nand ( n10080 , n10072 , n10079 );
xor ( n10081 , n10069 , n10080 );
not ( n10082 , n6095 );
xor ( n10083 , n549 , n9688 );
not ( n10084 , n10083 );
or ( n10085 , n10082 , n10084 );
nand ( n10086 , n9846 , n6667 );
nand ( n10087 , n10085 , n10086 );
xor ( n10088 , n10081 , n10087 );
xor ( n10089 , n10057 , n10088 );
not ( n10090 , n543 );
not ( n10091 , n7484 );
or ( n10092 , n10090 , n10091 );
nand ( n10093 , n7340 , n5146 );
nand ( n10094 , n10092 , n10093 );
nand ( n10095 , n10094 , n5330 );
not ( n10096 , n7396 );
nand ( n10097 , n10096 , n7016 );
nand ( n10098 , n7015 , n7402 );
nand ( n10099 , n10095 , n10097 , n10098 );
xor ( n10100 , n9988 , n9995 );
and ( n10101 , n10100 , n10011 );
and ( n10102 , n9988 , n9995 );
or ( n10103 , n10101 , n10102 );
xor ( n10104 , n10099 , n10103 );
not ( n10105 , n7026 );
not ( n10106 , n9871 );
or ( n10107 , n10105 , n10106 );
not ( n10108 , n8576 );
not ( n10109 , n7326 );
or ( n10110 , n10108 , n10109 );
or ( n10111 , n7326 , n8576 );
nand ( n10112 , n10110 , n10111 );
nand ( n10113 , n10112 , n6983 );
nand ( n10114 , n10107 , n10113 );
xor ( n10115 , n10104 , n10114 );
xor ( n10116 , n10089 , n10115 );
not ( n10117 , n6974 );
not ( n10118 , n9981 );
or ( n10119 , n10117 , n10118 );
not ( n10120 , n7491 );
nand ( n10121 , n10119 , n10120 );
not ( n10122 , n4660 );
not ( n10123 , n539 );
not ( n10124 , n5322 );
or ( n10125 , n10123 , n10124 );
nand ( n10126 , n5321 , n4477 );
nand ( n10127 , n10125 , n10126 );
not ( n10128 , n10127 );
or ( n10129 , n10122 , n10128 );
not ( n10130 , n5145 );
not ( n10131 , n5964 );
and ( n10132 , n10130 , n10131 );
and ( n10133 , n8090 , n5962 );
nor ( n10134 , n10132 , n10133 );
nand ( n10135 , n10129 , n10134 );
and ( n10136 , n10006 , n10000 );
nor ( n10137 , n10136 , n9998 );
xor ( n10138 , n10135 , n10137 );
and ( n10139 , n4655 , n537 );
not ( n10140 , n5697 );
not ( n10141 , n537 );
not ( n10142 , n7784 );
or ( n10143 , n10141 , n10142 );
nand ( n10144 , n7780 , n5605 );
nand ( n10145 , n10143 , n10144 );
not ( n10146 , n10145 );
or ( n10147 , n10140 , n10146 );
nand ( n10148 , n10005 , n5609 );
nand ( n10149 , n10147 , n10148 );
xor ( n10150 , n10139 , n10149 );
xor ( n10151 , n10138 , n10150 );
xor ( n10152 , n10121 , n10151 );
xor ( n10153 , n9857 , n9861 );
and ( n10154 , n10153 , n9873 );
and ( n10155 , n9857 , n9861 );
or ( n10156 , n10154 , n10155 );
xor ( n10157 , n10152 , n10156 );
xor ( n10158 , n9983 , n10012 );
and ( n10159 , n10158 , n10017 );
and ( n10160 , n9983 , n10012 );
or ( n10161 , n10159 , n10160 );
xor ( n10162 , n10157 , n10161 );
xor ( n10163 , n9820 , n9851 );
and ( n10164 , n10163 , n9874 );
and ( n10165 , n9820 , n9851 );
or ( n10166 , n10164 , n10165 );
xor ( n10167 , n10162 , n10166 );
xor ( n10168 , n10116 , n10167 );
xor ( n10169 , n9884 , n10018 );
and ( n10170 , n10169 , n10023 );
and ( n10171 , n9884 , n10018 );
or ( n10172 , n10170 , n10171 );
xor ( n10173 , n10168 , n10172 );
xor ( n10174 , n9875 , n9879 );
and ( n10175 , n10174 , n10024 );
and ( n10176 , n9875 , n9879 );
or ( n10177 , n10175 , n10176 );
nor ( n10178 , n10173 , n10177 );
not ( n10179 , n10178 );
nand ( n10180 , n10173 , n10177 );
buf ( n10181 , n10180 );
nand ( n10182 , n10179 , n10181 );
not ( n10183 , n10182 );
and ( n10184 , n10053 , n10183 );
not ( n10185 , n10053 );
and ( n10186 , n10185 , n10182 );
nor ( n10187 , n10184 , n10186 );
not ( n10188 , n10187 );
or ( n10189 , n4441 , n10188 );
not ( n10190 , n454 );
not ( n10191 , n504 );
not ( n10192 , n503 );
xor ( n10193 , n529 , n457 );
not ( n10194 , n10193 );
xor ( n10195 , n458 , n459 );
not ( n10196 , n10195 );
not ( n10197 , n10196 );
not ( n10198 , n10197 );
or ( n10199 , n10194 , n10198 );
xnor ( n10200 , n458 , n457 );
xor ( n10201 , n458 , n459 );
nor ( n10202 , n10200 , n10201 );
and ( n10203 , n530 , n457 );
not ( n10204 , n530 );
and ( n10205 , n10204 , n2984 );
nor ( n10206 , n10203 , n10205 );
nand ( n10207 , n10202 , n10206 );
nand ( n10208 , n10199 , n10207 );
xor ( n10209 , n528 , n459 );
not ( n10210 , n10209 );
not ( n10211 , n460 );
nand ( n10212 , n3352 , n10211 , n459 );
nand ( n10213 , n2624 , n460 , n461 );
nand ( n10214 , n10212 , n10213 );
not ( n10215 , n10214 );
not ( n10216 , n10215 );
not ( n10217 , n10216 );
or ( n10218 , n10210 , n10217 );
and ( n10219 , n461 , n460 );
not ( n10220 , n461 );
and ( n10221 , n10220 , n2801 );
nor ( n10222 , n10219 , n10221 );
buf ( n10223 , n10222 );
xor ( n10224 , n527 , n459 );
nand ( n10225 , n10223 , n10224 );
nand ( n10226 , n10218 , n10225 );
xor ( n10227 , n10208 , n10226 );
xor ( n10228 , n524 , n463 );
not ( n10229 , n10228 );
not ( n10230 , n465 );
and ( n10231 , n464 , n10230 );
not ( n10232 , n464 );
and ( n10233 , n10232 , n465 );
nor ( n10234 , n10231 , n10233 );
xor ( n10235 , n464 , n463 );
nand ( n10236 , n10234 , n10235 );
not ( n10237 , n10236 );
not ( n10238 , n10237 );
or ( n10239 , n10229 , n10238 );
xor ( n10240 , n464 , n465 );
buf ( n10241 , n10240 );
xor ( n10242 , n463 , n523 );
nand ( n10243 , n10241 , n10242 );
nand ( n10244 , n10239 , n10243 );
and ( n10245 , n10227 , n10244 );
and ( n10246 , n10208 , n10226 );
or ( n10247 , n10245 , n10246 );
not ( n10248 , n10224 );
not ( n10249 , n10214 );
or ( n10250 , n10248 , n10249 );
xor ( n10251 , n526 , n459 );
nand ( n10252 , n10223 , n10251 );
nand ( n10253 , n10250 , n10252 );
not ( n10254 , n10193 );
nor ( n10255 , n10200 , n10201 );
buf ( n10256 , n10255 );
not ( n10257 , n10256 );
or ( n10258 , n10254 , n10257 );
xor ( n10259 , n457 , n528 );
nand ( n10260 , n10197 , n10259 );
nand ( n10261 , n10258 , n10260 );
xor ( n10262 , n10253 , n10261 );
xor ( n10263 , n521 , n465 );
not ( n10264 , n10263 );
nand ( n10265 , n2827 , n467 );
not ( n10266 , n467 );
nand ( n10267 , n10266 , n466 );
nand ( n10268 , n10265 , n10267 );
not ( n10269 , n10268 );
xor ( n10270 , n466 , n465 );
and ( n10271 , n10269 , n10270 );
not ( n10272 , n10271 );
or ( n10273 , n10264 , n10272 );
xor ( n10274 , n466 , n467 );
nand ( n10275 , n10274 , n465 );
nand ( n10276 , n10273 , n10275 );
xor ( n10277 , n10262 , n10276 );
xor ( n10278 , n10247 , n10277 );
not ( n10279 , n468 );
and ( n10280 , n10279 , n469 );
not ( n10281 , n469 );
and ( n10282 , n10281 , n468 );
nor ( n10283 , n10280 , n10282 );
not ( n10284 , n10283 );
xnor ( n10285 , n468 , n469 );
xor ( n10286 , n468 , n467 );
nand ( n10287 , n10285 , n10286 );
not ( n10288 , n10287 );
buf ( n10289 , n10288 );
not ( n10290 , n10289 );
not ( n10291 , n10290 );
or ( n10292 , n10284 , n10291 );
nand ( n10293 , n10292 , n467 );
not ( n10294 , n10293 );
xor ( n10295 , n522 , n465 );
not ( n10296 , n10295 );
not ( n10297 , n10271 );
or ( n10298 , n10296 , n10297 );
nand ( n10299 , n10274 , n10263 );
nand ( n10300 , n10298 , n10299 );
not ( n10301 , n10300 );
or ( n10302 , n10294 , n10301 );
nor ( n10303 , n10293 , n10300 );
xor ( n10304 , n526 , n461 );
not ( n10305 , n10304 );
xor ( n10306 , n461 , n462 );
not ( n10307 , n10306 );
and ( n10308 , n462 , n463 );
not ( n10309 , n462 );
not ( n10310 , n463 );
and ( n10311 , n10309 , n10310 );
nor ( n10312 , n10308 , n10311 );
or ( n10313 , n10307 , n10312 );
not ( n10314 , n10313 );
not ( n10315 , n10314 );
or ( n10316 , n10305 , n10315 );
xor ( n10317 , n462 , n463 );
xor ( n10318 , n525 , n461 );
nand ( n10319 , n10317 , n10318 );
nand ( n10320 , n10316 , n10319 );
not ( n10321 , n10320 );
or ( n10322 , n10303 , n10321 );
nand ( n10323 , n10302 , n10322 );
and ( n10324 , n10278 , n10323 );
and ( n10325 , n10247 , n10277 );
or ( n10326 , n10324 , n10325 );
not ( n10327 , n10251 );
not ( n10328 , n10214 );
or ( n10329 , n10327 , n10328 );
xor ( n10330 , n525 , n459 );
nand ( n10331 , n10223 , n10330 );
nand ( n10332 , n10329 , n10331 );
xor ( n10333 , n522 , n463 );
not ( n10334 , n10333 );
not ( n10335 , n10237 );
or ( n10336 , n10334 , n10335 );
xor ( n10337 , n521 , n463 );
nand ( n10338 , n10241 , n10337 );
nand ( n10339 , n10336 , n10338 );
xor ( n10340 , n10332 , n10339 );
not ( n10341 , n10274 );
not ( n10342 , n10341 );
xnor ( n10343 , n466 , n467 );
nand ( n10344 , n10343 , n10270 );
not ( n10345 , n10344 );
or ( n10346 , n10342 , n10345 );
nand ( n10347 , n10346 , n465 );
xor ( n10348 , n10340 , n10347 );
not ( n10349 , n10348 );
nand ( n10350 , n530 , n457 );
not ( n10351 , n10350 );
not ( n10352 , n10351 );
not ( n10353 , n10242 );
not ( n10354 , n10237 );
or ( n10355 , n10353 , n10354 );
nand ( n10356 , n10241 , n10333 );
nand ( n10357 , n10355 , n10356 );
not ( n10358 , n10357 );
not ( n10359 , n10358 );
or ( n10360 , n10352 , n10359 );
not ( n10361 , n10350 );
not ( n10362 , n10357 );
or ( n10363 , n10361 , n10362 );
not ( n10364 , n463 );
nand ( n10365 , n10364 , n462 );
nand ( n10366 , n2224 , n463 );
nand ( n10367 , n10365 , n10366 );
xor ( n10368 , n524 , n461 );
nand ( n10369 , n10367 , n10368 );
and ( n10370 , n462 , n463 );
not ( n10371 , n462 );
and ( n10372 , n10371 , n10310 );
nor ( n10373 , n10370 , n10372 );
not ( n10374 , n10373 );
nand ( n10375 , n10374 , n10306 );
not ( n10376 , n10375 );
nand ( n10377 , n10318 , n10376 );
nand ( n10378 , n10369 , n10377 );
nand ( n10379 , n10363 , n10378 );
nand ( n10380 , n10360 , n10379 );
not ( n10381 , n10380 );
not ( n10382 , n10381 );
and ( n10383 , n10349 , n10382 );
and ( n10384 , n10348 , n10381 );
nor ( n10385 , n10383 , n10384 );
nand ( n10386 , n529 , n457 );
not ( n10387 , n10259 );
not ( n10388 , n10256 );
or ( n10389 , n10387 , n10388 );
xor ( n10390 , n457 , n527 );
nand ( n10391 , n10197 , n10390 );
nand ( n10392 , n10389 , n10391 );
xor ( n10393 , n10386 , n10392 );
not ( n10394 , n10368 );
not ( n10395 , n10314 );
or ( n10396 , n10394 , n10395 );
xor ( n10397 , n523 , n461 );
nand ( n10398 , n10317 , n10397 );
nand ( n10399 , n10396 , n10398 );
xnor ( n10400 , n10393 , n10399 );
xor ( n10401 , n10357 , n10400 );
or ( n10402 , n10253 , n10261 );
nand ( n10403 , n10402 , n10276 );
nand ( n10404 , n10253 , n10261 );
nand ( n10405 , n10403 , n10404 );
xor ( n10406 , n10401 , n10405 );
or ( n10407 , n10385 , n10406 );
nand ( n10408 , n10406 , n10385 );
nand ( n10409 , n10407 , n10408 );
xor ( n10410 , n10326 , n10409 );
xor ( n10411 , n10208 , n10226 );
xor ( n10412 , n10411 , n10244 );
not ( n10413 , n10412 );
and ( n10414 , n532 , n457 );
xnor ( n10415 , n458 , n457 );
nor ( n10416 , n10415 , n10201 );
not ( n10417 , n10416 );
xor ( n10418 , n531 , n457 );
not ( n10419 , n10418 );
or ( n10420 , n10417 , n10419 );
nand ( n10421 , n10195 , n10206 );
nand ( n10422 , n10420 , n10421 );
xor ( n10423 , n10414 , n10422 );
xor ( n10424 , n525 , n463 );
not ( n10425 , n10424 );
not ( n10426 , n10237 );
or ( n10427 , n10425 , n10426 );
nand ( n10428 , n10241 , n10228 );
nand ( n10429 , n10427 , n10428 );
and ( n10430 , n10423 , n10429 );
and ( n10431 , n10414 , n10422 );
or ( n10432 , n10430 , n10431 );
not ( n10433 , n10432 );
or ( n10434 , n10413 , n10433 );
nor ( n10435 , n10412 , n10432 );
xor ( n10436 , n10300 , n10293 );
and ( n10437 , n10436 , n10321 );
not ( n10438 , n10436 );
and ( n10439 , n10438 , n10320 );
nor ( n10440 , n10437 , n10439 );
or ( n10441 , n10435 , n10440 );
nand ( n10442 , n10434 , n10441 );
not ( n10443 , n10442 );
xor ( n10444 , n521 , n467 );
not ( n10445 , n10444 );
not ( n10446 , n10288 );
or ( n10447 , n10445 , n10446 );
not ( n10448 , n468 );
not ( n10449 , n10281 );
or ( n10450 , n10448 , n10449 );
nand ( n10451 , n10279 , n469 );
nand ( n10452 , n10450 , n10451 );
nand ( n10453 , n10452 , n467 );
nand ( n10454 , n10447 , n10453 );
not ( n10455 , n10454 );
nand ( n10456 , n531 , n457 );
nand ( n10457 , n10455 , n10456 );
not ( n10458 , n10457 );
not ( n10459 , n3352 );
not ( n10460 , n463 );
and ( n10461 , n10459 , n10460 );
nor ( n10462 , n10461 , n462 );
not ( n10463 , n10462 );
xor ( n10464 , n527 , n461 );
not ( n10465 , n462 );
not ( n10466 , n463 );
nor ( n10467 , n10466 , n461 );
nor ( n10468 , n10465 , n10467 );
not ( n10469 , n10468 );
nand ( n10470 , n10463 , n10464 , n10469 );
nand ( n10471 , n10365 , n10366 );
nand ( n10472 , n10471 , n10304 );
nand ( n10473 , n10470 , n10472 );
xor ( n10474 , n465 , n523 );
not ( n10475 , n10474 );
not ( n10476 , n10344 );
not ( n10477 , n10476 );
or ( n10478 , n10475 , n10477 );
xor ( n10479 , n467 , n466 );
buf ( n10480 , n10479 );
nand ( n10481 , n10480 , n10295 );
nand ( n10482 , n10478 , n10481 );
xor ( n10483 , n10473 , n10482 );
xor ( n10484 , n529 , n459 );
not ( n10485 , n10484 );
not ( n10486 , n10214 );
or ( n10487 , n10485 , n10486 );
nand ( n10488 , n10223 , n10209 );
nand ( n10489 , n10487 , n10488 );
and ( n10490 , n10483 , n10489 );
and ( n10491 , n10473 , n10482 );
or ( n10492 , n10490 , n10491 );
not ( n10493 , n10492 );
or ( n10494 , n10458 , n10493 );
not ( n10495 , n10456 );
nand ( n10496 , n10454 , n10495 );
nand ( n10497 , n10494 , n10496 );
not ( n10498 , n10497 );
xor ( n10499 , n10351 , n10358 );
xor ( n10500 , n10499 , n10378 );
not ( n10501 , n10500 );
nand ( n10502 , n10498 , n10501 );
not ( n10503 , n10502 );
or ( n10504 , n10443 , n10503 );
not ( n10505 , n10501 );
nand ( n10506 , n10505 , n10497 );
nand ( n10507 , n10504 , n10506 );
and ( n10508 , n10410 , n10507 );
and ( n10509 , n10326 , n10409 );
or ( n10510 , n10508 , n10509 );
not ( n10511 , n10510 );
not ( n10512 , n10348 );
nand ( n10513 , n10512 , n10381 );
not ( n10514 , n10513 );
not ( n10515 , n10406 );
or ( n10516 , n10514 , n10515 );
nand ( n10517 , n10348 , n10380 );
nand ( n10518 , n10516 , n10517 );
not ( n10519 , n10518 );
not ( n10520 , n10519 );
xor ( n10521 , n10357 , n10400 );
and ( n10522 , n10521 , n10405 );
and ( n10523 , n10357 , n10400 );
or ( n10524 , n10522 , n10523 );
not ( n10525 , n10524 );
not ( n10526 , n10525 );
xor ( n10527 , n10332 , n10339 );
and ( n10528 , n10527 , n10347 );
and ( n10529 , n10332 , n10339 );
or ( n10530 , n10528 , n10529 );
and ( n10531 , n457 , n528 );
not ( n10532 , n10390 );
not ( n10533 , n10256 );
or ( n10534 , n10532 , n10533 );
xor ( n10535 , n457 , n526 );
nand ( n10536 , n10197 , n10535 );
nand ( n10537 , n10534 , n10536 );
xor ( n10538 , n10531 , n10537 );
not ( n10539 , n10337 );
not ( n10540 , n10237 );
or ( n10541 , n10539 , n10540 );
nand ( n10542 , n463 , n10241 );
nand ( n10543 , n10541 , n10542 );
xor ( n10544 , n10538 , n10543 );
xor ( n10545 , n10530 , n10544 );
not ( n10546 , n10330 );
not ( n10547 , n10216 );
or ( n10548 , n10546 , n10547 );
xor ( n10549 , n459 , n524 );
nand ( n10550 , n10223 , n10549 );
nand ( n10551 , n10548 , n10550 );
not ( n10552 , n10551 );
not ( n10553 , n10397 );
not ( n10554 , n10376 );
or ( n10555 , n10553 , n10554 );
xor ( n10556 , n522 , n461 );
nand ( n10557 , n10556 , n10471 );
nand ( n10558 , n10555 , n10557 );
not ( n10559 , n10558 );
and ( n10560 , n10552 , n10559 );
and ( n10561 , n10551 , n10558 );
nor ( n10562 , n10560 , n10561 );
not ( n10563 , n10562 );
not ( n10564 , n10386 );
not ( n10565 , n10564 );
not ( n10566 , n10399 );
or ( n10567 , n10565 , n10566 );
or ( n10568 , n10399 , n10564 );
not ( n10569 , n10259 );
not ( n10570 , n10256 );
or ( n10571 , n10569 , n10570 );
nand ( n10572 , n10571 , n10391 );
nand ( n10573 , n10568 , n10572 );
nand ( n10574 , n10567 , n10573 );
not ( n10575 , n10574 );
or ( n10576 , n10563 , n10575 );
or ( n10577 , n10574 , n10562 );
nand ( n10578 , n10576 , n10577 );
xor ( n10579 , n10545 , n10578 );
not ( n10580 , n10579 );
or ( n10581 , n10526 , n10580 );
not ( n10582 , n10579 );
nand ( n10583 , n10582 , n10524 );
nand ( n10584 , n10581 , n10583 );
not ( n10585 , n10584 );
not ( n10586 , n10585 );
or ( n10587 , n10520 , n10586 );
nand ( n10588 , n10518 , n10584 );
nand ( n10589 , n10587 , n10588 );
nand ( n10590 , n10511 , n10589 );
not ( n10591 , n10590 );
xor ( n10592 , n468 , n469 );
not ( n10593 , n10592 );
not ( n10594 , n10444 );
or ( n10595 , n10593 , n10594 );
xor ( n10596 , n468 , n469 );
not ( n10597 , n10596 );
xor ( n10598 , n522 , n467 );
nand ( n10599 , n10597 , n10598 , n10286 );
nand ( n10600 , n10595 , n10599 );
xor ( n10601 , n526 , n463 );
not ( n10602 , n10601 );
and ( n10603 , n10234 , n10235 );
not ( n10604 , n10603 );
or ( n10605 , n10602 , n10604 );
nand ( n10606 , n10241 , n10424 );
nand ( n10607 , n10605 , n10606 );
xor ( n10608 , n10600 , n10607 );
xor ( n10609 , n470 , n471 );
not ( n10610 , n10609 );
not ( n10611 , n10610 );
xor ( n10612 , n470 , n469 );
not ( n10613 , n10612 );
xor ( n10614 , n470 , n471 );
nor ( n10615 , n10613 , n10614 );
not ( n10616 , n10615 );
not ( n10617 , n10616 );
or ( n10618 , n10611 , n10617 );
nand ( n10619 , n10618 , n469 );
and ( n10620 , n10608 , n10619 );
and ( n10621 , n10600 , n10607 );
or ( n10622 , n10620 , n10621 );
xor ( n10623 , n10455 , n10622 );
and ( n10624 , n524 , n465 );
not ( n10625 , n524 );
not ( n10626 , n465 );
and ( n10627 , n10625 , n10626 );
nor ( n10628 , n10624 , n10627 );
not ( n10629 , n10628 );
not ( n10630 , n10271 );
or ( n10631 , n10629 , n10630 );
nand ( n10632 , n10480 , n10474 );
nand ( n10633 , n10631 , n10632 );
and ( n10634 , n533 , n457 );
or ( n10635 , n10633 , n10634 );
xor ( n10636 , n528 , n461 );
not ( n10637 , n10636 );
not ( n10638 , n10376 );
or ( n10639 , n10637 , n10638 );
nand ( n10640 , n10367 , n10464 );
nand ( n10641 , n10639 , n10640 );
nand ( n10642 , n10635 , n10641 );
nand ( n10643 , n10633 , n10634 );
nand ( n10644 , n10642 , n10643 );
and ( n10645 , n10623 , n10644 );
and ( n10646 , n10455 , n10622 );
or ( n10647 , n10645 , n10646 );
not ( n10648 , n10492 );
not ( n10649 , n10455 );
not ( n10650 , n10495 );
and ( n10651 , n10649 , n10650 );
and ( n10652 , n10455 , n10495 );
nor ( n10653 , n10651 , n10652 );
not ( n10654 , n10653 );
or ( n10655 , n10648 , n10654 );
or ( n10656 , n10492 , n10653 );
nand ( n10657 , n10655 , n10656 );
xor ( n10658 , n10647 , n10657 );
xor ( n10659 , n10414 , n10422 );
xor ( n10660 , n10659 , n10429 );
xor ( n10661 , n532 , n457 );
not ( n10662 , n10661 );
not ( n10663 , n10256 );
or ( n10664 , n10662 , n10663 );
nand ( n10665 , n10197 , n10418 );
nand ( n10666 , n10664 , n10665 );
not ( n10667 , n10666 );
not ( n10668 , n10214 );
xor ( n10669 , n530 , n459 );
not ( n10670 , n10669 );
or ( n10671 , n10668 , n10670 );
nand ( n10672 , n10223 , n10484 );
nand ( n10673 , n10671 , n10672 );
not ( n10674 , n10673 );
or ( n10675 , n10667 , n10674 );
or ( n10676 , n10673 , n10666 );
xor ( n10677 , n521 , n469 );
not ( n10678 , n10677 );
not ( n10679 , n470 );
nand ( n10680 , n10679 , n471 );
not ( n10681 , n471 );
nand ( n10682 , n10681 , n470 );
and ( n10683 , n10680 , n10682 , n10612 );
not ( n10684 , n10683 );
or ( n10685 , n10678 , n10684 );
buf ( n10686 , n10609 );
nand ( n10687 , n469 , n10686 );
nand ( n10688 , n10685 , n10687 );
nand ( n10689 , n10676 , n10688 );
nand ( n10690 , n10675 , n10689 );
xor ( n10691 , n10660 , n10690 );
xor ( n10692 , n10473 , n10482 );
xor ( n10693 , n10692 , n10489 );
and ( n10694 , n10691 , n10693 );
and ( n10695 , n10660 , n10690 );
or ( n10696 , n10694 , n10695 );
xnor ( n10697 , n10658 , n10696 );
not ( n10698 , n10697 );
not ( n10699 , n10698 );
not ( n10700 , n10440 );
not ( n10701 , n10700 );
not ( n10702 , n10701 );
xor ( n10703 , n10412 , n10432 );
not ( n10704 , n10703 );
not ( n10705 , n10704 );
or ( n10706 , n10702 , n10705 );
nand ( n10707 , n10703 , n10700 );
nand ( n10708 , n10706 , n10707 );
not ( n10709 , n10708 );
not ( n10710 , n10709 );
or ( n10711 , n10699 , n10710 );
not ( n10712 , n10708 );
not ( n10713 , n10697 );
or ( n10714 , n10712 , n10713 );
xor ( n10715 , n527 , n463 );
not ( n10716 , n10715 );
not ( n10717 , n10603 );
or ( n10718 , n10716 , n10717 );
nand ( n10719 , n10241 , n10601 );
nand ( n10720 , n10718 , n10719 );
not ( n10721 , n10720 );
not ( n10722 , n10592 );
and ( n10723 , n467 , n523 );
not ( n10724 , n467 );
not ( n10725 , n523 );
and ( n10726 , n10724 , n10725 );
nor ( n10727 , n10723 , n10726 );
nand ( n10728 , n10727 , n10286 );
and ( n10729 , n10722 , n10728 );
not ( n10730 , n10722 );
not ( n10731 , n10598 );
and ( n10732 , n10730 , n10731 );
nor ( n10733 , n10729 , n10732 );
nand ( n10734 , n534 , n457 );
not ( n10735 , n10734 );
nor ( n10736 , n10733 , n10735 );
not ( n10737 , n10736 );
not ( n10738 , n10737 );
or ( n10739 , n10721 , n10738 );
not ( n10740 , n10734 );
nand ( n10741 , n10740 , n10733 );
nand ( n10742 , n10739 , n10741 );
not ( n10743 , n10268 );
not ( n10744 , n10628 );
or ( n10745 , n10743 , n10744 );
xor ( n10746 , n525 , n465 );
nand ( n10747 , n10746 , n10270 );
or ( n10748 , n10747 , n10479 );
nand ( n10749 , n10745 , n10748 );
xor ( n10750 , n529 , n461 );
not ( n10751 , n10750 );
not ( n10752 , n10376 );
or ( n10753 , n10751 , n10752 );
nand ( n10754 , n10471 , n10636 );
nand ( n10755 , n10753 , n10754 );
xor ( n10756 , n10749 , n10755 );
xor ( n10757 , n531 , n459 );
not ( n10758 , n10757 );
not ( n10759 , n10214 );
or ( n10760 , n10758 , n10759 );
nand ( n10761 , n10222 , n10669 );
nand ( n10762 , n10760 , n10761 );
and ( n10763 , n10756 , n10762 );
and ( n10764 , n10749 , n10755 );
or ( n10765 , n10763 , n10764 );
xor ( n10766 , n10742 , n10765 );
xor ( n10767 , n10600 , n10607 );
xor ( n10768 , n10767 , n10619 );
and ( n10769 , n10766 , n10768 );
and ( n10770 , n10742 , n10765 );
or ( n10771 , n10769 , n10770 );
xor ( n10772 , n10455 , n10622 );
xor ( n10773 , n10772 , n10644 );
xor ( n10774 , n10771 , n10773 );
xor ( n10775 , n10660 , n10690 );
xor ( n10776 , n10775 , n10693 );
and ( n10777 , n10774 , n10776 );
and ( n10778 , n10771 , n10773 );
or ( n10779 , n10777 , n10778 );
nand ( n10780 , n10714 , n10779 );
nand ( n10781 , n10711 , n10780 );
not ( n10782 , n10781 );
xor ( n10783 , n10247 , n10277 );
xor ( n10784 , n10783 , n10323 );
not ( n10785 , n10501 );
not ( n10786 , n10497 );
or ( n10787 , n10785 , n10786 );
or ( n10788 , n10497 , n10501 );
nand ( n10789 , n10787 , n10788 );
xor ( n10790 , n10789 , n10442 );
xor ( n10791 , n10784 , n10790 );
buf ( n10792 , n10647 );
not ( n10793 , n10792 );
not ( n10794 , n10657 );
or ( n10795 , n10793 , n10794 );
or ( n10796 , n10657 , n10792 );
nand ( n10797 , n10796 , n10696 );
nand ( n10798 , n10795 , n10797 );
xor ( n10799 , n10791 , n10798 );
not ( n10800 , n10799 );
and ( n10801 , n10782 , n10800 );
xor ( n10802 , n10784 , n10790 );
and ( n10803 , n10802 , n10798 );
and ( n10804 , n10784 , n10790 );
or ( n10805 , n10803 , n10804 );
xor ( n10806 , n10326 , n10409 );
xor ( n10807 , n10806 , n10507 );
nor ( n10808 , n10805 , n10807 );
nor ( n10809 , n10801 , n10808 );
buf ( n10810 , n10809 );
not ( n10811 , n10810 );
nor ( n10812 , n10591 , n10811 );
not ( n10813 , n10812 );
xor ( n10814 , n524 , n467 );
not ( n10815 , n10814 );
not ( n10816 , n10286 );
nor ( n10817 , n10816 , n10592 );
not ( n10818 , n10817 );
or ( n10819 , n10815 , n10818 );
nand ( n10820 , n10596 , n10727 );
nand ( n10821 , n10819 , n10820 );
xor ( n10822 , n528 , n463 );
not ( n10823 , n10822 );
not ( n10824 , n10237 );
or ( n10825 , n10823 , n10824 );
nand ( n10826 , n10241 , n10715 );
nand ( n10827 , n10825 , n10826 );
xor ( n10828 , n10821 , n10827 );
xor ( n10829 , n522 , n469 );
not ( n10830 , n10829 );
buf ( n10831 , n10683 );
not ( n10832 , n10831 );
or ( n10833 , n10830 , n10832 );
nand ( n10834 , n10686 , n10677 );
nand ( n10835 , n10833 , n10834 );
xor ( n10836 , n10828 , n10835 );
not ( n10837 , n10836 );
and ( n10838 , n534 , n2984 );
not ( n10839 , n534 );
and ( n10840 , n10839 , n457 );
nor ( n10841 , n10838 , n10840 );
not ( n10842 , n10841 );
not ( n10843 , n10842 );
not ( n10844 , n10202 );
or ( n10845 , n10843 , n10844 );
xor ( n10846 , n533 , n457 );
nand ( n10847 , n10195 , n10846 );
nand ( n10848 , n10845 , n10847 );
nand ( n10849 , n535 , n457 );
not ( n10850 , n10849 );
not ( n10851 , n471 );
and ( n10852 , n10850 , n10851 );
not ( n10853 , n10850 );
not ( n10854 , n10681 );
and ( n10855 , n10853 , n10854 );
or ( n10856 , n10852 , n10855 );
and ( n10857 , n10848 , n10856 );
not ( n10858 , n10848 );
not ( n10859 , n471 );
and ( n10860 , n10849 , n10859 );
not ( n10861 , n10849 );
not ( n10862 , n10681 );
and ( n10863 , n10861 , n10862 );
or ( n10864 , n10860 , n10863 );
and ( n10865 , n10858 , n10864 );
or ( n10866 , n10857 , n10865 );
not ( n10867 , n10866 );
nand ( n10868 , n10837 , n10867 );
nand ( n10869 , n10836 , n10866 );
nand ( n10870 , n10868 , n10869 );
xor ( n10871 , n461 , n532 );
not ( n10872 , n10871 );
not ( n10873 , n10376 );
or ( n10874 , n10872 , n10873 );
and ( n10875 , n461 , n531 );
not ( n10876 , n461 );
not ( n10877 , n531 );
and ( n10878 , n10876 , n10877 );
nor ( n10879 , n10875 , n10878 );
nand ( n10880 , n10317 , n10879 );
nand ( n10881 , n10874 , n10880 );
not ( n10882 , n10881 );
not ( n10883 , n10596 );
xor ( n10884 , n525 , n467 );
not ( n10885 , n10884 );
or ( n10886 , n10883 , n10885 );
xor ( n10887 , n526 , n467 );
nand ( n10888 , n10283 , n10286 , n10887 );
nand ( n10889 , n10886 , n10888 );
xor ( n10890 , n529 , n463 );
not ( n10891 , n10890 );
not ( n10892 , n10234 );
not ( n10893 , n10892 );
or ( n10894 , n10891 , n10893 );
and ( n10895 , n530 , n463 );
not ( n10896 , n530 );
and ( n10897 , n10896 , n2650 );
nor ( n10898 , n10895 , n10897 );
and ( n10899 , n10235 , n10898 );
not ( n10900 , n10240 );
nand ( n10901 , n10899 , n10900 );
nand ( n10902 , n10894 , n10901 );
or ( n10903 , n10889 , n10902 );
not ( n10904 , n10903 );
or ( n10905 , n10882 , n10904 );
nand ( n10906 , n10889 , n10902 );
nand ( n10907 , n10905 , n10906 );
not ( n10908 , n10907 );
or ( n10909 , n536 , n458 );
nand ( n10910 , n10909 , n459 );
nand ( n10911 , n536 , n458 );
and ( n10912 , n10910 , n10911 , n457 );
and ( n10913 , n522 , n471 );
not ( n10914 , n522 );
not ( n10915 , n471 );
and ( n10916 , n10914 , n10915 );
nor ( n10917 , n10913 , n10916 );
not ( n10918 , n10917 );
not ( n10919 , n471 );
nor ( n10920 , n10919 , n472 );
not ( n10921 , n10920 );
or ( n10922 , n10918 , n10921 );
xor ( n10923 , n521 , n471 );
nand ( n10924 , n10923 , n472 );
nand ( n10925 , n10922 , n10924 );
and ( n10926 , n10912 , n10925 );
not ( n10927 , n10926 );
not ( n10928 , n10610 );
and ( n10929 , n523 , n469 );
not ( n10930 , n523 );
and ( n10931 , n10930 , n10281 );
nor ( n10932 , n10929 , n10931 );
nand ( n10933 , n10928 , n10932 );
and ( n10934 , n524 , n10281 );
not ( n10935 , n524 );
and ( n10936 , n10935 , n469 );
or ( n10937 , n10934 , n10936 );
nand ( n10938 , n10610 , n10612 , n10937 );
nor ( n10939 , n10415 , n10201 );
xor ( n10940 , n536 , n457 );
nand ( n10941 , n10939 , n10940 );
buf ( n10942 , n10195 );
not ( n10943 , n535 );
not ( n10944 , n10943 );
not ( n10945 , n457 );
or ( n10946 , n10944 , n10945 );
nand ( n10947 , n2984 , n535 );
nand ( n10948 , n10946 , n10947 );
nand ( n10949 , n10942 , n10948 );
nand ( n10950 , n10933 , n10938 , n10941 , n10949 );
xor ( n10951 , n528 , n465 );
and ( n10952 , n10270 , n10951 );
not ( n10953 , n10952 );
not ( n10954 , n10480 );
not ( n10955 , n10954 );
or ( n10956 , n10953 , n10955 );
xor ( n10957 , n527 , n465 );
nand ( n10958 , n10957 , n10480 );
nand ( n10959 , n10956 , n10958 );
nand ( n10960 , n10950 , n10959 );
nand ( n10961 , n10941 , n10949 );
nand ( n10962 , n10937 , n10612 );
not ( n10963 , n10962 );
not ( n10964 , n10686 );
and ( n10965 , n10963 , n10964 );
or ( n10966 , n10725 , n469 );
or ( n10967 , n10281 , n523 );
nand ( n10968 , n10966 , n10967 );
and ( n10969 , n10968 , n10609 );
nor ( n10970 , n10965 , n10969 );
not ( n10971 , n10970 );
nand ( n10972 , n10961 , n10971 );
nand ( n10973 , n10927 , n10960 , n10972 );
not ( n10974 , n10973 );
or ( n10975 , n10908 , n10974 );
nand ( n10976 , n10960 , n10972 );
nand ( n10977 , n10926 , n10976 );
nand ( n10978 , n10975 , n10977 );
xor ( n10979 , n10870 , n10978 );
xor ( n10980 , n534 , n459 );
not ( n10981 , n10980 );
not ( n10982 , n10216 );
or ( n10983 , n10981 , n10982 );
xor ( n10984 , n459 , n533 );
nand ( n10985 , n10223 , n10984 );
nand ( n10986 , n10983 , n10985 );
xor ( n10987 , n10912 , n10925 );
xor ( n10988 , n10986 , n10987 );
xor ( n10989 , n525 , n469 );
not ( n10990 , n10989 );
not ( n10991 , n10683 );
or ( n10992 , n10990 , n10991 );
nand ( n10993 , n10686 , n10937 );
nand ( n10994 , n10992 , n10993 );
not ( n10995 , n10994 );
and ( n10996 , n471 , n523 );
not ( n10997 , n471 );
and ( n10998 , n10997 , n10725 );
nor ( n10999 , n10996 , n10998 );
not ( n11000 , n10999 );
not ( n11001 , n471 );
nor ( n11002 , n11001 , n472 );
not ( n11003 , n11002 );
or ( n11004 , n11000 , n11003 );
nand ( n11005 , n10917 , n472 );
nand ( n11006 , n11004 , n11005 );
not ( n11007 , n11006 );
nand ( n11008 , n536 , n10195 );
nand ( n11009 , n11007 , n11008 );
not ( n11010 , n11009 );
or ( n11011 , n10995 , n11010 );
not ( n11012 , n11008 );
nand ( n11013 , n11012 , n11006 );
nand ( n11014 , n11011 , n11013 );
and ( n11015 , n10988 , n11014 );
and ( n11016 , n10986 , n10987 );
or ( n11017 , n11015 , n11016 );
xor ( n11018 , n10926 , n10976 );
xor ( n11019 , n11018 , n10907 );
xor ( n11020 , n11017 , n11019 );
not ( n11021 , n10902 );
xor ( n11022 , n10889 , n11021 );
xor ( n11023 , n11022 , n10881 );
not ( n11024 , n11023 );
not ( n11025 , n11024 );
not ( n11026 , n10959 );
not ( n11027 , n10961 );
and ( n11028 , n11027 , n10970 );
not ( n11029 , n11027 );
or ( n11030 , n10962 , n10928 );
nand ( n11031 , n11030 , n10933 );
and ( n11032 , n11029 , n11031 );
nor ( n11033 , n11028 , n11032 );
not ( n11034 , n11033 );
not ( n11035 , n11034 );
or ( n11036 , n11026 , n11035 );
not ( n11037 , n10959 );
nand ( n11038 , n11037 , n11033 );
nand ( n11039 , n11036 , n11038 );
not ( n11040 , n11039 );
or ( n11041 , n11025 , n11040 );
or ( n11042 , n11039 , n11024 );
xor ( n11043 , n531 , n463 );
not ( n11044 , n11043 );
not ( n11045 , n10603 );
or ( n11046 , n11044 , n11045 );
nand ( n11047 , n10241 , n10898 );
nand ( n11048 , n11046 , n11047 );
xor ( n11049 , n529 , n465 );
not ( n11050 , n11049 );
not ( n11051 , n10270 );
buf ( n11052 , n10479 );
nor ( n11053 , n11051 , n11052 );
not ( n11054 , n11053 );
or ( n11055 , n11050 , n11054 );
nand ( n11056 , n11052 , n10951 );
nand ( n11057 , n11055 , n11056 );
xor ( n11058 , n11048 , n11057 );
not ( n11059 , n10596 );
not ( n11060 , n11059 );
not ( n11061 , n11060 );
not ( n11062 , n10887 );
or ( n11063 , n11061 , n11062 );
xor ( n11064 , n467 , n527 );
nand ( n11065 , n10288 , n11064 );
nand ( n11066 , n11063 , n11065 );
and ( n11067 , n11058 , n11066 );
and ( n11068 , n11048 , n11057 );
or ( n11069 , n11067 , n11068 );
nand ( n11070 , n11042 , n11069 );
nand ( n11071 , n11041 , n11070 );
and ( n11072 , n11020 , n11071 );
and ( n11073 , n11017 , n11019 );
or ( n11074 , n11072 , n11073 );
not ( n11075 , n11074 );
xor ( n11076 , n10979 , n11075 );
xor ( n11077 , n461 , n530 );
not ( n11078 , n11077 );
not ( n11079 , n10376 );
or ( n11080 , n11078 , n11079 );
nand ( n11081 , n10367 , n10750 );
nand ( n11082 , n11080 , n11081 );
xor ( n11083 , n532 , n459 );
not ( n11084 , n11083 );
not ( n11085 , n10216 );
or ( n11086 , n11084 , n11085 );
nand ( n11087 , n10223 , n10757 );
nand ( n11088 , n11086 , n11087 );
xor ( n11089 , n11082 , n11088 );
and ( n11090 , n526 , n465 );
not ( n11091 , n526 );
and ( n11092 , n11091 , n10626 );
nor ( n11093 , n11090 , n11092 );
not ( n11094 , n11093 );
not ( n11095 , n10476 );
or ( n11096 , n11094 , n11095 );
nand ( n11097 , n10274 , n10746 );
nand ( n11098 , n11096 , n11097 );
not ( n11099 , n11098 );
xor ( n11100 , n11089 , n11099 );
not ( n11101 , n10932 );
not ( n11102 , n10831 );
or ( n11103 , n11101 , n11102 );
nand ( n11104 , n10686 , n10829 );
nand ( n11105 , n11103 , n11104 );
not ( n11106 , n11105 );
not ( n11107 , n11106 );
nand ( n11108 , n536 , n457 );
not ( n11109 , n10923 );
not ( n11110 , n10920 );
or ( n11111 , n11109 , n11110 );
nand ( n11112 , n471 , n472 );
nand ( n11113 , n11111 , n11112 );
and ( n11114 , n11108 , n11113 );
not ( n11115 , n11108 );
not ( n11116 , n11113 );
and ( n11117 , n11115 , n11116 );
nor ( n11118 , n11114 , n11117 );
not ( n11119 , n11118 );
and ( n11120 , n11107 , n11119 );
and ( n11121 , n11106 , n11118 );
nor ( n11122 , n11120 , n11121 );
not ( n11123 , n11122 );
not ( n11124 , n10196 );
not ( n11125 , n10841 );
and ( n11126 , n11124 , n11125 );
and ( n11127 , n10416 , n10948 );
nor ( n11128 , n11126 , n11127 );
not ( n11129 , n11128 );
not ( n11130 , n11129 );
nand ( n11131 , n10957 , n10270 );
not ( n11132 , n11131 );
not ( n11133 , n10268 );
and ( n11134 , n11132 , n11133 );
and ( n11135 , n11093 , n10479 );
nor ( n11136 , n11134 , n11135 );
not ( n11137 , n11136 );
not ( n11138 , n11137 );
or ( n11139 , n11130 , n11138 );
nand ( n11140 , n11136 , n11128 );
nand ( n11141 , n11139 , n11140 );
not ( n11142 , n10890 );
not ( n11143 , n10603 );
or ( n11144 , n11142 , n11143 );
nand ( n11145 , n10241 , n10822 );
nand ( n11146 , n11144 , n11145 );
buf ( n11147 , n11146 );
not ( n11148 , n11147 );
and ( n11149 , n11141 , n11148 );
not ( n11150 , n11141 );
and ( n11151 , n11150 , n11147 );
nor ( n11152 , n11149 , n11151 );
not ( n11153 , n11152 );
or ( n11154 , n11123 , n11153 );
not ( n11155 , n11152 );
not ( n11156 , n11155 );
not ( n11157 , n11122 );
not ( n11158 , n11157 );
or ( n11159 , n11156 , n11158 );
and ( n11160 , n460 , n461 );
not ( n11161 , n460 );
not ( n11162 , n461 );
and ( n11163 , n11161 , n11162 );
nor ( n11164 , n11160 , n11163 );
not ( n11165 , n11164 );
and ( n11166 , n459 , n460 );
not ( n11167 , n459 );
and ( n11168 , n11167 , n10211 );
nor ( n11169 , n11166 , n11168 );
nand ( n11170 , n11165 , n10984 , n11169 );
nand ( n11171 , n3352 , n460 );
not ( n11172 , n11171 );
nand ( n11173 , n10211 , n461 );
not ( n11174 , n11173 );
or ( n11175 , n11172 , n11174 );
nand ( n11176 , n11175 , n11083 );
nand ( n11177 , n11170 , n11176 );
not ( n11178 , n10817 );
not ( n11179 , n10884 );
or ( n11180 , n11178 , n11179 );
nand ( n11181 , n10596 , n10814 );
nand ( n11182 , n11180 , n11181 );
xor ( n11183 , n11177 , n11182 );
not ( n11184 , n11077 );
not ( n11185 , n10471 );
or ( n11186 , n11184 , n11185 );
nand ( n11187 , n10469 , n10463 , n10879 );
nand ( n11188 , n11186 , n11187 );
xor ( n11189 , n11183 , n11188 );
nand ( n11190 , n11159 , n11189 );
nand ( n11191 , n11154 , n11190 );
xor ( n11192 , n11100 , n11191 );
not ( n11193 , n11146 );
not ( n11194 , n11140 );
or ( n11195 , n11193 , n11194 );
nand ( n11196 , n11137 , n11129 );
nand ( n11197 , n11195 , n11196 );
not ( n11198 , n11197 );
not ( n11199 , n11198 );
xor ( n11200 , n11177 , n11182 );
and ( n11201 , n11200 , n11188 );
and ( n11202 , n11177 , n11182 );
or ( n11203 , n11201 , n11202 );
not ( n11204 , n11203 );
not ( n11205 , n11204 );
or ( n11206 , n11199 , n11205 );
nand ( n11207 , n11203 , n11197 );
nand ( n11208 , n11206 , n11207 );
not ( n11209 , n11108 );
not ( n11210 , n11116 );
or ( n11211 , n11209 , n11210 );
nand ( n11212 , n11211 , n11105 );
not ( n11213 , n11108 );
nand ( n11214 , n11213 , n11113 );
nand ( n11215 , n11212 , n11214 );
not ( n11216 , n11215 );
and ( n11217 , n11208 , n11216 );
not ( n11218 , n11208 );
and ( n11219 , n11218 , n11215 );
nor ( n11220 , n11217 , n11219 );
xnor ( n11221 , n11192 , n11220 );
xor ( n11222 , n11076 , n11221 );
xor ( n11223 , n11189 , n11157 );
xor ( n11224 , n11223 , n11155 );
xor ( n11225 , n461 , n533 );
not ( n11226 , n11225 );
nor ( n11227 , n10462 , n10468 );
not ( n11228 , n11227 );
or ( n11229 , n11226 , n11228 );
not ( n11230 , n10365 );
not ( n11231 , n10366 );
or ( n11232 , n11230 , n11231 );
nand ( n11233 , n11232 , n10871 );
nand ( n11234 , n11229 , n11233 );
not ( n11235 , n10980 );
not ( n11236 , n10222 );
or ( n11237 , n11235 , n11236 );
and ( n11238 , n459 , n535 );
not ( n11239 , n459 );
and ( n11240 , n11239 , n10943 );
nor ( n11241 , n11238 , n11240 );
nand ( n11242 , n10214 , n11241 );
nand ( n11243 , n11237 , n11242 );
or ( n11244 , n11234 , n11243 );
xor ( n11245 , n523 , n471 );
nand ( n11246 , n11245 , n472 );
not ( n11247 , n11246 );
nand ( n11248 , n10681 , n524 );
not ( n11249 , n11248 );
not ( n11250 , n524 );
nand ( n11251 , n11250 , n471 );
not ( n11252 , n11251 );
or ( n11253 , n11249 , n11252 );
nor ( n11254 , n10681 , n472 );
nand ( n11255 , n11253 , n11254 );
not ( n11256 , n11255 );
or ( n11257 , n11247 , n11256 );
and ( n11258 , n536 , n460 );
nor ( n11259 , n11258 , n2624 );
or ( n11260 , n536 , n460 );
nand ( n11261 , n11260 , n461 );
nand ( n11262 , n11259 , n11261 );
not ( n11263 , n11262 );
nand ( n11264 , n11257 , n11263 );
not ( n11265 , n11264 );
nand ( n11266 , n11244 , n11265 );
nand ( n11267 , n11234 , n11243 );
nand ( n11268 , n11266 , n11267 );
not ( n11269 , n11268 );
xor ( n11270 , n10986 , n10987 );
xor ( n11271 , n11270 , n11014 );
buf ( n11272 , n11271 );
not ( n11273 , n11272 );
or ( n11274 , n11269 , n11273 );
or ( n11275 , n11271 , n11268 );
nor ( n11276 , n10283 , n11064 );
not ( n11277 , n11276 );
xor ( n11278 , n467 , n528 );
not ( n11279 , n11278 );
not ( n11280 , n10286 );
or ( n11281 , n11279 , n11280 );
nand ( n11282 , n11281 , n10283 );
nand ( n11283 , n11277 , n11282 );
not ( n11284 , n10471 );
not ( n11285 , n11225 );
or ( n11286 , n11284 , n11285 );
not ( n11287 , n10373 );
xor ( n11288 , n461 , n534 );
nand ( n11289 , n11287 , n10306 , n11288 );
nand ( n11290 , n11286 , n11289 );
not ( n11291 , n11290 );
nand ( n11292 , n11283 , n11291 );
not ( n11293 , n11292 );
xor ( n11294 , n536 , n459 );
not ( n11295 , n11294 );
not ( n11296 , n10216 );
or ( n11297 , n11295 , n11296 );
nand ( n11298 , n10223 , n11241 );
nand ( n11299 , n11297 , n11298 );
not ( n11300 , n11299 );
or ( n11301 , n11293 , n11300 );
not ( n11302 , n11283 );
nand ( n11303 , n11302 , n11290 );
nand ( n11304 , n11301 , n11303 );
not ( n11305 , n11304 );
not ( n11306 , n11305 );
not ( n11307 , n11006 );
not ( n11308 , n11008 );
and ( n11309 , n11307 , n11308 );
and ( n11310 , n11006 , n11008 );
nor ( n11311 , n11309 , n11310 );
not ( n11312 , n11311 );
not ( n11313 , n11312 );
not ( n11314 , n10994 );
or ( n11315 , n11313 , n11314 );
not ( n11316 , n10994 );
nand ( n11317 , n11316 , n11311 );
nand ( n11318 , n11315 , n11317 );
not ( n11319 , n11318 );
or ( n11320 , n11306 , n11319 );
xor ( n11321 , n530 , n465 );
not ( n11322 , n11321 );
not ( n11323 , n10476 );
or ( n11324 , n11322 , n11323 );
nand ( n11325 , n10480 , n11049 );
nand ( n11326 , n11324 , n11325 );
and ( n11327 , n532 , n463 );
not ( n11328 , n532 );
and ( n11329 , n11328 , n2650 );
nor ( n11330 , n11327 , n11329 );
not ( n11331 , n11330 );
not ( n11332 , n10237 );
or ( n11333 , n11331 , n11332 );
nand ( n11334 , n10241 , n11043 );
nand ( n11335 , n11333 , n11334 );
xor ( n11336 , n11326 , n11335 );
xor ( n11337 , n526 , n469 );
not ( n11338 , n11337 );
not ( n11339 , n10831 );
or ( n11340 , n11338 , n11339 );
nand ( n11341 , n10928 , n10989 );
nand ( n11342 , n11340 , n11341 );
and ( n11343 , n11336 , n11342 );
and ( n11344 , n11326 , n11335 );
or ( n11345 , n11343 , n11344 );
nand ( n11346 , n11320 , n11345 );
not ( n11347 , n11318 );
nand ( n11348 , n11347 , n11304 );
nand ( n11349 , n11346 , n11348 );
nand ( n11350 , n11275 , n11349 );
nand ( n11351 , n11274 , n11350 );
xor ( n11352 , n11224 , n11351 );
xor ( n11353 , n11017 , n11019 );
xor ( n11354 , n11353 , n11071 );
and ( n11355 , n11352 , n11354 );
and ( n11356 , n11224 , n11351 );
or ( n11357 , n11355 , n11356 );
not ( n11358 , n11357 );
nand ( n11359 , n11222 , n11358 );
xor ( n11360 , n11304 , n11318 );
xor ( n11361 , n11360 , n11345 );
not ( n11362 , n11361 );
not ( n11363 , n11362 );
xor ( n11364 , n529 , n467 );
not ( n11365 , n11364 );
not ( n11366 , n10289 );
or ( n11367 , n11365 , n11366 );
nand ( n11368 , n11060 , n11278 );
nand ( n11369 , n11367 , n11368 );
not ( n11370 , n11369 );
nand ( n11371 , n536 , n462 );
or ( n11372 , n536 , n462 );
nand ( n11373 , n11372 , n463 );
nand ( n11374 , n11371 , n461 , n11373 );
not ( n11375 , n11374 );
xor ( n11376 , n528 , n469 );
not ( n11377 , n11376 );
not ( n11378 , n10831 );
or ( n11379 , n11377 , n11378 );
xor ( n11380 , n527 , n469 );
nand ( n11381 , n10686 , n11380 );
nand ( n11382 , n11379 , n11381 );
nand ( n11383 , n11375 , n11382 );
nand ( n11384 , n11370 , n11383 );
not ( n11385 , n11384 );
not ( n11386 , n10920 );
xor ( n11387 , n471 , n526 );
not ( n11388 , n11387 );
or ( n11389 , n11386 , n11388 );
and ( n11390 , n471 , n525 );
not ( n11391 , n471 );
not ( n11392 , n525 );
and ( n11393 , n11391 , n11392 );
nor ( n11394 , n11390 , n11393 );
nand ( n11395 , n11394 , n472 );
nand ( n11396 , n11389 , n11395 );
xor ( n11397 , n532 , n465 );
not ( n11398 , n11397 );
not ( n11399 , n10271 );
or ( n11400 , n11398 , n11399 );
and ( n11401 , n465 , n531 );
not ( n11402 , n465 );
and ( n11403 , n11402 , n10877 );
nor ( n11404 , n11401 , n11403 );
nand ( n11405 , n10274 , n11404 );
nand ( n11406 , n11400 , n11405 );
xor ( n11407 , n11396 , n11406 );
xor ( n11408 , n534 , n463 );
not ( n11409 , n11408 );
not ( n11410 , n10237 );
or ( n11411 , n11409 , n11410 );
xor ( n11412 , n533 , n463 );
nand ( n11413 , n10241 , n11412 );
nand ( n11414 , n11411 , n11413 );
and ( n11415 , n11407 , n11414 );
and ( n11416 , n11396 , n11406 );
or ( n11417 , n11415 , n11416 );
not ( n11418 , n11417 );
or ( n11419 , n11385 , n11418 );
not ( n11420 , n11383 );
nand ( n11421 , n11420 , n11369 );
nand ( n11422 , n11419 , n11421 );
not ( n11423 , n11422 );
xor ( n11424 , n11326 , n11335 );
xor ( n11425 , n11424 , n11342 );
not ( n11426 , n11425 );
xor ( n11427 , n11290 , n11283 );
xor ( n11428 , n11427 , n11299 );
nand ( n11429 , n11426 , n11428 );
not ( n11430 , n11429 );
or ( n11431 , n11423 , n11430 );
not ( n11432 , n11428 );
nand ( n11433 , n11432 , n11425 );
nand ( n11434 , n11431 , n11433 );
not ( n11435 , n11434 );
nand ( n11436 , n11363 , n11435 );
not ( n11437 , n11436 );
xor ( n11438 , n11264 , n11234 );
xnor ( n11439 , n11438 , n11243 );
xor ( n11440 , n11048 , n11057 );
xor ( n11441 , n11440 , n11066 );
xor ( n11442 , n11439 , n11441 );
buf ( n11443 , n11262 );
not ( n11444 , n11443 );
nand ( n11445 , n11255 , n11246 );
not ( n11446 , n11445 );
or ( n11447 , n11444 , n11446 );
or ( n11448 , n11445 , n11443 );
nand ( n11449 , n11447 , n11448 );
not ( n11450 , n11394 );
not ( n11451 , n11002 );
or ( n11452 , n11450 , n11451 );
not ( n11453 , n11248 );
not ( n11454 , n11251 );
or ( n11455 , n11453 , n11454 );
nand ( n11456 , n11455 , n472 );
nand ( n11457 , n11452 , n11456 );
not ( n11458 , n11457 );
nand ( n11459 , n11412 , n10900 , n10235 );
nand ( n11460 , n11330 , n10892 );
nand ( n11461 , n11459 , n11460 );
not ( n11462 , n11461 );
or ( n11463 , n11458 , n11462 );
not ( n11464 , n11457 );
nand ( n11465 , n11459 , n11460 , n11464 );
xor ( n11466 , n535 , n461 );
not ( n11467 , n11466 );
not ( n11468 , n10376 );
or ( n11469 , n11467 , n11468 );
nand ( n11470 , n10471 , n11288 );
nand ( n11471 , n11469 , n11470 );
nand ( n11472 , n11465 , n11471 );
nand ( n11473 , n11463 , n11472 );
xor ( n11474 , n11449 , n11473 );
not ( n11475 , n11321 );
not ( n11476 , n11052 );
or ( n11477 , n11475 , n11476 );
not ( n11478 , n10479 );
nand ( n11479 , n10270 , n11478 , n11404 );
nand ( n11480 , n11477 , n11479 );
not ( n11481 , n11480 );
nand ( n11482 , n11164 , n536 );
not ( n11483 , n11482 );
not ( n11484 , n11483 );
or ( n11485 , n11481 , n11484 );
or ( n11486 , n11480 , n11483 );
not ( n11487 , n11380 );
not ( n11488 , n10831 );
or ( n11489 , n11487 , n11488 );
nand ( n11490 , n10686 , n11337 );
nand ( n11491 , n11489 , n11490 );
nand ( n11492 , n11486 , n11491 );
nand ( n11493 , n11485 , n11492 );
and ( n11494 , n11474 , n11493 );
and ( n11495 , n11449 , n11473 );
or ( n11496 , n11494 , n11495 );
xor ( n11497 , n11442 , n11496 );
not ( n11498 , n11497 );
or ( n11499 , n11437 , n11498 );
nand ( n11500 , n11434 , n11362 );
nand ( n11501 , n11499 , n11500 );
xor ( n11502 , n11439 , n11441 );
and ( n11503 , n11502 , n11496 );
and ( n11504 , n11439 , n11441 );
or ( n11505 , n11503 , n11504 );
and ( n11506 , n11069 , n11023 );
not ( n11507 , n11069 );
and ( n11508 , n11507 , n11024 );
nor ( n11509 , n11506 , n11508 );
not ( n11510 , n11039 );
and ( n11511 , n11509 , n11510 );
not ( n11512 , n11509 );
and ( n11513 , n11512 , n11039 );
nor ( n11514 , n11511 , n11513 );
xor ( n11515 , n11505 , n11514 );
not ( n11516 , n11271 );
xor ( n11517 , n11268 , n11516 );
xnor ( n11518 , n11517 , n11349 );
xor ( n11519 , n11515 , n11518 );
nor ( n11520 , n11501 , n11519 );
not ( n11521 , n11520 );
xor ( n11522 , n11224 , n11351 );
xor ( n11523 , n11522 , n11354 );
not ( n11524 , n11523 );
xor ( n11525 , n11505 , n11514 );
and ( n11526 , n11525 , n11518 );
and ( n11527 , n11505 , n11514 );
or ( n11528 , n11526 , n11527 );
not ( n11529 , n11528 );
nand ( n11530 , n11524 , n11529 );
and ( n11531 , n11359 , n11521 , n11530 );
not ( n11532 , n11531 );
xor ( n11533 , n532 , n467 );
not ( n11534 , n11533 );
not ( n11535 , n10288 );
or ( n11536 , n11534 , n11535 );
xor ( n11537 , n531 , n467 );
nand ( n11538 , n11060 , n11537 );
nand ( n11539 , n11536 , n11538 );
not ( n11540 , n11539 );
not ( n11541 , n11540 );
xor ( n11542 , n530 , n469 );
not ( n11543 , n11542 );
not ( n11544 , n10615 );
or ( n11545 , n11543 , n11544 );
xor ( n11546 , n529 , n469 );
nand ( n11547 , n10686 , n11546 );
nand ( n11548 , n11545 , n11547 );
or ( n11549 , n536 , n464 );
nand ( n11550 , n11549 , n465 );
nand ( n11551 , n536 , n464 );
and ( n11552 , n11550 , n11551 , n463 );
nor ( n11553 , n11548 , n11552 );
not ( n11554 , n11553 );
nand ( n11555 , n11552 , n11548 );
nand ( n11556 , n11554 , n11555 );
not ( n11557 , n11556 );
or ( n11558 , n11541 , n11557 );
and ( n11559 , n10240 , n536 );
not ( n11560 , n472 );
xor ( n11561 , n471 , n528 );
not ( n11562 , n11561 );
or ( n11563 , n11560 , n11562 );
and ( n11564 , n471 , n529 );
not ( n11565 , n471 );
not ( n11566 , n529 );
and ( n11567 , n11565 , n11566 );
nor ( n11568 , n11564 , n11567 );
not ( n11569 , n471 );
nor ( n11570 , n11569 , n472 );
nand ( n11571 , n11568 , n11570 );
nand ( n11572 , n11563 , n11571 );
xor ( n11573 , n11559 , n11572 );
xor ( n11574 , n535 , n465 );
not ( n11575 , n11574 );
not ( n11576 , n10476 );
or ( n11577 , n11575 , n11576 );
xor ( n11578 , n534 , n465 );
nand ( n11579 , n11578 , n10274 );
nand ( n11580 , n11577 , n11579 );
and ( n11581 , n11573 , n11580 );
and ( n11582 , n11559 , n11572 );
or ( n11583 , n11581 , n11582 );
nand ( n11584 , n11558 , n11583 );
not ( n11585 , n11556 );
nand ( n11586 , n11585 , n11539 );
nand ( n11587 , n11584 , n11586 );
not ( n11588 , n11587 );
xor ( n11589 , n471 , n527 );
not ( n11590 , n11589 );
not ( n11591 , n10920 );
or ( n11592 , n11590 , n11591 );
nand ( n11593 , n11387 , n472 );
nand ( n11594 , n11592 , n11593 );
xor ( n11595 , n535 , n463 );
not ( n11596 , n11595 );
not ( n11597 , n10237 );
or ( n11598 , n11596 , n11597 );
nand ( n11599 , n10241 , n11408 );
nand ( n11600 , n11598 , n11599 );
xor ( n11601 , n11594 , n11600 );
not ( n11602 , n11537 );
not ( n11603 , n10288 );
or ( n11604 , n11602 , n11603 );
xor ( n11605 , n467 , n530 );
nand ( n11606 , n10596 , n11605 );
nand ( n11607 , n11604 , n11606 );
buf ( n11608 , n11607 );
xor ( n11609 , n11601 , n11608 );
not ( n11610 , n11609 );
or ( n11611 , n11588 , n11610 );
not ( n11612 , n11587 );
not ( n11613 , n11609 );
nand ( n11614 , n11612 , n11613 );
nand ( n11615 , n11611 , n11614 );
not ( n11616 , n11615 );
not ( n11617 , n11561 );
not ( n11618 , n11570 );
or ( n11619 , n11617 , n11618 );
nand ( n11620 , n11589 , n472 );
nand ( n11621 , n11619 , n11620 );
not ( n11622 , n11621 );
not ( n11623 , n11578 );
not ( n11624 , n10476 );
or ( n11625 , n11623 , n11624 );
xor ( n11626 , n533 , n465 );
nand ( n11627 , n10480 , n11626 );
nand ( n11628 , n11625 , n11627 );
not ( n11629 , n11628 );
or ( n11630 , n11622 , n11629 );
or ( n11631 , n11628 , n11621 );
xor ( n11632 , n536 , n463 );
not ( n11633 , n11632 );
not ( n11634 , n10237 );
or ( n11635 , n11633 , n11634 );
nand ( n11636 , n10241 , n11595 );
nand ( n11637 , n11635 , n11636 );
nand ( n11638 , n11631 , n11637 );
nand ( n11639 , n11630 , n11638 );
xor ( n11640 , n11555 , n11639 );
and ( n11641 , n10471 , n536 );
not ( n11642 , n11626 );
not ( n11643 , n11053 );
or ( n11644 , n11642 , n11643 );
nand ( n11645 , n11052 , n11397 );
nand ( n11646 , n11644 , n11645 );
not ( n11647 , n11646 );
xor ( n11648 , n11641 , n11647 );
not ( n11649 , n10831 );
not ( n11650 , n11546 );
or ( n11651 , n11649 , n11650 );
nand ( n11652 , n10686 , n11376 );
nand ( n11653 , n11651 , n11652 );
xnor ( n11654 , n11648 , n11653 );
xnor ( n11655 , n11640 , n11654 );
not ( n11656 , n11655 );
not ( n11657 , n11656 );
or ( n11658 , n11616 , n11657 );
or ( n11659 , n11615 , n11656 );
nand ( n11660 , n11658 , n11659 );
not ( n11661 , n11660 );
buf ( n11662 , n11556 );
xor ( n11663 , n11540 , n11662 );
xnor ( n11664 , n11663 , n11583 );
or ( n11665 , n536 , n466 );
nand ( n11666 , n11665 , n467 );
nand ( n11667 , n536 , n466 );
and ( n11668 , n11666 , n11667 , n465 );
nor ( n11669 , n530 , n472 );
nand ( n11670 , n11669 , n471 );
not ( n11671 , n471 );
nand ( n11672 , n11671 , n472 , n529 );
nand ( n11673 , n11566 , n471 , n472 );
nand ( n11674 , n11670 , n11672 , n11673 );
nand ( n11675 , n11668 , n11674 );
xor ( n11676 , n531 , n469 );
not ( n11677 , n11676 );
not ( n11678 , n10615 );
or ( n11679 , n11677 , n11678 );
nand ( n11680 , n11542 , n10686 );
nand ( n11681 , n11679 , n11680 );
not ( n11682 , n11681 );
xor ( n11683 , n11675 , n11682 );
xor ( n11684 , n533 , n467 );
not ( n11685 , n11684 );
not ( n11686 , n10288 );
or ( n11687 , n11685 , n11686 );
nand ( n11688 , n10452 , n11533 );
nand ( n11689 , n11687 , n11688 );
not ( n11690 , n11689 );
and ( n11691 , n11683 , n11690 );
and ( n11692 , n11675 , n11682 );
or ( n11693 , n11691 , n11692 );
xor ( n11694 , n11621 , n11637 );
xnor ( n11695 , n11694 , n11628 );
and ( n11696 , n11693 , n11695 );
or ( n11697 , n11664 , n11696 );
or ( n11698 , n11695 , n11693 );
nand ( n11699 , n11697 , n11698 );
nand ( n11700 , n11661 , n11699 );
not ( n11701 , n11700 );
xor ( n11702 , n11559 , n11572 );
xor ( n11703 , n11702 , n11580 );
not ( n11704 , n11703 );
xor ( n11705 , n11675 , n11682 );
xor ( n11706 , n11705 , n11690 );
or ( n11707 , n11704 , n11706 );
not ( n11708 , n11706 );
not ( n11709 , n11704 );
or ( n11710 , n11708 , n11709 );
xor ( n11711 , n536 , n465 );
not ( n11712 , n11711 );
not ( n11713 , n10271 );
or ( n11714 , n11712 , n11713 );
nand ( n11715 , n10274 , n11574 );
nand ( n11716 , n11714 , n11715 );
xor ( n11717 , n534 , n467 );
not ( n11718 , n11717 );
not ( n11719 , n10289 );
or ( n11720 , n11718 , n11719 );
nand ( n11721 , n11060 , n11684 );
nand ( n11722 , n11720 , n11721 );
xor ( n11723 , n11716 , n11722 );
xor ( n11724 , n532 , n469 );
not ( n11725 , n11724 );
not ( n11726 , n10831 );
or ( n11727 , n11725 , n11726 );
nand ( n11728 , n10686 , n11676 );
nand ( n11729 , n11727 , n11728 );
and ( n11730 , n11723 , n11729 );
and ( n11731 , n11716 , n11722 );
or ( n11732 , n11730 , n11731 );
nand ( n11733 , n11710 , n11732 );
nand ( n11734 , n11707 , n11733 );
not ( n11735 , n11734 );
xor ( n11736 , n11539 , n11583 );
xnor ( n11737 , n11736 , n11662 );
xor ( n11738 , n11693 , n11695 );
xnor ( n11739 , n11737 , n11738 );
nand ( n11740 , n11735 , n11739 );
not ( n11741 , n11704 );
not ( n11742 , n11706 );
not ( n11743 , n11742 );
or ( n11744 , n11741 , n11743 );
nand ( n11745 , n11706 , n11703 );
nand ( n11746 , n11744 , n11745 );
not ( n11747 , n11746 );
not ( n11748 , n11732 );
nand ( n11749 , n11747 , n11748 );
not ( n11750 , n11748 );
nand ( n11751 , n11750 , n11746 );
nand ( n11752 , n10480 , n536 );
not ( n11753 , n11752 );
not ( n11754 , n11753 );
xor ( n11755 , n531 , n471 );
not ( n11756 , n11755 );
not ( n11757 , n10920 );
or ( n11758 , n11756 , n11757 );
xor ( n11759 , n471 , n530 );
nand ( n11760 , n11759 , n472 );
nand ( n11761 , n11758 , n11760 );
not ( n11762 , n11761 );
or ( n11763 , n11754 , n11762 );
not ( n11764 , n11752 );
not ( n11765 , n11761 );
not ( n11766 , n11765 );
or ( n11767 , n11764 , n11766 );
xor ( n11768 , n533 , n469 );
not ( n11769 , n11768 );
not ( n11770 , n10831 );
or ( n11771 , n11769 , n11770 );
nand ( n11772 , n10686 , n11724 );
nand ( n11773 , n11771 , n11772 );
nand ( n11774 , n11767 , n11773 );
nand ( n11775 , n11763 , n11774 );
not ( n11776 , n11775 );
not ( n11777 , n11674 );
not ( n11778 , n11777 );
not ( n11779 , n11668 );
not ( n11780 , n11779 );
or ( n11781 , n11778 , n11780 );
nand ( n11782 , n11781 , n11675 );
nand ( n11783 , n11776 , n11782 );
not ( n11784 , n11783 );
xor ( n11785 , n11716 , n11722 );
xor ( n11786 , n11785 , n11729 );
not ( n11787 , n11786 );
or ( n11788 , n11784 , n11787 );
not ( n11789 , n11782 );
nand ( n11790 , n11789 , n11775 );
nand ( n11791 , n11788 , n11790 );
and ( n11792 , n11749 , n11751 , n11791 );
nand ( n11793 , n11740 , n11792 );
not ( n11794 , n11739 );
nand ( n11795 , n11794 , n11734 );
and ( n11796 , n11793 , n11795 );
xor ( n11797 , n536 , n467 );
nand ( n11798 , n10286 , n11797 );
not ( n11799 , n11798 );
not ( n11800 , n10452 );
and ( n11801 , n11799 , n11800 );
xor ( n11802 , n535 , n467 );
and ( n11803 , n11060 , n11802 );
nor ( n11804 , n11801 , n11803 );
not ( n11805 , n11804 );
xor ( n11806 , n534 , n469 );
not ( n11807 , n11806 );
not ( n11808 , n10831 );
or ( n11809 , n11807 , n11808 );
nand ( n11810 , n10686 , n11768 );
nand ( n11811 , n11809 , n11810 );
and ( n11812 , n11805 , n11811 );
not ( n11813 , n11805 );
not ( n11814 , n11811 );
and ( n11815 , n11813 , n11814 );
nor ( n11816 , n11812 , n11815 );
or ( n11817 , n536 , n468 );
nand ( n11818 , n11817 , n469 );
nand ( n11819 , n536 , n468 );
nand ( n11820 , n11818 , n11819 , n467 );
xor ( n11821 , n471 , n532 );
not ( n11822 , n11821 );
not ( n11823 , n11570 );
or ( n11824 , n11822 , n11823 );
nand ( n11825 , n11755 , n472 );
nand ( n11826 , n11824 , n11825 );
xor ( n11827 , n11820 , n11826 );
and ( n11828 , n11816 , n11827 );
not ( n11829 , n11816 );
not ( n11830 , n11827 );
and ( n11831 , n11829 , n11830 );
nor ( n11832 , n11828 , n11831 );
xor ( n11833 , n535 , n469 );
not ( n11834 , n11833 );
not ( n11835 , n10831 );
or ( n11836 , n11834 , n11835 );
nand ( n11837 , n10686 , n11806 );
nand ( n11838 , n11836 , n11837 );
not ( n11839 , n11838 );
xor ( n11840 , n471 , n533 );
not ( n11841 , n11840 );
not ( n11842 , n10920 );
or ( n11843 , n11841 , n11842 );
nand ( n11844 , n11821 , n472 );
nand ( n11845 , n11843 , n11844 );
not ( n11846 , n11845 );
not ( n11847 , n536 );
not ( n11848 , n11847 );
nand ( n11849 , n11848 , n10452 );
nand ( n11850 , n11846 , n11849 );
not ( n11851 , n11850 );
or ( n11852 , n11839 , n11851 );
not ( n11853 , n11849 );
nand ( n11854 , n11853 , n11845 );
nand ( n11855 , n11852 , n11854 );
not ( n11856 , n11855 );
nand ( n11857 , n11832 , n11856 );
not ( n11858 , n11857 );
not ( n11859 , n11570 );
xor ( n11860 , n534 , n471 );
not ( n11861 , n11860 );
or ( n11862 , n11859 , n11861 );
nand ( n11863 , n11840 , n472 );
nand ( n11864 , n11862 , n11863 );
not ( n11865 , n11864 );
or ( n11866 , n536 , n470 );
nand ( n11867 , n11866 , n471 );
nand ( n11868 , n536 , n470 );
nand ( n11869 , n11867 , n11868 , n469 );
not ( n11870 , n11869 );
and ( n11871 , n11865 , n11870 );
and ( n11872 , n11864 , n11869 );
nor ( n11873 , n11871 , n11872 );
xor ( n11874 , n536 , n469 );
not ( n11875 , n11874 );
not ( n11876 , n10831 );
or ( n11877 , n11875 , n11876 );
nand ( n11878 , n10686 , n11833 );
nand ( n11879 , n11877 , n11878 );
not ( n11880 , n11879 );
nand ( n11881 , n11873 , n11880 );
not ( n11882 , n11881 );
not ( n11883 , n11847 );
not ( n11884 , n11570 );
or ( n11885 , n11883 , n11884 );
xor ( n11886 , n471 , n535 );
nand ( n11887 , n11886 , n472 );
nand ( n11888 , n11885 , n11887 );
and ( n11889 , n536 , n472 );
nor ( n11890 , n11889 , n10681 );
nand ( n11891 , n11888 , n11890 );
nand ( n11892 , n10686 , n536 );
not ( n11893 , n11892 );
not ( n11894 , n11886 );
not ( n11895 , n10920 );
or ( n11896 , n11894 , n11895 );
nand ( n11897 , n11860 , n472 );
nand ( n11898 , n11896 , n11897 );
nor ( n11899 , n11893 , n11898 );
or ( n11900 , n11891 , n11899 );
not ( n11901 , n11892 );
nand ( n11902 , n11901 , n11898 );
nand ( n11903 , n11900 , n11902 );
not ( n11904 , n11903 );
or ( n11905 , n11882 , n11904 );
not ( n11906 , n11873 );
nand ( n11907 , n11906 , n11879 );
nand ( n11908 , n11905 , n11907 );
not ( n11909 , n11908 );
not ( n11910 , n11845 );
not ( n11911 , n11849 );
and ( n11912 , n11910 , n11911 );
and ( n11913 , n11845 , n11849 );
nor ( n11914 , n11912 , n11913 );
not ( n11915 , n11914 );
not ( n11916 , n11838 );
and ( n11917 , n11915 , n11916 );
and ( n11918 , n11838 , n11914 );
nor ( n11919 , n11917 , n11918 );
not ( n11920 , n11869 );
nand ( n11921 , n11920 , n11864 );
nand ( n11922 , n11919 , n11921 );
not ( n11923 , n11922 );
or ( n11924 , n11909 , n11923 );
not ( n11925 , n11919 );
not ( n11926 , n11921 );
nand ( n11927 , n11925 , n11926 );
nand ( n11928 , n11924 , n11927 );
not ( n11929 , n11928 );
or ( n11930 , n11858 , n11929 );
not ( n11931 , n11832 );
nand ( n11932 , n11931 , n11855 );
nand ( n11933 , n11930 , n11932 );
not ( n11934 , n11827 );
not ( n11935 , n11804 );
or ( n11936 , n11934 , n11935 );
nand ( n11937 , n11936 , n11811 );
nand ( n11938 , n11830 , n11805 );
nand ( n11939 , n11937 , n11938 );
not ( n11940 , n11939 );
not ( n11941 , n11761 );
not ( n11942 , n11752 );
or ( n11943 , n11941 , n11942 );
or ( n11944 , n11761 , n11752 );
nand ( n11945 , n11943 , n11944 );
xor ( n11946 , n11945 , n11773 );
not ( n11947 , n11946 );
not ( n11948 , n11826 );
nor ( n11949 , n11948 , n11820 );
not ( n11950 , n11949 );
not ( n11951 , n11802 );
not ( n11952 , n10288 );
or ( n11953 , n11951 , n11952 );
nand ( n11954 , n11060 , n11717 );
nand ( n11955 , n11953 , n11954 );
not ( n11956 , n11955 );
not ( n11957 , n11956 );
and ( n11958 , n11950 , n11957 );
and ( n11959 , n11949 , n11956 );
nor ( n11960 , n11958 , n11959 );
not ( n11961 , n11960 );
and ( n11962 , n11947 , n11961 );
and ( n11963 , n11946 , n11960 );
nor ( n11964 , n11962 , n11963 );
nand ( n11965 , n11940 , n11964 );
nand ( n11966 , n11933 , n11965 );
xor ( n11967 , n11782 , n11775 );
xnor ( n11968 , n11967 , n11786 );
or ( n11969 , n11949 , n11955 );
nand ( n11970 , n11969 , n11946 );
nand ( n11971 , n11949 , n11955 );
nand ( n11972 , n11970 , n11971 );
nand ( n11973 , n11968 , n11972 );
not ( n11974 , n11964 );
nand ( n11975 , n11974 , n11939 );
nand ( n11976 , n11966 , n11973 , n11975 );
nand ( n11977 , n11747 , n11748 );
and ( n11978 , n11977 , n11751 );
nor ( n11979 , n11978 , n11791 );
nor ( n11980 , n11968 , n11972 );
nor ( n11981 , n11979 , n11980 );
nand ( n11982 , n11740 , n11976 , n11981 );
nand ( n11983 , n11796 , n11982 );
not ( n11984 , n11699 );
nand ( n11985 , n11984 , n11660 );
nand ( n11986 , n11983 , n11985 );
not ( n11987 , n11986 );
or ( n11988 , n11701 , n11987 );
not ( n11989 , n11383 );
not ( n11990 , n11369 );
and ( n11991 , n11989 , n11990 );
and ( n11992 , n11383 , n11369 );
nor ( n11993 , n11991 , n11992 );
not ( n11994 , n11993 );
not ( n11995 , n11417 );
and ( n11996 , n11994 , n11995 );
and ( n11997 , n11417 , n11993 );
nor ( n11998 , n11996 , n11997 );
not ( n11999 , n11998 );
xor ( n12000 , n11457 , n11471 );
xor ( n12001 , n12000 , n11461 );
not ( n12002 , n12001 );
xor ( n12003 , n11483 , n11480 );
xnor ( n12004 , n12003 , n11491 );
nand ( n12005 , n12002 , n12004 );
not ( n12006 , n12005 );
not ( n12007 , n11364 );
not ( n12008 , n11060 );
or ( n12009 , n12007 , n12008 );
nand ( n12010 , n11605 , n10286 , n10722 );
nand ( n12011 , n12009 , n12010 );
buf ( n12012 , n12011 );
not ( n12013 , n12012 );
not ( n12014 , n10313 );
xnor ( n12015 , n536 , n461 );
not ( n12016 , n12015 );
and ( n12017 , n12014 , n12016 );
and ( n12018 , n10317 , n11466 );
nor ( n12019 , n12017 , n12018 );
nand ( n12020 , n12013 , n12019 );
not ( n12021 , n11374 );
not ( n12022 , n12021 );
not ( n12023 , n11382 );
not ( n12024 , n12023 );
or ( n12025 , n12022 , n12024 );
nand ( n12026 , n11382 , n11374 );
nand ( n12027 , n12025 , n12026 );
and ( n12028 , n12020 , n12027 );
not ( n12029 , n12019 );
and ( n12030 , n12029 , n12012 );
nor ( n12031 , n12028 , n12030 );
not ( n12032 , n12001 );
nor ( n12033 , n12032 , n12004 );
nor ( n12034 , n12031 , n12033 );
not ( n12035 , n12034 );
or ( n12036 , n12006 , n12035 );
not ( n12037 , n12004 );
nor ( n12038 , n12037 , n12001 );
or ( n12039 , n12038 , n12033 );
nand ( n12040 , n12039 , n12031 );
nand ( n12041 , n12036 , n12040 );
not ( n12042 , n12041 );
or ( n12043 , n11999 , n12042 );
not ( n12044 , n11594 );
not ( n12045 , n11600 );
or ( n12046 , n12044 , n12045 );
or ( n12047 , n11594 , n11600 );
nand ( n12048 , n12047 , n11607 );
nand ( n12049 , n12046 , n12048 );
not ( n12050 , n12049 );
xor ( n12051 , n11396 , n11406 );
xor ( n12052 , n12051 , n11414 );
not ( n12053 , n12052 );
or ( n12054 , n12050 , n12053 );
or ( n12055 , n12049 , n12052 );
not ( n12056 , n11641 );
not ( n12057 , n11646 );
or ( n12058 , n12056 , n12057 );
not ( n12059 , n11647 );
not ( n12060 , n11641 );
not ( n12061 , n12060 );
or ( n12062 , n12059 , n12061 );
nand ( n12063 , n12062 , n11653 );
nand ( n12064 , n12058 , n12063 );
nand ( n12065 , n12055 , n12064 );
nand ( n12066 , n12054 , n12065 );
nand ( n12067 , n12043 , n12066 );
not ( n12068 , n11998 );
not ( n12069 , n12041 );
nand ( n12070 , n12068 , n12069 );
nand ( n12071 , n12067 , n12070 );
not ( n12072 , n12071 );
xor ( n12073 , n11449 , n11473 );
xor ( n12074 , n12073 , n11493 );
not ( n12075 , n12074 );
not ( n12076 , n12001 );
not ( n12077 , n12037 );
or ( n12078 , n12076 , n12077 );
not ( n12079 , n12032 );
not ( n12080 , n12004 );
or ( n12081 , n12079 , n12080 );
not ( n12082 , n12031 );
nand ( n12083 , n12081 , n12082 );
nand ( n12084 , n12078 , n12083 );
xor ( n12085 , n12075 , n12084 );
and ( n12086 , n11425 , n11428 );
not ( n12087 , n11425 );
and ( n12088 , n12087 , n11432 );
nor ( n12089 , n12086 , n12088 );
and ( n12090 , n12089 , n11422 );
not ( n12091 , n12089 );
not ( n12092 , n11422 );
and ( n12093 , n12091 , n12092 );
nor ( n12094 , n12090 , n12093 );
xnor ( n12095 , n12085 , n12094 );
nand ( n12096 , n12072 , n12095 );
or ( n12097 , n11998 , n12066 );
nand ( n12098 , n12066 , n11998 );
nand ( n12099 , n12097 , n12098 );
xnor ( n12100 , n12099 , n12069 );
not ( n12101 , n11654 );
not ( n12102 , n11555 );
not ( n12103 , n12102 );
or ( n12104 , n12101 , n12103 );
or ( n12105 , n11654 , n12102 );
nand ( n12106 , n12105 , n11639 );
nand ( n12107 , n12104 , n12106 );
not ( n12108 , n12107 );
not ( n12109 , n12108 );
not ( n12110 , n12052 );
xor ( n12111 , n12049 , n12064 );
xor ( n12112 , n12110 , n12111 );
not ( n12113 , n12112 );
or ( n12114 , n12109 , n12113 );
xor ( n12115 , n12012 , n12029 );
xnor ( n12116 , n12115 , n12027 );
not ( n12117 , n12116 );
nand ( n12118 , n12114 , n12117 );
not ( n12119 , n12112 );
nand ( n12120 , n12119 , n12107 );
nand ( n12121 , n12118 , n12120 );
not ( n12122 , n12121 );
nand ( n12123 , n12100 , n12122 );
nor ( n12124 , n12107 , n12117 );
and ( n12125 , n12124 , n12112 );
nor ( n12126 , n12107 , n12116 );
not ( n12127 , n12112 );
and ( n12128 , n12126 , n12127 );
nor ( n12129 , n12125 , n12128 );
not ( n12130 , n12129 );
and ( n12131 , n12116 , n12112 );
not ( n12132 , n12116 );
and ( n12133 , n12132 , n12127 );
nor ( n12134 , n12131 , n12133 );
not ( n12135 , n12108 );
nand ( n12136 , n12134 , n12135 );
not ( n12137 , n12136 );
or ( n12138 , n12130 , n12137 );
not ( n12139 , n11655 );
nand ( n12140 , n11612 , n11613 );
not ( n12141 , n12140 );
or ( n12142 , n12139 , n12141 );
not ( n12143 , n11612 );
nand ( n12144 , n12143 , n11609 );
nand ( n12145 , n12142 , n12144 );
not ( n12146 , n12145 );
nand ( n12147 , n12138 , n12146 );
nand ( n12148 , n12096 , n12123 , n12147 );
not ( n12149 , n12094 );
not ( n12150 , n12149 );
not ( n12151 , n12075 );
not ( n12152 , n12151 );
or ( n12153 , n12150 , n12152 );
not ( n12154 , n12075 );
not ( n12155 , n12094 );
or ( n12156 , n12154 , n12155 );
buf ( n12157 , n12084 );
nand ( n12158 , n12156 , n12157 );
nand ( n12159 , n12153 , n12158 );
not ( n12160 , n12159 );
and ( n12161 , n11497 , n11362 );
not ( n12162 , n11497 );
and ( n12163 , n12162 , n11361 );
nor ( n12164 , n12161 , n12163 );
and ( n12165 , n12164 , n11435 );
not ( n12166 , n12164 );
and ( n12167 , n12166 , n11434 );
nor ( n12168 , n12165 , n12167 );
nand ( n12169 , n12160 , n12168 );
not ( n12170 , n12169 );
nor ( n12171 , n12148 , n12170 );
nand ( n12172 , n11988 , n12171 );
buf ( n12173 , n12096 );
nand ( n12174 , n12136 , n12129 );
nor ( n12175 , n12174 , n12146 );
not ( n12176 , n12175 );
not ( n12177 , n12123 );
or ( n12178 , n12176 , n12177 );
not ( n12179 , n12100 );
nand ( n12180 , n12179 , n12121 );
nand ( n12181 , n12178 , n12180 );
not ( n12182 , n12170 );
nand ( n12183 , n12173 , n12181 , n12182 );
not ( n12184 , n12169 );
nor ( n12185 , n12072 , n12095 );
not ( n12186 , n12185 );
or ( n12187 , n12184 , n12186 );
not ( n12188 , n12168 );
nand ( n12189 , n12188 , n12159 );
nand ( n12190 , n12187 , n12189 );
not ( n12191 , n12190 );
nand ( n12192 , n12172 , n12183 , n12191 );
not ( n12193 , n12192 );
or ( n12194 , n11532 , n12193 );
not ( n12195 , n11529 );
not ( n12196 , n11524 );
or ( n12197 , n12195 , n12196 );
nand ( n12198 , n11523 , n11528 );
nand ( n12199 , n11519 , n11501 );
nand ( n12200 , n12198 , n12199 );
nand ( n12201 , n12197 , n12200 );
not ( n12202 , n11359 );
or ( n12203 , n12201 , n12202 );
not ( n12204 , n11222 );
nand ( n12205 , n12204 , n11357 );
nand ( n12206 , n12203 , n12205 );
not ( n12207 , n12206 );
nand ( n12208 , n12194 , n12207 );
not ( n12209 , n12208 );
xor ( n12210 , n10742 , n10765 );
xor ( n12211 , n12210 , n10768 );
or ( n12212 , n10681 , n10850 );
nand ( n12213 , n12212 , n10848 );
nand ( n12214 , n10681 , n10850 );
nand ( n12215 , n12213 , n12214 );
xor ( n12216 , n10749 , n10755 );
xor ( n12217 , n12216 , n10762 );
xor ( n12218 , n12215 , n12217 );
xor ( n12219 , n10821 , n10827 );
and ( n12220 , n12219 , n10835 );
and ( n12221 , n10821 , n10827 );
or ( n12222 , n12220 , n12221 );
and ( n12223 , n12218 , n12222 );
and ( n12224 , n12215 , n12217 );
or ( n12225 , n12223 , n12224 );
xor ( n12226 , n12211 , n12225 );
or ( n12227 , n11203 , n11197 );
nand ( n12228 , n12227 , n11215 );
nand ( n12229 , n11203 , n11197 );
nand ( n12230 , n12228 , n12229 );
not ( n12231 , n12230 );
not ( n12232 , n10846 );
not ( n12233 , n10255 );
or ( n12234 , n12232 , n12233 );
nand ( n12235 , n10195 , n10661 );
nand ( n12236 , n12234 , n12235 );
not ( n12237 , n12236 );
not ( n12238 , n12237 );
not ( n12239 , n10688 );
not ( n12240 , n12239 );
or ( n12241 , n12238 , n12240 );
nand ( n12242 , n10688 , n12236 );
nand ( n12243 , n12241 , n12242 );
and ( n12244 , n12243 , n11099 );
not ( n12245 , n12243 );
and ( n12246 , n12245 , n11098 );
nor ( n12247 , n12244 , n12246 );
not ( n12248 , n10720 );
not ( n12249 , n10736 );
nand ( n12250 , n12249 , n10741 );
not ( n12251 , n12250 );
not ( n12252 , n12251 );
or ( n12253 , n12248 , n12252 );
not ( n12254 , n10720 );
nand ( n12255 , n12254 , n12250 );
nand ( n12256 , n12253 , n12255 );
nand ( n12257 , n12247 , n12256 );
not ( n12258 , n12257 );
or ( n12259 , n12231 , n12258 );
not ( n12260 , n12256 );
not ( n12261 , n12247 );
nand ( n12262 , n12260 , n12261 );
nand ( n12263 , n12259 , n12262 );
xor ( n12264 , n12226 , n12263 );
not ( n12265 , n12264 );
not ( n12266 , n10641 );
not ( n12267 , n10633 );
not ( n12268 , n10634 );
and ( n12269 , n12267 , n12268 );
and ( n12270 , n10633 , n10634 );
nor ( n12271 , n12269 , n12270 );
xor ( n12272 , n12266 , n12271 );
not ( n12273 , n12272 );
xor ( n12274 , n12239 , n10673 );
xnor ( n12275 , n12274 , n10666 );
not ( n12276 , n12275 );
xor ( n12277 , n12273 , n12276 );
not ( n12278 , n12237 );
not ( n12279 , n11099 );
or ( n12280 , n12278 , n12279 );
nand ( n12281 , n12280 , n12239 );
nand ( n12282 , n11098 , n12236 );
nand ( n12283 , n12281 , n12282 );
xor ( n12284 , n12277 , n12283 );
not ( n12285 , n12284 );
or ( n12286 , n12265 , n12285 );
not ( n12287 , n12264 );
not ( n12288 , n12275 );
not ( n12289 , n12283 );
not ( n12290 , n12272 );
or ( n12291 , n12289 , n12290 );
or ( n12292 , n12283 , n12272 );
nand ( n12293 , n12291 , n12292 );
not ( n12294 , n12293 );
not ( n12295 , n12294 );
or ( n12296 , n12288 , n12295 );
not ( n12297 , n12275 );
nand ( n12298 , n12297 , n12293 );
nand ( n12299 , n12296 , n12298 );
nand ( n12300 , n12287 , n12299 );
nand ( n12301 , n12286 , n12300 );
xor ( n12302 , n11082 , n11088 );
and ( n12303 , n12302 , n11099 );
and ( n12304 , n11082 , n11088 );
or ( n12305 , n12303 , n12304 );
not ( n12306 , n12305 );
xor ( n12307 , n12215 , n12217 );
xor ( n12308 , n12307 , n12222 );
not ( n12309 , n12308 );
or ( n12310 , n12306 , n12309 );
or ( n12311 , n12305 , n12308 );
not ( n12312 , n10868 );
not ( n12313 , n10978 );
or ( n12314 , n12312 , n12313 );
nand ( n12315 , n12314 , n10869 );
nand ( n12316 , n12311 , n12315 );
nand ( n12317 , n12310 , n12316 );
not ( n12318 , n12317 );
and ( n12319 , n12301 , n12318 );
not ( n12320 , n12301 );
and ( n12321 , n12320 , n12317 );
nor ( n12322 , n12319 , n12321 );
buf ( n12323 , n12230 );
and ( n12324 , n12261 , n12256 );
not ( n12325 , n12261 );
and ( n12326 , n12325 , n12260 );
nor ( n12327 , n12324 , n12326 );
xor ( n12328 , n12323 , n12327 );
not ( n12329 , n12328 );
xor ( n12330 , n12305 , n12308 );
xnor ( n12331 , n12330 , n12315 );
not ( n12332 , n12331 );
or ( n12333 , n12329 , n12332 );
not ( n12334 , n11100 );
not ( n12335 , n11220 );
or ( n12336 , n12334 , n12335 );
or ( n12337 , n11220 , n11100 );
nand ( n12338 , n12337 , n11191 );
nand ( n12339 , n12336 , n12338 );
nand ( n12340 , n12333 , n12339 );
not ( n12341 , n12331 );
not ( n12342 , n12328 );
nand ( n12343 , n12341 , n12342 );
nand ( n12344 , n12340 , n12343 );
not ( n12345 , n12344 );
nand ( n12346 , n12322 , n12345 );
and ( n12347 , n12339 , n12328 );
not ( n12348 , n12339 );
and ( n12349 , n12348 , n12342 );
nor ( n12350 , n12347 , n12349 );
and ( n12351 , n12350 , n12341 );
not ( n12352 , n12350 );
not ( n12353 , n12341 );
and ( n12354 , n12352 , n12353 );
nor ( n12355 , n12351 , n12354 );
xor ( n12356 , n10979 , n11075 );
and ( n12357 , n12356 , n11221 );
and ( n12358 , n10979 , n11075 );
or ( n12359 , n12357 , n12358 );
nand ( n12360 , n12355 , n12359 );
and ( n12361 , n12346 , n12360 );
not ( n12362 , n12361 );
not ( n12363 , n12272 );
not ( n12364 , n12276 );
or ( n12365 , n12363 , n12364 );
nand ( n12366 , n12365 , n12283 );
nand ( n12367 , n12275 , n12273 );
nand ( n12368 , n12366 , n12367 );
not ( n12369 , n12368 );
not ( n12370 , n12369 );
xor ( n12371 , n10771 , n10773 );
xor ( n12372 , n12371 , n10776 );
nand ( n12373 , n12370 , n12372 );
or ( n12374 , n12372 , n12368 );
xor ( n12375 , n12211 , n12225 );
and ( n12376 , n12375 , n12263 );
and ( n12377 , n12211 , n12225 );
or ( n12378 , n12376 , n12377 );
nand ( n12379 , n12374 , n12378 );
nand ( n12380 , n12373 , n12379 );
not ( n12381 , n12380 );
not ( n12382 , n12381 );
xor ( n12383 , n10708 , n10779 );
xor ( n12384 , n12383 , n10698 );
not ( n12385 , n12384 );
or ( n12386 , n12382 , n12385 );
not ( n12387 , n12378 );
not ( n12388 , n12369 );
not ( n12389 , n12372 );
or ( n12390 , n12388 , n12389 );
or ( n12391 , n12372 , n12369 );
nand ( n12392 , n12390 , n12391 );
xor ( n12393 , n12387 , n12392 );
not ( n12394 , n12299 );
not ( n12395 , n12287 );
not ( n12396 , n12395 );
or ( n12397 , n12394 , n12396 );
not ( n12398 , n12284 );
not ( n12399 , n12287 );
or ( n12400 , n12398 , n12399 );
nand ( n12401 , n12400 , n12317 );
nand ( n12402 , n12397 , n12401 );
not ( n12403 , n12402 );
nand ( n12404 , n12393 , n12403 );
nand ( n12405 , n12386 , n12404 );
nor ( n12406 , n12362 , n12405 );
not ( n12407 , n12406 );
or ( n12408 , n12209 , n12407 );
not ( n12409 , n12405 );
not ( n12410 , n12409 );
nor ( n12411 , n12355 , n12359 );
not ( n12412 , n12411 );
not ( n12413 , n12346 );
or ( n12414 , n12412 , n12413 );
not ( n12415 , n12322 );
nand ( n12416 , n12415 , n12344 );
nand ( n12417 , n12414 , n12416 );
not ( n12418 , n12417 );
not ( n12419 , n12418 );
not ( n12420 , n12419 );
or ( n12421 , n12410 , n12420 );
not ( n12422 , n12384 );
nand ( n12423 , n12422 , n12380 );
not ( n12424 , n12402 );
nor ( n12425 , n12424 , n12393 );
nand ( n12426 , n12381 , n12384 );
nand ( n12427 , n12425 , n12426 );
nand ( n12428 , n12423 , n12427 );
not ( n12429 , n12428 );
nand ( n12430 , n12421 , n12429 );
not ( n12431 , n12430 );
nand ( n12432 , n12408 , n12431 );
not ( n12433 , n12432 );
or ( n12434 , n10813 , n12433 );
not ( n12435 , n10590 );
nand ( n12436 , n10799 , n10781 );
or ( n12437 , n10808 , n12436 );
nand ( n12438 , n10805 , n10807 );
nand ( n12439 , n12437 , n12438 );
not ( n12440 , n12439 );
or ( n12441 , n12435 , n12440 );
not ( n12442 , n10510 );
nor ( n12443 , n12442 , n10589 );
not ( n12444 , n12443 );
nand ( n12445 , n12441 , n12444 );
not ( n12446 , n12445 );
nand ( n12447 , n12434 , n12446 );
not ( n12448 , n12447 );
not ( n12449 , n10551 );
nand ( n12450 , n12449 , n10558 );
not ( n12451 , n12450 );
not ( n12452 , n10574 );
or ( n12453 , n12451 , n12452 );
not ( n12454 , n10558 );
nand ( n12455 , n12454 , n10551 );
nand ( n12456 , n12453 , n12455 );
not ( n12457 , n12456 );
xor ( n12458 , n10531 , n10537 );
and ( n12459 , n12458 , n10543 );
and ( n12460 , n10531 , n10537 );
or ( n12461 , n12459 , n12460 );
and ( n12462 , n457 , n527 );
not ( n12463 , n10558 );
xor ( n12464 , n12462 , n12463 );
not ( n12465 , n10549 );
not ( n12466 , n10216 );
or ( n12467 , n12465 , n12466 );
xor ( n12468 , n523 , n459 );
nand ( n12469 , n10223 , n12468 );
nand ( n12470 , n12467 , n12469 );
xnor ( n12471 , n12464 , n12470 );
xor ( n12472 , n12461 , n12471 );
not ( n12473 , n10535 );
not ( n12474 , n10256 );
or ( n12475 , n12473 , n12474 );
xor ( n12476 , n457 , n525 );
nand ( n12477 , n10197 , n12476 );
nand ( n12478 , n12475 , n12477 );
not ( n12479 , n10556 );
not ( n12480 , n10314 );
or ( n12481 , n12479 , n12480 );
xor ( n12482 , n461 , n521 );
nand ( n12483 , n10317 , n12482 );
nand ( n12484 , n12481 , n12483 );
xor ( n12485 , n12478 , n12484 );
or ( n12486 , n10603 , n10241 );
nand ( n12487 , n12486 , n463 );
xor ( n12488 , n12485 , n12487 );
xor ( n12489 , n12472 , n12488 );
xor ( n12490 , n12457 , n12489 );
xor ( n12491 , n10530 , n10544 );
and ( n12492 , n12491 , n10578 );
and ( n12493 , n10530 , n10544 );
or ( n12494 , n12492 , n12493 );
xor ( n12495 , n12490 , n12494 );
not ( n12496 , n12495 );
nand ( n12497 , n10582 , n10525 );
not ( n12498 , n12497 );
not ( n12499 , n10518 );
or ( n12500 , n12498 , n12499 );
nand ( n12501 , n10579 , n10524 );
nand ( n12502 , n12500 , n12501 );
nand ( n12503 , n12496 , n12502 );
not ( n12504 , n12502 );
nand ( n12505 , n12504 , n12495 );
nand ( n12506 , n12503 , n12505 );
not ( n12507 , n12506 );
and ( n12508 , n12448 , n12507 );
and ( n12509 , n12447 , n12506 );
nor ( n12510 , n12508 , n12509 );
not ( n12511 , n12510 );
not ( n12512 , n12511 );
not ( n12513 , n12512 );
or ( n12514 , n10192 , n12513 );
not ( n12515 , n12512 );
not ( n12516 , n503 );
nand ( n12517 , n12515 , n12516 );
nand ( n12518 , n12514 , n12517 );
not ( n12519 , n12518 );
or ( n12520 , n10191 , n12519 );
not ( n12521 , n503 );
nor ( n12522 , n10811 , n12405 );
not ( n12523 , n12522 );
not ( n12524 , n12206 );
not ( n12525 , n12361 );
or ( n12526 , n12524 , n12525 );
nand ( n12527 , n12526 , n12418 );
not ( n12528 , n12527 );
not ( n12529 , n12202 );
and ( n12530 , n11521 , n11530 );
and ( n12531 , n12529 , n12530 , n12346 , n12360 );
nand ( n12532 , n12531 , n12192 );
nand ( n12533 , n12528 , n12532 );
not ( n12534 , n12533 );
or ( n12535 , n12523 , n12534 );
and ( n12536 , n10810 , n12428 );
nor ( n12537 , n12536 , n12439 );
nand ( n12538 , n12535 , n12537 );
not ( n12539 , n12443 );
nand ( n12540 , n12539 , n10590 );
not ( n12541 , n12540 );
and ( n12542 , n12538 , n12541 );
not ( n12543 , n12538 );
and ( n12544 , n12543 , n12540 );
nor ( n12545 , n12542 , n12544 );
not ( n12546 , n12545 );
not ( n12547 , n12546 );
or ( n12548 , n12521 , n12547 );
not ( n12549 , n12546 );
buf ( n12550 , n12516 );
nand ( n12551 , n12549 , n12550 );
nand ( n12552 , n12548 , n12551 );
not ( n12553 , n504 );
nand ( n12554 , n12553 , n503 );
not ( n12555 , n12554 );
nand ( n12556 , n12552 , n12555 );
nand ( n12557 , n12520 , n12556 );
and ( n12558 , n498 , n499 );
not ( n12559 , n498 );
not ( n12560 , n499 );
and ( n12561 , n12559 , n12560 );
or ( n12562 , n12558 , n12561 );
not ( n12563 , n12562 );
not ( n12564 , n12563 );
not ( n12565 , n497 );
or ( n12566 , n12359 , n12355 );
nand ( n12567 , n12360 , n12566 );
not ( n12568 , n12567 );
not ( n12569 , n12208 );
or ( n12570 , n12568 , n12569 );
not ( n12571 , n12208 );
not ( n12572 , n12567 );
nand ( n12573 , n12571 , n12572 );
nand ( n12574 , n12570 , n12573 );
not ( n12575 , n12574 );
buf ( n12576 , n12575 );
not ( n12577 , n12576 );
or ( n12578 , n12565 , n12577 );
not ( n12579 , n497 );
nand ( n12580 , n12574 , n12579 );
nand ( n12581 , n12578 , n12580 );
not ( n12582 , n12581 );
or ( n12583 , n12564 , n12582 );
not ( n12584 , n497 );
nand ( n12585 , n12529 , n12205 );
not ( n12586 , n12585 );
not ( n12587 , n12586 );
not ( n12588 , n12530 );
nand ( n12589 , n12191 , n12172 , n12183 );
not ( n12590 , n12589 );
or ( n12591 , n12588 , n12590 );
buf ( n12592 , n12201 );
nand ( n12593 , n12591 , n12592 );
not ( n12594 , n12593 );
not ( n12595 , n12594 );
or ( n12596 , n12587 , n12595 );
nand ( n12597 , n12593 , n12585 );
nand ( n12598 , n12596 , n12597 );
not ( n12599 , n12598 );
not ( n12600 , n12599 );
or ( n12601 , n12584 , n12600 );
buf ( n12602 , n12598 );
nand ( n12603 , n12602 , n12579 );
nand ( n12604 , n12601 , n12603 );
and ( n12605 , n498 , n497 );
not ( n12606 , n498 );
and ( n12607 , n12606 , n12579 );
nor ( n12608 , n12605 , n12607 );
and ( n12609 , n12562 , n12608 );
buf ( n12610 , n12609 );
nand ( n12611 , n12604 , n12610 );
nand ( n12612 , n12583 , n12611 );
not ( n12613 , n489 );
buf ( n12614 , n11979 );
not ( n12615 , n12614 );
buf ( n12616 , n11792 );
not ( n12617 , n12616 );
nand ( n12618 , n12615 , n12617 );
or ( n12619 , n11968 , n11972 );
not ( n12620 , n12619 );
not ( n12621 , n12620 );
buf ( n12622 , n11976 );
nand ( n12623 , n12621 , n12622 );
xor ( n12624 , n12618 , n12623 );
not ( n12625 , n12624 );
nor ( n12626 , n12613 , n12625 );
not ( n12627 , n12626 );
and ( n12628 , n490 , n491 );
not ( n12629 , n490 );
and ( n12630 , n12629 , n1993 );
nor ( n12631 , n12628 , n12630 );
not ( n12632 , n12631 );
xor ( n12633 , n489 , n490 );
nand ( n12634 , n12632 , n12633 );
not ( n12635 , n12634 );
not ( n12636 , n12635 );
not ( n12637 , n489 );
nand ( n12638 , n11795 , n11740 );
not ( n12639 , n12638 );
nor ( n12640 , n12614 , n12620 );
and ( n12641 , n12622 , n12640 );
nor ( n12642 , n12641 , n12616 );
not ( n12643 , n12642 );
not ( n12644 , n12643 );
or ( n12645 , n12639 , n12644 );
not ( n12646 , n12638 );
nand ( n12647 , n12646 , n12642 );
nand ( n12648 , n12645 , n12647 );
not ( n12649 , n12648 );
not ( n12650 , n12649 );
or ( n12651 , n12637 , n12650 );
buf ( n12652 , n12648 );
not ( n12653 , n489 );
nand ( n12654 , n12652 , n12653 );
nand ( n12655 , n12651 , n12654 );
not ( n12656 , n12655 );
or ( n12657 , n12636 , n12656 );
not ( n12658 , n11983 );
not ( n12659 , n12658 );
nand ( n12660 , n11700 , n11985 );
not ( n12661 , n12660 );
not ( n12662 , n12661 );
or ( n12663 , n12659 , n12662 );
nand ( n12664 , n12660 , n11983 );
nand ( n12665 , n12663 , n12664 );
buf ( n12666 , n12665 );
not ( n12667 , n12666 );
not ( n12668 , n12653 );
or ( n12669 , n12667 , n12668 );
not ( n12670 , n12665 );
nand ( n12671 , n12670 , n489 );
nand ( n12672 , n12669 , n12671 );
buf ( n12673 , n12631 );
nand ( n12674 , n12672 , n12673 );
nand ( n12675 , n12657 , n12674 );
not ( n12676 , n12675 );
or ( n12677 , n12627 , n12676 );
or ( n12678 , n12675 , n12626 );
nand ( n12679 , n12677 , n12678 );
and ( n12680 , n491 , n492 );
nor ( n12681 , n491 , n492 );
nor ( n12682 , n12680 , n12681 );
and ( n12683 , n492 , n493 );
not ( n12684 , n492 );
and ( n12685 , n12684 , n2264 );
or ( n12686 , n12683 , n12685 );
nand ( n12687 , n12682 , n12686 );
not ( n12688 , n12687 );
not ( n12689 , n12688 );
not ( n12690 , n491 );
not ( n12691 , n11985 );
not ( n12692 , n11983 );
or ( n12693 , n12691 , n12692 );
nand ( n12694 , n12693 , n11700 );
not ( n12695 , n12175 );
nand ( n12696 , n12146 , n12174 );
nand ( n12697 , n12695 , n12696 );
xnor ( n12698 , n12694 , n12697 );
buf ( n12699 , n12698 );
not ( n12700 , n12699 );
not ( n12701 , n12700 );
or ( n12702 , n12690 , n12701 );
not ( n12703 , n491 );
nand ( n12704 , n12699 , n12703 );
nand ( n12705 , n12702 , n12704 );
not ( n12706 , n12705 );
or ( n12707 , n12689 , n12706 );
not ( n12708 , n491 );
and ( n12709 , n12123 , n12180 );
not ( n12710 , n12709 );
not ( n12711 , n12696 );
nand ( n12712 , n11986 , n11700 );
not ( n12713 , n12712 );
or ( n12714 , n12711 , n12713 );
nand ( n12715 , n12714 , n12695 );
not ( n12716 , n12715 );
not ( n12717 , n12716 );
or ( n12718 , n12710 , n12717 );
not ( n12719 , n12709 );
nand ( n12720 , n12719 , n12715 );
nand ( n12721 , n12718 , n12720 );
not ( n12722 , n12721 );
not ( n12723 , n12722 );
or ( n12724 , n12708 , n12723 );
and ( n12725 , n12709 , n12716 );
not ( n12726 , n12709 );
and ( n12727 , n12726 , n12715 );
or ( n12728 , n12725 , n12727 );
nand ( n12729 , n12703 , n12728 );
nand ( n12730 , n12724 , n12729 );
not ( n12731 , n12686 );
nand ( n12732 , n12730 , n12731 );
nand ( n12733 , n12707 , n12732 );
and ( n12734 , n12679 , n12733 );
not ( n12735 , n12679 );
not ( n12736 , n12733 );
and ( n12737 , n12735 , n12736 );
or ( n12738 , n12734 , n12737 );
xor ( n12739 , n12612 , n12738 );
xor ( n12740 , n500 , n501 );
buf ( n12741 , n12740 );
not ( n12742 , n12741 );
not ( n12743 , n12742 );
not ( n12744 , n12743 );
not ( n12745 , n499 );
not ( n12746 , n12425 );
nand ( n12747 , n12393 , n12403 );
nand ( n12748 , n12746 , n12747 );
not ( n12749 , n12748 );
not ( n12750 , n12749 );
not ( n12751 , n12192 );
not ( n12752 , n12531 );
or ( n12753 , n12751 , n12752 );
not ( n12754 , n12527 );
nand ( n12755 , n12753 , n12754 );
not ( n12756 , n12755 );
not ( n12757 , n12756 );
or ( n12758 , n12750 , n12757 );
nand ( n12759 , n12755 , n12748 );
nand ( n12760 , n12758 , n12759 );
not ( n12761 , n12760 );
not ( n12762 , n12761 );
or ( n12763 , n12745 , n12762 );
not ( n12764 , n12761 );
nand ( n12765 , n12764 , n12560 );
nand ( n12766 , n12763 , n12765 );
not ( n12767 , n12766 );
or ( n12768 , n12744 , n12767 );
nand ( n12769 , n12416 , n12346 );
not ( n12770 , n12769 );
not ( n12771 , n12770 );
not ( n12772 , n12360 );
not ( n12773 , n12208 );
or ( n12774 , n12772 , n12773 );
nand ( n12775 , n12774 , n12566 );
not ( n12776 , n12775 );
not ( n12777 , n12776 );
or ( n12778 , n12771 , n12777 );
nand ( n12779 , n12775 , n12769 );
nand ( n12780 , n12778 , n12779 );
not ( n12781 , n12780 );
and ( n12782 , n12781 , n499 );
not ( n12783 , n12781 );
and ( n12784 , n12783 , n12560 );
or ( n12785 , n12782 , n12784 );
not ( n12786 , n12740 );
xor ( n12787 , n500 , n499 );
nand ( n12788 , n12786 , n12787 );
not ( n12789 , n12788 );
nand ( n12790 , n12785 , n12789 );
nand ( n12791 , n12768 , n12790 );
and ( n12792 , n12739 , n12791 );
and ( n12793 , n12612 , n12738 );
or ( n12794 , n12792 , n12793 );
xor ( n12795 , n12557 , n12794 );
not ( n12796 , n12673 );
and ( n12797 , n12625 , n489 );
not ( n12798 , n12625 );
and ( n12799 , n12798 , n12653 );
or ( n12800 , n12797 , n12799 );
not ( n12801 , n12800 );
or ( n12802 , n12796 , n12801 );
nand ( n12803 , n11966 , n11975 );
not ( n12804 , n12803 );
not ( n12805 , n12804 );
nand ( n12806 , n11973 , n12619 );
not ( n12807 , n12806 );
not ( n12808 , n12807 );
or ( n12809 , n12805 , n12808 );
nand ( n12810 , n12806 , n12803 );
nand ( n12811 , n12809 , n12810 );
buf ( n12812 , n12811 );
xor ( n12813 , n489 , n12812 );
nand ( n12814 , n12635 , n12813 );
nand ( n12815 , n12802 , n12814 );
not ( n12816 , n11939 );
not ( n12817 , n12816 );
not ( n12818 , n11964 );
or ( n12819 , n12817 , n12818 );
nand ( n12820 , n12819 , n11975 );
not ( n12821 , n11933 );
xor ( n12822 , n12820 , n12821 );
and ( n12823 , n489 , n12822 );
xor ( n12824 , n12815 , n12823 );
not ( n12825 , n12731 );
not ( n12826 , n491 );
not ( n12827 , n12670 );
or ( n12828 , n12826 , n12827 );
nand ( n12829 , n12666 , n12703 );
nand ( n12830 , n12828 , n12829 );
not ( n12831 , n12830 );
or ( n12832 , n12825 , n12831 );
not ( n12833 , n491 );
not ( n12834 , n12649 );
or ( n12835 , n12833 , n12834 );
nand ( n12836 , n12652 , n12703 );
nand ( n12837 , n12835 , n12836 );
nand ( n12838 , n12837 , n12688 );
nand ( n12839 , n12832 , n12838 );
and ( n12840 , n12824 , n12839 );
and ( n12841 , n12815 , n12823 );
or ( n12842 , n12840 , n12841 );
xor ( n12843 , n494 , n495 );
not ( n12844 , n12843 );
not ( n12845 , n12844 );
not ( n12846 , n12845 );
and ( n12847 , n12123 , n12147 );
not ( n12848 , n12847 );
not ( n12849 , n12712 );
or ( n12850 , n12848 , n12849 );
not ( n12851 , n12181 );
nand ( n12852 , n12850 , n12851 );
buf ( n12853 , n12852 );
not ( n12854 , n12185 );
nand ( n12855 , n12854 , n12173 );
not ( n12856 , n12855 );
and ( n12857 , n12853 , n12856 );
not ( n12858 , n12853 );
and ( n12859 , n12858 , n12855 );
nor ( n12860 , n12857 , n12859 );
buf ( n12861 , n12860 );
not ( n12862 , n493 );
and ( n12863 , n12861 , n12862 );
not ( n12864 , n12861 );
and ( n12865 , n12864 , n493 );
or ( n12866 , n12863 , n12865 );
not ( n12867 , n12866 );
or ( n12868 , n12846 , n12867 );
not ( n12869 , n493 );
buf ( n12870 , n12722 );
not ( n12871 , n12870 );
or ( n12872 , n12869 , n12871 );
nand ( n12873 , n12862 , n12728 );
nand ( n12874 , n12872 , n12873 );
and ( n12875 , n493 , n494 );
nor ( n12876 , n493 , n494 );
nor ( n12877 , n12875 , n12876 );
and ( n12878 , n12844 , n12877 );
nand ( n12879 , n12874 , n12878 );
nand ( n12880 , n12868 , n12879 );
xor ( n12881 , n12842 , n12880 );
buf ( n12882 , n12631 );
not ( n12883 , n12882 );
not ( n12884 , n12655 );
or ( n12885 , n12883 , n12884 );
nand ( n12886 , n12800 , n12635 );
nand ( n12887 , n12885 , n12886 );
and ( n12888 , n489 , n12812 );
xor ( n12889 , n12887 , n12888 );
not ( n12890 , n12731 );
not ( n12891 , n12705 );
or ( n12892 , n12890 , n12891 );
nand ( n12893 , n12830 , n12688 );
nand ( n12894 , n12892 , n12893 );
xor ( n12895 , n12889 , n12894 );
and ( n12896 , n12881 , n12895 );
and ( n12897 , n12842 , n12880 );
or ( n12898 , n12896 , n12897 );
not ( n12899 , n502 );
nand ( n12900 , n12899 , n501 );
not ( n12901 , n501 );
nand ( n12902 , n12901 , n502 );
and ( n12903 , n12900 , n12902 );
and ( n12904 , n502 , n3291 );
not ( n12905 , n502 );
and ( n12906 , n12905 , n503 );
or ( n12907 , n12904 , n12906 );
nor ( n12908 , n12903 , n12907 );
buf ( n12909 , n12908 );
not ( n12910 , n12909 );
nand ( n12911 , n12426 , n12423 );
not ( n12912 , n12911 );
not ( n12913 , n12747 );
not ( n12914 , n12533 );
or ( n12915 , n12913 , n12914 );
nand ( n12916 , n12915 , n12746 );
not ( n12917 , n12916 );
or ( n12918 , n12912 , n12917 );
not ( n12919 , n12911 );
nand ( n12920 , n12533 , n12747 );
nand ( n12921 , n12919 , n12920 , n12746 );
nand ( n12922 , n12918 , n12921 );
not ( n12923 , n12922 );
and ( n12924 , n755 , n12923 );
not ( n12925 , n755 );
and ( n12926 , n12925 , n12922 );
nor ( n12927 , n12924 , n12926 );
not ( n12928 , n12927 );
or ( n12929 , n12910 , n12928 );
buf ( n12930 , n12907 );
not ( n12931 , n501 );
or ( n12932 , n10799 , n10781 );
nand ( n12933 , n12436 , n12932 );
not ( n12934 , n12933 );
not ( n12935 , n12432 );
or ( n12936 , n12934 , n12935 );
or ( n12937 , n12933 , n12432 );
nand ( n12938 , n12936 , n12937 );
not ( n12939 , n12938 );
not ( n12940 , n12939 );
or ( n12941 , n12931 , n12940 );
not ( n12942 , n12939 );
not ( n12943 , n501 );
nand ( n12944 , n12942 , n12943 );
nand ( n12945 , n12941 , n12944 );
nand ( n12946 , n12930 , n12945 );
nand ( n12947 , n12929 , n12946 );
xor ( n12948 , n12898 , n12947 );
not ( n12949 , n12555 );
not ( n12950 , n10808 );
nand ( n12951 , n12950 , n12438 );
not ( n12952 , n12951 );
not ( n12953 , n12532 );
not ( n12954 , n12207 );
nand ( n12955 , n12954 , n12361 );
not ( n12956 , n12955 );
or ( n12957 , n12953 , n12956 );
and ( n12958 , n12409 , n12932 );
nand ( n12959 , n12957 , n12958 );
and ( n12960 , n12428 , n12932 );
not ( n12961 , n12436 );
nor ( n12962 , n12960 , n12961 );
nand ( n12963 , n12419 , n12932 );
not ( n12964 , n12963 );
nand ( n12965 , n12964 , n12409 );
nand ( n12966 , n12959 , n12962 , n12965 );
not ( n12967 , n12966 );
or ( n12968 , n12952 , n12967 );
not ( n12969 , n12960 );
nor ( n12970 , n12951 , n12961 );
nand ( n12971 , n12969 , n12959 , n12965 , n12970 );
nand ( n12972 , n12968 , n12971 );
not ( n12973 , n12972 );
not ( n12974 , n12973 );
or ( n12975 , n12949 , n12974 );
nand ( n12976 , n12552 , n504 );
nand ( n12977 , n12975 , n12976 );
and ( n12978 , n12948 , n12977 );
and ( n12979 , n12898 , n12947 );
or ( n12980 , n12978 , n12979 );
and ( n12981 , n12795 , n12980 );
and ( n12982 , n12557 , n12794 );
or ( n12983 , n12981 , n12982 );
and ( n12984 , n12675 , n12626 );
not ( n12985 , n12731 );
not ( n12986 , n491 );
not ( n12987 , n12861 );
not ( n12988 , n12987 );
or ( n12989 , n12986 , n12988 );
nand ( n12990 , n12861 , n12703 );
nand ( n12991 , n12989 , n12990 );
not ( n12992 , n12991 );
or ( n12993 , n12985 , n12992 );
nand ( n12994 , n12730 , n12688 );
nand ( n12995 , n12993 , n12994 );
xor ( n12996 , n12984 , n12995 );
and ( n12997 , n12652 , n489 );
not ( n12998 , n12882 );
not ( n12999 , n489 );
not ( n13000 , n12700 );
or ( n13001 , n12999 , n13000 );
nand ( n13002 , n12699 , n12653 );
nand ( n13003 , n13001 , n13002 );
not ( n13004 , n13003 );
or ( n13005 , n12998 , n13004 );
nand ( n13006 , n12672 , n12635 );
nand ( n13007 , n13005 , n13006 );
xor ( n13008 , n12997 , n13007 );
xor ( n13009 , n12996 , n13008 );
not ( n13010 , n12563 );
not ( n13011 , n497 );
not ( n13012 , n12781 );
or ( n13013 , n13011 , n13012 );
nand ( n13014 , n12780 , n12579 );
nand ( n13015 , n13013 , n13014 );
not ( n13016 , n13015 );
or ( n13017 , n13010 , n13016 );
nand ( n13018 , n12581 , n12610 );
nand ( n13019 , n13017 , n13018 );
xor ( n13020 , n13009 , n13019 );
not ( n13021 , n12878 );
not ( n13022 , n12866 );
or ( n13023 , n13021 , n13022 );
not ( n13024 , n493 );
not ( n13025 , n12173 );
not ( n13026 , n12852 );
or ( n13027 , n13025 , n13026 );
buf ( n13028 , n12854 );
nand ( n13029 , n13027 , n13028 );
nand ( n13030 , n12182 , n12189 );
not ( n13031 , n13030 );
and ( n13032 , n13029 , n13031 );
not ( n13033 , n13029 );
and ( n13034 , n13033 , n13030 );
nor ( n13035 , n13032 , n13034 );
buf ( n13036 , n13035 );
not ( n13037 , n13036 );
not ( n13038 , n13037 );
or ( n13039 , n13024 , n13038 );
nand ( n13040 , n13036 , n12862 );
nand ( n13041 , n13039 , n13040 );
nand ( n13042 , n13041 , n12845 );
nand ( n13043 , n13023 , n13042 );
xor ( n13044 , n12887 , n12888 );
and ( n13045 , n13044 , n12894 );
and ( n13046 , n12887 , n12888 );
or ( n13047 , n13045 , n13046 );
xor ( n13048 , n13043 , n13047 );
and ( n13049 , n496 , n497 );
not ( n13050 , n496 );
and ( n13051 , n13050 , n12579 );
or ( n13052 , n13049 , n13051 );
and ( n13053 , n496 , n495 );
nor ( n13054 , n495 , n496 );
nor ( n13055 , n13053 , n13054 );
and ( n13056 , n13052 , n13055 );
not ( n13057 , n13056 );
not ( n13058 , n495 );
nand ( n13059 , n12199 , n11521 );
not ( n13060 , n13059 );
buf ( n13061 , n12589 );
not ( n13062 , n13061 );
or ( n13063 , n13060 , n13062 );
not ( n13064 , n13061 );
not ( n13065 , n13059 );
nand ( n13066 , n13064 , n13065 );
nand ( n13067 , n13063 , n13066 );
not ( n13068 , n13067 );
not ( n13069 , n13068 );
or ( n13070 , n13058 , n13069 );
not ( n13071 , n495 );
buf ( n13072 , n13067 );
nand ( n13073 , n13071 , n13072 );
nand ( n13074 , n13070 , n13073 );
not ( n13075 , n13074 );
or ( n13076 , n13057 , n13075 );
not ( n13077 , n12852 );
not ( n13078 , n12170 );
nand ( n13079 , n13078 , n12173 );
nor ( n13080 , n13079 , n11520 );
not ( n13081 , n13080 );
or ( n13082 , n13077 , n13081 );
not ( n13083 , n12190 );
not ( n13084 , n11521 );
or ( n13085 , n13083 , n13084 );
nand ( n13086 , n13085 , n12199 );
not ( n13087 , n13086 );
nand ( n13088 , n13082 , n13087 );
nand ( n13089 , n11530 , n12198 );
not ( n13090 , n13089 );
and ( n13091 , n13088 , n13090 );
not ( n13092 , n13088 );
and ( n13093 , n13092 , n13089 );
nor ( n13094 , n13091 , n13093 );
buf ( n13095 , n13094 );
not ( n13096 , n13095 );
and ( n13097 , n495 , n13096 );
not ( n13098 , n495 );
and ( n13099 , n13098 , n13095 );
or ( n13100 , n13097 , n13099 );
not ( n13101 , n13100 );
or ( n13102 , n13101 , n13052 );
nand ( n13103 , n13076 , n13102 );
and ( n13104 , n13048 , n13103 );
and ( n13105 , n13043 , n13047 );
or ( n13106 , n13104 , n13105 );
xor ( n13107 , n13020 , n13106 );
nor ( n13108 , n12679 , n12736 );
not ( n13109 , n12845 );
and ( n13110 , n13072 , n493 );
not ( n13111 , n13072 );
and ( n13112 , n13111 , n2264 );
nor ( n13113 , n13110 , n13112 );
not ( n13114 , n13113 );
or ( n13115 , n13109 , n13114 );
nand ( n13116 , n13041 , n12878 );
nand ( n13117 , n13115 , n13116 );
xor ( n13118 , n13108 , n13117 );
not ( n13119 , n13052 );
not ( n13120 , n13119 );
and ( n13121 , n495 , n12599 );
not ( n13122 , n495 );
and ( n13123 , n13122 , n12598 );
or ( n13124 , n13121 , n13123 );
not ( n13125 , n13124 );
or ( n13126 , n13120 , n13125 );
nand ( n13127 , n13100 , n13056 );
nand ( n13128 , n13126 , n13127 );
xor ( n13129 , n13118 , n13128 );
not ( n13130 , n12930 );
and ( n13131 , n501 , n12973 );
not ( n13132 , n501 );
not ( n13133 , n12973 );
and ( n13134 , n13132 , n13133 );
or ( n13135 , n13131 , n13134 );
not ( n13136 , n13135 );
or ( n13137 , n13130 , n13136 );
nand ( n13138 , n12945 , n12908 );
nand ( n13139 , n13137 , n13138 );
xor ( n13140 , n13129 , n13139 );
not ( n13141 , n12743 );
and ( n13142 , n12922 , n12560 );
not ( n13143 , n12922 );
and ( n13144 , n13143 , n499 );
or ( n13145 , n13142 , n13144 );
not ( n13146 , n13145 );
or ( n13147 , n13141 , n13146 );
nand ( n13148 , n12766 , n12789 );
nand ( n13149 , n13147 , n13148 );
xor ( n13150 , n13140 , n13149 );
xor ( n13151 , n13107 , n13150 );
xor ( n13152 , n13043 , n13047 );
xor ( n13153 , n13152 , n13103 );
not ( n13154 , n13119 );
not ( n13155 , n13074 );
or ( n13156 , n13154 , n13155 );
not ( n13157 , n495 );
not ( n13158 , n13037 );
or ( n13159 , n13157 , n13158 );
not ( n13160 , n13036 );
not ( n13161 , n13160 );
nand ( n13162 , n13161 , n3583 );
nand ( n13163 , n13159 , n13162 );
nand ( n13164 , n13163 , n13056 );
nand ( n13165 , n13156 , n13164 );
not ( n13166 , n12563 );
not ( n13167 , n12604 );
or ( n13168 , n13166 , n13167 );
and ( n13169 , n12579 , n13096 );
not ( n13170 , n12579 );
and ( n13171 , n13170 , n13095 );
or ( n13172 , n13169 , n13171 );
not ( n13173 , n13172 );
nand ( n13174 , n13173 , n12610 );
nand ( n13175 , n13168 , n13174 );
xor ( n13176 , n13165 , n13175 );
not ( n13177 , n12845 );
not ( n13178 , n12874 );
or ( n13179 , n13177 , n13178 );
not ( n13180 , n493 );
not ( n13181 , n12698 );
not ( n13182 , n13181 );
or ( n13183 , n13180 , n13182 );
nand ( n13184 , n12862 , n12699 );
nand ( n13185 , n13183 , n13184 );
nand ( n13186 , n13185 , n12878 );
nand ( n13187 , n13179 , n13186 );
not ( n13188 , n12673 );
not ( n13189 , n12813 );
or ( n13190 , n13188 , n13189 );
xor ( n13191 , n489 , n12822 );
nand ( n13192 , n13191 , n12635 );
nand ( n13193 , n13190 , n13192 );
nand ( n13194 , n11932 , n11857 );
xnor ( n13195 , n11928 , n13194 );
and ( n13196 , n489 , n13195 );
xor ( n13197 , n13193 , n13196 );
not ( n13198 , n12731 );
not ( n13199 , n12837 );
or ( n13200 , n13198 , n13199 );
and ( n13201 , n12624 , n12703 );
not ( n13202 , n12624 );
and ( n13203 , n13202 , n491 );
or ( n13204 , n13201 , n13203 );
nand ( n13205 , n13204 , n12688 );
nand ( n13206 , n13200 , n13205 );
and ( n13207 , n13197 , n13206 );
and ( n13208 , n13193 , n13196 );
or ( n13209 , n13207 , n13208 );
xor ( n13210 , n13187 , n13209 );
not ( n13211 , n13119 );
not ( n13212 , n13163 );
or ( n13213 , n13211 , n13212 );
and ( n13214 , n495 , n12987 );
not ( n13215 , n495 );
and ( n13216 , n13215 , n12861 );
or ( n13217 , n13214 , n13216 );
nand ( n13218 , n13217 , n13056 );
nand ( n13219 , n13213 , n13218 );
and ( n13220 , n13210 , n13219 );
and ( n13221 , n13187 , n13209 );
or ( n13222 , n13220 , n13221 );
and ( n13223 , n13176 , n13222 );
and ( n13224 , n13165 , n13175 );
or ( n13225 , n13223 , n13224 );
xor ( n13226 , n13153 , n13225 );
xor ( n13227 , n12612 , n12738 );
xor ( n13228 , n13227 , n12791 );
and ( n13229 , n13226 , n13228 );
and ( n13230 , n13153 , n13225 );
or ( n13231 , n13229 , n13230 );
and ( n13232 , n13151 , n13231 );
and ( n13233 , n13107 , n13150 );
or ( n13234 , n13232 , n13233 );
xor ( n13235 , n12983 , n13234 );
xor ( n13236 , n13129 , n13139 );
and ( n13237 , n13236 , n13149 );
and ( n13238 , n13129 , n13139 );
or ( n13239 , n13237 , n13238 );
not ( n13240 , n12909 );
not ( n13241 , n13135 );
or ( n13242 , n13240 , n13241 );
not ( n13243 , n501 );
not ( n13244 , n12546 );
or ( n13245 , n13243 , n13244 );
nand ( n13246 , n12549 , n12943 );
nand ( n13247 , n13245 , n13246 );
nand ( n13248 , n13247 , n12930 );
nand ( n13249 , n13242 , n13248 );
not ( n13250 , n12789 );
not ( n13251 , n13145 );
or ( n13252 , n13250 , n13251 );
and ( n13253 , n499 , n12942 );
not ( n13254 , n499 );
and ( n13255 , n13254 , n12939 );
nor ( n13256 , n13253 , n13255 );
nand ( n13257 , n12743 , n13256 );
nand ( n13258 , n13252 , n13257 );
xor ( n13259 , n13249 , n13258 );
not ( n13260 , n12555 );
not ( n13261 , n12518 );
or ( n13262 , n13260 , n13261 );
not ( n13263 , n503 );
not ( n13264 , n10809 );
nand ( n13265 , n10590 , n12505 );
nor ( n13266 , n13264 , n13265 );
and ( n13267 , n13266 , n12409 );
not ( n13268 , n13267 );
not ( n13269 , n12755 );
or ( n13270 , n13268 , n13269 );
not ( n13271 , n12428 );
not ( n13272 , n13266 );
or ( n13273 , n13271 , n13272 );
nand ( n13274 , n13273 , n12503 );
nand ( n13275 , n12445 , n12505 );
not ( n13276 , n13275 );
nor ( n13277 , n13274 , n13276 );
nand ( n13278 , n13270 , n13277 );
not ( n13279 , n12462 );
not ( n13280 , n12470 );
or ( n13281 , n13279 , n13280 );
or ( n13282 , n12462 , n12470 );
nand ( n13283 , n13282 , n10558 );
nand ( n13284 , n13281 , n13283 );
xor ( n13285 , n12461 , n12471 );
and ( n13286 , n13285 , n12488 );
and ( n13287 , n12461 , n12471 );
or ( n13288 , n13286 , n13287 );
xor ( n13289 , n13284 , n13288 );
not ( n13290 , n12482 );
not ( n13291 , n10314 );
or ( n13292 , n13290 , n13291 );
nand ( n13293 , n10317 , n461 );
nand ( n13294 , n13292 , n13293 );
not ( n13295 , n13294 );
and ( n13296 , n457 , n526 );
not ( n13297 , n12476 );
not ( n13298 , n10256 );
or ( n13299 , n13297 , n13298 );
xor ( n13300 , n457 , n524 );
nand ( n13301 , n10197 , n13300 );
nand ( n13302 , n13299 , n13301 );
xor ( n13303 , n13296 , n13302 );
not ( n13304 , n12468 );
not ( n13305 , n10216 );
or ( n13306 , n13304 , n13305 );
xor ( n13307 , n459 , n522 );
nand ( n13308 , n10223 , n13307 );
nand ( n13309 , n13306 , n13308 );
xor ( n13310 , n13303 , n13309 );
xor ( n13311 , n13295 , n13310 );
xor ( n13312 , n12478 , n12484 );
and ( n13313 , n13312 , n12487 );
and ( n13314 , n12478 , n12484 );
or ( n13315 , n13313 , n13314 );
xor ( n13316 , n13311 , n13315 );
xor ( n13317 , n13289 , n13316 );
not ( n13318 , n12456 );
not ( n13319 , n12489 );
or ( n13320 , n13318 , n13319 );
not ( n13321 , n12457 );
not ( n13322 , n12489 );
not ( n13323 , n13322 );
or ( n13324 , n13321 , n13323 );
nand ( n13325 , n13324 , n12494 );
nand ( n13326 , n13320 , n13325 );
nor ( n13327 , n13317 , n13326 );
not ( n13328 , n13327 );
nand ( n13329 , n13326 , n13317 );
nand ( n13330 , n13328 , n13329 );
and ( n13331 , n13278 , n13330 );
not ( n13332 , n13278 );
not ( n13333 , n13330 );
and ( n13334 , n13332 , n13333 );
nor ( n13335 , n13331 , n13334 );
buf ( n13336 , n13335 );
not ( n13337 , n13336 );
or ( n13338 , n13263 , n13337 );
not ( n13339 , n13335 );
nand ( n13340 , n13339 , n12516 );
nand ( n13341 , n13338 , n13340 );
nand ( n13342 , n13341 , n504 );
nand ( n13343 , n13262 , n13342 );
xor ( n13344 , n13259 , n13343 );
xor ( n13345 , n13239 , n13344 );
not ( n13346 , n12878 );
not ( n13347 , n13113 );
or ( n13348 , n13346 , n13347 );
and ( n13349 , n493 , n13095 );
not ( n13350 , n493 );
and ( n13351 , n13350 , n13096 );
nor ( n13352 , n13349 , n13351 );
nand ( n13353 , n13352 , n12845 );
nand ( n13354 , n13348 , n13353 );
not ( n13355 , n13056 );
not ( n13356 , n13124 );
or ( n13357 , n13355 , n13356 );
and ( n13358 , n495 , n12574 );
not ( n13359 , n495 );
and ( n13360 , n13359 , n12575 );
nor ( n13361 , n13358 , n13360 );
nand ( n13362 , n13361 , n13119 );
nand ( n13363 , n13357 , n13362 );
xor ( n13364 , n13354 , n13363 );
xor ( n13365 , n12984 , n12995 );
and ( n13366 , n13365 , n13008 );
and ( n13367 , n12984 , n12995 );
or ( n13368 , n13366 , n13367 );
xor ( n13369 , n13364 , n13368 );
xor ( n13370 , n13009 , n13019 );
and ( n13371 , n13370 , n13106 );
and ( n13372 , n13009 , n13019 );
or ( n13373 , n13371 , n13372 );
xor ( n13374 , n13369 , n13373 );
not ( n13375 , n12610 );
not ( n13376 , n13015 );
or ( n13377 , n13375 , n13376 );
not ( n13378 , n497 );
not ( n13379 , n12761 );
or ( n13380 , n13378 , n13379 );
nand ( n13381 , n12764 , n12579 );
nand ( n13382 , n13380 , n13381 );
nand ( n13383 , n13382 , n12563 );
nand ( n13384 , n13377 , n13383 );
and ( n13385 , n13036 , n12703 );
not ( n13386 , n13036 );
and ( n13387 , n13386 , n491 );
or ( n13388 , n13385 , n13387 );
not ( n13389 , n13388 );
not ( n13390 , n12731 );
or ( n13391 , n13389 , n13390 );
nand ( n13392 , n12991 , n12688 );
nand ( n13393 , n13391 , n13392 );
and ( n13394 , n12997 , n13007 );
xor ( n13395 , n13393 , n13394 );
not ( n13396 , n12635 );
not ( n13397 , n13003 );
or ( n13398 , n13396 , n13397 );
not ( n13399 , n489 );
not ( n13400 , n12722 );
or ( n13401 , n13399 , n13400 );
nand ( n13402 , n12721 , n12653 );
nand ( n13403 , n13401 , n13402 );
nand ( n13404 , n13403 , n12882 );
nand ( n13405 , n13398 , n13404 );
and ( n13406 , n12666 , n489 );
xor ( n13407 , n13405 , n13406 );
xor ( n13408 , n13395 , n13407 );
xor ( n13409 , n13384 , n13408 );
xor ( n13410 , n13108 , n13117 );
and ( n13411 , n13410 , n13128 );
and ( n13412 , n13108 , n13117 );
or ( n13413 , n13411 , n13412 );
xor ( n13414 , n13409 , n13413 );
xor ( n13415 , n13374 , n13414 );
xor ( n13416 , n13345 , n13415 );
xor ( n13417 , n13235 , n13416 );
not ( n13418 , n13417 );
xor ( n13419 , n12557 , n12794 );
xor ( n13420 , n13419 , n12980 );
not ( n13421 , n12743 );
not ( n13422 , n12785 );
or ( n13423 , n13421 , n13422 );
and ( n13424 , n499 , n12575 );
not ( n13425 , n499 );
and ( n13426 , n13425 , n12574 );
nor ( n13427 , n13424 , n13426 );
not ( n13428 , n13427 );
nand ( n13429 , n13428 , n12789 );
nand ( n13430 , n13423 , n13429 );
xor ( n13431 , n12842 , n12880 );
xor ( n13432 , n13431 , n12895 );
xor ( n13433 , n13430 , n13432 );
not ( n13434 , n12930 );
not ( n13435 , n12927 );
or ( n13436 , n13434 , n13435 );
not ( n13437 , n501 );
not ( n13438 , n12760 );
not ( n13439 , n13438 );
or ( n13440 , n13437 , n13439 );
or ( n13441 , n13438 , n501 );
nand ( n13442 , n13440 , n13441 );
nand ( n13443 , n13442 , n12909 );
nand ( n13444 , n13436 , n13443 );
and ( n13445 , n13433 , n13444 );
and ( n13446 , n13430 , n13432 );
or ( n13447 , n13445 , n13446 );
not ( n13448 , n699 );
nand ( n13449 , n13448 , n12973 );
buf ( n13450 , n12938 );
not ( n13451 , n13450 );
nand ( n13452 , n13451 , n12555 );
buf ( n13453 , n12972 );
nand ( n13454 , n13453 , n4208 );
nand ( n13455 , n13449 , n13452 , n13454 );
xor ( n13456 , n12815 , n12823 );
xor ( n13457 , n13456 , n12839 );
not ( n13458 , n497 );
not ( n13459 , n13072 );
not ( n13460 , n13459 );
or ( n13461 , n13458 , n13460 );
nand ( n13462 , n13072 , n12579 );
nand ( n13463 , n13461 , n13462 );
not ( n13464 , n13463 );
not ( n13465 , n12610 );
or ( n13466 , n13464 , n13465 );
or ( n13467 , n13172 , n12562 );
nand ( n13468 , n13466 , n13467 );
xor ( n13469 , n13457 , n13468 );
and ( n13470 , n12560 , n12602 );
not ( n13471 , n12560 );
and ( n13472 , n13471 , n12599 );
nor ( n13473 , n13470 , n13472 );
or ( n13474 , n13473 , n12788 );
or ( n13475 , n13427 , n12742 );
nand ( n13476 , n13474 , n13475 );
and ( n13477 , n13469 , n13476 );
and ( n13478 , n13457 , n13468 );
or ( n13479 , n13477 , n13478 );
xor ( n13480 , n13455 , n13479 );
xor ( n13481 , n13165 , n13175 );
xor ( n13482 , n13481 , n13222 );
and ( n13483 , n13480 , n13482 );
and ( n13484 , n13455 , n13479 );
or ( n13485 , n13483 , n13484 );
xor ( n13486 , n13447 , n13485 );
xor ( n13487 , n12898 , n12947 );
xor ( n13488 , n13487 , n12977 );
and ( n13489 , n13486 , n13488 );
and ( n13490 , n13447 , n13485 );
or ( n13491 , n13489 , n13490 );
xor ( n13492 , n13420 , n13491 );
xor ( n13493 , n13107 , n13150 );
xor ( n13494 , n13493 , n13231 );
and ( n13495 , n13492 , n13494 );
and ( n13496 , n13420 , n13491 );
or ( n13497 , n13495 , n13496 );
not ( n13498 , n13497 );
nand ( n13499 , n13418 , n13498 );
xor ( n13500 , n13420 , n13491 );
xor ( n13501 , n13500 , n13494 );
xor ( n13502 , n13153 , n13225 );
xor ( n13503 , n13502 , n13228 );
not ( n13504 , n12882 );
not ( n13505 , n13191 );
or ( n13506 , n13504 , n13505 );
xor ( n13507 , n489 , n13195 );
nand ( n13508 , n13507 , n12635 );
nand ( n13509 , n13506 , n13508 );
not ( n13510 , n11908 );
not ( n13511 , n11926 );
not ( n13512 , n11925 );
or ( n13513 , n13511 , n13512 );
nand ( n13514 , n13513 , n11922 );
not ( n13515 , n13514 );
or ( n13516 , n13510 , n13515 );
or ( n13517 , n13514 , n11908 );
nand ( n13518 , n13516 , n13517 );
buf ( n13519 , n13518 );
and ( n13520 , n489 , n13519 );
xor ( n13521 , n13509 , n13520 );
not ( n13522 , n12731 );
not ( n13523 , n13204 );
or ( n13524 , n13522 , n13523 );
not ( n13525 , n491 );
not ( n13526 , n12811 );
not ( n13527 , n13526 );
or ( n13528 , n13525 , n13527 );
nand ( n13529 , n12812 , n12703 );
nand ( n13530 , n13528 , n13529 );
nand ( n13531 , n13530 , n12688 );
nand ( n13532 , n13524 , n13531 );
and ( n13533 , n13521 , n13532 );
and ( n13534 , n13509 , n13520 );
or ( n13535 , n13533 , n13534 );
not ( n13536 , n12845 );
not ( n13537 , n13185 );
or ( n13538 , n13536 , n13537 );
not ( n13539 , n493 );
not ( n13540 , n12665 );
or ( n13541 , n13539 , n13540 );
or ( n13542 , n12665 , n493 );
nand ( n13543 , n13541 , n13542 );
not ( n13544 , n13543 );
nand ( n13545 , n13544 , n12878 );
nand ( n13546 , n13538 , n13545 );
xor ( n13547 , n13535 , n13546 );
xor ( n13548 , n13193 , n13196 );
xor ( n13549 , n13548 , n13206 );
and ( n13550 , n13547 , n13549 );
and ( n13551 , n13535 , n13546 );
or ( n13552 , n13550 , n13551 );
xor ( n13553 , n13187 , n13209 );
xor ( n13554 , n13553 , n13219 );
xor ( n13555 , n13552 , n13554 );
not ( n13556 , n12909 );
not ( n13557 , n501 );
buf ( n13558 , n12780 );
not ( n13559 , n13558 );
not ( n13560 , n13559 );
or ( n13561 , n13557 , n13560 );
nand ( n13562 , n13558 , n12943 );
nand ( n13563 , n13561 , n13562 );
not ( n13564 , n13563 );
or ( n13565 , n13556 , n13564 );
nand ( n13566 , n13442 , n12930 );
nand ( n13567 , n13565 , n13566 );
and ( n13568 , n13555 , n13567 );
and ( n13569 , n13552 , n13554 );
or ( n13570 , n13568 , n13569 );
not ( n13571 , n13119 );
not ( n13572 , n13217 );
or ( n13573 , n13571 , n13572 );
and ( n13574 , n495 , n12722 );
not ( n13575 , n495 );
and ( n13576 , n13575 , n12721 );
nor ( n13577 , n13574 , n13576 );
not ( n13578 , n13577 );
nand ( n13579 , n13578 , n13056 );
nand ( n13580 , n13573 , n13579 );
and ( n13581 , n11907 , n11881 );
buf ( n13582 , n11903 );
and ( n13583 , n13581 , n13582 );
not ( n13584 , n13581 );
not ( n13585 , n13582 );
and ( n13586 , n13584 , n13585 );
nor ( n13587 , n13583 , n13586 );
and ( n13588 , n489 , n13587 );
xor ( n13589 , n489 , n13519 );
not ( n13590 , n13589 );
not ( n13591 , n12635 );
or ( n13592 , n13590 , n13591 );
not ( n13593 , n13507 );
or ( n13594 , n13593 , n12632 );
nand ( n13595 , n13592 , n13594 );
xor ( n13596 , n13588 , n13595 );
not ( n13597 , n12688 );
not ( n13598 , n491 );
not ( n13599 , n12822 );
not ( n13600 , n13599 );
or ( n13601 , n13598 , n13600 );
nand ( n13602 , n12822 , n12703 );
nand ( n13603 , n13601 , n13602 );
not ( n13604 , n13603 );
or ( n13605 , n13597 , n13604 );
nand ( n13606 , n13530 , n12731 );
nand ( n13607 , n13605 , n13606 );
and ( n13608 , n13596 , n13607 );
and ( n13609 , n13588 , n13595 );
or ( n13610 , n13608 , n13609 );
and ( n13611 , n12862 , n12649 );
not ( n13612 , n12862 );
and ( n13613 , n13612 , n12652 );
or ( n13614 , n13611 , n13613 );
not ( n13615 , n12878 );
or ( n13616 , n13614 , n13615 );
or ( n13617 , n13543 , n12844 );
nand ( n13618 , n13616 , n13617 );
xor ( n13619 , n13610 , n13618 );
xor ( n13620 , n13509 , n13520 );
xor ( n13621 , n13620 , n13532 );
and ( n13622 , n13619 , n13621 );
and ( n13623 , n13610 , n13618 );
or ( n13624 , n13622 , n13623 );
xor ( n13625 , n13580 , n13624 );
not ( n13626 , n12563 );
not ( n13627 , n13463 );
or ( n13628 , n13626 , n13627 );
and ( n13629 , n12579 , n13036 );
not ( n13630 , n12579 );
and ( n13631 , n13630 , n13160 );
nor ( n13632 , n13629 , n13631 );
not ( n13633 , n13632 );
nand ( n13634 , n13633 , n12610 );
nand ( n13635 , n13628 , n13634 );
and ( n13636 , n13625 , n13635 );
and ( n13637 , n13580 , n13624 );
or ( n13638 , n13636 , n13637 );
not ( n13639 , n499 );
not ( n13640 , n13096 );
or ( n13641 , n13639 , n13640 );
nand ( n13642 , n13095 , n12560 );
nand ( n13643 , n13641 , n13642 );
nand ( n13644 , n13643 , n12789 );
nand ( n13645 , n12741 , n499 );
or ( n13646 , n12598 , n13645 );
nor ( n13647 , n12742 , n499 );
nand ( n13648 , n12598 , n13647 );
nand ( n13649 , n13644 , n13646 , n13648 );
xor ( n13650 , n13535 , n13546 );
xor ( n13651 , n13650 , n13549 );
xor ( n13652 , n13649 , n13651 );
and ( n13653 , n495 , n13181 );
not ( n13654 , n495 );
and ( n13655 , n13654 , n12699 );
nor ( n13656 , n13653 , n13655 );
not ( n13657 , n13056 );
or ( n13658 , n13656 , n13657 );
or ( n13659 , n13577 , n13052 );
nand ( n13660 , n13658 , n13659 );
xor ( n13661 , n12579 , n12861 );
or ( n13662 , n13661 , n13465 );
or ( n13663 , n13632 , n12562 );
nand ( n13664 , n13662 , n13663 );
xor ( n13665 , n13660 , n13664 );
not ( n13666 , n11891 );
not ( n13667 , n13666 );
not ( n13668 , n13667 );
not ( n13669 , n11899 );
nand ( n13670 , n13669 , n11902 );
not ( n13671 , n13670 );
not ( n13672 , n13671 );
or ( n13673 , n13668 , n13672 );
nand ( n13674 , n13670 , n13666 );
nand ( n13675 , n13673 , n13674 );
and ( n13676 , n13675 , n489 );
not ( n13677 , n12882 );
not ( n13678 , n13589 );
or ( n13679 , n13677 , n13678 );
xor ( n13680 , n489 , n13587 );
nand ( n13681 , n13680 , n12635 );
nand ( n13682 , n13679 , n13681 );
xor ( n13683 , n13676 , n13682 );
not ( n13684 , n12731 );
not ( n13685 , n13603 );
or ( n13686 , n13684 , n13685 );
not ( n13687 , n13195 );
not ( n13688 , n13687 );
and ( n13689 , n491 , n13688 );
not ( n13690 , n491 );
and ( n13691 , n13690 , n13687 );
nor ( n13692 , n13689 , n13691 );
nand ( n13693 , n13692 , n12688 );
nand ( n13694 , n13686 , n13693 );
and ( n13695 , n13683 , n13694 );
and ( n13696 , n13676 , n13682 );
or ( n13697 , n13695 , n13696 );
not ( n13698 , n493 );
not ( n13699 , n12625 );
or ( n13700 , n13698 , n13699 );
nand ( n13701 , n12624 , n12862 );
nand ( n13702 , n13700 , n13701 );
not ( n13703 , n13702 );
not ( n13704 , n12878 );
or ( n13705 , n13703 , n13704 );
or ( n13706 , n13614 , n12844 );
nand ( n13707 , n13705 , n13706 );
xor ( n13708 , n13697 , n13707 );
xor ( n13709 , n13588 , n13595 );
xor ( n13710 , n13709 , n13607 );
and ( n13711 , n13708 , n13710 );
and ( n13712 , n13697 , n13707 );
or ( n13713 , n13711 , n13712 );
and ( n13714 , n13665 , n13713 );
and ( n13715 , n13660 , n13664 );
or ( n13716 , n13714 , n13715 );
and ( n13717 , n13652 , n13716 );
and ( n13718 , n13649 , n13651 );
or ( n13719 , n13717 , n13718 );
xor ( n13720 , n13638 , n13719 );
not ( n13721 , n12555 );
not ( n13722 , n503 );
not ( n13723 , n12923 );
or ( n13724 , n13722 , n13723 );
not ( n13725 , n12923 );
nand ( n13726 , n13725 , n12550 );
nand ( n13727 , n13724 , n13726 );
not ( n13728 , n13727 );
or ( n13729 , n13721 , n13728 );
nand ( n13730 , n12942 , n12550 );
not ( n13731 , n13730 );
nand ( n13732 , n12939 , n503 );
not ( n13733 , n13732 );
or ( n13734 , n13731 , n13733 );
nand ( n13735 , n13734 , n504 );
nand ( n13736 , n13729 , n13735 );
and ( n13737 , n13720 , n13736 );
and ( n13738 , n13638 , n13719 );
or ( n13739 , n13737 , n13738 );
xor ( n13740 , n13570 , n13739 );
xor ( n13741 , n13430 , n13432 );
xor ( n13742 , n13741 , n13444 );
and ( n13743 , n13740 , n13742 );
and ( n13744 , n13570 , n13739 );
or ( n13745 , n13743 , n13744 );
xor ( n13746 , n13503 , n13745 );
xor ( n13747 , n13447 , n13485 );
xor ( n13748 , n13747 , n13488 );
and ( n13749 , n13746 , n13748 );
and ( n13750 , n13503 , n13745 );
or ( n13751 , n13749 , n13750 );
and ( n13752 , n13501 , n13751 );
and ( n13753 , n13499 , n13752 );
and ( n13754 , n13417 , n13497 );
nor ( n13755 , n13753 , n13754 );
not ( n13756 , n13755 );
xor ( n13757 , n13503 , n13745 );
xor ( n13758 , n13757 , n13748 );
xor ( n13759 , n13455 , n13479 );
xor ( n13760 , n13759 , n13482 );
xor ( n13761 , n13457 , n13468 );
xor ( n13762 , n13761 , n13476 );
xor ( n13763 , n13552 , n13554 );
xor ( n13764 , n13763 , n13567 );
xor ( n13765 , n13762 , n13764 );
xor ( n13766 , n13580 , n13624 );
xor ( n13767 , n13766 , n13635 );
not ( n13768 , n12930 );
not ( n13769 , n13563 );
or ( n13770 , n13768 , n13769 );
not ( n13771 , n501 );
not ( n13772 , n12576 );
or ( n13773 , n13771 , n13772 );
not ( n13774 , n12576 );
nand ( n13775 , n13774 , n12943 );
nand ( n13776 , n13773 , n13775 );
nand ( n13777 , n13776 , n12909 );
nand ( n13778 , n13770 , n13777 );
xor ( n13779 , n13767 , n13778 );
not ( n13780 , n13727 );
not ( n13781 , n504 );
or ( n13782 , n13780 , n13781 );
not ( n13783 , n503 );
not ( n13784 , n12761 );
or ( n13785 , n13783 , n13784 );
nand ( n13786 , n12764 , n12550 );
nand ( n13787 , n13785 , n13786 );
nand ( n13788 , n13787 , n12555 );
nand ( n13789 , n13782 , n13788 );
and ( n13790 , n13779 , n13789 );
and ( n13791 , n13767 , n13778 );
or ( n13792 , n13790 , n13791 );
and ( n13793 , n13765 , n13792 );
and ( n13794 , n13762 , n13764 );
or ( n13795 , n13793 , n13794 );
xor ( n13796 , n13760 , n13795 );
xor ( n13797 , n13570 , n13739 );
xor ( n13798 , n13797 , n13742 );
and ( n13799 , n13796 , n13798 );
and ( n13800 , n13760 , n13795 );
or ( n13801 , n13799 , n13800 );
nor ( n13802 , n13758 , n13801 );
not ( n13803 , n13802 );
not ( n13804 , n12845 );
not ( n13805 , n12822 );
not ( n13806 , n13805 );
and ( n13807 , n493 , n13806 );
not ( n13808 , n493 );
and ( n13809 , n13808 , n13599 );
nor ( n13810 , n13807 , n13809 );
not ( n13811 , n13810 );
or ( n13812 , n13804 , n13811 );
and ( n13813 , n493 , n13688 );
not ( n13814 , n493 );
and ( n13815 , n13814 , n13687 );
nor ( n13816 , n13813 , n13815 );
nand ( n13817 , n13816 , n12878 );
nand ( n13818 , n13812 , n13817 );
not ( n13819 , n13119 );
and ( n13820 , n495 , n12625 );
not ( n13821 , n495 );
and ( n13822 , n13821 , n12624 );
or ( n13823 , n13820 , n13822 );
not ( n13824 , n13823 );
or ( n13825 , n13819 , n13824 );
and ( n13826 , n495 , n12812 );
not ( n13827 , n495 );
and ( n13828 , n13827 , n13526 );
nor ( n13829 , n13826 , n13828 );
nand ( n13830 , n13829 , n13056 );
nand ( n13831 , n13825 , n13830 );
xor ( n13832 , n13818 , n13831 );
not ( n13833 , n12731 );
not ( n13834 , n491 );
not ( n13835 , n13519 );
not ( n13836 , n13835 );
or ( n13837 , n13834 , n13836 );
nand ( n13838 , n13519 , n12703 );
nand ( n13839 , n13837 , n13838 );
not ( n13840 , n13839 );
or ( n13841 , n13833 , n13840 );
buf ( n13842 , n13587 );
and ( n13843 , n491 , n13842 );
not ( n13844 , n491 );
not ( n13845 , n13587 );
and ( n13846 , n13844 , n13845 );
nor ( n13847 , n13843 , n13846 );
nand ( n13848 , n13847 , n12688 );
nand ( n13849 , n13841 , n13848 );
nand ( n13850 , n536 , n472 );
not ( n13851 , n13850 );
and ( n13852 , n489 , n13851 );
not ( n13853 , n12882 );
not ( n13854 , n489 );
not ( n13855 , n11891 );
not ( n13856 , n13670 );
or ( n13857 , n13855 , n13856 );
nand ( n13858 , n13671 , n13666 );
nand ( n13859 , n13857 , n13858 );
not ( n13860 , n13859 );
or ( n13861 , n13854 , n13860 );
or ( n13862 , n13859 , n489 );
nand ( n13863 , n13861 , n13862 );
not ( n13864 , n13863 );
or ( n13865 , n13853 , n13864 );
not ( n13866 , n11890 );
not ( n13867 , n11888 );
or ( n13868 , n13866 , n13867 );
or ( n13869 , n11888 , n11890 );
nand ( n13870 , n13868 , n13869 );
not ( n13871 , n13870 );
xor ( n13872 , n489 , n13871 );
nand ( n13873 , n13872 , n12635 );
nand ( n13874 , n13865 , n13873 );
xor ( n13875 , n13852 , n13874 );
or ( n13876 , n13851 , n490 );
nand ( n13877 , n13876 , n491 );
nand ( n13878 , n13851 , n490 );
and ( n13879 , n13877 , n13878 , n489 );
not ( n13880 , n12882 );
not ( n13881 , n13872 );
or ( n13882 , n13880 , n13881 );
xor ( n13883 , n489 , n13851 );
nand ( n13884 , n13883 , n12635 );
nand ( n13885 , n13882 , n13884 );
and ( n13886 , n13879 , n13885 );
xor ( n13887 , n13875 , n13886 );
xor ( n13888 , n13849 , n13887 );
xor ( n13889 , n13879 , n13885 );
not ( n13890 , n12731 );
not ( n13891 , n13847 );
or ( n13892 , n13890 , n13891 );
or ( n13893 , n13675 , n1993 );
nand ( n13894 , n13675 , n12703 );
nand ( n13895 , n13893 , n13894 );
nand ( n13896 , n12688 , n13895 );
nand ( n13897 , n13892 , n13896 );
xor ( n13898 , n13889 , n13897 );
nor ( n13899 , n13850 , n12632 );
not ( n13900 , n12731 );
not ( n13901 , n13895 );
or ( n13902 , n13900 , n13901 );
and ( n13903 , n491 , n13871 );
not ( n13904 , n491 );
and ( n13905 , n13904 , n13870 );
nor ( n13906 , n13903 , n13905 );
nand ( n13907 , n13906 , n12688 );
nand ( n13908 , n13902 , n13907 );
xor ( n13909 , n13899 , n13908 );
or ( n13910 , n13851 , n492 );
nand ( n13911 , n13910 , n493 );
and ( n13912 , n13851 , n492 );
nor ( n13913 , n13912 , n12703 );
and ( n13914 , n13911 , n13913 );
not ( n13915 , n12731 );
not ( n13916 , n13906 );
or ( n13917 , n13915 , n13916 );
or ( n13918 , n13850 , n491 );
or ( n13919 , n13851 , n12703 );
nand ( n13920 , n13918 , n13919 );
nand ( n13921 , n13920 , n12688 );
nand ( n13922 , n13917 , n13921 );
and ( n13923 , n13914 , n13922 );
and ( n13924 , n13909 , n13923 );
and ( n13925 , n13899 , n13908 );
or ( n13926 , n13924 , n13925 );
and ( n13927 , n13898 , n13926 );
and ( n13928 , n13889 , n13897 );
or ( n13929 , n13927 , n13928 );
xor ( n13930 , n13888 , n13929 );
and ( n13931 , n13832 , n13930 );
and ( n13932 , n13818 , n13831 );
or ( n13933 , n13931 , n13932 );
not ( n13934 , n12563 );
and ( n13935 , n497 , n12699 );
not ( n13936 , n497 );
and ( n13937 , n13936 , n12700 );
nor ( n13938 , n13935 , n13937 );
not ( n13939 , n13938 );
or ( n13940 , n13934 , n13939 );
not ( n13941 , n497 );
not ( n13942 , n12670 );
or ( n13943 , n13941 , n13942 );
nand ( n13944 , n12666 , n12579 );
nand ( n13945 , n13943 , n13944 );
nand ( n13946 , n12610 , n13945 );
nand ( n13947 , n13940 , n13946 );
xor ( n13948 , n13933 , n13947 );
not ( n13949 , n12743 );
not ( n13950 , n499 );
not ( n13951 , n12987 );
or ( n13952 , n13950 , n13951 );
nand ( n13953 , n12861 , n12560 );
nand ( n13954 , n13952 , n13953 );
not ( n13955 , n13954 );
or ( n13956 , n13949 , n13955 );
not ( n13957 , n499 );
not ( n13958 , n12722 );
or ( n13959 , n13957 , n13958 );
nand ( n13960 , n12560 , n12721 );
nand ( n13961 , n13959 , n13960 );
nand ( n13962 , n13961 , n12789 );
nand ( n13963 , n13956 , n13962 );
xor ( n13964 , n13948 , n13963 );
not ( n13965 , n12555 );
not ( n13966 , n503 );
not ( n13967 , n13096 );
or ( n13968 , n13966 , n13967 );
nand ( n13969 , n13095 , n12516 );
nand ( n13970 , n13968 , n13969 );
not ( n13971 , n13970 );
or ( n13972 , n13965 , n13971 );
and ( n13973 , n12599 , n503 );
not ( n13974 , n12599 );
and ( n13975 , n13974 , n12550 );
or ( n13976 , n13973 , n13975 );
nand ( n13977 , n13976 , n504 );
nand ( n13978 , n13972 , n13977 );
xor ( n13979 , n13964 , n13978 );
xor ( n13980 , n13818 , n13831 );
xor ( n13981 , n13980 , n13930 );
not ( n13982 , n12845 );
and ( n13983 , n12862 , n13835 );
not ( n13984 , n12862 );
and ( n13985 , n13984 , n13519 );
nor ( n13986 , n13983 , n13985 );
not ( n13987 , n13986 );
or ( n13988 , n13982 , n13987 );
and ( n13989 , n493 , n13587 );
not ( n13990 , n493 );
and ( n13991 , n13990 , n13845 );
nor ( n13992 , n13989 , n13991 );
nand ( n13993 , n13992 , n12878 );
nand ( n13994 , n13988 , n13993 );
xor ( n13995 , n13899 , n13908 );
xor ( n13996 , n13995 , n13923 );
xor ( n13997 , n13994 , n13996 );
xor ( n13998 , n13914 , n13922 );
not ( n13999 , n12845 );
not ( n14000 , n13992 );
or ( n14001 , n13999 , n14000 );
not ( n14002 , n493 );
not ( n14003 , n13859 );
or ( n14004 , n14002 , n14003 );
or ( n14005 , n13859 , n493 );
nand ( n14006 , n14004 , n14005 );
nand ( n14007 , n14006 , n12878 );
nand ( n14008 , n14001 , n14007 );
xor ( n14009 , n13998 , n14008 );
nor ( n14010 , n12686 , n13850 );
not ( n14011 , n12843 );
and ( n14012 , n493 , n13871 );
not ( n14013 , n493 );
and ( n14014 , n14013 , n13870 );
nor ( n14015 , n14012 , n14014 );
not ( n14016 , n14015 );
or ( n14017 , n14011 , n14016 );
or ( n14018 , n13850 , n493 );
or ( n14019 , n13851 , n12862 );
nand ( n14020 , n14018 , n14019 );
nand ( n14021 , n14020 , n12878 );
nand ( n14022 , n14017 , n14021 );
or ( n14023 , n13851 , n494 );
nand ( n14024 , n14023 , n495 );
and ( n14025 , n13851 , n494 );
nor ( n14026 , n14025 , n12862 );
nand ( n14027 , n14024 , n14026 );
not ( n14028 , n14027 );
and ( n14029 , n14022 , n14028 );
xor ( n14030 , n14010 , n14029 );
not ( n14031 , n12845 );
not ( n14032 , n14006 );
or ( n14033 , n14031 , n14032 );
nand ( n14034 , n14015 , n12878 );
nand ( n14035 , n14033 , n14034 );
and ( n14036 , n14030 , n14035 );
or ( n14037 , n14036 , C0 );
and ( n14038 , n14009 , n14037 );
and ( n14039 , n13998 , n14008 );
or ( n14040 , n14038 , n14039 );
and ( n14041 , n13997 , n14040 );
and ( n14042 , n13994 , n13996 );
or ( n14043 , n14041 , n14042 );
not ( n14044 , n12563 );
not ( n14045 , n497 );
not ( n14046 , n12649 );
or ( n14047 , n14045 , n14046 );
nand ( n14048 , n12652 , n12579 );
nand ( n14049 , n14047 , n14048 );
not ( n14050 , n14049 );
or ( n14051 , n14044 , n14050 );
and ( n14052 , n12624 , n12579 );
not ( n14053 , n12624 );
and ( n14054 , n14053 , n497 );
or ( n14055 , n14052 , n14054 );
nand ( n14056 , n14055 , n12610 );
nand ( n14057 , n14051 , n14056 );
xor ( n14058 , n14043 , n14057 );
not ( n14059 , n12845 );
not ( n14060 , n13816 );
or ( n14061 , n14059 , n14060 );
nand ( n14062 , n13986 , n12878 );
nand ( n14063 , n14061 , n14062 );
xor ( n14064 , n13889 , n13897 );
xor ( n14065 , n14064 , n13926 );
xor ( n14066 , n14063 , n14065 );
not ( n14067 , n13119 );
not ( n14068 , n13829 );
or ( n14069 , n14067 , n14068 );
and ( n14070 , n495 , n13805 );
not ( n14071 , n495 );
and ( n14072 , n14071 , n13806 );
or ( n14073 , n14070 , n14072 );
nand ( n14074 , n14073 , n13056 );
nand ( n14075 , n14069 , n14074 );
xor ( n14076 , n14066 , n14075 );
and ( n14077 , n14058 , n14076 );
and ( n14078 , n14043 , n14057 );
or ( n14079 , n14077 , n14078 );
xor ( n14080 , n13981 , n14079 );
not ( n14081 , n12930 );
not ( n14082 , n501 );
not ( n14083 , n13037 );
or ( n14084 , n14082 , n14083 );
nand ( n14085 , n13161 , n12943 );
nand ( n14086 , n14084 , n14085 );
not ( n14087 , n14086 );
or ( n14088 , n14081 , n14087 );
not ( n14089 , n501 );
not ( n14090 , n12987 );
or ( n14091 , n14089 , n14090 );
nand ( n14092 , n12861 , n12943 );
nand ( n14093 , n14091 , n14092 );
nand ( n14094 , n14093 , n12908 );
nand ( n14095 , n14088 , n14094 );
and ( n14096 , n14080 , n14095 );
and ( n14097 , n13981 , n14079 );
or ( n14098 , n14096 , n14097 );
and ( n14099 , n13979 , n14098 );
and ( n14100 , n13964 , n13978 );
or ( n14101 , n14099 , n14100 );
not ( n14102 , n12731 );
not ( n14103 , n13692 );
or ( n14104 , n14102 , n14103 );
nand ( n14105 , n13839 , n12688 );
nand ( n14106 , n14104 , n14105 );
and ( n14107 , n489 , n13871 );
not ( n14108 , n12635 );
not ( n14109 , n13863 );
or ( n14110 , n14108 , n14109 );
nand ( n14111 , n13680 , n12882 );
nand ( n14112 , n14110 , n14111 );
xor ( n14113 , n14107 , n14112 );
xor ( n14114 , n13852 , n13874 );
and ( n14115 , n14114 , n13886 );
and ( n14116 , n13852 , n13874 );
or ( n14117 , n14115 , n14116 );
xor ( n14118 , n14113 , n14117 );
xor ( n14119 , n14106 , n14118 );
not ( n14120 , n12878 );
not ( n14121 , n13810 );
or ( n14122 , n14120 , n14121 );
not ( n14123 , n493 );
not ( n14124 , n13526 );
or ( n14125 , n14123 , n14124 );
nand ( n14126 , n12812 , n12862 );
nand ( n14127 , n14125 , n14126 );
nand ( n14128 , n14127 , n12845 );
nand ( n14129 , n14122 , n14128 );
and ( n14130 , n14119 , n14129 );
and ( n14131 , n14106 , n14118 );
or ( n14132 , n14130 , n14131 );
not ( n14133 , n13119 );
and ( n14134 , n495 , n12670 );
not ( n14135 , n495 );
and ( n14136 , n14135 , n12666 );
or ( n14137 , n14134 , n14136 );
not ( n14138 , n14137 );
or ( n14139 , n14133 , n14138 );
not ( n14140 , n495 );
not ( n14141 , n12652 );
not ( n14142 , n14141 );
or ( n14143 , n14140 , n14142 );
not ( n14144 , n495 );
not ( n14145 , n12649 );
nand ( n14146 , n14144 , n14145 );
nand ( n14147 , n14143 , n14146 );
nand ( n14148 , n14147 , n13056 );
nand ( n14149 , n14139 , n14148 );
xor ( n14150 , n14132 , n14149 );
not ( n14151 , n12610 );
not ( n14152 , n13938 );
or ( n14153 , n14151 , n14152 );
not ( n14154 , n497 );
not ( n14155 , n12722 );
or ( n14156 , n14154 , n14155 );
not ( n14157 , n12870 );
nand ( n14158 , n14157 , n12579 );
nand ( n14159 , n14156 , n14158 );
nand ( n14160 , n14159 , n12563 );
nand ( n14161 , n14153 , n14160 );
xor ( n14162 , n14150 , n14161 );
not ( n14163 , n12908 );
not ( n14164 , n501 );
not ( n14165 , n13068 );
or ( n14166 , n14164 , n14165 );
not ( n14167 , n13068 );
nand ( n14168 , n14167 , n12943 );
nand ( n14169 , n14166 , n14168 );
not ( n14170 , n14169 );
or ( n14171 , n14163 , n14170 );
not ( n14172 , n501 );
not ( n14173 , n13096 );
or ( n14174 , n14172 , n14173 );
nand ( n14175 , n13095 , n12943 );
nand ( n14176 , n14174 , n14175 );
nand ( n14177 , n14176 , n12930 );
nand ( n14178 , n14171 , n14177 );
xor ( n14179 , n14162 , n14178 );
not ( n14180 , n504 );
not ( n14181 , n503 );
not ( n14182 , n12576 );
or ( n14183 , n14181 , n14182 );
nand ( n14184 , n13774 , n12550 );
nand ( n14185 , n14183 , n14184 );
not ( n14186 , n14185 );
or ( n14187 , n14180 , n14186 );
nand ( n14188 , n13976 , n12555 );
nand ( n14189 , n14187 , n14188 );
xor ( n14190 , n14179 , n14189 );
xor ( n14191 , n14101 , n14190 );
xor ( n14192 , n13933 , n13947 );
and ( n14193 , n14192 , n13963 );
and ( n14194 , n13933 , n13947 );
or ( n14195 , n14193 , n14194 );
xor ( n14196 , n14107 , n14112 );
and ( n14197 , n14196 , n14117 );
and ( n14198 , n14107 , n14112 );
or ( n14199 , n14197 , n14198 );
not ( n14200 , n12845 );
not ( n14201 , n13702 );
or ( n14202 , n14200 , n14201 );
nand ( n14203 , n14127 , n12878 );
nand ( n14204 , n14202 , n14203 );
xor ( n14205 , n14199 , n14204 );
xor ( n14206 , n13676 , n13682 );
xor ( n14207 , n14206 , n13694 );
xor ( n14208 , n14205 , n14207 );
not ( n14209 , n12789 );
not ( n14210 , n13954 );
or ( n14211 , n14209 , n14210 );
and ( n14212 , n13036 , n12560 );
not ( n14213 , n13036 );
and ( n14214 , n14213 , n499 );
or ( n14215 , n14212 , n14214 );
nand ( n14216 , n14215 , n12741 );
nand ( n14217 , n14211 , n14216 );
xor ( n14218 , n14208 , n14217 );
xor ( n14219 , n13849 , n13887 );
and ( n14220 , n14219 , n13929 );
and ( n14221 , n13849 , n13887 );
or ( n14222 , n14220 , n14221 );
not ( n14223 , n13119 );
not ( n14224 , n14147 );
or ( n14225 , n14223 , n14224 );
nand ( n14226 , n13823 , n13056 );
nand ( n14227 , n14225 , n14226 );
xor ( n14228 , n14222 , n14227 );
xor ( n14229 , n14106 , n14118 );
xor ( n14230 , n14229 , n14129 );
and ( n14231 , n14228 , n14230 );
and ( n14232 , n14222 , n14227 );
or ( n14233 , n14231 , n14232 );
xor ( n14234 , n14218 , n14233 );
xor ( n14235 , n14195 , n14234 );
xor ( n14236 , n14222 , n14227 );
xor ( n14237 , n14236 , n14230 );
not ( n14238 , n12610 );
not ( n14239 , n14049 );
or ( n14240 , n14238 , n14239 );
nand ( n14241 , n13945 , n12563 );
nand ( n14242 , n14240 , n14241 );
xor ( n14243 , n14063 , n14065 );
and ( n14244 , n14243 , n14075 );
and ( n14245 , n14063 , n14065 );
or ( n14246 , n14244 , n14245 );
xor ( n14247 , n14242 , n14246 );
not ( n14248 , n12789 );
not ( n14249 , n499 );
not ( n14250 , n13181 );
or ( n14251 , n14249 , n14250 );
nand ( n14252 , n12560 , n12699 );
nand ( n14253 , n14251 , n14252 );
not ( n14254 , n14253 );
or ( n14255 , n14248 , n14254 );
nand ( n14256 , n13961 , n12741 );
nand ( n14257 , n14255 , n14256 );
and ( n14258 , n14247 , n14257 );
and ( n14259 , n14242 , n14246 );
or ( n14260 , n14258 , n14259 );
xor ( n14261 , n14237 , n14260 );
not ( n14262 , n12930 );
not ( n14263 , n14169 );
or ( n14264 , n14262 , n14263 );
nand ( n14265 , n14086 , n12908 );
nand ( n14266 , n14264 , n14265 );
and ( n14267 , n14261 , n14266 );
and ( n14268 , n14237 , n14260 );
or ( n14269 , n14267 , n14268 );
xor ( n14270 , n14235 , n14269 );
xor ( n14271 , n14191 , n14270 );
xor ( n14272 , n14237 , n14260 );
xor ( n14273 , n14272 , n14266 );
xor ( n14274 , n14242 , n14246 );
xor ( n14275 , n14274 , n14257 );
not ( n14276 , n12555 );
not ( n14277 , n503 );
not ( n14278 , n13459 );
or ( n14279 , n14277 , n14278 );
not ( n14280 , n503 );
nand ( n14281 , n14280 , n14167 );
nand ( n14282 , n14279 , n14281 );
not ( n14283 , n14282 );
or ( n14284 , n14276 , n14283 );
nand ( n14285 , n13970 , n504 );
nand ( n14286 , n14284 , n14285 );
xor ( n14287 , n14275 , n14286 );
not ( n14288 , n13119 );
not ( n14289 , n14073 );
or ( n14290 , n14288 , n14289 );
and ( n14291 , n495 , n13195 );
not ( n14292 , n495 );
and ( n14293 , n14292 , n13687 );
nor ( n14294 , n14291 , n14293 );
nand ( n14295 , n14294 , n13056 );
nand ( n14296 , n14290 , n14295 );
not ( n14297 , n12563 );
not ( n14298 , n14055 );
or ( n14299 , n14297 , n14298 );
not ( n14300 , n497 );
not ( n14301 , n13526 );
or ( n14302 , n14300 , n14301 );
nand ( n14303 , n12812 , n12579 );
nand ( n14304 , n14302 , n14303 );
nand ( n14305 , n14304 , n12610 );
nand ( n14306 , n14299 , n14305 );
xor ( n14307 , n14296 , n14306 );
xor ( n14308 , n13994 , n13996 );
xor ( n14309 , n14308 , n14040 );
and ( n14310 , n14307 , n14309 );
and ( n14311 , n14296 , n14306 );
or ( n14312 , n14310 , n14311 );
not ( n14313 , n12743 );
not ( n14314 , n14253 );
or ( n14315 , n14313 , n14314 );
not ( n14316 , n499 );
not ( n14317 , n12670 );
or ( n14318 , n14316 , n14317 );
nand ( n14319 , n12666 , n12560 );
nand ( n14320 , n14318 , n14319 );
nand ( n14321 , n14320 , n12789 );
nand ( n14322 , n14315 , n14321 );
xor ( n14323 , n14312 , n14322 );
not ( n14324 , n12930 );
not ( n14325 , n14093 );
or ( n14326 , n14324 , n14325 );
and ( n14327 , n12722 , n501 );
not ( n14328 , n12722 );
and ( n14329 , n14328 , n12943 );
or ( n14330 , n14327 , n14329 );
nand ( n14331 , n14330 , n12908 );
nand ( n14332 , n14326 , n14331 );
and ( n14333 , n14323 , n14332 );
and ( n14334 , n14312 , n14322 );
or ( n14335 , n14333 , n14334 );
and ( n14336 , n14287 , n14335 );
and ( n14337 , n14275 , n14286 );
or ( n14338 , n14336 , n14337 );
xor ( n14339 , n14273 , n14338 );
xor ( n14340 , n13964 , n13978 );
xor ( n14341 , n14340 , n14098 );
and ( n14342 , n14339 , n14341 );
and ( n14343 , n14273 , n14338 );
or ( n14344 , n14342 , n14343 );
or ( n14345 , n14271 , n14344 );
not ( n14346 , n14345 );
xor ( n14347 , n14273 , n14338 );
xor ( n14348 , n14347 , n14341 );
xor ( n14349 , n13981 , n14079 );
xor ( n14350 , n14349 , n14095 );
xor ( n14351 , n14043 , n14057 );
xor ( n14352 , n14351 , n14076 );
not ( n14353 , n13119 );
not ( n14354 , n14294 );
or ( n14355 , n14353 , n14354 );
and ( n14356 , n495 , n13519 );
not ( n14357 , n495 );
and ( n14358 , n14357 , n13835 );
nor ( n14359 , n14356 , n14358 );
nand ( n14360 , n14359 , n13056 );
nand ( n14361 , n14355 , n14360 );
xor ( n14362 , n13998 , n14008 );
xor ( n14363 , n14362 , n14037 );
xor ( n14364 , n14361 , n14363 );
not ( n14365 , n12563 );
not ( n14366 , n14304 );
or ( n14367 , n14365 , n14366 );
buf ( n14368 , n12822 );
and ( n14369 , n497 , n14368 );
not ( n14370 , n497 );
and ( n14371 , n14370 , n13805 );
nor ( n14372 , n14369 , n14371 );
nand ( n14373 , n14372 , n12609 );
nand ( n14374 , n14367 , n14373 );
and ( n14375 , n14364 , n14374 );
and ( n14376 , n14361 , n14363 );
or ( n14377 , n14375 , n14376 );
not ( n14378 , n12789 );
and ( n14379 , n499 , n14145 );
not ( n14380 , n499 );
and ( n14381 , n14380 , n12649 );
nor ( n14382 , n14379 , n14381 );
not ( n14383 , n14382 );
or ( n14384 , n14378 , n14383 );
nand ( n14385 , n14320 , n12741 );
nand ( n14386 , n14384 , n14385 );
xor ( n14387 , n14377 , n14386 );
xor ( n14388 , n14296 , n14306 );
xor ( n14389 , n14388 , n14309 );
and ( n14390 , n14387 , n14389 );
and ( n14391 , n14377 , n14386 );
or ( n14392 , n14390 , n14391 );
xor ( n14393 , n14352 , n14392 );
not ( n14394 , n12555 );
not ( n14395 , n503 );
not ( n14396 , n13160 );
or ( n14397 , n14395 , n14396 );
nand ( n14398 , n13161 , n12516 );
nand ( n14399 , n14397 , n14398 );
not ( n14400 , n14399 );
or ( n14401 , n14394 , n14400 );
nand ( n14402 , n14282 , n504 );
nand ( n14403 , n14401 , n14402 );
and ( n14404 , n14393 , n14403 );
and ( n14405 , n14352 , n14392 );
or ( n14406 , n14404 , n14405 );
xor ( n14407 , n14350 , n14406 );
xor ( n14408 , n14275 , n14286 );
xor ( n14409 , n14408 , n14335 );
and ( n14410 , n14407 , n14409 );
and ( n14411 , n14350 , n14406 );
or ( n14412 , n14410 , n14411 );
or ( n14413 , n14348 , n14412 );
not ( n14414 , n14413 );
xor ( n14415 , n14350 , n14406 );
xor ( n14416 , n14415 , n14409 );
not ( n14417 , n14416 );
not ( n14418 , n12908 );
and ( n14419 , n501 , n12699 );
not ( n14420 , n501 );
and ( n14421 , n14420 , n12700 );
nor ( n14422 , n14419 , n14421 );
not ( n14423 , n14422 );
or ( n14424 , n14418 , n14423 );
nand ( n14425 , n14330 , n12930 );
nand ( n14426 , n14424 , n14425 );
not ( n14427 , n13056 );
and ( n14428 , n495 , n13842 );
not ( n14429 , n495 );
and ( n14430 , n14429 , n13845 );
nor ( n14431 , n14428 , n14430 );
not ( n14432 , n14431 );
or ( n14433 , n14427 , n14432 );
nand ( n14434 , n14359 , n13119 );
nand ( n14435 , n14433 , n14434 );
xor ( n14436 , n14010 , n14029 );
xor ( n14437 , n14436 , n14035 );
xor ( n14438 , n14435 , n14437 );
and ( n14439 , n14022 , n14028 );
not ( n14440 , n14022 );
and ( n14441 , n14440 , n14027 );
nor ( n14442 , n14439 , n14441 );
not ( n14443 , n13119 );
not ( n14444 , n14431 );
or ( n14445 , n14443 , n14444 );
not ( n14446 , n495 );
not ( n14447 , n13859 );
or ( n14448 , n14446 , n14447 );
or ( n14449 , n13859 , n495 );
nand ( n14450 , n14448 , n14449 );
nand ( n14451 , n14450 , n13056 );
nand ( n14452 , n14445 , n14451 );
xor ( n14453 , n14442 , n14452 );
nor ( n14454 , n13850 , n12844 );
not ( n14455 , n13119 );
not ( n14456 , n14450 );
or ( n14457 , n14455 , n14456 );
and ( n14458 , n495 , n13871 );
not ( n14459 , n495 );
and ( n14460 , n14459 , n13870 );
nor ( n14461 , n14458 , n14460 );
nand ( n14462 , n14461 , n13056 );
nand ( n14463 , n14457 , n14462 );
xor ( n14464 , n14454 , n14463 );
or ( n14465 , n13851 , n496 );
nand ( n14466 , n14465 , n497 );
and ( n14467 , n13851 , n496 );
nor ( n14468 , n14467 , n3583 );
and ( n14469 , n14466 , n14468 );
not ( n14470 , n13056 );
and ( n14471 , n495 , n13851 );
not ( n14472 , n495 );
and ( n14473 , n14472 , n13850 );
nor ( n14474 , n14471 , n14473 );
not ( n14475 , n14474 );
or ( n14476 , n14470 , n14475 );
nand ( n14477 , n14461 , n13119 );
nand ( n14478 , n14476 , n14477 );
and ( n14479 , n14469 , n14478 );
and ( n14480 , n14464 , n14479 );
and ( n14481 , n14454 , n14463 );
or ( n14482 , n14480 , n14481 );
and ( n14483 , n14453 , n14482 );
and ( n14484 , n14442 , n14452 );
or ( n14485 , n14483 , n14484 );
and ( n14486 , n14438 , n14485 );
and ( n14487 , n14435 , n14437 );
or ( n14488 , n14486 , n14487 );
xor ( n14489 , n14361 , n14363 );
xor ( n14490 , n14489 , n14374 );
xor ( n14491 , n14488 , n14490 );
not ( n14492 , n14382 );
or ( n14493 , n14492 , n12742 );
and ( n14494 , n12624 , n12560 );
not ( n14495 , n12624 );
and ( n14496 , n14495 , n499 );
or ( n14497 , n14494 , n14496 );
nand ( n14498 , n14497 , n12789 );
nand ( n14499 , n14493 , n14498 );
and ( n14500 , n14491 , n14499 );
and ( n14501 , n14488 , n14490 );
or ( n14502 , n14500 , n14501 );
xor ( n14503 , n14426 , n14502 );
not ( n14504 , n12555 );
not ( n14505 , n503 );
not ( n14506 , n12987 );
or ( n14507 , n14505 , n14506 );
nand ( n14508 , n12861 , n12516 );
nand ( n14509 , n14507 , n14508 );
not ( n14510 , n14509 );
or ( n14511 , n14504 , n14510 );
nand ( n14512 , n14399 , n504 );
nand ( n14513 , n14511 , n14512 );
and ( n14514 , n14503 , n14513 );
and ( n14515 , n14426 , n14502 );
or ( n14516 , n14514 , n14515 );
xor ( n14517 , n14312 , n14322 );
xor ( n14518 , n14517 , n14332 );
xor ( n14519 , n14516 , n14518 );
xor ( n14520 , n14352 , n14392 );
xor ( n14521 , n14520 , n14403 );
and ( n14522 , n14519 , n14521 );
and ( n14523 , n14516 , n14518 );
or ( n14524 , n14522 , n14523 );
not ( n14525 , n14524 );
and ( n14526 , n14417 , n14525 );
xor ( n14527 , n14516 , n14518 );
xor ( n14528 , n14527 , n14521 );
xor ( n14529 , n14377 , n14386 );
xor ( n14530 , n14529 , n14389 );
not ( n14531 , n12563 );
not ( n14532 , n14372 );
or ( n14533 , n14531 , n14532 );
and ( n14534 , n497 , n13688 );
not ( n14535 , n497 );
and ( n14536 , n14535 , n13687 );
nor ( n14537 , n14534 , n14536 );
nand ( n14538 , n14537 , n12609 );
nand ( n14539 , n14533 , n14538 );
not ( n14540 , n12741 );
not ( n14541 , n14497 );
or ( n14542 , n14540 , n14541 );
not ( n14543 , n499 );
not ( n14544 , n13526 );
or ( n14545 , n14543 , n14544 );
nand ( n14546 , n12812 , n12560 );
nand ( n14547 , n14545 , n14546 );
nand ( n14548 , n14547 , n12789 );
nand ( n14549 , n14542 , n14548 );
xor ( n14550 , n14539 , n14549 );
xor ( n14551 , n14435 , n14437 );
xor ( n14552 , n14551 , n14485 );
and ( n14553 , n14550 , n14552 );
and ( n14554 , n14539 , n14549 );
or ( n14555 , n14553 , n14554 );
not ( n14556 , n12930 );
not ( n14557 , n14422 );
or ( n14558 , n14556 , n14557 );
not ( n14559 , n501 );
not ( n14560 , n12670 );
or ( n14561 , n14559 , n14560 );
nand ( n14562 , n12666 , n12943 );
nand ( n14563 , n14561 , n14562 );
nand ( n14564 , n14563 , n12909 );
nand ( n14565 , n14558 , n14564 );
xor ( n14566 , n14555 , n14565 );
not ( n14567 , n504 );
not ( n14568 , n14509 );
or ( n14569 , n14567 , n14568 );
not ( n14570 , n503 );
not ( n14571 , n12870 );
or ( n14572 , n14570 , n14571 );
nand ( n14573 , n12550 , n12721 );
nand ( n14574 , n14572 , n14573 );
nand ( n14575 , n14574 , n12555 );
nand ( n14576 , n14569 , n14575 );
and ( n14577 , n14566 , n14576 );
and ( n14578 , n14555 , n14565 );
or ( n14579 , n14577 , n14578 );
xor ( n14580 , n14530 , n14579 );
xor ( n14581 , n14426 , n14502 );
xor ( n14582 , n14581 , n14513 );
and ( n14583 , n14580 , n14582 );
and ( n14584 , n14530 , n14579 );
or ( n14585 , n14583 , n14584 );
nor ( n14586 , n14528 , n14585 );
nor ( n14587 , n14526 , n14586 );
not ( n14588 , n14587 );
xor ( n14589 , n14530 , n14579 );
xor ( n14590 , n14589 , n14582 );
not ( n14591 , n14590 );
xor ( n14592 , n14488 , n14490 );
xor ( n14593 , n14592 , n14499 );
not ( n14594 , n12930 );
not ( n14595 , n14563 );
or ( n14596 , n14594 , n14595 );
and ( n14597 , n501 , n12652 );
not ( n14598 , n501 );
and ( n14599 , n14598 , n12649 );
nor ( n14600 , n14597 , n14599 );
nand ( n14601 , n14600 , n12908 );
nand ( n14602 , n14596 , n14601 );
not ( n14603 , n12609 );
and ( n14604 , n497 , n13519 );
not ( n14605 , n497 );
and ( n14606 , n14605 , n13835 );
nor ( n14607 , n14604 , n14606 );
not ( n14608 , n14607 );
or ( n14609 , n14603 , n14608 );
nand ( n14610 , n14537 , n12563 );
nand ( n14611 , n14609 , n14610 );
xor ( n14612 , n14442 , n14452 );
xor ( n14613 , n14612 , n14482 );
xor ( n14614 , n14611 , n14613 );
not ( n14615 , n12741 );
not ( n14616 , n14547 );
or ( n14617 , n14615 , n14616 );
and ( n14618 , n499 , n13806 );
not ( n14619 , n499 );
and ( n14620 , n14619 , n13599 );
nor ( n14621 , n14618 , n14620 );
nand ( n14622 , n14621 , n12789 );
nand ( n14623 , n14617 , n14622 );
and ( n14624 , n14614 , n14623 );
and ( n14625 , n14611 , n14613 );
or ( n14626 , n14624 , n14625 );
xor ( n14627 , n14602 , n14626 );
not ( n14628 , n504 );
not ( n14629 , n14574 );
or ( n14630 , n14628 , n14629 );
and ( n14631 , n503 , n12699 );
not ( n14632 , n503 );
and ( n14633 , n14632 , n12700 );
nor ( n14634 , n14631 , n14633 );
nand ( n14635 , n14634 , n12555 );
nand ( n14636 , n14630 , n14635 );
and ( n14637 , n14627 , n14636 );
and ( n14638 , n14602 , n14626 );
or ( n14639 , n14637 , n14638 );
xor ( n14640 , n14593 , n14639 );
xor ( n14641 , n14555 , n14565 );
xor ( n14642 , n14641 , n14576 );
and ( n14643 , n14640 , n14642 );
and ( n14644 , n14593 , n14639 );
or ( n14645 , n14643 , n14644 );
not ( n14646 , n14645 );
and ( n14647 , n14591 , n14646 );
xor ( n14648 , n14593 , n14639 );
xor ( n14649 , n14648 , n14642 );
xor ( n14650 , n14539 , n14549 );
xor ( n14651 , n14650 , n14552 );
not ( n14652 , n12563 );
not ( n14653 , n14607 );
or ( n14654 , n14652 , n14653 );
not ( n14655 , n497 );
not ( n14656 , n13845 );
or ( n14657 , n14655 , n14656 );
nand ( n14658 , n13842 , n12579 );
nand ( n14659 , n14657 , n14658 );
nand ( n14660 , n14659 , n12609 );
nand ( n14661 , n14654 , n14660 );
xor ( n14662 , n14454 , n14463 );
xor ( n14663 , n14662 , n14479 );
xor ( n14664 , n14661 , n14663 );
xor ( n14665 , n14469 , n14478 );
not ( n14666 , n12563 );
not ( n14667 , n14659 );
or ( n14668 , n14666 , n14667 );
not ( n14669 , n12579 );
not ( n14670 , n13675 );
or ( n14671 , n14669 , n14670 );
nand ( n14672 , n13859 , n497 );
nand ( n14673 , n14671 , n14672 );
nand ( n14674 , n14673 , n12609 );
nand ( n14675 , n14668 , n14674 );
xor ( n14676 , n14665 , n14675 );
nor ( n14677 , n13850 , n13052 );
not ( n14678 , n12563 );
not ( n14679 , n14673 );
or ( n14680 , n14678 , n14679 );
or ( n14681 , n13871 , n497 );
nand ( n14682 , n13871 , n497 );
nand ( n14683 , n14681 , n14682 );
not ( n14684 , n14683 );
nand ( n14685 , n14684 , n12609 );
nand ( n14686 , n14680 , n14685 );
xor ( n14687 , n14677 , n14686 );
or ( n14688 , n13851 , n498 );
nand ( n14689 , n14688 , n499 );
and ( n14690 , n13851 , n498 );
nor ( n14691 , n14690 , n12579 );
and ( n14692 , n14689 , n14691 );
not ( n14693 , n12609 );
or ( n14694 , n13850 , n497 );
or ( n14695 , n13851 , n12579 );
nand ( n14696 , n14694 , n14695 );
not ( n14697 , n14696 );
or ( n14698 , n14693 , n14697 );
or ( n14699 , n14683 , n12562 );
nand ( n14700 , n14698 , n14699 );
and ( n14701 , n14692 , n14700 );
and ( n14702 , n14687 , n14701 );
and ( n14703 , n14677 , n14686 );
or ( n14704 , n14702 , n14703 );
and ( n14705 , n14676 , n14704 );
and ( n14706 , n14665 , n14675 );
or ( n14707 , n14705 , n14706 );
and ( n14708 , n14664 , n14707 );
and ( n14709 , n14661 , n14663 );
or ( n14710 , n14708 , n14709 );
xor ( n14711 , n14611 , n14613 );
xor ( n14712 , n14711 , n14623 );
xor ( n14713 , n14710 , n14712 );
not ( n14714 , n12909 );
xor ( n14715 , n501 , n12624 );
not ( n14716 , n14715 );
or ( n14717 , n14714 , n14716 );
nand ( n14718 , n14600 , n12930 );
nand ( n14719 , n14717 , n14718 );
and ( n14720 , n14713 , n14719 );
and ( n14721 , n14710 , n14712 );
or ( n14722 , n14720 , n14721 );
xor ( n14723 , n14651 , n14722 );
xor ( n14724 , n14602 , n14626 );
xor ( n14725 , n14724 , n14636 );
and ( n14726 , n14723 , n14725 );
and ( n14727 , n14651 , n14722 );
or ( n14728 , n14726 , n14727 );
nor ( n14729 , n14649 , n14728 );
nor ( n14730 , n14647 , n14729 );
not ( n14731 , n14730 );
not ( n14732 , n12789 );
and ( n14733 , n499 , n13687 );
not ( n14734 , n499 );
and ( n14735 , n14734 , n13195 );
or ( n14736 , n14733 , n14735 );
not ( n14737 , n14736 );
or ( n14738 , n14732 , n14737 );
nand ( n14739 , n14621 , n12741 );
nand ( n14740 , n14738 , n14739 );
xor ( n14741 , n14661 , n14663 );
xor ( n14742 , n14741 , n14707 );
xor ( n14743 , n14740 , n14742 );
not ( n14744 , n12930 );
not ( n14745 , n14715 );
or ( n14746 , n14744 , n14745 );
and ( n14747 , n12908 , n12943 );
and ( n14748 , n12812 , n14747 );
not ( n14749 , n12812 );
not ( n14750 , n12516 );
nor ( n14751 , n14750 , n12900 );
and ( n14752 , n14749 , n14751 );
nor ( n14753 , n14748 , n14752 );
nand ( n14754 , n14746 , n14753 );
and ( n14755 , n14743 , n14754 );
and ( n14756 , n14740 , n14742 );
or ( n14757 , n14755 , n14756 );
not ( n14758 , n504 );
not ( n14759 , n14634 );
or ( n14760 , n14758 , n14759 );
and ( n14761 , n503 , n12666 );
not ( n14762 , n503 );
and ( n14763 , n14762 , n12670 );
nor ( n14764 , n14761 , n14763 );
nand ( n14765 , n14764 , n12555 );
nand ( n14766 , n14760 , n14765 );
xor ( n14767 , n14757 , n14766 );
xor ( n14768 , n14710 , n14712 );
xor ( n14769 , n14768 , n14719 );
and ( n14770 , n14767 , n14769 );
and ( n14771 , n14757 , n14766 );
or ( n14772 , n14770 , n14771 );
not ( n14773 , n14772 );
xor ( n14774 , n14651 , n14722 );
xor ( n14775 , n14774 , n14725 );
not ( n14776 , n14775 );
nand ( n14777 , n14773 , n14776 );
not ( n14778 , n14777 );
xor ( n14779 , n14757 , n14766 );
xor ( n14780 , n14779 , n14769 );
not ( n14781 , n12555 );
not ( n14782 , n503 );
not ( n14783 , n12649 );
or ( n14784 , n14782 , n14783 );
nand ( n14785 , n12652 , n12516 );
nand ( n14786 , n14784 , n14785 );
not ( n14787 , n14786 );
or ( n14788 , n14781 , n14787 );
nand ( n14789 , n14764 , n504 );
nand ( n14790 , n14788 , n14789 );
not ( n14791 , n12741 );
not ( n14792 , n14736 );
or ( n14793 , n14791 , n14792 );
and ( n14794 , n13835 , n1407 );
not ( n14795 , n13835 );
and ( n14796 , n14795 , n499 );
nor ( n14797 , n14794 , n14796 );
nand ( n14798 , n14797 , n12789 );
nand ( n14799 , n14793 , n14798 );
xor ( n14800 , n14665 , n14675 );
xor ( n14801 , n14800 , n14704 );
xor ( n14802 , n14799 , n14801 );
not ( n14803 , n501 );
not ( n14804 , n13526 );
or ( n14805 , n14803 , n14804 );
nand ( n14806 , n12812 , n12943 );
nand ( n14807 , n14805 , n14806 );
not ( n14808 , n14807 );
not ( n14809 , n12930 );
or ( n14810 , n14808 , n14809 );
not ( n14811 , n14368 );
not ( n14812 , n14751 );
not ( n14813 , n14812 );
and ( n14814 , n14811 , n14813 );
not ( n14815 , n13599 );
and ( n14816 , n14815 , n14747 );
nor ( n14817 , n14814 , n14816 );
nand ( n14818 , n14810 , n14817 );
and ( n14819 , n14802 , n14818 );
and ( n14820 , n14799 , n14801 );
or ( n14821 , n14819 , n14820 );
xor ( n14822 , n14790 , n14821 );
xor ( n14823 , n14740 , n14742 );
xor ( n14824 , n14823 , n14754 );
and ( n14825 , n14822 , n14824 );
and ( n14826 , n14790 , n14821 );
or ( n14827 , n14825 , n14826 );
or ( n14828 , n14780 , n14827 );
not ( n14829 , n14828 );
xor ( n14830 , n14692 , n14700 );
not ( n14831 , n12740 );
and ( n14832 , n499 , n13842 );
not ( n14833 , n499 );
and ( n14834 , n14833 , n13845 );
nor ( n14835 , n14832 , n14834 );
not ( n14836 , n14835 );
or ( n14837 , n14831 , n14836 );
not ( n14838 , n499 );
not ( n14839 , n13859 );
or ( n14840 , n14838 , n14839 );
nand ( n14841 , n13675 , n12560 );
nand ( n14842 , n14840 , n14841 );
nand ( n14843 , n14842 , n12789 );
nand ( n14844 , n14837 , n14843 );
xor ( n14845 , n14830 , n14844 );
nor ( n14846 , n13850 , n12562 );
not ( n14847 , n12740 );
not ( n14848 , n14842 );
or ( n14849 , n14847 , n14848 );
and ( n14850 , n499 , n13871 );
not ( n14851 , n499 );
and ( n14852 , n14851 , n13870 );
nor ( n14853 , n14850 , n14852 );
nand ( n14854 , n14853 , n12789 );
nand ( n14855 , n14849 , n14854 );
xor ( n14856 , n14846 , n14855 );
or ( n14857 , n13851 , n500 );
nand ( n14858 , n14857 , n501 );
and ( n14859 , n13851 , n500 );
nor ( n14860 , n14859 , n12560 );
and ( n14861 , n14858 , n14860 );
not ( n14862 , n12740 );
not ( n14863 , n14853 );
or ( n14864 , n14862 , n14863 );
or ( n14865 , n13850 , n499 );
or ( n14866 , n13851 , n12560 );
nand ( n14867 , n14865 , n14866 );
nand ( n14868 , n14867 , n12789 );
nand ( n14869 , n14864 , n14868 );
and ( n14870 , n14861 , n14869 );
and ( n14871 , n14856 , n14870 );
and ( n14872 , n14846 , n14855 );
or ( n14873 , n14871 , n14872 );
and ( n14874 , n14845 , n14873 );
and ( n14875 , n14830 , n14844 );
or ( n14876 , n14874 , n14875 );
not ( n14877 , n12741 );
not ( n14878 , n14797 );
or ( n14879 , n14877 , n14878 );
nand ( n14880 , n14835 , n12789 );
nand ( n14881 , n14879 , n14880 );
xor ( n14882 , n14677 , n14686 );
xor ( n14883 , n14882 , n14701 );
xor ( n14884 , n14881 , n14883 );
not ( n14885 , n12907 );
xor ( n14886 , n501 , n12822 );
not ( n14887 , n14886 );
or ( n14888 , n14885 , n14887 );
and ( n14889 , n501 , n13195 );
not ( n14890 , n501 );
and ( n14891 , n14890 , n13687 );
nor ( n14892 , n14889 , n14891 );
nand ( n14893 , n14892 , n12908 );
nand ( n14894 , n14888 , n14893 );
xor ( n14895 , n14884 , n14894 );
xor ( n14896 , n14876 , n14895 );
not ( n14897 , n699 );
nand ( n14898 , n14897 , n12625 );
nand ( n14899 , n12624 , n4208 );
not ( n14900 , n503 );
not ( n14901 , n13526 );
or ( n14902 , n14900 , n14901 );
or ( n14903 , n13526 , n503 );
nand ( n14904 , n14902 , n14903 );
nand ( n14905 , n14904 , n12555 );
nand ( n14906 , n14898 , n14899 , n14905 );
xor ( n14907 , n14896 , n14906 );
not ( n14908 , n12908 );
or ( n14909 , n13519 , n12943 );
nand ( n14910 , n13519 , n3378 );
nand ( n14911 , n14909 , n14910 );
not ( n14912 , n14911 );
or ( n14913 , n14908 , n14912 );
nand ( n14914 , n14892 , n12907 );
nand ( n14915 , n14913 , n14914 );
xor ( n14916 , n14830 , n14844 );
xor ( n14917 , n14916 , n14873 );
xor ( n14918 , n14915 , n14917 );
not ( n14919 , n12555 );
xor ( n14920 , n503 , n12822 );
not ( n14921 , n14920 );
or ( n14922 , n14919 , n14921 );
nand ( n14923 , n14904 , n504 );
nand ( n14924 , n14922 , n14923 );
and ( n14925 , n14918 , n14924 );
and ( n14926 , n14915 , n14917 );
or ( n14927 , n14925 , n14926 );
or ( n14928 , n14907 , n14927 );
not ( n14929 , n14928 );
not ( n14930 , n12908 );
and ( n14931 , n13587 , n501 );
not ( n14932 , n13587 );
and ( n14933 , n14932 , n12943 );
nor ( n14934 , n14931 , n14933 );
not ( n14935 , n14934 );
or ( n14936 , n14930 , n14935 );
nand ( n14937 , n14911 , n12907 );
nand ( n14938 , n14936 , n14937 );
xor ( n14939 , n14846 , n14855 );
xor ( n14940 , n14939 , n14870 );
xor ( n14941 , n14938 , n14940 );
not ( n14942 , n12555 );
and ( n14943 , n13195 , n12516 );
not ( n14944 , n13195 );
and ( n14945 , n14944 , n503 );
or ( n14946 , n14943 , n14945 );
not ( n14947 , n14946 );
or ( n14948 , n14942 , n14947 );
nand ( n14949 , n14920 , n504 );
nand ( n14950 , n14948 , n14949 );
and ( n14951 , n14941 , n14950 );
and ( n14952 , n14938 , n14940 );
or ( n14953 , n14951 , n14952 );
xor ( n14954 , n14915 , n14917 );
xor ( n14955 , n14954 , n14924 );
xor ( n14956 , n14953 , n14955 );
xor ( n14957 , n14861 , n14869 );
not ( n14958 , n12907 );
not ( n14959 , n14934 );
or ( n14960 , n14958 , n14959 );
not ( n14961 , n501 );
not ( n14962 , n13859 );
or ( n14963 , n14961 , n14962 );
nand ( n14964 , n13675 , n12943 );
nand ( n14965 , n14963 , n14964 );
nand ( n14966 , n14965 , n12908 );
nand ( n14967 , n14960 , n14966 );
xor ( n14968 , n14957 , n14967 );
and ( n14969 , n13851 , n12740 );
and ( n14970 , n13870 , n3378 );
not ( n14971 , n13870 );
and ( n14972 , n14971 , n501 );
nor ( n14973 , n14970 , n14972 );
nand ( n14974 , n14973 , n12907 );
nand ( n14975 , n14747 , n13851 );
nand ( n14976 , n14751 , n13850 );
and ( n14977 , n14974 , n14975 , n14976 );
or ( n14978 , n13851 , n502 );
nand ( n14979 , n14978 , n503 );
and ( n14980 , n13851 , n502 );
nor ( n14981 , n14980 , n12943 );
nand ( n14982 , n14979 , n14981 );
nor ( n14983 , n14977 , n14982 );
xor ( n14984 , n14969 , n14983 );
not ( n14985 , n12907 );
not ( n14986 , n14965 );
or ( n14987 , n14985 , n14986 );
nand ( n14988 , n14973 , n12908 );
nand ( n14989 , n14987 , n14988 );
and ( n14990 , n14984 , n14989 );
or ( n14991 , n14990 , C0 );
and ( n14992 , n14968 , n14991 );
and ( n14993 , n14957 , n14967 );
or ( n14994 , n14992 , n14993 );
xor ( n14995 , n14957 , n14967 );
xor ( n14996 , n14995 , n14991 );
not ( n14997 , n14946 );
not ( n14998 , n504 );
or ( n14999 , n14997 , n14998 );
not ( n15000 , n13519 );
not ( n15001 , n503 );
and ( n15002 , n15000 , n15001 );
and ( n15003 , n13519 , n503 );
nor ( n15004 , n15002 , n15003 );
nand ( n15005 , n15004 , n12555 );
nand ( n15006 , n14999 , n15005 );
or ( n15007 , n14996 , n15006 );
xor ( n15008 , n14969 , n14983 );
xor ( n15009 , n15008 , n14989 );
not ( n15010 , n13587 );
not ( n15011 , n12516 );
or ( n15012 , n15010 , n15011 );
or ( n15013 , n13587 , n12516 );
nand ( n15014 , n15012 , n15013 );
not ( n15015 , n15014 );
not ( n15016 , n12555 );
or ( n15017 , n15015 , n15016 );
not ( n15018 , n15004 );
or ( n15019 , n15018 , n1939 );
nand ( n15020 , n15017 , n15019 );
nor ( n15021 , n15009 , n15020 );
not ( n15022 , n14982 );
nand ( n15023 , n14974 , n14975 , n14976 );
not ( n15024 , n15023 );
or ( n15025 , n15022 , n15024 );
or ( n15026 , n15023 , n14982 );
nand ( n15027 , n15025 , n15026 );
not ( n15028 , n504 );
not ( n15029 , n15014 );
or ( n15030 , n15028 , n15029 );
not ( n15031 , n13675 );
not ( n15032 , n503 );
and ( n15033 , n15031 , n15032 );
and ( n15034 , n13675 , n503 );
nor ( n15035 , n15033 , n15034 );
nand ( n15036 , n15035 , n12555 );
nand ( n15037 , n15030 , n15036 );
xor ( n15038 , n15027 , n15037 );
not ( n15039 , n504 );
or ( n15040 , n13871 , n12516 , n15039 );
nor ( n15041 , n503 , n15039 );
and ( n15042 , n13871 , n15041 );
and ( n15043 , n12555 , n13850 );
nor ( n15044 , n15042 , n15043 );
nand ( n15045 , n15040 , n15044 );
not ( n15046 , n504 );
nor ( n15047 , n15046 , n13850 );
nor ( n15048 , n15047 , n12516 );
nand ( n15049 , n15045 , n15048 );
not ( n15050 , n15049 );
not ( n15051 , n12907 );
nor ( n15052 , n15051 , n13850 );
nor ( n15053 , n15050 , n15052 );
not ( n15054 , n503 );
not ( n15055 , n13871 );
or ( n15056 , n15054 , n15055 );
or ( n15057 , n13871 , n503 );
nand ( n15058 , n15056 , n15057 );
not ( n15059 , n15058 );
not ( n15060 , n12554 );
and ( n15061 , n15059 , n15060 );
and ( n15062 , n15035 , n504 );
nor ( n15063 , n15061 , n15062 );
or ( n15064 , n15053 , n15063 );
nand ( n15065 , n15064 , C1 );
and ( n15066 , n15038 , n15065 );
and ( n15067 , n15027 , n15037 );
or ( n15068 , n15066 , n15067 );
not ( n15069 , n15068 );
or ( n15070 , n15021 , n15069 );
nand ( n15071 , n15020 , n15009 );
nand ( n15072 , n15070 , n15071 );
nand ( n15073 , n15007 , n15072 );
nand ( n15074 , n14996 , n15006 );
nand ( n15075 , n15073 , n15074 );
xor ( n15076 , n14994 , n15075 );
xor ( n15077 , n14938 , n14940 );
xor ( n15078 , n15077 , n14950 );
and ( n15079 , n15076 , n15078 );
and ( n15080 , n14994 , n15075 );
or ( n15081 , n15079 , n15080 );
and ( n15082 , n14956 , n15081 );
and ( n15083 , n14953 , n14955 );
or ( n15084 , n15082 , n15083 );
not ( n15085 , n15084 );
or ( n15086 , n14929 , n15085 );
nand ( n15087 , n14907 , n14927 );
nand ( n15088 , n15086 , n15087 );
not ( n15089 , n15088 );
xor ( n15090 , n14881 , n14883 );
and ( n15091 , n15090 , n14894 );
and ( n15092 , n14881 , n14883 );
or ( n15093 , n15091 , n15092 );
xor ( n15094 , n14799 , n14801 );
xor ( n15095 , n15094 , n14818 );
xor ( n15096 , n15093 , n15095 );
not ( n15097 , n504 );
not ( n15098 , n14786 );
or ( n15099 , n15097 , n15098 );
nand ( n15100 , n12625 , n12555 );
nand ( n15101 , n15099 , n15100 );
xor ( n15102 , n15096 , n15101 );
not ( n15103 , n15102 );
xor ( n15104 , n14876 , n14895 );
and ( n15105 , n15104 , n14906 );
and ( n15106 , n14876 , n14895 );
or ( n15107 , n15105 , n15106 );
not ( n15108 , n15107 );
nand ( n15109 , n15103 , n15108 );
not ( n15110 , n15109 );
or ( n15111 , n15089 , n15110 );
nand ( n15112 , n15102 , n15107 );
nand ( n15113 , n15111 , n15112 );
not ( n15114 , n15113 );
xor ( n15115 , n14790 , n14821 );
xor ( n15116 , n15115 , n14824 );
not ( n15117 , n15116 );
xor ( n15118 , n15093 , n15095 );
and ( n15119 , n15118 , n15101 );
and ( n15120 , n15093 , n15095 );
or ( n15121 , n15119 , n15120 );
not ( n15122 , n15121 );
nand ( n15123 , n15117 , n15122 );
not ( n15124 , n15123 );
or ( n15125 , n15114 , n15124 );
nand ( n15126 , n15116 , n15121 );
nand ( n15127 , n15125 , n15126 );
not ( n15128 , n15127 );
or ( n15129 , n14829 , n15128 );
nand ( n15130 , n14780 , n14827 );
nand ( n15131 , n15129 , n15130 );
not ( n15132 , n15131 );
or ( n15133 , n14778 , n15132 );
nand ( n15134 , n14775 , n14772 );
nand ( n15135 , n15133 , n15134 );
not ( n15136 , n15135 );
or ( n15137 , n14731 , n15136 );
or ( n15138 , n14645 , n14590 );
and ( n15139 , n14649 , n14728 );
and ( n15140 , n15138 , n15139 );
and ( n15141 , n14590 , n14645 );
nor ( n15142 , n15140 , n15141 );
nand ( n15143 , n15137 , n15142 );
not ( n15144 , n15143 );
or ( n15145 , n14588 , n15144 );
not ( n15146 , n14416 );
not ( n15147 , n14524 );
nand ( n15148 , n15146 , n15147 );
nand ( n15149 , n14528 , n14585 );
not ( n15150 , n15149 );
and ( n15151 , n15148 , n15150 );
nand ( n15152 , n14416 , n14524 );
not ( n15153 , n15152 );
nor ( n15154 , n15151 , n15153 );
nand ( n15155 , n15145 , n15154 );
not ( n15156 , n15155 );
or ( n15157 , n14414 , n15156 );
nand ( n15158 , n14348 , n14412 );
nand ( n15159 , n15157 , n15158 );
not ( n15160 , n15159 );
or ( n15161 , n14346 , n15160 );
nand ( n15162 , n14344 , n14271 );
nand ( n15163 , n15161 , n15162 );
not ( n15164 , n15163 );
xor ( n15165 , n14199 , n14204 );
and ( n15166 , n15165 , n14207 );
and ( n15167 , n14199 , n14204 );
or ( n15168 , n15166 , n15167 );
not ( n15169 , n13119 );
not ( n15170 , n13656 );
not ( n15171 , n15170 );
or ( n15172 , n15169 , n15171 );
nand ( n15173 , n14137 , n13056 );
nand ( n15174 , n15172 , n15173 );
xor ( n15175 , n15168 , n15174 );
not ( n15176 , n14159 );
not ( n15177 , n12610 );
or ( n15178 , n15176 , n15177 );
not ( n15179 , n13661 );
nand ( n15180 , n15179 , n12563 );
nand ( n15181 , n15178 , n15180 );
and ( n15182 , n15175 , n15181 );
and ( n15183 , n15168 , n15174 );
or ( n15184 , n15182 , n15183 );
xor ( n15185 , n13660 , n13664 );
xor ( n15186 , n15185 , n13713 );
xor ( n15187 , n15184 , n15186 );
xor ( n15188 , n13697 , n13707 );
xor ( n15189 , n15188 , n13710 );
not ( n15190 , n12743 );
not ( n15191 , n499 );
not ( n15192 , n13459 );
or ( n15193 , n15191 , n15192 );
not ( n15194 , n499 );
nand ( n15195 , n15194 , n14167 );
nand ( n15196 , n15193 , n15195 );
not ( n15197 , n15196 );
or ( n15198 , n15190 , n15197 );
nand ( n15199 , n12789 , n14215 );
nand ( n15200 , n15198 , n15199 );
xor ( n15201 , n15189 , n15200 );
xor ( n15202 , n14132 , n14149 );
and ( n15203 , n15202 , n14161 );
and ( n15204 , n14132 , n14149 );
or ( n15205 , n15203 , n15204 );
and ( n15206 , n15201 , n15205 );
and ( n15207 , n15189 , n15200 );
or ( n15208 , n15206 , n15207 );
xor ( n15209 , n15187 , n15208 );
not ( n15210 , n12555 );
not ( n15211 , n14185 );
or ( n15212 , n15210 , n15211 );
not ( n15213 , n503 );
not ( n15214 , n13559 );
or ( n15215 , n15213 , n15214 );
nand ( n15216 , n13558 , n12550 );
nand ( n15217 , n15215 , n15216 );
nand ( n15218 , n15217 , n504 );
nand ( n15219 , n15212 , n15218 );
xor ( n15220 , n15189 , n15200 );
xor ( n15221 , n15220 , n15205 );
xor ( n15222 , n15219 , n15221 );
xor ( n15223 , n14162 , n14178 );
and ( n15224 , n15223 , n14189 );
and ( n15225 , n14162 , n14178 );
or ( n15226 , n15224 , n15225 );
and ( n15227 , n15222 , n15226 );
and ( n15228 , n15219 , n15221 );
or ( n15229 , n15227 , n15228 );
xor ( n15230 , n15209 , n15229 );
not ( n15231 , n12555 );
not ( n15232 , n15217 );
or ( n15233 , n15231 , n15232 );
nand ( n15234 , n13787 , n504 );
nand ( n15235 , n15233 , n15234 );
xor ( n15236 , n14208 , n14217 );
and ( n15237 , n15236 , n14233 );
and ( n15238 , n14208 , n14217 );
or ( n15239 , n15237 , n15238 );
xor ( n15240 , n15168 , n15174 );
xor ( n15241 , n15240 , n15181 );
xor ( n15242 , n15239 , n15241 );
not ( n15243 , n14176 );
not ( n15244 , n12909 );
or ( n15245 , n15243 , n15244 );
not ( n15246 , n501 );
not ( n15247 , n12599 );
or ( n15248 , n15246 , n15247 );
nand ( n15249 , n12602 , n12943 );
nand ( n15250 , n15248 , n15249 );
not ( n15251 , n15250 );
not ( n15252 , n12930 );
or ( n15253 , n15251 , n15252 );
nand ( n15254 , n15245 , n15253 );
and ( n15255 , n15242 , n15254 );
and ( n15256 , n15239 , n15241 );
or ( n15257 , n15255 , n15256 );
xor ( n15258 , n15235 , n15257 );
xor ( n15259 , n13610 , n13618 );
xor ( n15260 , n15259 , n13621 );
not ( n15261 , n12789 );
not ( n15262 , n15196 );
or ( n15263 , n15261 , n15262 );
nand ( n15264 , n13643 , n12743 );
nand ( n15265 , n15263 , n15264 );
xor ( n15266 , n15260 , n15265 );
not ( n15267 , n12909 );
not ( n15268 , n15250 );
or ( n15269 , n15267 , n15268 );
nand ( n15270 , n13776 , n12930 );
nand ( n15271 , n15269 , n15270 );
xor ( n15272 , n15266 , n15271 );
xor ( n15273 , n15258 , n15272 );
xor ( n15274 , n15230 , n15273 );
xor ( n15275 , n15239 , n15241 );
xor ( n15276 , n15275 , n15254 );
xor ( n15277 , n14195 , n14234 );
and ( n15278 , n15277 , n14269 );
and ( n15279 , n14195 , n14234 );
or ( n15280 , n15278 , n15279 );
xor ( n15281 , n15276 , n15280 );
xor ( n15282 , n15219 , n15221 );
xor ( n15283 , n15282 , n15226 );
and ( n15284 , n15281 , n15283 );
and ( n15285 , n15276 , n15280 );
or ( n15286 , n15284 , n15285 );
nor ( n15287 , n15274 , n15286 );
xor ( n15288 , n15276 , n15280 );
xor ( n15289 , n15288 , n15283 );
xor ( n15290 , n14101 , n14190 );
and ( n15291 , n15290 , n14270 );
and ( n15292 , n14101 , n14190 );
or ( n15293 , n15291 , n15292 );
nor ( n15294 , n15289 , n15293 );
nor ( n15295 , n15287 , n15294 );
not ( n15296 , n15295 );
or ( n15297 , n15164 , n15296 );
not ( n15298 , n15287 );
nand ( n15299 , n15289 , n15293 );
not ( n15300 , n15299 );
and ( n15301 , n15298 , n15300 );
and ( n15302 , n15274 , n15286 );
nor ( n15303 , n15301 , n15302 );
nand ( n15304 , n15297 , n15303 );
xor ( n15305 , n15235 , n15257 );
and ( n15306 , n15305 , n15272 );
and ( n15307 , n15235 , n15257 );
or ( n15308 , n15306 , n15307 );
xor ( n15309 , n13767 , n13778 );
xor ( n15310 , n15309 , n13789 );
xor ( n15311 , n15308 , n15310 );
xor ( n15312 , n15260 , n15265 );
and ( n15313 , n15312 , n15271 );
and ( n15314 , n15260 , n15265 );
or ( n15315 , n15313 , n15314 );
xor ( n15316 , n13649 , n13651 );
xor ( n15317 , n15316 , n13716 );
xor ( n15318 , n15315 , n15317 );
xor ( n15319 , n15184 , n15186 );
and ( n15320 , n15319 , n15208 );
and ( n15321 , n15184 , n15186 );
or ( n15322 , n15320 , n15321 );
xor ( n15323 , n15318 , n15322 );
and ( n15324 , n15311 , n15323 );
and ( n15325 , n15308 , n15310 );
or ( n15326 , n15324 , n15325 );
xor ( n15327 , n13638 , n13719 );
xor ( n15328 , n15327 , n13736 );
xor ( n15329 , n15315 , n15317 );
and ( n15330 , n15329 , n15322 );
and ( n15331 , n15315 , n15317 );
or ( n15332 , n15330 , n15331 );
xor ( n15333 , n15328 , n15332 );
xor ( n15334 , n13762 , n13764 );
xor ( n15335 , n15334 , n13792 );
xor ( n15336 , n15333 , n15335 );
nor ( n15337 , n15326 , n15336 );
xor ( n15338 , n15308 , n15310 );
xor ( n15339 , n15338 , n15323 );
xor ( n15340 , n15209 , n15229 );
and ( n15341 , n15340 , n15273 );
and ( n15342 , n15209 , n15229 );
or ( n15343 , n15341 , n15342 );
nor ( n15344 , n15339 , n15343 );
nor ( n15345 , n15337 , n15344 );
xor ( n15346 , n13760 , n13795 );
xor ( n15347 , n15346 , n13798 );
xor ( n15348 , n15328 , n15332 );
and ( n15349 , n15348 , n15335 );
and ( n15350 , n15328 , n15332 );
or ( n15351 , n15349 , n15350 );
nor ( n15352 , n15347 , n15351 );
not ( n15353 , n15352 );
and ( n15354 , n13803 , n15304 , n15345 , n15353 );
nand ( n15355 , n15339 , n15343 );
or ( n15356 , n15337 , n15355 );
nand ( n15357 , n15326 , n15336 );
nand ( n15358 , n15356 , n15357 );
not ( n15359 , n15358 );
nor ( n15360 , n13802 , n15352 );
not ( n15361 , n15360 );
or ( n15362 , n15359 , n15361 );
not ( n15363 , n13802 );
nand ( n15364 , n15347 , n15351 );
not ( n15365 , n15364 );
and ( n15366 , n15363 , n15365 );
and ( n15367 , n13758 , n13801 );
nor ( n15368 , n15366 , n15367 );
nand ( n15369 , n15362 , n15368 );
or ( n15370 , n15354 , n15369 );
nand ( n15371 , n13418 , n13498 );
not ( n15372 , n13501 );
not ( n15373 , n13751 );
nand ( n15374 , n15372 , n15373 );
and ( n15375 , n15371 , n15374 );
nand ( n15376 , n15370 , n15375 );
not ( n15377 , n15376 );
or ( n15378 , n13756 , n15377 );
not ( n15379 , n12845 );
and ( n15380 , n493 , n12602 );
not ( n15381 , n493 );
and ( n15382 , n15381 , n12599 );
nor ( n15383 , n15380 , n15382 );
not ( n15384 , n15383 );
or ( n15385 , n15379 , n15384 );
buf ( n15386 , n12878 );
nand ( n15387 , n13352 , n15386 );
nand ( n15388 , n15385 , n15387 );
xor ( n15389 , n13393 , n13394 );
and ( n15390 , n15389 , n13407 );
and ( n15391 , n13393 , n13394 );
or ( n15392 , n15390 , n15391 );
xor ( n15393 , n15388 , n15392 );
and ( n15394 , n495 , n13559 );
not ( n15395 , n495 );
and ( n15396 , n15395 , n13558 );
or ( n15397 , n15394 , n15396 );
not ( n15398 , n15397 );
not ( n15399 , n13119 );
or ( n15400 , n15398 , n15399 );
nand ( n15401 , n13361 , n13056 );
nand ( n15402 , n15400 , n15401 );
xor ( n15403 , n15393 , n15402 );
xor ( n15404 , n13384 , n13408 );
and ( n15405 , n15404 , n13413 );
and ( n15406 , n13384 , n13408 );
or ( n15407 , n15405 , n15406 );
xor ( n15408 , n15403 , n15407 );
xor ( n15409 , n13249 , n13258 );
and ( n15410 , n15409 , n13343 );
and ( n15411 , n13249 , n13258 );
or ( n15412 , n15410 , n15411 );
and ( n15413 , n15408 , n15412 );
and ( n15414 , n15403 , n15407 );
or ( n15415 , n15413 , n15414 );
not ( n15416 , n12789 );
not ( n15417 , n13256 );
or ( n15418 , n15416 , n15417 );
not ( n15419 , n499 );
not ( n15420 , n12973 );
or ( n15421 , n15419 , n15420 );
nand ( n15422 , n13453 , n12560 );
nand ( n15423 , n15421 , n15422 );
nand ( n15424 , n15423 , n12743 );
nand ( n15425 , n15418 , n15424 );
not ( n15426 , n12563 );
not ( n15427 , n497 );
not ( n15428 , n12923 );
or ( n15429 , n15427 , n15428 );
nand ( n15430 , n13725 , n12579 );
nand ( n15431 , n15429 , n15430 );
not ( n15432 , n15431 );
or ( n15433 , n15426 , n15432 );
nand ( n15434 , n13382 , n12610 );
nand ( n15435 , n15433 , n15434 );
xor ( n15436 , n15425 , n15435 );
and ( n15437 , n13405 , n13406 );
not ( n15438 , n12731 );
not ( n15439 , n491 );
not ( n15440 , n13068 );
or ( n15441 , n15439 , n15440 );
not ( n15442 , n491 );
nand ( n15443 , n15442 , n13067 );
nand ( n15444 , n15441 , n15443 );
not ( n15445 , n15444 );
or ( n15446 , n15438 , n15445 );
nand ( n15447 , n13388 , n12688 );
nand ( n15448 , n15446 , n15447 );
xor ( n15449 , n15437 , n15448 );
nand ( n15450 , n12699 , n489 );
not ( n15451 , n15450 );
not ( n15452 , n15451 );
not ( n15453 , n12882 );
not ( n15454 , n489 );
not ( n15455 , n12987 );
or ( n15456 , n15454 , n15455 );
nand ( n15457 , n12861 , n12653 );
nand ( n15458 , n15456 , n15457 );
not ( n15459 , n15458 );
or ( n15460 , n15453 , n15459 );
nand ( n15461 , n13403 , n12635 );
nand ( n15462 , n15460 , n15461 );
not ( n15463 , n15462 );
not ( n15464 , n15463 );
or ( n15465 , n15452 , n15464 );
or ( n15466 , n15463 , n15451 );
nand ( n15467 , n15465 , n15466 );
xor ( n15468 , n15449 , n15467 );
xor ( n15469 , n15436 , n15468 );
not ( n15470 , n12907 );
not ( n15471 , n501 );
not ( n15472 , n12512 );
or ( n15473 , n15471 , n15472 );
not ( n15474 , n12511 );
not ( n15475 , n15474 );
nand ( n15476 , n15475 , n12943 );
nand ( n15477 , n15473 , n15476 );
not ( n15478 , n15477 );
or ( n15479 , n15470 , n15478 );
nand ( n15480 , n13247 , n12909 );
nand ( n15481 , n15479 , n15480 );
xor ( n15482 , n13354 , n13363 );
and ( n15483 , n15482 , n13368 );
and ( n15484 , n13354 , n13363 );
or ( n15485 , n15483 , n15484 );
xor ( n15486 , n15481 , n15485 );
not ( n15487 , n12555 );
not ( n15488 , n13341 );
or ( n15489 , n15487 , n15488 );
not ( n15490 , n503 );
not ( n15491 , n13329 );
xor ( n15492 , n13284 , n13288 );
and ( n15493 , n15492 , n13316 );
and ( n15494 , n13284 , n13288 );
or ( n15495 , n15493 , n15494 );
not ( n15496 , n15495 );
xor ( n15497 , n13295 , n13310 );
and ( n15498 , n15497 , n13315 );
and ( n15499 , n13295 , n13310 );
or ( n15500 , n15498 , n15499 );
not ( n15501 , n15500 );
nand ( n15502 , n525 , n457 );
not ( n15503 , n13307 );
not ( n15504 , n10216 );
or ( n15505 , n15503 , n15504 );
not ( n15506 , n459 );
nor ( n15507 , n15506 , n521 );
not ( n15508 , n521 );
nor ( n15509 , n15508 , n459 );
nor ( n15510 , n15507 , n15509 );
not ( n15511 , n15510 );
nand ( n15512 , n15511 , n10223 );
nand ( n15513 , n15505 , n15512 );
xor ( n15514 , n15502 , n15513 );
and ( n15515 , n462 , n463 );
not ( n15516 , n462 );
and ( n15517 , n15516 , n2650 );
nor ( n15518 , n15515 , n15517 );
or ( n15519 , n10307 , n15518 );
not ( n15520 , n10317 );
nand ( n15521 , n15519 , n15520 );
nand ( n15522 , n15521 , n461 );
xor ( n15523 , n15514 , n15522 );
not ( n15524 , n15523 );
not ( n15525 , n13300 );
not ( n15526 , n10256 );
or ( n15527 , n15525 , n15526 );
xor ( n15528 , n457 , n523 );
nand ( n15529 , n10197 , n15528 );
nand ( n15530 , n15527 , n15529 );
xor ( n15531 , n13294 , n15530 );
xor ( n15532 , n13296 , n13302 );
and ( n15533 , n15532 , n13309 );
and ( n15534 , n13296 , n13302 );
or ( n15535 , n15533 , n15534 );
xor ( n15536 , n15531 , n15535 );
not ( n15537 , n15536 );
or ( n15538 , n15524 , n15537 );
or ( n15539 , n15536 , n15523 );
nand ( n15540 , n15538 , n15539 );
not ( n15541 , n15540 );
or ( n15542 , n15501 , n15541 );
or ( n15543 , n15540 , n15500 );
nand ( n15544 , n15542 , n15543 );
nand ( n15545 , n15496 , n15544 );
not ( n15546 , n15545 );
not ( n15547 , n15546 );
not ( n15548 , n15544 );
nand ( n15549 , n15548 , n15495 );
nand ( n15550 , n15547 , n15549 );
nor ( n15551 , n15491 , n15550 );
not ( n15552 , n15551 );
nand ( n15553 , n12427 , n12423 , n12503 );
nor ( n15554 , n13276 , n15553 );
not ( n15555 , n15554 );
nand ( n15556 , n12755 , n12409 );
not ( n15557 , n15556 );
or ( n15558 , n15555 , n15557 );
not ( n15559 , n13265 );
not ( n15560 , n15559 );
not ( n15561 , n10809 );
or ( n15562 , n15560 , n15561 );
nand ( n15563 , n15562 , n12503 );
not ( n15564 , n15563 );
and ( n15565 , n15564 , n13275 );
nor ( n15566 , n15565 , n13327 );
nand ( n15567 , n15558 , n15566 );
not ( n15568 , n15567 );
or ( n15569 , n15552 , n15568 );
not ( n15570 , n13329 );
not ( n15571 , n15567 );
or ( n15572 , n15570 , n15571 );
nand ( n15573 , n15572 , n15550 );
nand ( n15574 , n15569 , n15573 );
buf ( n15575 , n15574 );
not ( n15576 , n15575 );
not ( n15577 , n15576 );
or ( n15578 , n15490 , n15577 );
not ( n15579 , n15574 );
not ( n15580 , n15579 );
nand ( n15581 , n15580 , n12516 );
nand ( n15582 , n15578 , n15581 );
nand ( n15583 , n15582 , n504 );
nand ( n15584 , n15489 , n15583 );
xor ( n15585 , n15486 , n15584 );
xor ( n15586 , n15469 , n15585 );
xor ( n15587 , n13369 , n13373 );
and ( n15588 , n15587 , n13414 );
and ( n15589 , n13369 , n13373 );
or ( n15590 , n15588 , n15589 );
and ( n15591 , n15586 , n15590 );
and ( n15592 , n15469 , n15585 );
or ( n15593 , n15591 , n15592 );
xor ( n15594 , n15415 , n15593 );
not ( n15595 , n12789 );
not ( n15596 , n15423 );
or ( n15597 , n15595 , n15596 );
not ( n15598 , n499 );
not ( n15599 , n12545 );
not ( n15600 , n15599 );
or ( n15601 , n15598 , n15600 );
buf ( n15602 , n12545 );
nand ( n15603 , n15602 , n12560 );
nand ( n15604 , n15601 , n15603 );
nand ( n15605 , n15604 , n12743 );
nand ( n15606 , n15597 , n15605 );
not ( n15607 , n12563 );
nand ( n15608 , n13450 , n12579 );
nand ( n15609 , n13451 , n497 );
nand ( n15610 , n15608 , n15609 );
not ( n15611 , n15610 );
or ( n15612 , n15607 , n15611 );
nand ( n15613 , n15431 , n12610 );
nand ( n15614 , n15612 , n15613 );
xor ( n15615 , n15606 , n15614 );
not ( n15616 , n15444 );
not ( n15617 , n12688 );
or ( n15618 , n15616 , n15617 );
not ( n15619 , n491 );
not ( n15620 , n13096 );
or ( n15621 , n15619 , n15620 );
or ( n15622 , n13096 , n491 );
nand ( n15623 , n15621 , n15622 );
nand ( n15624 , n15623 , n12731 );
nand ( n15625 , n15618 , n15624 );
not ( n15626 , n15462 );
nor ( n15627 , n15626 , n15450 );
xor ( n15628 , n15625 , n15627 );
not ( n15629 , n12722 );
and ( n15630 , n15629 , n489 );
not ( n15631 , n12635 );
not ( n15632 , n15458 );
or ( n15633 , n15631 , n15632 );
not ( n15634 , n489 );
not ( n15635 , n13160 );
or ( n15636 , n15634 , n15635 );
nand ( n15637 , n13036 , n12653 );
nand ( n15638 , n15636 , n15637 );
nand ( n15639 , n15638 , n12882 );
nand ( n15640 , n15633 , n15639 );
xor ( n15641 , n15630 , n15640 );
xor ( n15642 , n15628 , n15641 );
xor ( n15643 , n15615 , n15642 );
not ( n15644 , n12909 );
not ( n15645 , n15477 );
or ( n15646 , n15644 , n15645 );
not ( n15647 , n501 );
not ( n15648 , n13336 );
or ( n15649 , n15647 , n15648 );
nand ( n15650 , n13339 , n12943 );
nand ( n15651 , n15649 , n15650 );
nand ( n15652 , n15651 , n12930 );
nand ( n15653 , n15646 , n15652 );
not ( n15654 , n12555 );
not ( n15655 , n15582 );
or ( n15656 , n15654 , n15655 );
not ( n15657 , n15523 );
not ( n15658 , n15657 );
not ( n15659 , n15536 );
or ( n15660 , n15658 , n15659 );
not ( n15661 , n15536 );
nand ( n15662 , n15661 , n15523 );
nand ( n15663 , n15500 , n15662 );
nand ( n15664 , n15660 , n15663 );
not ( n15665 , n15502 );
or ( n15666 , n15513 , n15665 );
nand ( n15667 , n15666 , n15522 );
nand ( n15668 , n15513 , n15665 );
nand ( n15669 , n15667 , n15668 );
and ( n15670 , n457 , n524 );
not ( n15671 , n15528 );
not ( n15672 , n10256 );
or ( n15673 , n15671 , n15672 );
xnor ( n15674 , n457 , n522 );
not ( n15675 , n15674 );
nand ( n15676 , n15675 , n10197 );
nand ( n15677 , n15673 , n15676 );
xor ( n15678 , n15670 , n15677 );
not ( n15679 , n10215 );
not ( n15680 , n15510 );
and ( n15681 , n15679 , n15680 );
and ( n15682 , n10223 , n459 );
nor ( n15683 , n15681 , n15682 );
xor ( n15684 , n15678 , n15683 );
xor ( n15685 , n15669 , n15684 );
xor ( n15686 , n13294 , n15530 );
and ( n15687 , n15686 , n15535 );
and ( n15688 , n13294 , n15530 );
or ( n15689 , n15687 , n15688 );
xor ( n15690 , n15685 , n15689 );
or ( n15691 , n15664 , n15690 );
nand ( n15692 , n15664 , n15690 );
nand ( n15693 , n15691 , n15692 );
not ( n15694 , n15693 );
not ( n15695 , n15694 );
not ( n15696 , n12533 );
not ( n15697 , n13267 );
or ( n15698 , n15696 , n15697 );
buf ( n15699 , n13275 );
nand ( n15700 , n15698 , n15699 );
nor ( n15701 , n13326 , n13317 );
nor ( n15702 , n15546 , n15701 );
buf ( n15703 , n15702 );
nand ( n15704 , n15700 , n15703 );
and ( n15705 , n13274 , n15702 );
not ( n15706 , n15545 );
not ( n15707 , n13329 );
not ( n15708 , n15707 );
or ( n15709 , n15706 , n15708 );
nand ( n15710 , n15709 , n15549 );
nor ( n15711 , n15705 , n15710 );
nand ( n15712 , n15704 , n15711 );
not ( n15713 , n15712 );
not ( n15714 , n15713 );
or ( n15715 , n15695 , n15714 );
not ( n15716 , n15711 );
not ( n15717 , n15704 );
or ( n15718 , n15716 , n15717 );
nand ( n15719 , n15718 , n15693 );
nand ( n15720 , n15715 , n15719 );
and ( n15721 , n12550 , n15720 );
not ( n15722 , n12550 );
not ( n15723 , n15694 );
not ( n15724 , n15713 );
or ( n15725 , n15723 , n15724 );
nand ( n15726 , n15725 , n15719 );
not ( n15727 , n15726 );
and ( n15728 , n15722 , n15727 );
nor ( n15729 , n15721 , n15728 );
not ( n15730 , n15729 );
nand ( n15731 , n15730 , n504 );
nand ( n15732 , n15656 , n15731 );
xor ( n15733 , n15653 , n15732 );
xor ( n15734 , n15388 , n15392 );
and ( n15735 , n15734 , n15402 );
and ( n15736 , n15388 , n15392 );
or ( n15737 , n15735 , n15736 );
xor ( n15738 , n15733 , n15737 );
xor ( n15739 , n15643 , n15738 );
not ( n15740 , n15386 );
not ( n15741 , n15383 );
or ( n15742 , n15740 , n15741 );
and ( n15743 , n12575 , n493 );
not ( n15744 , n12575 );
and ( n15745 , n15744 , n12862 );
or ( n15746 , n15743 , n15745 );
nand ( n15747 , n15746 , n12845 );
nand ( n15748 , n15742 , n15747 );
xor ( n15749 , n15437 , n15448 );
and ( n15750 , n15749 , n15467 );
and ( n15751 , n15437 , n15448 );
or ( n15752 , n15750 , n15751 );
xor ( n15753 , n15748 , n15752 );
not ( n15754 , n13056 );
not ( n15755 , n15397 );
or ( n15756 , n15754 , n15755 );
not ( n15757 , n495 );
not ( n15758 , n12761 );
or ( n15759 , n15757 , n15758 );
not ( n15760 , n495 );
nand ( n15761 , n15760 , n12764 );
nand ( n15762 , n15759 , n15761 );
nand ( n15763 , n15762 , n13119 );
nand ( n15764 , n15756 , n15763 );
xor ( n15765 , n15753 , n15764 );
xor ( n15766 , n15425 , n15435 );
and ( n15767 , n15766 , n15468 );
and ( n15768 , n15425 , n15435 );
or ( n15769 , n15767 , n15768 );
xor ( n15770 , n15765 , n15769 );
xor ( n15771 , n15481 , n15485 );
and ( n15772 , n15771 , n15584 );
and ( n15773 , n15481 , n15485 );
or ( n15774 , n15772 , n15773 );
xor ( n15775 , n15770 , n15774 );
xor ( n15776 , n15739 , n15775 );
xor ( n15777 , n15594 , n15776 );
not ( n15778 , n15777 );
xor ( n15779 , n15403 , n15407 );
xor ( n15780 , n15779 , n15412 );
xor ( n15781 , n15469 , n15585 );
xor ( n15782 , n15781 , n15590 );
xor ( n15783 , n15780 , n15782 );
xor ( n15784 , n13239 , n13344 );
and ( n15785 , n15784 , n13415 );
and ( n15786 , n13239 , n13344 );
or ( n15787 , n15785 , n15786 );
and ( n15788 , n15783 , n15787 );
and ( n15789 , n15780 , n15782 );
or ( n15790 , n15788 , n15789 );
not ( n15791 , n15790 );
and ( n15792 , n15778 , n15791 );
xor ( n15793 , n15780 , n15782 );
xor ( n15794 , n15793 , n15787 );
xor ( n15795 , n12983 , n13234 );
and ( n15796 , n15795 , n13416 );
and ( n15797 , n12983 , n13234 );
or ( n15798 , n15796 , n15797 );
nor ( n15799 , n15794 , n15798 );
nor ( n15800 , n15792 , n15799 );
nand ( n15801 , n15378 , n15800 );
or ( n15802 , n15777 , n15790 );
nand ( n15803 , n15794 , n15798 );
not ( n15804 , n15803 );
and ( n15805 , n15802 , n15804 );
and ( n15806 , n15777 , n15790 );
nor ( n15807 , n15805 , n15806 );
nand ( n15808 , n15801 , n15807 );
xor ( n15809 , n15606 , n15614 );
and ( n15810 , n15809 , n15642 );
and ( n15811 , n15606 , n15614 );
or ( n15812 , n15810 , n15811 );
xor ( n15813 , n15625 , n15627 );
and ( n15814 , n15813 , n15641 );
and ( n15815 , n15625 , n15627 );
or ( n15816 , n15814 , n15815 );
not ( n15817 , n12845 );
and ( n15818 , n12781 , n493 );
not ( n15819 , n12781 );
and ( n15820 , n15819 , n12862 );
or ( n15821 , n15818 , n15820 );
not ( n15822 , n15821 );
or ( n15823 , n15817 , n15822 );
nand ( n15824 , n15746 , n15386 );
nand ( n15825 , n15823 , n15824 );
xor ( n15826 , n15816 , n15825 );
not ( n15827 , n13119 );
and ( n15828 , n495 , n12922 );
not ( n15829 , n495 );
and ( n15830 , n15829 , n12923 );
nor ( n15831 , n15828 , n15830 );
not ( n15832 , n15831 );
or ( n15833 , n15827 , n15832 );
nand ( n15834 , n15762 , n13056 );
nand ( n15835 , n15833 , n15834 );
xor ( n15836 , n15826 , n15835 );
xor ( n15837 , n15812 , n15836 );
not ( n15838 , n12743 );
not ( n15839 , n12560 );
not ( n15840 , n12515 );
or ( n15841 , n15839 , n15840 );
nand ( n15842 , n12512 , n499 );
nand ( n15843 , n15841 , n15842 );
not ( n15844 , n15843 );
or ( n15845 , n15838 , n15844 );
nand ( n15846 , n15604 , n12789 );
nand ( n15847 , n15845 , n15846 );
and ( n15848 , n15630 , n15640 );
not ( n15849 , n12731 );
xor ( n15850 , n491 , n12585 );
xnor ( n15851 , n15850 , n12593 );
not ( n15852 , n15851 );
or ( n15853 , n15849 , n15852 );
nand ( n15854 , n15623 , n12688 );
nand ( n15855 , n15853 , n15854 );
xor ( n15856 , n15848 , n15855 );
and ( n15857 , n12861 , n489 );
not ( n15858 , n12882 );
not ( n15859 , n489 );
not ( n15860 , n13068 );
or ( n15861 , n15859 , n15860 );
nand ( n15862 , n13067 , n12653 );
nand ( n15863 , n15861 , n15862 );
not ( n15864 , n15863 );
or ( n15865 , n15858 , n15864 );
nand ( n15866 , n15638 , n12635 );
nand ( n15867 , n15865 , n15866 );
xor ( n15868 , n15857 , n15867 );
xor ( n15869 , n15856 , n15868 );
xor ( n15870 , n15847 , n15869 );
xor ( n15871 , n15748 , n15752 );
and ( n15872 , n15871 , n15764 );
and ( n15873 , n15748 , n15752 );
or ( n15874 , n15872 , n15873 );
xor ( n15875 , n15870 , n15874 );
xor ( n15876 , n15837 , n15875 );
xor ( n15877 , n15653 , n15732 );
and ( n15878 , n15877 , n15737 );
and ( n15879 , n15653 , n15732 );
or ( n15880 , n15878 , n15879 );
not ( n15881 , n12563 );
not ( n15882 , n497 );
not ( n15883 , n13453 );
not ( n15884 , n15883 );
or ( n15885 , n15882 , n15884 );
nand ( n15886 , n13133 , n12579 );
nand ( n15887 , n15885 , n15886 );
not ( n15888 , n15887 );
or ( n15889 , n15881 , n15888 );
nand ( n15890 , n15610 , n12610 );
nand ( n15891 , n15889 , n15890 );
nand ( n15892 , n15575 , n12943 , n12930 );
nand ( n15893 , n15651 , n12909 );
nand ( n15894 , n15579 , n12930 , n501 );
nand ( n15895 , n15892 , n15893 , n15894 );
xor ( n15896 , n15891 , n15895 );
or ( n15897 , n15729 , n12554 );
xor ( n15898 , n15669 , n15684 );
and ( n15899 , n15898 , n15689 );
and ( n15900 , n15669 , n15684 );
or ( n15901 , n15899 , n15900 );
xor ( n15902 , n15670 , n15677 );
and ( n15903 , n15902 , n15683 );
and ( n15904 , n15670 , n15677 );
or ( n15905 , n15903 , n15904 );
not ( n15906 , n15683 );
xor ( n15907 , n15905 , n15906 );
not ( n15908 , n10256 );
or ( n15909 , n15908 , n15674 );
xnor ( n15910 , n457 , n521 );
or ( n15911 , n10196 , n15910 );
nand ( n15912 , n15909 , n15911 );
and ( n15913 , n457 , n523 );
xor ( n15914 , n15912 , n15913 );
not ( n15915 , n10223 );
not ( n15916 , n15915 );
not ( n15917 , n10215 );
or ( n15918 , n15916 , n15917 );
nand ( n15919 , n15918 , n459 );
xor ( n15920 , n15914 , n15919 );
xor ( n15921 , n15907 , n15920 );
nor ( n15922 , n15901 , n15921 );
not ( n15923 , n15922 );
nand ( n15924 , n15901 , n15921 );
nand ( n15925 , n15923 , n15924 );
nand ( n15926 , n15545 , n15691 );
nor ( n15927 , n15926 , n15701 );
nand ( n15928 , n12409 , n15927 );
not ( n15929 , n15928 );
buf ( n15930 , n12527 );
nand ( n15931 , n15929 , n15930 );
or ( n15932 , n15931 , n15564 );
not ( n15933 , n12505 );
not ( n15934 , n15927 );
nor ( n15935 , n15933 , n15934 );
and ( n15936 , n15935 , n12445 );
not ( n15937 , n15691 );
not ( n15938 , n15710 );
or ( n15939 , n15937 , n15938 );
nand ( n15940 , n15939 , n15692 );
nor ( n15941 , n15936 , n15940 );
nand ( n15942 , n15932 , n15941 );
not ( n15943 , n15563 );
nor ( n15944 , n12532 , n15928 );
not ( n15945 , n15944 );
or ( n15946 , n15943 , n15945 );
and ( n15947 , n12429 , n12503 );
nor ( n15948 , n15947 , n15934 );
nand ( n15949 , n15563 , n15948 );
nand ( n15950 , n15946 , n15949 );
nor ( n15951 , n15942 , n15950 );
xor ( n15952 , n15925 , n15951 );
and ( n15953 , n12550 , n15952 );
not ( n15954 , n12550 );
not ( n15955 , n15952 );
and ( n15956 , n15954 , n15955 );
nor ( n15957 , n15953 , n15956 );
or ( n15958 , n15957 , n15039 );
nand ( n15959 , n15897 , n15958 );
xor ( n15960 , n15896 , n15959 );
xor ( n15961 , n15880 , n15960 );
xor ( n15962 , n15765 , n15769 );
and ( n15963 , n15962 , n15774 );
and ( n15964 , n15765 , n15769 );
or ( n15965 , n15963 , n15964 );
xor ( n15966 , n15961 , n15965 );
xor ( n15967 , n15876 , n15966 );
xor ( n15968 , n15643 , n15738 );
and ( n15969 , n15968 , n15775 );
and ( n15970 , n15643 , n15738 );
or ( n15971 , n15969 , n15970 );
xor ( n15972 , n15967 , n15971 );
xor ( n15973 , n15415 , n15593 );
and ( n15974 , n15973 , n15776 );
and ( n15975 , n15415 , n15593 );
or ( n15976 , n15974 , n15975 );
or ( n15977 , n15972 , n15976 );
nand ( n15978 , n15972 , n15976 );
nand ( n15979 , n15977 , n15978 );
xnor ( n15980 , n15808 , n15979 );
nand ( n15981 , n10190 , n15980 );
nand ( n15982 , n10189 , n15981 );
and ( n15983 , n15982 , n471 );
not ( n15984 , n9401 );
not ( n15985 , n10040 );
buf ( n15986 , n10044 );
not ( n15987 , n15986 );
or ( n15988 , n15985 , n15987 );
nand ( n15989 , n15988 , n454 );
and ( n15990 , n15984 , n15989 );
not ( n15991 , n15984 );
nand ( n15992 , n454 , n10040 , n15986 );
and ( n15993 , n15991 , n15992 );
nor ( n15994 , n15990 , n15993 );
not ( n15995 , n15994 );
not ( n15996 , n15374 );
not ( n15997 , n15360 );
not ( n15998 , n15345 );
not ( n15999 , n15304 );
or ( n16000 , n15998 , n15999 );
not ( n16001 , n15358 );
nand ( n16002 , n16000 , n16001 );
not ( n16003 , n16002 );
or ( n16004 , n15997 , n16003 );
buf ( n16005 , n15368 );
nand ( n16006 , n16004 , n16005 );
not ( n16007 , n16006 );
or ( n16008 , n15996 , n16007 );
not ( n16009 , n13752 );
nand ( n16010 , n16008 , n16009 );
not ( n16011 , n13754 );
nand ( n16012 , n16011 , n13499 );
not ( n16013 , n16012 );
and ( n16014 , n16010 , n16013 );
not ( n16015 , n16010 );
and ( n16016 , n16015 , n16012 );
nor ( n16017 , n16014 , n16016 );
nand ( n16018 , n16017 , n10190 );
nand ( n16019 , n15995 , n16018 );
and ( n16020 , n16019 , n469 );
not ( n16021 , n10190 );
not ( n16022 , n15799 );
not ( n16023 , n16022 );
not ( n16024 , n15375 );
not ( n16025 , n16006 );
or ( n16026 , n16024 , n16025 );
nand ( n16027 , n16026 , n13755 );
not ( n16028 , n16027 );
or ( n16029 , n16023 , n16028 );
nand ( n16030 , n16029 , n15803 );
not ( n16031 , n15802 );
nor ( n16032 , n16031 , n15806 );
and ( n16033 , n16030 , n16032 );
not ( n16034 , n16030 );
not ( n16035 , n16032 );
and ( n16036 , n16034 , n16035 );
nor ( n16037 , n16033 , n16036 );
not ( n16038 , n16037 );
or ( n16039 , n16021 , n16038 );
buf ( n16040 , n10046 );
not ( n16041 , n16040 );
nor ( n16042 , n9802 , n9814 );
not ( n16043 , n16042 );
not ( n16044 , n16043 );
or ( n16045 , n16041 , n16044 );
not ( n16046 , n10040 );
nor ( n16047 , n16046 , n16042 );
nand ( n16048 , n15984 , n16047 );
nand ( n16049 , n16045 , n16048 );
nand ( n16050 , n10031 , n10048 );
not ( n16051 , n16050 );
and ( n16052 , n16049 , n16051 );
not ( n16053 , n16049 );
and ( n16054 , n16053 , n16050 );
nor ( n16055 , n16052 , n16054 );
nand ( n16056 , n16055 , n454 );
nand ( n16057 , n16039 , n16056 );
and ( n16058 , n16057 , n471 );
xor ( n16059 , n16020 , n16058 );
not ( n16060 , n454 );
not ( n16061 , n10040 );
not ( n16062 , n15984 );
or ( n16063 , n16061 , n16062 );
nand ( n16064 , n16063 , n15986 );
and ( n16065 , n16043 , n10045 );
xor ( n16066 , n16064 , n16065 );
not ( n16067 , n16066 );
or ( n16068 , n16060 , n16067 );
nand ( n16069 , n16022 , n15803 );
xnor ( n16070 , n16027 , n16069 );
nand ( n16071 , n16070 , n10190 );
nand ( n16072 , n16068 , n16071 );
and ( n16073 , n16072 , n470 );
and ( n16074 , n16059 , n16073 );
and ( n16075 , n16020 , n16058 );
or ( n16076 , n16074 , n16075 );
xor ( n16077 , n15983 , n16076 );
and ( n16078 , n16057 , n470 );
not ( n16079 , n16072 );
not ( n16080 , n469 );
nor ( n16081 , n16079 , n16080 );
xor ( n16082 , n16078 , n16081 );
buf ( n16083 , n10178 );
not ( n16084 , n16083 );
not ( n16085 , n16084 );
not ( n16086 , n10052 );
or ( n16087 , n16085 , n16086 );
nand ( n16088 , n16087 , n10181 );
xor ( n16089 , n10116 , n10167 );
and ( n16090 , n16089 , n10172 );
and ( n16091 , n10116 , n10167 );
or ( n16092 , n16090 , n16091 );
xor ( n16093 , n10069 , n10080 );
and ( n16094 , n16093 , n10087 );
and ( n16095 , n10069 , n10080 );
or ( n16096 , n16094 , n16095 );
not ( n16097 , n9730 );
and ( n16098 , n6618 , n5146 );
not ( n16099 , n6618 );
and ( n16100 , n16099 , n543 );
or ( n16101 , n16098 , n16100 );
not ( n16102 , n16101 );
or ( n16103 , n16097 , n16102 );
nand ( n16104 , n10094 , n4671 );
nand ( n16105 , n16103 , n16104 );
not ( n16106 , n541 );
not ( n16107 , n7019 );
or ( n16108 , n16106 , n16107 );
nand ( n16109 , n7015 , n5734 );
nand ( n16110 , n16108 , n16109 );
not ( n16111 , n16110 );
not ( n16112 , n5786 );
or ( n16113 , n16111 , n16112 );
nand ( n16114 , n10064 , n10067 );
nand ( n16115 , n16113 , n16114 );
xor ( n16116 , n16105 , n16115 );
xor ( n16117 , n10135 , n10137 );
and ( n16118 , n16117 , n10150 );
and ( n16119 , n10135 , n10137 );
or ( n16120 , n16118 , n16119 );
xor ( n16121 , n16116 , n16120 );
xor ( n16122 , n16096 , n16121 );
not ( n16123 , n4659 );
not ( n16124 , n539 );
not ( n16125 , n5467 );
or ( n16126 , n16124 , n16125 );
nand ( n16127 , n5466 , n4477 );
nand ( n16128 , n16126 , n16127 );
not ( n16129 , n16128 );
or ( n16130 , n16123 , n16129 );
nand ( n16131 , n10127 , n4450 );
nand ( n16132 , n16130 , n16131 );
not ( n16133 , n5595 );
not ( n16134 , n545 );
not ( n16135 , n9867 );
or ( n16136 , n16134 , n16135 );
nand ( n16137 , n9866 , n4666 );
nand ( n16138 , n16136 , n16137 );
not ( n16139 , n16138 );
or ( n16140 , n16133 , n16139 );
nand ( n16141 , n10078 , n5339 );
nand ( n16142 , n16140 , n16141 );
xor ( n16143 , n16132 , n16142 );
not ( n16144 , n6667 );
not ( n16145 , n10083 );
or ( n16146 , n16144 , n16145 );
not ( n16147 , n7190 );
not ( n16148 , n9976 );
or ( n16149 , n16147 , n16148 );
nand ( n16150 , n9977 , n549 );
nand ( n16151 , n16149 , n16150 );
nand ( n16152 , n16151 , n6095 );
nand ( n16153 , n16146 , n16152 );
xor ( n16154 , n16143 , n16153 );
xor ( n16155 , n16122 , n16154 );
not ( n16156 , n6983 );
and ( n16157 , n547 , n9692 );
not ( n16158 , n547 );
not ( n16159 , n9692 );
and ( n16160 , n16158 , n16159 );
or ( n16161 , n16157 , n16160 );
not ( n16162 , n16161 );
or ( n16163 , n16156 , n16162 );
nand ( n16164 , n10112 , n7026 );
nand ( n16165 , n16163 , n16164 );
not ( n16166 , n5697 );
and ( n16167 , n5145 , n5605 );
not ( n16168 , n5145 );
and ( n16169 , n16168 , n537 );
or ( n16170 , n16167 , n16169 );
not ( n16171 , n16170 );
or ( n16172 , n16166 , n16171 );
buf ( n16173 , n5609 );
nand ( n16174 , n10145 , n16173 );
nand ( n16175 , n16172 , n16174 );
and ( n16176 , n10139 , n10149 );
xor ( n16177 , n16175 , n16176 );
nand ( n16178 , n7946 , n537 );
nand ( n16179 , n9020 , n10120 );
or ( n16180 , n16178 , n16179 );
nand ( n16181 , n16178 , n16179 );
nand ( n16182 , n16180 , n16181 );
xor ( n16183 , n16177 , n16182 );
xor ( n16184 , n16165 , n16183 );
xor ( n16185 , n10099 , n10103 );
and ( n16186 , n16185 , n10114 );
and ( n16187 , n10099 , n10103 );
or ( n16188 , n16186 , n16187 );
xor ( n16189 , n16184 , n16188 );
xor ( n16190 , n10121 , n10151 );
and ( n16191 , n16190 , n10156 );
and ( n16192 , n10121 , n10151 );
or ( n16193 , n16191 , n16192 );
xor ( n16194 , n16189 , n16193 );
xor ( n16195 , n10057 , n10088 );
and ( n16196 , n16195 , n10115 );
and ( n16197 , n10057 , n10088 );
or ( n16198 , n16196 , n16197 );
xor ( n16199 , n16194 , n16198 );
xor ( n16200 , n16155 , n16199 );
xor ( n16201 , n10157 , n10161 );
and ( n16202 , n16201 , n10166 );
and ( n16203 , n10157 , n10161 );
or ( n16204 , n16202 , n16203 );
xor ( n16205 , n16200 , n16204 );
nand ( n16206 , n16092 , n16205 );
not ( n16207 , n16205 );
not ( n16208 , n16092 );
nand ( n16209 , n16207 , n16208 );
nand ( n16210 , n16206 , n16209 );
not ( n16211 , n16210 );
and ( n16212 , n16088 , n16211 );
not ( n16213 , n16088 );
and ( n16214 , n16213 , n16210 );
nor ( n16215 , n16212 , n16214 );
nand ( n16216 , n16215 , n454 );
not ( n16217 , n15977 );
not ( n16218 , n15808 );
or ( n16219 , n16217 , n16218 );
not ( n16220 , n15386 );
not ( n16221 , n15821 );
or ( n16222 , n16220 , n16221 );
not ( n16223 , n493 );
not ( n16224 , n13438 );
or ( n16225 , n16223 , n16224 );
nand ( n16226 , n12764 , n12862 );
nand ( n16227 , n16225 , n16226 );
nand ( n16228 , n16227 , n12845 );
nand ( n16229 , n16222 , n16228 );
not ( n16230 , n13056 );
not ( n16231 , n15831 );
or ( n16232 , n16230 , n16231 );
not ( n16233 , n495 );
nand ( n16234 , n16233 , n13450 );
not ( n16235 , n16234 );
nand ( n16236 , n13451 , n495 );
not ( n16237 , n16236 );
or ( n16238 , n16235 , n16237 );
nand ( n16239 , n16238 , n13119 );
nand ( n16240 , n16232 , n16239 );
xor ( n16241 , n16229 , n16240 );
not ( n16242 , n12610 );
not ( n16243 , n15887 );
or ( n16244 , n16242 , n16243 );
not ( n16245 , n12579 );
not ( n16246 , n15602 );
or ( n16247 , n16245 , n16246 );
nand ( n16248 , n15599 , n497 );
nand ( n16249 , n16247 , n16248 );
nand ( n16250 , n16249 , n12563 );
nand ( n16251 , n16244 , n16250 );
xor ( n16252 , n16241 , n16251 );
xor ( n16253 , n15891 , n15895 );
and ( n16254 , n16253 , n15959 );
and ( n16255 , n15891 , n15895 );
or ( n16256 , n16254 , n16255 );
xor ( n16257 , n16252 , n16256 );
xor ( n16258 , n15847 , n15869 );
and ( n16259 , n16258 , n15874 );
and ( n16260 , n15847 , n15869 );
or ( n16261 , n16259 , n16260 );
xor ( n16262 , n16257 , n16261 );
xor ( n16263 , n15880 , n15960 );
and ( n16264 , n16263 , n15965 );
and ( n16265 , n15880 , n15960 );
or ( n16266 , n16264 , n16265 );
xor ( n16267 , n16262 , n16266 );
not ( n16268 , n15694 );
not ( n16269 , n15713 );
or ( n16270 , n16268 , n16269 );
nand ( n16271 , n16270 , n15719 );
nand ( n16272 , n12930 , n501 );
or ( n16273 , n16271 , n16272 );
not ( n16274 , n15575 );
not ( n16275 , n12908 );
nor ( n16276 , n16275 , n12943 );
nand ( n16277 , n16274 , n16276 );
nor ( n16278 , n15252 , n501 );
nand ( n16279 , n15726 , n16278 );
nand ( n16280 , n15575 , n14747 );
nand ( n16281 , n16273 , n16277 , n16279 , n16280 );
xor ( n16282 , n15848 , n15855 );
and ( n16283 , n16282 , n15868 );
and ( n16284 , n15848 , n15855 );
or ( n16285 , n16283 , n16284 );
xor ( n16286 , n16281 , n16285 );
not ( n16287 , n12789 );
not ( n16288 , n15843 );
or ( n16289 , n16287 , n16288 );
and ( n16290 , n13339 , n12560 );
not ( n16291 , n13339 );
and ( n16292 , n16291 , n499 );
nor ( n16293 , n16290 , n16292 );
or ( n16294 , n16293 , n12742 );
nand ( n16295 , n16289 , n16294 );
xor ( n16296 , n16286 , n16295 );
not ( n16297 , n504 );
not ( n16298 , n503 );
or ( n16299 , n15942 , n15950 );
xor ( n16300 , n15905 , n15906 );
and ( n16301 , n16300 , n15920 );
and ( n16302 , n15905 , n15906 );
or ( n16303 , n16301 , n16302 );
or ( n16304 , n15908 , n15910 );
or ( n16305 , n10196 , n2984 );
nand ( n16306 , n16304 , n16305 );
nand ( n16307 , n522 , n457 );
xor ( n16308 , n16306 , n16307 );
xor ( n16309 , n15912 , n15913 );
and ( n16310 , n16309 , n15919 );
and ( n16311 , n15912 , n15913 );
or ( n16312 , n16310 , n16311 );
xor ( n16313 , n16308 , n16312 );
nor ( n16314 , n16303 , n16313 );
not ( n16315 , n16314 );
not ( n16316 , n16315 );
and ( n16317 , n16303 , n16313 );
nor ( n16318 , n16316 , n16317 );
not ( n16319 , n16318 );
not ( n16320 , n15924 );
and ( n16321 , n16319 , n16320 );
and ( n16322 , n16318 , n15924 , n15922 );
nor ( n16323 , n16321 , n16322 );
or ( n16324 , n16318 , n15922 );
nand ( n16325 , n16299 , n16323 , n16324 );
not ( n16326 , n15942 );
not ( n16327 , n15924 );
not ( n16328 , n16318 );
or ( n16329 , n16327 , n16328 );
nand ( n16330 , n16329 , n16323 );
nor ( n16331 , n15950 , n16330 );
nand ( n16332 , n16326 , n16331 );
nand ( n16333 , n16325 , n16332 );
not ( n16334 , n16333 );
or ( n16335 , n16298 , n16334 );
not ( n16336 , n16333 );
nand ( n16337 , n16336 , n12550 );
nand ( n16338 , n16335 , n16337 );
not ( n16339 , n16338 );
or ( n16340 , n16297 , n16339 );
not ( n16341 , n15957 );
nand ( n16342 , n16341 , n12555 );
nand ( n16343 , n16340 , n16342 );
not ( n16344 , n12688 );
not ( n16345 , n15851 );
or ( n16346 , n16344 , n16345 );
xor ( n16347 , n12574 , n12703 );
or ( n16348 , n16347 , n12686 );
nand ( n16349 , n16346 , n16348 );
and ( n16350 , n15867 , n15857 );
xor ( n16351 , n16349 , n16350 );
not ( n16352 , n489 );
nor ( n16353 , n16352 , n13037 );
not ( n16354 , n12882 );
xor ( n16355 , n13095 , n12653 );
not ( n16356 , n16355 );
not ( n16357 , n16356 );
or ( n16358 , n16354 , n16357 );
nand ( n16359 , n15863 , n12635 );
nand ( n16360 , n16358 , n16359 );
xor ( n16361 , n16353 , n16360 );
xor ( n16362 , n16351 , n16361 );
xor ( n16363 , n16343 , n16362 );
xor ( n16364 , n15816 , n15825 );
and ( n16365 , n16364 , n15835 );
and ( n16366 , n15816 , n15825 );
or ( n16367 , n16365 , n16366 );
xor ( n16368 , n16363 , n16367 );
xor ( n16369 , n16296 , n16368 );
xor ( n16370 , n15812 , n15836 );
and ( n16371 , n16370 , n15875 );
and ( n16372 , n15812 , n15836 );
or ( n16373 , n16371 , n16372 );
xor ( n16374 , n16369 , n16373 );
xor ( n16375 , n16267 , n16374 );
xor ( n16376 , n15876 , n15966 );
and ( n16377 , n16376 , n15971 );
and ( n16378 , n15876 , n15966 );
or ( n16379 , n16377 , n16378 );
nand ( n16380 , n16375 , n16379 );
buf ( n16381 , n16380 );
not ( n16382 , n16381 );
nor ( n16383 , n16375 , n16379 );
buf ( n16384 , n16383 );
nor ( n16385 , n16382 , n16384 );
not ( n16386 , n15978 );
nor ( n16387 , n16385 , n16386 );
nand ( n16388 , n16219 , n16387 );
and ( n16389 , n16385 , n16386 );
nor ( n16390 , n16389 , n454 );
nand ( n16391 , n15977 , n15808 , n16385 );
nand ( n16392 , n16388 , n16390 , n16391 );
nand ( n16393 , n16216 , n16392 );
not ( n16394 , n16393 );
not ( n16395 , n472 );
nor ( n16396 , n16394 , n16395 );
xor ( n16397 , n16082 , n16396 );
and ( n16398 , n16077 , n16397 );
and ( n16399 , n15983 , n16076 );
or ( n16400 , n16398 , n16399 );
not ( n16401 , n16400 );
nor ( n16402 , n16205 , n16092 );
nor ( n16403 , n16402 , n10178 );
not ( n16404 , n16403 );
not ( n16405 , n10052 );
or ( n16406 , n16404 , n16405 );
nand ( n16407 , n16206 , n10180 );
nand ( n16408 , n16407 , n16209 );
buf ( n16409 , n16408 );
nand ( n16410 , n16406 , n16409 );
xor ( n16411 , n16155 , n16199 );
and ( n16412 , n16411 , n16204 );
and ( n16413 , n16155 , n16199 );
or ( n16414 , n16412 , n16413 );
xor ( n16415 , n16132 , n16142 );
and ( n16416 , n16415 , n16153 );
and ( n16417 , n16132 , n16142 );
or ( n16418 , n16416 , n16417 );
not ( n16419 , n10067 );
not ( n16420 , n16110 );
or ( n16421 , n16419 , n16420 );
not ( n16422 , n541 );
not ( n16423 , n6657 );
or ( n16424 , n16422 , n16423 );
nand ( n16425 , n6656 , n5734 );
nand ( n16426 , n16424 , n16425 );
nand ( n16427 , n16426 , n5786 );
nand ( n16428 , n16421 , n16427 );
not ( n16429 , n5595 );
and ( n16430 , n9517 , n545 );
not ( n16431 , n9517 );
and ( n16432 , n16431 , n4666 );
or ( n16433 , n16430 , n16432 );
not ( n16434 , n16433 );
or ( n16435 , n16429 , n16434 );
nand ( n16436 , n16138 , n5341 );
nand ( n16437 , n16435 , n16436 );
xor ( n16438 , n16428 , n16437 );
not ( n16439 , n6667 );
not ( n16440 , n16151 );
or ( n16441 , n16439 , n16440 );
nand ( n16442 , n16441 , n7192 );
xor ( n16443 , n16438 , n16442 );
xor ( n16444 , n16418 , n16443 );
not ( n16445 , n4450 );
not ( n16446 , n16128 );
or ( n16447 , n16445 , n16446 );
nand ( n16448 , n539 , n10060 );
not ( n16449 , n16448 );
not ( n16450 , n10060 );
nand ( n16451 , n16450 , n4477 );
not ( n16452 , n16451 );
or ( n16453 , n16449 , n16452 );
nand ( n16454 , n16453 , n4447 );
nand ( n16455 , n16447 , n16454 );
not ( n16456 , n5330 );
not ( n16457 , n543 );
not ( n16458 , n6968 );
or ( n16459 , n16457 , n16458 );
nand ( n16460 , n6967 , n5146 );
nand ( n16461 , n16459 , n16460 );
not ( n16462 , n16461 );
or ( n16463 , n16456 , n16462 );
nand ( n16464 , n4671 , n16101 );
nand ( n16465 , n16463 , n16464 );
xor ( n16466 , n16455 , n16465 );
not ( n16467 , n7026 );
not ( n16468 , n16161 );
or ( n16469 , n16467 , n16468 );
xor ( n16470 , n547 , n9688 );
nand ( n16471 , n16470 , n6983 );
nand ( n16472 , n16469 , n16471 );
xor ( n16473 , n16466 , n16472 );
xor ( n16474 , n16444 , n16473 );
not ( n16475 , n16173 );
not ( n16476 , n16170 );
or ( n16477 , n16475 , n16476 );
not ( n16478 , n537 );
not ( n16479 , n8068 );
or ( n16480 , n16478 , n16479 );
nand ( n16481 , n7109 , n5605 );
nand ( n16482 , n16480 , n16481 );
nand ( n16483 , n16482 , n5697 );
nand ( n16484 , n16477 , n16483 );
nand ( n16485 , n7781 , n537 );
xor ( n16486 , n16484 , n16485 );
xor ( n16487 , n16486 , n16181 );
xor ( n16488 , n16175 , n16176 );
and ( n16489 , n16488 , n16182 );
and ( n16490 , n16175 , n16176 );
or ( n16491 , n16489 , n16490 );
xor ( n16492 , n16487 , n16491 );
xor ( n16493 , n16105 , n16115 );
and ( n16494 , n16493 , n16120 );
and ( n16495 , n16105 , n16115 );
or ( n16496 , n16494 , n16495 );
xor ( n16497 , n16492 , n16496 );
xor ( n16498 , n16165 , n16183 );
and ( n16499 , n16498 , n16188 );
and ( n16500 , n16165 , n16183 );
or ( n16501 , n16499 , n16500 );
xor ( n16502 , n16497 , n16501 );
xor ( n16503 , n16096 , n16121 );
and ( n16504 , n16503 , n16154 );
and ( n16505 , n16096 , n16121 );
or ( n16506 , n16504 , n16505 );
xor ( n16507 , n16502 , n16506 );
xor ( n16508 , n16474 , n16507 );
xor ( n16509 , n16189 , n16193 );
and ( n16510 , n16509 , n16198 );
and ( n16511 , n16189 , n16193 );
or ( n16512 , n16510 , n16511 );
xor ( n16513 , n16508 , n16512 );
nor ( n16514 , n16414 , n16513 );
buf ( n16515 , n16514 );
not ( n16516 , n16515 );
buf ( n16517 , n16513 );
nand ( n16518 , n16414 , n16517 );
nand ( n16519 , n16516 , n16518 );
not ( n16520 , n16519 );
and ( n16521 , n16410 , n16520 );
not ( n16522 , n16410 );
and ( n16523 , n16522 , n16519 );
nor ( n16524 , n16521 , n16523 );
not ( n16525 , n16524 );
not ( n16526 , n454 );
or ( n16527 , n16525 , n16526 );
not ( n16528 , n15977 );
nor ( n16529 , n16528 , n16384 );
not ( n16530 , n16529 );
not ( n16531 , n15808 );
or ( n16532 , n16530 , n16531 );
nor ( n16533 , n16383 , n15978 );
not ( n16534 , n16533 );
and ( n16535 , n16381 , n16534 );
nand ( n16536 , n16532 , n16535 );
not ( n16537 , n13119 );
and ( n16538 , n495 , n12973 );
not ( n16539 , n495 );
and ( n16540 , n16539 , n13453 );
or ( n16541 , n16538 , n16540 );
not ( n16542 , n16541 );
or ( n16543 , n16537 , n16542 );
not ( n16544 , n16236 );
not ( n16545 , n16234 );
or ( n16546 , n16544 , n16545 );
nand ( n16547 , n16546 , n13056 );
nand ( n16548 , n16543 , n16547 );
not ( n16549 , n12845 );
not ( n16550 , n493 );
not ( n16551 , n12923 );
or ( n16552 , n16550 , n16551 );
or ( n16553 , n12923 , n493 );
nand ( n16554 , n16552 , n16553 );
not ( n16555 , n16554 );
or ( n16556 , n16549 , n16555 );
nand ( n16557 , n16227 , n15386 );
nand ( n16558 , n16556 , n16557 );
xor ( n16559 , n16548 , n16558 );
not ( n16560 , n12909 );
and ( n16561 , n501 , n15720 );
not ( n16562 , n501 );
and ( n16563 , n16562 , n15727 );
nor ( n16564 , n16561 , n16563 );
not ( n16565 , n16564 );
or ( n16566 , n16560 , n16565 );
and ( n16567 , n15952 , n12943 );
not ( n16568 , n15952 );
and ( n16569 , n16568 , n501 );
or ( n16570 , n16567 , n16569 );
nand ( n16571 , n16570 , n12930 );
nand ( n16572 , n16566 , n16571 );
xor ( n16573 , n16559 , n16572 );
xor ( n16574 , n16281 , n16285 );
and ( n16575 , n16574 , n16295 );
and ( n16576 , n16281 , n16285 );
or ( n16577 , n16575 , n16576 );
xor ( n16578 , n16573 , n16577 );
not ( n16579 , n15474 );
nor ( n16580 , n12562 , n497 );
nand ( n16581 , n16579 , n16580 );
nand ( n16582 , n16249 , n12610 );
nand ( n16583 , n12563 , n497 );
or ( n16584 , n12511 , n16583 );
nand ( n16585 , n16581 , n16582 , n16584 );
xor ( n16586 , n16349 , n16350 );
and ( n16587 , n16586 , n16361 );
and ( n16588 , n16349 , n16350 );
or ( n16589 , n16587 , n16588 );
xor ( n16590 , n16585 , n16589 );
not ( n16591 , n12742 );
not ( n16592 , n499 );
not ( n16593 , n16274 );
or ( n16594 , n16592 , n16593 );
nand ( n16595 , n15575 , n1407 );
nand ( n16596 , n16594 , n16595 );
nand ( n16597 , n16591 , n16596 );
not ( n16598 , n16293 );
nand ( n16599 , n16598 , n12789 );
nand ( n16600 , n16597 , n16599 );
xor ( n16601 , n16590 , n16600 );
xor ( n16602 , n16578 , n16601 );
xor ( n16603 , n16343 , n16362 );
and ( n16604 , n16603 , n16367 );
and ( n16605 , n16343 , n16362 );
or ( n16606 , n16604 , n16605 );
not ( n16607 , n504 );
not ( n16608 , n503 );
or ( n16609 , n15692 , n15922 );
nand ( n16610 , n16609 , n15924 );
and ( n16611 , n16610 , n16315 );
nor ( n16612 , n16611 , n16317 );
not ( n16613 , n16612 );
xor ( n16614 , n16306 , n16307 );
and ( n16615 , n16614 , n16312 );
and ( n16616 , n16306 , n16307 );
or ( n16617 , n16615 , n16616 );
not ( n16618 , n16307 );
nand ( n16619 , n521 , n457 );
not ( n16620 , n16619 );
or ( n16621 , n10256 , n10197 );
nand ( n16622 , n16621 , n457 );
not ( n16623 , n16622 );
or ( n16624 , n16620 , n16623 );
or ( n16625 , n16622 , n16619 );
nand ( n16626 , n16624 , n16625 );
not ( n16627 , n16626 );
or ( n16628 , n16618 , n16627 );
or ( n16629 , n16626 , n16307 );
nand ( n16630 , n16628 , n16629 );
xnor ( n16631 , n16617 , n16630 );
nor ( n16632 , n16613 , n16631 );
not ( n16633 , n16632 );
not ( n16634 , n15711 );
not ( n16635 , n15704 );
or ( n16636 , n16634 , n16635 );
not ( n16637 , n15691 );
nor ( n16638 , n16637 , n16314 , n15922 );
nand ( n16639 , n16636 , n16638 );
not ( n16640 , n16639 );
or ( n16641 , n16633 , n16640 );
not ( n16642 , n16612 );
not ( n16643 , n16639 );
or ( n16644 , n16642 , n16643 );
xor ( n16645 , n16617 , n16307 );
xor ( n16646 , n16645 , n16626 );
nand ( n16647 , n16644 , n16646 );
nand ( n16648 , n16641 , n16647 );
not ( n16649 , n16648 );
not ( n16650 , n16649 );
or ( n16651 , n16608 , n16650 );
nand ( n16652 , n12516 , n16648 );
nand ( n16653 , n16651 , n16652 );
not ( n16654 , n16653 );
or ( n16655 , n16607 , n16654 );
nand ( n16656 , n16338 , n12555 );
nand ( n16657 , n16655 , n16656 );
xor ( n16658 , n16229 , n16240 );
and ( n16659 , n16658 , n16251 );
and ( n16660 , n16229 , n16240 );
or ( n16661 , n16659 , n16660 );
xor ( n16662 , n16657 , n16661 );
and ( n16663 , n16353 , n16360 );
xor ( n16664 , n491 , n12780 );
not ( n16665 , n16664 );
or ( n16666 , n16665 , n12686 );
not ( n16667 , n16347 );
nand ( n16668 , n16667 , n12688 );
nand ( n16669 , n16666 , n16668 );
xor ( n16670 , n16663 , n16669 );
and ( n16671 , n14167 , n489 );
not ( n16672 , n12673 );
and ( n16673 , n12598 , n12653 );
not ( n16674 , n12598 );
and ( n16675 , n16674 , n489 );
or ( n16676 , n16673 , n16675 );
not ( n16677 , n16676 );
or ( n16678 , n16672 , n16677 );
not ( n16679 , n16355 );
nand ( n16680 , n16679 , n12635 );
nand ( n16681 , n16678 , n16680 );
xor ( n16682 , n16671 , n16681 );
xor ( n16683 , n16670 , n16682 );
xor ( n16684 , n16662 , n16683 );
xor ( n16685 , n16606 , n16684 );
xor ( n16686 , n16252 , n16256 );
and ( n16687 , n16686 , n16261 );
and ( n16688 , n16252 , n16256 );
or ( n16689 , n16687 , n16688 );
xor ( n16690 , n16685 , n16689 );
xor ( n16691 , n16602 , n16690 );
xor ( n16692 , n16296 , n16368 );
and ( n16693 , n16692 , n16373 );
and ( n16694 , n16296 , n16368 );
or ( n16695 , n16693 , n16694 );
xor ( n16696 , n16691 , n16695 );
xor ( n16697 , n16262 , n16266 );
and ( n16698 , n16697 , n16374 );
and ( n16699 , n16262 , n16266 );
or ( n16700 , n16698 , n16699 );
or ( n16701 , n16696 , n16700 );
nand ( n16702 , n16696 , n16700 );
nand ( n16703 , n16701 , n16702 );
not ( n16704 , n16703 );
and ( n16705 , n16536 , n16704 );
not ( n16706 , n16536 );
and ( n16707 , n16706 , n16703 );
nor ( n16708 , n16705 , n16707 );
nand ( n16709 , n16708 , n10190 );
nand ( n16710 , n16527 , n16709 );
and ( n16711 , n16710 , n472 );
xor ( n16712 , n16078 , n16081 );
and ( n16713 , n16712 , n16396 );
and ( n16714 , n16078 , n16081 );
or ( n16715 , n16713 , n16714 );
xor ( n16716 , n16711 , n16715 );
and ( n16717 , n16057 , n469 );
nand ( n16718 , n16216 , n16392 );
and ( n16719 , n16718 , n471 );
xor ( n16720 , n16717 , n16719 );
and ( n16721 , n15982 , n470 );
xor ( n16722 , n16720 , n16721 );
xor ( n16723 , n16716 , n16722 );
not ( n16724 , n16723 );
and ( n16725 , n16401 , n16724 );
xor ( n16726 , n15983 , n16076 );
xor ( n16727 , n16726 , n16397 );
and ( n16728 , n15982 , n472 );
and ( n16729 , n16019 , n470 );
nor ( n16730 , n8323 , n8318 );
not ( n16731 , n454 );
nor ( n16732 , n16730 , n16731 );
or ( n16733 , n7540 , n7760 );
not ( n16734 , n16733 );
buf ( n16735 , n8304 );
not ( n16736 , n16735 );
not ( n16737 , n9399 );
not ( n16738 , n8339 );
not ( n16739 , n16738 );
or ( n16740 , n16737 , n16739 );
not ( n16741 , n8280 );
nand ( n16742 , n16740 , n16741 );
not ( n16743 , n16742 );
or ( n16744 , n16736 , n16743 );
buf ( n16745 , n8314 );
nand ( n16746 , n16744 , n16745 );
not ( n16747 , n16746 );
or ( n16748 , n16734 , n16747 );
nand ( n16749 , n16748 , n8320 );
and ( n16750 , n16732 , n16749 );
nand ( n16751 , n16009 , n15374 );
xnor ( n16752 , n16006 , n16751 );
and ( n16753 , n16752 , n10190 );
nor ( n16754 , n16750 , n16753 );
not ( n16755 , n16749 );
and ( n16756 , n16730 , n454 );
nand ( n16757 , n16755 , n16756 );
nand ( n16758 , n16754 , n16757 );
and ( n16759 , n16758 , n469 );
xor ( n16760 , n16729 , n16759 );
and ( n16761 , n16057 , n472 );
and ( n16762 , n16760 , n16761 );
and ( n16763 , n16729 , n16759 );
or ( n16764 , n16762 , n16763 );
xor ( n16765 , n16728 , n16764 );
xor ( n16766 , n16020 , n16058 );
xor ( n16767 , n16766 , n16073 );
and ( n16768 , n16765 , n16767 );
and ( n16769 , n16728 , n16764 );
or ( n16770 , n16768 , n16769 );
nor ( n16771 , n16727 , n16770 );
nor ( n16772 , n16725 , n16771 );
not ( n16773 , n15294 );
nand ( n16774 , n15299 , n16773 );
xnor ( n16775 , n15163 , n16774 );
nand ( n16776 , n16775 , n10190 );
buf ( n16777 , n9330 );
not ( n16778 , n9376 );
nand ( n16779 , n16777 , n16778 );
not ( n16780 , n9394 );
nand ( n16781 , n16779 , n16780 );
nand ( n16782 , n9396 , n9389 );
nand ( n16783 , n16781 , n16782 , n454 );
not ( n16784 , n16782 );
nand ( n16785 , n16784 , n16779 , n16780 , n454 );
nand ( n16786 , n16776 , n16783 , n16785 );
and ( n16787 , n16786 , n471 );
not ( n16788 , n8767 );
not ( n16789 , n16788 );
not ( n16790 , n8832 );
not ( n16791 , n9314 );
or ( n16792 , n16790 , n16791 );
nand ( n16793 , n16792 , n9318 );
buf ( n16794 , n16793 );
not ( n16795 , n16794 );
or ( n16796 , n16789 , n16795 );
buf ( n16797 , n9322 );
nand ( n16798 , n16796 , n16797 );
not ( n16799 , n16798 );
not ( n16800 , n454 );
not ( n16801 , n8674 );
nand ( n16802 , n16801 , n9327 );
nor ( n16803 , n16800 , n16802 );
nand ( n16804 , n16799 , n16803 );
and ( n16805 , n16802 , n454 );
and ( n16806 , n16798 , n16805 );
nand ( n16807 , n15148 , n15152 );
not ( n16808 , n14586 );
not ( n16809 , n16808 );
buf ( n16810 , n15143 );
not ( n16811 , n16810 );
or ( n16812 , n16809 , n16811 );
nand ( n16813 , n16812 , n15149 );
xnor ( n16814 , n16807 , n16813 );
and ( n16815 , n16814 , n10190 );
nor ( n16816 , n16806 , n16815 );
nand ( n16817 , n16804 , n16816 );
and ( n16818 , n16817 , n469 );
not ( n16819 , n9390 );
nand ( n16820 , n16819 , n9393 );
not ( n16821 , n16820 );
nor ( n16822 , n16821 , n16731 );
not ( n16823 , n16822 );
nand ( n16824 , n16777 , n9375 );
nand ( n16825 , n16824 , n9391 );
not ( n16826 , n16825 );
or ( n16827 , n16823 , n16826 );
nand ( n16828 , n9391 , n454 );
nor ( n16829 , n16820 , n16828 );
and ( n16830 , n16829 , n16824 );
nand ( n16831 , n14345 , n15162 );
xnor ( n16832 , n15159 , n16831 );
and ( n16833 , n16832 , n10190 );
nor ( n16834 , n16830 , n16833 );
nand ( n16835 , n16827 , n16834 );
and ( n16836 , n16835 , n471 );
xor ( n16837 , n16818 , n16836 );
not ( n16838 , n454 );
nand ( n16839 , n9375 , n9391 );
xnor ( n16840 , n16839 , n16777 );
not ( n16841 , n16840 );
or ( n16842 , n16838 , n16841 );
nand ( n16843 , n14413 , n15158 );
xnor ( n16844 , n15155 , n16843 );
nand ( n16845 , n16844 , n10190 );
nand ( n16846 , n16842 , n16845 );
and ( n16847 , n16846 , n470 );
and ( n16848 , n16837 , n16847 );
and ( n16849 , n16818 , n16836 );
or ( n16850 , n16848 , n16849 );
xor ( n16851 , n16787 , n16850 );
and ( n16852 , n16835 , n470 );
and ( n16853 , n16846 , n469 );
xor ( n16854 , n16852 , n16853 );
not ( n16855 , n15274 );
not ( n16856 , n15286 );
or ( n16857 , n16855 , n16856 );
or ( n16858 , n15286 , n15274 );
nand ( n16859 , n16857 , n16858 );
not ( n16860 , n16773 );
not ( n16861 , n15163 );
or ( n16862 , n16860 , n16861 );
nand ( n16863 , n16862 , n15299 );
xnor ( n16864 , n16859 , n16863 );
not ( n16865 , n16864 );
not ( n16866 , n10190 );
or ( n16867 , n16865 , n16866 );
buf ( n16868 , n8338 );
buf ( n16869 , n8277 );
nand ( n16870 , n16868 , n16869 );
not ( n16871 , n454 );
nor ( n16872 , n16870 , n16871 );
buf ( n16873 , n9399 );
or ( n16874 , n16872 , n16873 );
not ( n16875 , n454 );
not ( n16876 , n16870 );
or ( n16877 , n16875 , n16876 );
nand ( n16878 , n16877 , n16873 );
nand ( n16879 , n16874 , n16878 );
nand ( n16880 , n16867 , n16879 );
and ( n16881 , n16880 , n472 );
xor ( n16882 , n16854 , n16881 );
xor ( n16883 , n16851 , n16882 );
and ( n16884 , n16786 , n472 );
nand ( n16885 , n16788 , n16797 );
not ( n16886 , n16885 );
and ( n16887 , n16794 , n16886 );
not ( n16888 , n16794 );
and ( n16889 , n16888 , n16885 );
nor ( n16890 , n16887 , n16889 );
nand ( n16891 , n16890 , n454 );
nand ( n16892 , n16808 , n15149 );
xnor ( n16893 , n16810 , n16892 );
nand ( n16894 , n16893 , n10190 );
nand ( n16895 , n16891 , n16894 );
and ( n16896 , n16895 , n469 );
and ( n16897 , n16817 , n470 );
xor ( n16898 , n16896 , n16897 );
and ( n16899 , n16835 , n472 );
and ( n16900 , n16898 , n16899 );
and ( n16901 , n16896 , n16897 );
or ( n16902 , n16900 , n16901 );
xor ( n16903 , n16884 , n16902 );
xor ( n16904 , n16818 , n16836 );
xor ( n16905 , n16904 , n16847 );
and ( n16906 , n16903 , n16905 );
and ( n16907 , n16884 , n16902 );
or ( n16908 , n16906 , n16907 );
nor ( n16909 , n16883 , n16908 );
xor ( n16910 , n16884 , n16902 );
xor ( n16911 , n16910 , n16905 );
and ( n16912 , n16846 , n471 );
nand ( n16913 , n9318 , n8832 );
not ( n16914 , n16913 );
buf ( n16915 , n9314 );
not ( n16916 , n16915 );
or ( n16917 , n16914 , n16916 );
or ( n16918 , n16915 , n16913 );
nand ( n16919 , n16917 , n16918 );
nand ( n16920 , n16919 , n454 );
not ( n16921 , n15141 );
nand ( n16922 , n16921 , n15138 );
not ( n16923 , n16922 );
not ( n16924 , n14729 );
not ( n16925 , n16924 );
buf ( n16926 , n15135 );
not ( n16927 , n16926 );
or ( n16928 , n16925 , n16927 );
not ( n16929 , n15139 );
nand ( n16930 , n16928 , n16929 );
not ( n16931 , n16930 );
or ( n16932 , n16923 , n16931 );
or ( n16933 , n16922 , n16930 );
nand ( n16934 , n16932 , n16933 );
nand ( n16935 , n10190 , n16934 );
nand ( n16936 , n16920 , n16935 );
and ( n16937 , n16936 , n469 );
and ( n16938 , n16895 , n470 );
xor ( n16939 , n16937 , n16938 );
and ( n16940 , n16817 , n471 );
and ( n16941 , n16939 , n16940 );
and ( n16942 , n16937 , n16938 );
or ( n16943 , n16941 , n16942 );
xor ( n16944 , n16912 , n16943 );
xor ( n16945 , n16896 , n16897 );
xor ( n16946 , n16945 , n16899 );
and ( n16947 , n16944 , n16946 );
and ( n16948 , n16912 , n16943 );
or ( n16949 , n16947 , n16948 );
nor ( n16950 , n16911 , n16949 );
nor ( n16951 , n16909 , n16950 );
not ( n16952 , n16951 );
not ( n16953 , n16952 );
xor ( n16954 , n16912 , n16943 );
xor ( n16955 , n16954 , n16946 );
and ( n16956 , n16846 , n472 );
not ( n16957 , n8893 );
not ( n16958 , n8948 );
nand ( n16959 , n16957 , n16958 );
not ( n16960 , n16959 );
buf ( n16961 , n9303 );
not ( n16962 , n16961 );
or ( n16963 , n16960 , n16962 );
nand ( n16964 , n8893 , n8948 );
nand ( n16965 , n16963 , n16964 );
not ( n16966 , n16965 );
not ( n16967 , n9312 );
nand ( n16968 , n16967 , n9308 );
nor ( n16969 , n16968 , n16731 );
nand ( n16970 , n16966 , n16969 );
and ( n16971 , n16968 , n454 );
and ( n16972 , n16965 , n16971 );
nand ( n16973 , n16929 , n16924 );
xnor ( n16974 , n16926 , n16973 );
and ( n16975 , n16974 , n10190 );
nor ( n16976 , n16972 , n16975 );
nand ( n16977 , n16970 , n16976 );
and ( n16978 , n16977 , n469 );
and ( n16979 , n16936 , n470 );
xor ( n16980 , n16978 , n16979 );
and ( n16981 , n16895 , n471 );
and ( n16982 , n16980 , n16981 );
and ( n16983 , n16978 , n16979 );
or ( n16984 , n16982 , n16983 );
xor ( n16985 , n16956 , n16984 );
xor ( n16986 , n16937 , n16938 );
xor ( n16987 , n16986 , n16940 );
and ( n16988 , n16985 , n16987 );
and ( n16989 , n16956 , n16984 );
or ( n16990 , n16988 , n16989 );
or ( n16991 , n16955 , n16990 );
not ( n16992 , n16991 );
not ( n16993 , n10190 );
not ( n16994 , n14777 );
and ( n16995 , n15131 , n16994 );
not ( n16996 , n15134 );
and ( n16997 , n15131 , n16996 );
nor ( n16998 , n16995 , n16997 );
not ( n16999 , n14772 );
not ( n17000 , n15131 );
nand ( n17001 , n16999 , n17000 , n14775 );
not ( n17002 , n14775 );
nand ( n17003 , n17002 , n17000 , n14772 );
nand ( n17004 , n16998 , n17001 , n17003 );
not ( n17005 , n17004 );
or ( n17006 , n16993 , n17005 );
nand ( n17007 , n16959 , n16964 );
not ( n17008 , n9303 );
and ( n17009 , n17007 , n17008 );
not ( n17010 , n17007 );
and ( n17011 , n17010 , n16961 );
nor ( n17012 , n17009 , n17011 );
nand ( n17013 , n17012 , n454 );
nand ( n17014 , n17006 , n17013 );
and ( n17015 , n17014 , n469 );
and ( n17016 , n16977 , n470 );
xor ( n17017 , n17015 , n17016 );
and ( n17018 , n16936 , n471 );
and ( n17019 , n17017 , n17018 );
and ( n17020 , n17015 , n17016 );
or ( n17021 , n17019 , n17020 );
and ( n17022 , n16817 , n472 );
xor ( n17023 , n17021 , n17022 );
xor ( n17024 , n16978 , n16979 );
xor ( n17025 , n17024 , n16981 );
and ( n17026 , n17023 , n17025 );
and ( n17027 , n17021 , n17022 );
or ( n17028 , n17026 , n17027 );
not ( n17029 , n17028 );
xor ( n17030 , n16956 , n16984 );
xor ( n17031 , n17030 , n16987 );
not ( n17032 , n17031 );
nand ( n17033 , n17029 , n17032 );
not ( n17034 , n17033 );
xor ( n17035 , n17021 , n17022 );
xor ( n17036 , n17035 , n17025 );
and ( n17037 , n16895 , n472 );
nand ( n17038 , n9302 , n9013 );
buf ( n17039 , n9299 );
not ( n17040 , n17039 );
and ( n17041 , n17038 , n17040 );
not ( n17042 , n17038 );
and ( n17043 , n17042 , n17039 );
nor ( n17044 , n17041 , n17043 );
nand ( n17045 , n17044 , n454 );
nand ( n17046 , n14828 , n15130 );
xnor ( n17047 , n15127 , n17046 );
nand ( n17048 , n17047 , n10190 );
nand ( n17049 , n17045 , n17048 );
and ( n17050 , n17049 , n469 );
and ( n17051 , n17014 , n470 );
xor ( n17052 , n17050 , n17051 );
and ( n17053 , n16977 , n471 );
and ( n17054 , n17052 , n17053 );
and ( n17055 , n17050 , n17051 );
or ( n17056 , n17054 , n17055 );
xor ( n17057 , n17037 , n17056 );
xor ( n17058 , n17015 , n17016 );
xor ( n17059 , n17058 , n17018 );
and ( n17060 , n17057 , n17059 );
and ( n17061 , n17037 , n17056 );
or ( n17062 , n17060 , n17061 );
or ( n17063 , n17036 , n17062 );
not ( n17064 , n17063 );
and ( n17065 , n16936 , n472 );
not ( n17066 , n10190 );
nand ( n17067 , n15123 , n15126 );
xnor ( n17068 , n17067 , n15113 );
not ( n17069 , n17068 );
or ( n17070 , n17066 , n17069 );
not ( n17071 , n9016 );
not ( n17072 , n9052 );
nand ( n17073 , n17071 , n17072 );
nand ( n17074 , n17073 , n9298 );
not ( n17075 , n9116 );
not ( n17076 , n9292 );
or ( n17077 , n17075 , n17076 );
not ( n17078 , n9295 );
nand ( n17079 , n17077 , n17078 );
not ( n17080 , n17079 );
and ( n17081 , n17074 , n17080 );
not ( n17082 , n17074 );
and ( n17083 , n17082 , n17079 );
nor ( n17084 , n17081 , n17083 );
nand ( n17085 , n17084 , n454 );
nand ( n17086 , n17070 , n17085 );
and ( n17087 , n17086 , n469 );
and ( n17088 , n17049 , n470 );
xor ( n17089 , n17087 , n17088 );
and ( n17090 , n17014 , n471 );
and ( n17091 , n17089 , n17090 );
and ( n17092 , n17087 , n17088 );
or ( n17093 , n17091 , n17092 );
xor ( n17094 , n17065 , n17093 );
xor ( n17095 , n17050 , n17051 );
xor ( n17096 , n17095 , n17053 );
and ( n17097 , n17094 , n17096 );
and ( n17098 , n17065 , n17093 );
or ( n17099 , n17097 , n17098 );
not ( n17100 , n17099 );
xor ( n17101 , n17037 , n17056 );
xor ( n17102 , n17101 , n17059 );
not ( n17103 , n17102 );
nand ( n17104 , n17100 , n17103 );
not ( n17105 , n17104 );
xor ( n17106 , n17065 , n17093 );
xor ( n17107 , n17106 , n17096 );
not ( n17108 , n17107 );
and ( n17109 , n16977 , n472 );
nand ( n17110 , n9116 , n9294 );
not ( n17111 , n17110 );
xor ( n17112 , n9292 , n17111 );
not ( n17113 , n17112 );
not ( n17114 , n454 );
or ( n17115 , n17113 , n17114 );
not ( n17116 , n15088 );
nand ( n17117 , n15109 , n15112 );
not ( n17118 , n17117 );
or ( n17119 , n17116 , n17118 );
or ( n17120 , n17117 , n15088 );
nand ( n17121 , n17119 , n17120 );
nand ( n17122 , n17121 , n10190 );
nand ( n17123 , n17115 , n17122 );
and ( n17124 , n17123 , n469 );
and ( n17125 , n17086 , n470 );
xor ( n17126 , n17124 , n17125 );
and ( n17127 , n17049 , n471 );
and ( n17128 , n17126 , n17127 );
and ( n17129 , n17124 , n17125 );
or ( n17130 , n17128 , n17129 );
xor ( n17131 , n17109 , n17130 );
xor ( n17132 , n17087 , n17088 );
xor ( n17133 , n17132 , n17090 );
and ( n17134 , n17131 , n17133 );
and ( n17135 , n17109 , n17130 );
or ( n17136 , n17134 , n17135 );
not ( n17137 , n17136 );
nand ( n17138 , n17108 , n17137 );
not ( n17139 , n17138 );
xor ( n17140 , n17109 , n17130 );
xor ( n17141 , n17140 , n17133 );
not ( n17142 , n17141 );
and ( n17143 , n17014 , n472 );
not ( n17144 , n10190 );
not ( n17145 , n15084 );
nand ( n17146 , n14928 , n15087 );
not ( n17147 , n17146 );
or ( n17148 , n17145 , n17147 );
or ( n17149 , n17146 , n15084 );
nand ( n17150 , n17148 , n17149 );
not ( n17151 , n17150 );
or ( n17152 , n17144 , n17151 );
xnor ( n17153 , n9138 , n9118 );
buf ( n17154 , n9289 );
and ( n17155 , n17153 , n17154 );
not ( n17156 , n17153 );
not ( n17157 , n17154 );
and ( n17158 , n17156 , n17157 );
nor ( n17159 , n17155 , n17158 );
nand ( n17160 , n17159 , n454 );
nand ( n17161 , n17152 , n17160 );
and ( n17162 , n17161 , n469 );
and ( n17163 , n17123 , n470 );
xor ( n17164 , n17162 , n17163 );
and ( n17165 , n17086 , n471 );
and ( n17166 , n17164 , n17165 );
and ( n17167 , n17162 , n17163 );
or ( n17168 , n17166 , n17167 );
xor ( n17169 , n17143 , n17168 );
xor ( n17170 , n17124 , n17125 );
xor ( n17171 , n17170 , n17127 );
and ( n17172 , n17169 , n17171 );
and ( n17173 , n17143 , n17168 );
or ( n17174 , n17172 , n17173 );
not ( n17175 , n17174 );
nand ( n17176 , n17142 , n17175 );
not ( n17177 , n17176 );
xor ( n17178 , n17143 , n17168 );
xor ( n17179 , n17178 , n17171 );
not ( n17180 , n17179 );
and ( n17181 , n17049 , n472 );
not ( n17182 , n10190 );
xor ( n17183 , n14953 , n14955 );
xor ( n17184 , n17183 , n15081 );
not ( n17185 , n17184 );
or ( n17186 , n17182 , n17185 );
not ( n17187 , n9160 );
nand ( n17188 , n17187 , n9164 );
and ( n17189 , n17188 , n9287 );
and ( n17190 , n17189 , n9285 );
not ( n17191 , n17189 );
not ( n17192 , n9285 );
and ( n17193 , n17191 , n17192 );
nor ( n17194 , n17190 , n17193 );
nand ( n17195 , n454 , n17194 );
nand ( n17196 , n17186 , n17195 );
and ( n17197 , n17196 , n469 );
and ( n17198 , n17161 , n470 );
xor ( n17199 , n17197 , n17198 );
and ( n17200 , n17123 , n471 );
and ( n17201 , n17199 , n17200 );
and ( n17202 , n17197 , n17198 );
or ( n17203 , n17201 , n17202 );
xor ( n17204 , n17181 , n17203 );
xor ( n17205 , n17162 , n17163 );
xor ( n17206 , n17205 , n17165 );
and ( n17207 , n17204 , n17206 );
and ( n17208 , n17181 , n17203 );
or ( n17209 , n17207 , n17208 );
not ( n17210 , n17209 );
nand ( n17211 , n17180 , n17210 );
not ( n17212 , n17211 );
xor ( n17213 , n17181 , n17203 );
xor ( n17214 , n17213 , n17206 );
not ( n17215 , n17214 );
nand ( n17216 , n9281 , n9284 );
not ( n17217 , n9271 );
and ( n17218 , n17216 , n17217 );
not ( n17219 , n17216 );
and ( n17220 , n17219 , n9271 );
nor ( n17221 , n17218 , n17220 );
not ( n17222 , n17221 );
not ( n17223 , n454 );
or ( n17224 , n17222 , n17223 );
xor ( n17225 , n14994 , n15075 );
xor ( n17226 , n17225 , n15078 );
nand ( n17227 , n17226 , n10190 );
nand ( n17228 , n17224 , n17227 );
and ( n17229 , n17228 , n469 );
and ( n17230 , n17196 , n470 );
xor ( n17231 , n17229 , n17230 );
nand ( n17232 , n17228 , n470 );
not ( n17233 , n454 );
not ( n17234 , n9268 );
nand ( n17235 , n17234 , n9270 );
xor ( n17236 , n9251 , n17235 );
not ( n17237 , n17236 );
or ( n17238 , n17233 , n17237 );
not ( n17239 , n15072 );
or ( n17240 , n14996 , n15006 );
nand ( n17241 , n17240 , n15074 );
not ( n17242 , n17241 );
or ( n17243 , n17239 , n17242 );
or ( n17244 , n17241 , n15072 );
nand ( n17245 , n17243 , n17244 );
nand ( n17246 , n17245 , n10190 );
nand ( n17247 , n17238 , n17246 );
nand ( n17248 , n17247 , n469 );
nor ( n17249 , n17232 , n17248 );
and ( n17250 , n17231 , n17249 );
and ( n17251 , n17229 , n17230 );
or ( n17252 , n17250 , n17251 );
and ( n17253 , n17086 , n472 );
xor ( n17254 , n17252 , n17253 );
and ( n17255 , n17161 , n471 );
not ( n17256 , n17196 );
not ( n17257 , n471 );
nor ( n17258 , n17256 , n17257 );
not ( n17259 , n17248 );
not ( n17260 , n17259 );
not ( n17261 , n17232 );
or ( n17262 , n17260 , n17261 );
nand ( n17263 , n17248 , n470 , n17228 );
nand ( n17264 , n17262 , n17263 );
xor ( n17265 , n17258 , n17264 );
and ( n17266 , n17228 , n471 );
not ( n17267 , n17266 );
nand ( n17268 , n470 , n17247 );
nor ( n17269 , n17267 , n17268 );
and ( n17270 , n17265 , n17269 );
and ( n17271 , n17258 , n17264 );
or ( n17272 , n17270 , n17271 );
xor ( n17273 , n17255 , n17272 );
and ( n17274 , n17123 , n472 );
and ( n17275 , n17273 , n17274 );
and ( n17276 , n17255 , n17272 );
or ( n17277 , n17275 , n17276 );
and ( n17278 , n17254 , n17277 );
and ( n17279 , n17252 , n17253 );
or ( n17280 , n17278 , n17279 );
not ( n17281 , n17280 );
nand ( n17282 , n17215 , n17281 );
not ( n17283 , n17282 );
xor ( n17284 , n17252 , n17253 );
xor ( n17285 , n17284 , n17277 );
xor ( n17286 , n17197 , n17198 );
xor ( n17287 , n17286 , n17200 );
nor ( n17288 , n17285 , n17287 );
and ( n17289 , n17161 , n472 );
xor ( n17290 , n17258 , n17264 );
xor ( n17291 , n17290 , n17269 );
xor ( n17292 , n17289 , n17291 );
not ( n17293 , n17266 );
not ( n17294 , n17268 );
or ( n17295 , n17293 , n17294 );
or ( n17296 , n17268 , n17266 );
nand ( n17297 , n17295 , n17296 );
not ( n17298 , n17297 );
not ( n17299 , n472 );
nor ( n17300 , n17299 , n17256 );
not ( n17301 , n17300 );
nand ( n17302 , n17228 , n17247 , n471 , n472 );
nand ( n17303 , n17301 , n17302 );
not ( n17304 , n17303 );
or ( n17305 , n17298 , n17304 );
not ( n17306 , n17302 );
nand ( n17307 , n17306 , n17300 );
nand ( n17308 , n17305 , n17307 );
and ( n17309 , n17292 , n17308 );
and ( n17310 , n17289 , n17291 );
or ( n17311 , n17309 , n17310 );
xor ( n17312 , n17255 , n17272 );
xor ( n17313 , n17312 , n17274 );
not ( n17314 , n17313 );
xor ( n17315 , n17229 , n17230 );
xor ( n17316 , n17315 , n17249 );
not ( n17317 , n17316 );
nand ( n17318 , n17314 , n17317 );
and ( n17319 , n17311 , n17318 );
nor ( n17320 , n17314 , n17317 );
nor ( n17321 , n17319 , n17320 );
or ( n17322 , n17288 , n17321 );
nand ( n17323 , n17285 , n17287 );
nand ( n17324 , n17322 , n17323 );
not ( n17325 , n17324 );
or ( n17326 , n17283 , n17325 );
nand ( n17327 , n17214 , n17280 );
nand ( n17328 , n17326 , n17327 );
not ( n17329 , n17328 );
or ( n17330 , n17212 , n17329 );
nand ( n17331 , n17179 , n17209 );
nand ( n17332 , n17330 , n17331 );
not ( n17333 , n17332 );
or ( n17334 , n17177 , n17333 );
nand ( n17335 , n17141 , n17174 );
nand ( n17336 , n17334 , n17335 );
not ( n17337 , n17336 );
or ( n17338 , n17139 , n17337 );
nand ( n17339 , n17107 , n17136 );
nand ( n17340 , n17338 , n17339 );
not ( n17341 , n17340 );
or ( n17342 , n17105 , n17341 );
nand ( n17343 , n17102 , n17099 );
nand ( n17344 , n17342 , n17343 );
not ( n17345 , n17344 );
or ( n17346 , n17064 , n17345 );
nand ( n17347 , n17036 , n17062 );
nand ( n17348 , n17346 , n17347 );
not ( n17349 , n17348 );
or ( n17350 , n17034 , n17349 );
not ( n17351 , n17032 );
nand ( n17352 , n17351 , n17028 );
nand ( n17353 , n17350 , n17352 );
not ( n17354 , n17353 );
or ( n17355 , n16992 , n17354 );
nand ( n17356 , n16955 , n16990 );
nand ( n17357 , n17355 , n17356 );
and ( n17358 , n16758 , n472 );
buf ( n17359 , n8308 );
nand ( n17360 , n17359 , n8330 );
not ( n17361 , n17360 );
not ( n17362 , n9399 );
not ( n17363 , n16738 );
or ( n17364 , n17362 , n17363 );
nand ( n17365 , n17364 , n16741 );
not ( n17366 , n17365 );
or ( n17367 , n17361 , n17366 );
or ( n17368 , n17360 , n16742 );
nand ( n17369 , n17367 , n17368 );
nand ( n17370 , n17369 , n454 );
not ( n17371 , n15337 );
nand ( n17372 , n17371 , n15357 );
not ( n17373 , n17372 );
not ( n17374 , n17373 );
not ( n17375 , n15163 );
not ( n17376 , n15295 );
or ( n17377 , n17375 , n17376 );
not ( n17378 , n15287 );
not ( n17379 , n15299 );
and ( n17380 , n17378 , n17379 );
nor ( n17381 , n17380 , n15302 );
nand ( n17382 , n17377 , n17381 );
not ( n17383 , n17382 );
not ( n17384 , n15344 );
buf ( n17385 , n17384 );
not ( n17386 , n17385 );
or ( n17387 , n17383 , n17386 );
buf ( n17388 , n15355 );
nand ( n17389 , n17387 , n17388 );
not ( n17390 , n17389 );
or ( n17391 , n17374 , n17390 );
nand ( n17392 , n17382 , n17385 );
and ( n17393 , n17392 , n17372 , n17388 );
nor ( n17394 , n17393 , n454 );
nand ( n17395 , n17391 , n17394 );
and ( n17396 , n17370 , n17395 );
not ( n17397 , n470 );
nor ( n17398 , n17396 , n17397 );
nand ( n17399 , n17384 , n15355 );
not ( n17400 , n17399 );
not ( n17401 , n17382 );
or ( n17402 , n17400 , n17401 );
or ( n17403 , n17382 , n17399 );
nand ( n17404 , n17402 , n17403 );
nand ( n17405 , n17404 , n10190 );
not ( n17406 , n17405 );
nand ( n17407 , n8335 , n8279 );
not ( n17408 , n17407 );
not ( n17409 , n16868 );
not ( n17410 , n9399 );
or ( n17411 , n17409 , n17410 );
nand ( n17412 , n17411 , n16869 );
not ( n17413 , n17412 );
or ( n17414 , n17408 , n17413 );
or ( n17415 , n17407 , n17412 );
nand ( n17416 , n17414 , n17415 );
nand ( n17417 , n17416 , n454 );
not ( n17418 , n17417 );
or ( n17419 , n17406 , n17418 );
nand ( n17420 , n17419 , n469 );
not ( n17421 , n17420 );
xor ( n17422 , n17398 , n17421 );
buf ( n17423 , n8313 );
not ( n17424 , n8327 );
nor ( n17425 , n17423 , n17424 );
not ( n17426 , n17359 );
nor ( n17427 , n17425 , n17426 );
buf ( n17428 , n8330 );
nand ( n17429 , n17365 , n17428 );
and ( n17430 , n17427 , n17429 );
nor ( n17431 , n17430 , n16731 );
not ( n17432 , n17431 );
not ( n17433 , n17359 );
not ( n17434 , n17429 );
or ( n17435 , n17433 , n17434 );
buf ( n17436 , n17425 );
nand ( n17437 , n17435 , n17436 );
not ( n17438 , n17437 );
or ( n17439 , n17432 , n17438 );
nand ( n17440 , n15353 , n15364 );
not ( n17441 , n17440 );
not ( n17442 , n16002 );
or ( n17443 , n17441 , n17442 );
or ( n17444 , n16002 , n17440 );
nand ( n17445 , n17443 , n17444 );
nand ( n17446 , n17445 , n10190 );
nand ( n17447 , n17439 , n17446 );
and ( n17448 , n17447 , n471 );
and ( n17449 , n17422 , n17448 );
and ( n17450 , n17398 , n17421 );
or ( n17451 , n17449 , n17450 );
xor ( n17452 , n17358 , n17451 );
nand ( n17453 , n17370 , n17395 );
and ( n17454 , n17453 , n469 );
and ( n17455 , n17447 , n470 );
xor ( n17456 , n17454 , n17455 );
not ( n17457 , n454 );
nand ( n17458 , n16733 , n8320 );
not ( n17459 , n17458 );
and ( n17460 , n16746 , n17459 );
not ( n17461 , n16746 );
and ( n17462 , n17461 , n17458 );
nor ( n17463 , n17460 , n17462 );
not ( n17464 , n17463 );
or ( n17465 , n17457 , n17464 );
not ( n17466 , n15353 );
not ( n17467 , n16002 );
or ( n17468 , n17466 , n17467 );
nand ( n17469 , n17468 , n15364 );
not ( n17470 , n13803 );
nor ( n17471 , n17470 , n15367 );
xor ( n17472 , n17469 , n17471 );
nand ( n17473 , n17472 , n10190 );
nand ( n17474 , n17465 , n17473 );
and ( n17475 , n17474 , n471 );
xor ( n17476 , n17456 , n17475 );
xor ( n17477 , n17452 , n17476 );
not ( n17478 , n17477 );
and ( n17479 , n17474 , n472 );
and ( n17480 , n16880 , n469 );
not ( n17481 , n17453 );
nor ( n17482 , n17481 , n17257 );
xor ( n17483 , n17480 , n17482 );
nand ( n17484 , n17417 , n17405 );
and ( n17485 , n17484 , n470 );
and ( n17486 , n17483 , n17485 );
and ( n17487 , n17480 , n17482 );
or ( n17488 , n17486 , n17487 );
xor ( n17489 , n17479 , n17488 );
xor ( n17490 , n17398 , n17421 );
xor ( n17491 , n17490 , n17448 );
and ( n17492 , n17489 , n17491 );
and ( n17493 , n17479 , n17488 );
or ( n17494 , n17492 , n17493 );
not ( n17495 , n17494 );
nand ( n17496 , n17478 , n17495 );
and ( n17497 , n17484 , n471 );
and ( n17498 , n16835 , n469 );
and ( n17499 , n16880 , n471 );
xor ( n17500 , n17498 , n17499 );
not ( n17501 , n16786 );
nor ( n17502 , n17501 , n17397 );
and ( n17503 , n17500 , n17502 );
and ( n17504 , n17498 , n17499 );
or ( n17505 , n17503 , n17504 );
xor ( n17506 , n17497 , n17505 );
and ( n17507 , n16880 , n470 );
and ( n17508 , n16786 , n469 );
xor ( n17509 , n17507 , n17508 );
and ( n17510 , n17453 , n472 );
xor ( n17511 , n17509 , n17510 );
xor ( n17512 , n17506 , n17511 );
not ( n17513 , n17512 );
and ( n17514 , n17484 , n472 );
xor ( n17515 , n16852 , n16853 );
and ( n17516 , n17515 , n16881 );
and ( n17517 , n16852 , n16853 );
or ( n17518 , n17516 , n17517 );
xor ( n17519 , n17514 , n17518 );
xor ( n17520 , n17498 , n17499 );
xor ( n17521 , n17520 , n17502 );
and ( n17522 , n17519 , n17521 );
and ( n17523 , n17514 , n17518 );
or ( n17524 , n17522 , n17523 );
not ( n17525 , n17524 );
and ( n17526 , n17513 , n17525 );
xor ( n17527 , n17514 , n17518 );
xor ( n17528 , n17527 , n17521 );
xor ( n17529 , n16787 , n16850 );
and ( n17530 , n17529 , n16882 );
and ( n17531 , n16787 , n16850 );
or ( n17532 , n17530 , n17531 );
nor ( n17533 , n17528 , n17532 );
nor ( n17534 , n17526 , n17533 );
nand ( n17535 , n16953 , n17357 , n17496 , n17534 );
not ( n17536 , n17535 );
and ( n17537 , n16758 , n471 );
xor ( n17538 , n17454 , n17455 );
and ( n17539 , n17538 , n17475 );
and ( n17540 , n17454 , n17455 );
or ( n17541 , n17539 , n17540 );
xor ( n17542 , n17537 , n17541 );
not ( n17543 , n17431 );
not ( n17544 , n17437 );
or ( n17545 , n17543 , n17544 );
nand ( n17546 , n17545 , n17446 );
and ( n17547 , n17546 , n469 );
and ( n17548 , n17474 , n470 );
xor ( n17549 , n17547 , n17548 );
and ( n17550 , n16019 , n472 );
xor ( n17551 , n17549 , n17550 );
xor ( n17552 , n17542 , n17551 );
not ( n17553 , n17552 );
xor ( n17554 , n17358 , n17451 );
and ( n17555 , n17554 , n17476 );
and ( n17556 , n17358 , n17451 );
or ( n17557 , n17555 , n17556 );
not ( n17558 , n17557 );
and ( n17559 , n17553 , n17558 );
and ( n17560 , n17546 , n472 );
xor ( n17561 , n17507 , n17508 );
and ( n17562 , n17561 , n17510 );
and ( n17563 , n17507 , n17508 );
or ( n17564 , n17562 , n17563 );
xor ( n17565 , n17560 , n17564 );
xor ( n17566 , n17480 , n17482 );
xor ( n17567 , n17566 , n17485 );
and ( n17568 , n17565 , n17567 );
and ( n17569 , n17560 , n17564 );
or ( n17570 , n17568 , n17569 );
not ( n17571 , n17570 );
not ( n17572 , n17571 );
xor ( n17573 , n17479 , n17488 );
xor ( n17574 , n17573 , n17491 );
not ( n17575 , n17574 );
not ( n17576 , n17575 );
or ( n17577 , n17572 , n17576 );
xor ( n17578 , n17560 , n17564 );
xor ( n17579 , n17578 , n17567 );
not ( n17580 , n17579 );
xor ( n17581 , n17497 , n17505 );
and ( n17582 , n17581 , n17511 );
and ( n17583 , n17497 , n17505 );
or ( n17584 , n17582 , n17583 );
not ( n17585 , n17584 );
nand ( n17586 , n17580 , n17585 );
nand ( n17587 , n17577 , n17586 );
nor ( n17588 , n17559 , n17587 );
nand ( n17589 , n17536 , n17588 );
nand ( n17590 , n17553 , n17558 );
and ( n17591 , n17477 , n17494 );
nand ( n17592 , n17590 , n17591 );
buf ( n17593 , n17552 );
nand ( n17594 , n17593 , n17557 );
buf ( n17595 , n17496 );
not ( n17596 , n17571 );
not ( n17597 , n17575 );
or ( n17598 , n17596 , n17597 );
nand ( n17599 , n17598 , n17586 );
not ( n17600 , n17599 );
not ( n17601 , n17600 );
nand ( n17602 , n16911 , n16949 );
or ( n17603 , n16909 , n17602 );
nand ( n17604 , n16883 , n16908 );
nand ( n17605 , n17603 , n17604 );
not ( n17606 , n17605 );
not ( n17607 , n17534 );
or ( n17608 , n17606 , n17607 );
not ( n17609 , n17512 );
not ( n17610 , n17524 );
nand ( n17611 , n17609 , n17610 );
and ( n17612 , n17528 , n17532 );
and ( n17613 , n17611 , n17612 );
not ( n17614 , n17512 );
nor ( n17615 , n17614 , n17610 );
nor ( n17616 , n17613 , n17615 );
nand ( n17617 , n17608 , n17616 );
not ( n17618 , n17617 );
or ( n17619 , n17601 , n17618 );
nand ( n17620 , n17575 , n17571 );
and ( n17621 , n17579 , n17584 );
and ( n17622 , n17620 , n17621 );
and ( n17623 , n17574 , n17570 );
nor ( n17624 , n17622 , n17623 );
nand ( n17625 , n17619 , n17624 );
nand ( n17626 , n17595 , n17625 , n17590 );
nand ( n17627 , n17589 , n17592 , n17594 , n17626 );
xor ( n17628 , n16728 , n16764 );
xor ( n17629 , n17628 , n16767 );
not ( n17630 , n17629 );
and ( n17631 , n16072 , n471 );
and ( n17632 , n17474 , n469 );
not ( n17633 , n16019 );
nor ( n17634 , n17633 , n17257 );
xor ( n17635 , n17632 , n17634 );
and ( n17636 , n16758 , n470 );
and ( n17637 , n17635 , n17636 );
and ( n17638 , n17632 , n17634 );
or ( n17639 , n17637 , n17638 );
xor ( n17640 , n17631 , n17639 );
xor ( n17641 , n16729 , n16759 );
xor ( n17642 , n17641 , n16761 );
and ( n17643 , n17640 , n17642 );
and ( n17644 , n17631 , n17639 );
or ( n17645 , n17643 , n17644 );
not ( n17646 , n17645 );
nand ( n17647 , n17630 , n17646 );
not ( n17648 , n17647 );
xor ( n17649 , n17631 , n17639 );
xor ( n17650 , n17649 , n17642 );
and ( n17651 , n16072 , n472 );
xor ( n17652 , n17547 , n17548 );
and ( n17653 , n17652 , n17550 );
and ( n17654 , n17547 , n17548 );
or ( n17655 , n17653 , n17654 );
xor ( n17656 , n17651 , n17655 );
xor ( n17657 , n17632 , n17634 );
xor ( n17658 , n17657 , n17636 );
and ( n17659 , n17656 , n17658 );
and ( n17660 , n17651 , n17655 );
or ( n17661 , n17659 , n17660 );
nor ( n17662 , n17650 , n17661 );
xor ( n17663 , n17651 , n17655 );
xor ( n17664 , n17663 , n17658 );
xor ( n17665 , n17537 , n17541 );
and ( n17666 , n17665 , n17551 );
and ( n17667 , n17537 , n17541 );
or ( n17668 , n17666 , n17667 );
nor ( n17669 , n17664 , n17668 );
nor ( n17670 , n17662 , n17669 );
not ( n17671 , n17670 );
nor ( n17672 , n17648 , n17671 );
nand ( n17673 , n16772 , n17627 , n17672 );
nand ( n17674 , n17664 , n17668 );
or ( n17675 , n17662 , n17674 );
nand ( n17676 , n17650 , n17661 );
nand ( n17677 , n17675 , n17676 );
and ( n17678 , n17647 , n17677 );
not ( n17679 , n17629 );
nor ( n17680 , n17679 , n17646 );
nor ( n17681 , n17678 , n17680 );
not ( n17682 , n17681 );
nand ( n17683 , n17682 , n16772 );
nand ( n17684 , n16727 , n16770 );
not ( n17685 , n17684 );
not ( n17686 , n16723 );
not ( n17687 , n16400 );
nand ( n17688 , n17686 , n17687 );
and ( n17689 , n17685 , n17688 );
and ( n17690 , n16723 , n16400 );
nor ( n17691 , n17689 , n17690 );
nand ( n17692 , n17673 , n17683 , n17691 );
and ( n17693 , n16710 , n471 );
xor ( n17694 , n16717 , n16719 );
and ( n17695 , n17694 , n16721 );
and ( n17696 , n16717 , n16719 );
or ( n17697 , n17695 , n17696 );
xor ( n17698 , n17693 , n17697 );
not ( n17699 , n454 );
not ( n17700 , n15807 );
not ( n17701 , n15801 );
or ( n17702 , n17700 , n17701 );
or ( n17703 , n16375 , n16379 );
nand ( n17704 , n16701 , n15977 , n17703 );
not ( n17705 , n17704 );
nand ( n17706 , n17702 , n17705 );
nand ( n17707 , n16380 , n16702 );
or ( n17708 , n17707 , n16533 );
nand ( n17709 , n17708 , n16701 );
buf ( n17710 , n17709 );
nand ( n17711 , n17706 , n17710 );
not ( n17712 , n13056 );
not ( n17713 , n16541 );
or ( n17714 , n17712 , n17713 );
and ( n17715 , n495 , n15599 );
not ( n17716 , n495 );
and ( n17717 , n17716 , n15602 );
or ( n17718 , n17715 , n17717 );
nand ( n17719 , n17718 , n13119 );
nand ( n17720 , n17714 , n17719 );
not ( n17721 , n15386 );
not ( n17722 , n16554 );
or ( n17723 , n17721 , n17722 );
not ( n17724 , n493 );
not ( n17725 , n12939 );
or ( n17726 , n17724 , n17725 );
nand ( n17727 , n13450 , n12862 );
nand ( n17728 , n17726 , n17727 );
nand ( n17729 , n17728 , n12845 );
nand ( n17730 , n17723 , n17729 );
xor ( n17731 , n17720 , n17730 );
not ( n17732 , n12789 );
not ( n17733 , n16596 );
or ( n17734 , n17732 , n17733 );
not ( n17735 , n499 );
not ( n17736 , n15727 );
or ( n17737 , n17735 , n17736 );
nand ( n17738 , n15720 , n12560 );
nand ( n17739 , n17737 , n17738 );
nand ( n17740 , n17739 , n12743 );
nand ( n17741 , n17734 , n17740 );
xor ( n17742 , n17731 , n17741 );
xor ( n17743 , n16548 , n16558 );
and ( n17744 , n17743 , n16572 );
and ( n17745 , n16548 , n16558 );
or ( n17746 , n17744 , n17745 );
xor ( n17747 , n17742 , n17746 );
xor ( n17748 , n16657 , n16661 );
and ( n17749 , n17748 , n16683 );
and ( n17750 , n16657 , n16661 );
or ( n17751 , n17749 , n17750 );
xor ( n17752 , n17747 , n17751 );
not ( n17753 , n12610 );
not ( n17754 , n497 );
not ( n17755 , n15474 );
or ( n17756 , n17754 , n17755 );
nand ( n17757 , n12511 , n12579 );
nand ( n17758 , n17756 , n17757 );
not ( n17759 , n17758 );
or ( n17760 , n17753 , n17759 );
not ( n17761 , n13339 );
not ( n17762 , n16583 );
and ( n17763 , n17761 , n17762 );
not ( n17764 , n13336 );
and ( n17765 , n17764 , n16580 );
nor ( n17766 , n17763 , n17765 );
nand ( n17767 , n17760 , n17766 );
not ( n17768 , n12909 );
not ( n17769 , n16570 );
or ( n17770 , n17768 , n17769 );
and ( n17771 , n16336 , n16278 );
not ( n17772 , n16336 );
and ( n17773 , n12930 , n501 );
and ( n17774 , n17772 , n17773 );
nor ( n17775 , n17771 , n17774 );
nand ( n17776 , n17770 , n17775 );
xor ( n17777 , n17767 , n17776 );
xor ( n17778 , n16663 , n16669 );
and ( n17779 , n17778 , n16682 );
and ( n17780 , n16663 , n16669 );
or ( n17781 , n17779 , n17780 );
xor ( n17782 , n17777 , n17781 );
not ( n17783 , n12555 );
not ( n17784 , n16653 );
or ( n17785 , n17783 , n17784 );
nand ( n17786 , n17785 , n699 );
not ( n17787 , n12688 );
not ( n17788 , n16664 );
or ( n17789 , n17787 , n17788 );
not ( n17790 , n491 );
not ( n17791 , n13438 );
or ( n17792 , n17790 , n17791 );
or ( n17793 , n491 , n13438 );
nand ( n17794 , n17792 , n17793 );
nand ( n17795 , n17794 , n12731 );
nand ( n17796 , n17789 , n17795 );
and ( n17797 , n16671 , n16681 );
xor ( n17798 , n17796 , n17797 );
nand ( n17799 , n489 , n13095 );
not ( n17800 , n17799 );
not ( n17801 , n12673 );
not ( n17802 , n489 );
not ( n17803 , n12575 );
or ( n17804 , n17802 , n17803 );
nand ( n17805 , n12574 , n12653 );
nand ( n17806 , n17804 , n17805 );
not ( n17807 , n17806 );
or ( n17808 , n17801 , n17807 );
nand ( n17809 , n16676 , n12635 );
nand ( n17810 , n17808 , n17809 );
not ( n17811 , n17810 );
or ( n17812 , n17800 , n17811 );
or ( n17813 , n17810 , n17799 );
nand ( n17814 , n17812 , n17813 );
xor ( n17815 , n17798 , n17814 );
xor ( n17816 , n17786 , n17815 );
xor ( n17817 , n16585 , n16589 );
and ( n17818 , n17817 , n16600 );
and ( n17819 , n16585 , n16589 );
or ( n17820 , n17818 , n17819 );
xor ( n17821 , n17816 , n17820 );
xor ( n17822 , n17782 , n17821 );
xor ( n17823 , n16573 , n16577 );
and ( n17824 , n17823 , n16601 );
and ( n17825 , n16573 , n16577 );
or ( n17826 , n17824 , n17825 );
xor ( n17827 , n17822 , n17826 );
xor ( n17828 , n17752 , n17827 );
xor ( n17829 , n16606 , n16684 );
and ( n17830 , n17829 , n16689 );
and ( n17831 , n16606 , n16684 );
or ( n17832 , n17830 , n17831 );
xor ( n17833 , n17828 , n17832 );
not ( n17834 , n17833 );
xor ( n17835 , n16602 , n16690 );
and ( n17836 , n17835 , n16695 );
and ( n17837 , n16602 , n16690 );
or ( n17838 , n17836 , n17837 );
not ( n17839 , n17838 );
nor ( n17840 , n17834 , n17839 );
not ( n17841 , n17840 );
not ( n17842 , n17833 );
nand ( n17843 , n17842 , n17839 );
buf ( n17844 , n17843 );
nand ( n17845 , n17841 , n17844 );
not ( n17846 , n17845 );
and ( n17847 , n17711 , n17846 );
not ( n17848 , n17711 );
and ( n17849 , n17848 , n17845 );
nor ( n17850 , n17847 , n17849 );
nand ( n17851 , n17699 , n17850 );
not ( n17852 , n16731 );
not ( n17853 , n16403 );
nor ( n17854 , n17853 , n16515 );
not ( n17855 , n17854 );
not ( n17856 , n10052 );
or ( n17857 , n17855 , n17856 );
buf ( n17858 , n16402 );
nor ( n17859 , n16515 , n17858 );
buf ( n17860 , n16407 );
and ( n17861 , n17859 , n17860 );
not ( n17862 , n16518 );
nor ( n17863 , n17861 , n17862 );
nand ( n17864 , n17857 , n17863 );
xor ( n17865 , n16428 , n16437 );
and ( n17866 , n17865 , n16442 );
and ( n17867 , n16428 , n16437 );
or ( n17868 , n17866 , n17867 );
not ( n17869 , n5786 );
not ( n17870 , n541 );
not ( n17871 , n7490 );
or ( n17872 , n17870 , n17871 );
nand ( n17873 , n6618 , n5734 );
nand ( n17874 , n17872 , n17873 );
not ( n17875 , n17874 );
or ( n17876 , n17869 , n17875 );
nand ( n17877 , n16426 , n10067 );
nand ( n17878 , n17876 , n17877 );
not ( n17879 , n4660 );
and ( n17880 , n7016 , n539 );
not ( n17881 , n7016 );
and ( n17882 , n17881 , n4477 );
or ( n17883 , n17880 , n17882 );
not ( n17884 , n17883 );
or ( n17885 , n17879 , n17884 );
and ( n17886 , n5588 , n4477 );
not ( n17887 , n5588 );
and ( n17888 , n17887 , n539 );
or ( n17889 , n17886 , n17888 );
nand ( n17890 , n17889 , n4450 );
nand ( n17891 , n17885 , n17890 );
xor ( n17892 , n17878 , n17891 );
not ( n17893 , n5595 );
not ( n17894 , n545 );
not ( n17895 , n9692 );
or ( n17896 , n17894 , n17895 );
nand ( n17897 , n16159 , n4666 );
nand ( n17898 , n17896 , n17897 );
not ( n17899 , n17898 );
or ( n17900 , n17893 , n17899 );
nand ( n17901 , n16433 , n5341 );
nand ( n17902 , n17900 , n17901 );
xor ( n17903 , n17892 , n17902 );
xor ( n17904 , n17868 , n17903 );
not ( n17905 , n5697 );
not ( n17906 , n537 );
not ( n17907 , n7544 );
or ( n17908 , n17906 , n17907 );
nand ( n17909 , n5466 , n5605 );
nand ( n17910 , n17908 , n17909 );
not ( n17911 , n17910 );
or ( n17912 , n17905 , n17911 );
nand ( n17913 , n16482 , n16173 );
nand ( n17914 , n17912 , n17913 );
not ( n17915 , n9730 );
not ( n17916 , n543 );
not ( n17917 , n9867 );
or ( n17918 , n17916 , n17917 );
nand ( n17919 , n9866 , n5146 );
nand ( n17920 , n17918 , n17919 );
not ( n17921 , n17920 );
or ( n17922 , n17915 , n17921 );
nand ( n17923 , n16461 , n4671 );
nand ( n17924 , n17922 , n17923 );
xor ( n17925 , n17914 , n17924 );
not ( n17926 , n6983 );
not ( n17927 , n547 );
not ( n17928 , n9977 );
or ( n17929 , n17927 , n17928 );
or ( n17930 , n9977 , n547 );
nand ( n17931 , n17929 , n17930 );
not ( n17932 , n17931 );
or ( n17933 , n17926 , n17932 );
nand ( n17934 , n16470 , n7026 );
nand ( n17935 , n17933 , n17934 );
xor ( n17936 , n17925 , n17935 );
xor ( n17937 , n17904 , n17936 );
or ( n17938 , n6667 , n6095 );
nand ( n17939 , n17938 , n549 );
and ( n17940 , n5145 , n537 );
xor ( n17941 , n17939 , n17940 );
not ( n17942 , n16485 );
xor ( n17943 , n17941 , n17942 );
xor ( n17944 , n16484 , n16485 );
and ( n17945 , n17944 , n16181 );
and ( n17946 , n16484 , n16485 );
or ( n17947 , n17945 , n17946 );
xor ( n17948 , n17943 , n17947 );
xor ( n17949 , n16455 , n16465 );
and ( n17950 , n17949 , n16472 );
and ( n17951 , n16455 , n16465 );
or ( n17952 , n17950 , n17951 );
xor ( n17953 , n17948 , n17952 );
xor ( n17954 , n16487 , n16491 );
and ( n17955 , n17954 , n16496 );
and ( n17956 , n16487 , n16491 );
or ( n17957 , n17955 , n17956 );
xor ( n17958 , n17953 , n17957 );
xor ( n17959 , n16418 , n16443 );
and ( n17960 , n17959 , n16473 );
and ( n17961 , n16418 , n16443 );
or ( n17962 , n17960 , n17961 );
xor ( n17963 , n17958 , n17962 );
xor ( n17964 , n17937 , n17963 );
xor ( n17965 , n16497 , n16501 );
and ( n17966 , n17965 , n16506 );
and ( n17967 , n16497 , n16501 );
or ( n17968 , n17966 , n17967 );
xor ( n17969 , n17964 , n17968 );
xor ( n17970 , n16474 , n16507 );
and ( n17971 , n17970 , n16512 );
and ( n17972 , n16474 , n16507 );
or ( n17973 , n17971 , n17972 );
nor ( n17974 , n17969 , n17973 );
not ( n17975 , n17974 );
buf ( n17976 , n17969 );
nand ( n17977 , n17976 , n17973 );
nand ( n17978 , n17975 , n17977 );
not ( n17979 , n17978 );
and ( n17980 , n17864 , n17979 );
not ( n17981 , n17864 );
and ( n17982 , n17981 , n17978 );
nor ( n17983 , n17980 , n17982 );
nand ( n17984 , n17852 , n17983 );
and ( n17985 , n17851 , n17984 );
nor ( n17986 , n17985 , n16395 );
and ( n17987 , n15982 , n469 );
xor ( n17988 , n17986 , n17987 );
nor ( n17989 , n16394 , n17397 );
xor ( n17990 , n17988 , n17989 );
xor ( n17991 , n17698 , n17990 );
xor ( n17992 , n16711 , n16715 );
and ( n17993 , n17992 , n16722 );
and ( n17994 , n16711 , n16715 );
or ( n17995 , n17993 , n17994 );
nor ( n17996 , n17991 , n17995 );
buf ( n17997 , n17996 );
not ( n17998 , n17997 );
nand ( n17999 , n17991 , n17995 );
nand ( n18000 , n17998 , n17999 );
not ( n18001 , n18000 );
and ( n18002 , n17692 , n18001 );
not ( n18003 , n17692 );
and ( n18004 , n18003 , n18000 );
or ( n18005 , n18002 , n18004 );
nor ( n18006 , n455 , n456 );
or ( n18007 , n18006 , n16871 );
or ( n18008 , n18005 , n18007 );
and ( n18009 , n536 , n6973 );
not ( n18010 , n536 );
and ( n18011 , n18010 , n552 );
or ( n18012 , n18009 , n18011 );
not ( n18013 , n18012 );
nand ( n18014 , n536 , n552 );
nand ( n18015 , n535 , n551 );
not ( n18016 , n18015 );
nor ( n18017 , n535 , n551 );
nor ( n18018 , n18016 , n18017 );
and ( n18019 , n18014 , n18018 );
not ( n18020 , n18014 );
not ( n18021 , n18018 );
and ( n18022 , n18020 , n18021 );
or ( n18023 , n18019 , n18022 );
nand ( n18024 , n18013 , n18023 );
not ( n18025 , n18024 );
not ( n18026 , n18025 );
not ( n18027 , n18023 );
buf ( n18028 , n18027 );
not ( n18029 , n18028 );
buf ( n18030 , n2373 );
xor ( n18031 , n2270 , n18030 );
not ( n18032 , n6206 );
not ( n18033 , n6303 );
or ( n18034 , n18032 , n18033 );
nand ( n18035 , n6304 , n2270 );
nand ( n18036 , n18034 , n18035 );
nor ( n18037 , n18031 , n18036 );
not ( n18038 , n18037 );
not ( n18039 , n18038 );
not ( n18040 , n18039 );
not ( n18041 , n6303 );
not ( n18042 , n18041 );
nor ( n18043 , n493 , n509 );
nor ( n18044 , n494 , n510 );
nor ( n18045 , n18043 , n18044 );
nor ( n18046 , n495 , n511 );
nor ( n18047 , n496 , n512 );
nor ( n18048 , n18046 , n18047 );
and ( n18049 , n18045 , n18048 );
not ( n18050 , n18049 );
nor ( n18051 , n498 , n514 );
not ( n18052 , n18051 );
not ( n18053 , n18052 );
or ( n18054 , n497 , n513 );
not ( n18055 , n18054 );
or ( n18056 , n18053 , n18055 );
nand ( n18057 , n497 , n513 );
nand ( n18058 , n18056 , n18057 );
not ( n18059 , n18058 );
nand ( n18060 , n500 , n516 );
nor ( n18061 , n499 , n515 );
or ( n18062 , n18060 , n18061 );
nand ( n18063 , n498 , n514 );
nand ( n18064 , n499 , n515 );
and ( n18065 , n18057 , n18063 , n18064 );
nand ( n18066 , n18062 , n18065 );
not ( n18067 , n18066 );
or ( n18068 , n18059 , n18067 );
nand ( n18069 , n501 , n517 );
nand ( n18070 , n502 , n518 );
and ( n18071 , n18069 , n18070 );
not ( n18072 , n18071 );
not ( n18073 , n504 );
not ( n18074 , n520 );
or ( n18075 , n18073 , n18074 );
nand ( n18076 , n503 , n519 );
nand ( n18077 , n18075 , n18076 );
nor ( n18078 , n503 , n519 );
not ( n18079 , n18078 );
not ( n18080 , n502 );
nand ( n18081 , n18080 , n758 );
nand ( n18082 , n18077 , n18079 , n18081 );
not ( n18083 , n18082 );
or ( n18084 , n18072 , n18083 );
or ( n18085 , n501 , n517 );
nand ( n18086 , n18054 , n18085 , n18052 );
or ( n18087 , n500 , n516 );
or ( n18088 , n499 , n515 );
nand ( n18089 , n18087 , n18088 );
nor ( n18090 , n18086 , n18089 );
nand ( n18091 , n18084 , n18090 );
nand ( n18092 , n18068 , n18091 );
not ( n18093 , n18092 );
or ( n18094 , n18050 , n18093 );
nor ( n18095 , n495 , n511 );
nand ( n18096 , n496 , n512 );
or ( n18097 , n18095 , n18096 );
nand ( n18098 , n495 , n511 );
nand ( n18099 , n18097 , n18098 );
not ( n18100 , n18099 );
not ( n18101 , n18045 );
or ( n18102 , n18100 , n18101 );
not ( n18103 , n18043 );
nand ( n18104 , n494 , n510 );
not ( n18105 , n18104 );
and ( n18106 , n18103 , n18105 );
nand ( n18107 , n493 , n509 );
not ( n18108 , n18107 );
nor ( n18109 , n18106 , n18108 );
nand ( n18110 , n18102 , n18109 );
not ( n18111 , n18110 );
nand ( n18112 , n18094 , n18111 );
nor ( n18113 , n492 , n508 );
not ( n18114 , n18113 );
nand ( n18115 , n492 , n508 );
nand ( n18116 , n18114 , n18115 );
xnor ( n18117 , n18112 , n18116 );
buf ( n18118 , n18117 );
not ( n18119 , n18118 );
not ( n18120 , n18119 );
or ( n18121 , n18042 , n18120 );
not ( n18122 , n18041 );
nand ( n18123 , n18118 , n18122 );
nand ( n18124 , n18121 , n18123 );
not ( n18125 , n18124 );
or ( n18126 , n18040 , n18125 );
not ( n18127 , n18041 );
not ( n18128 , n18049 );
nor ( n18129 , n18128 , n18113 );
not ( n18130 , n18129 );
not ( n18131 , n18092 );
or ( n18132 , n18130 , n18131 );
and ( n18133 , n18110 , n18114 );
not ( n18134 , n18115 );
nor ( n18135 , n18133 , n18134 );
nand ( n18136 , n18132 , n18135 );
nor ( n18137 , n491 , n507 );
not ( n18138 , n18137 );
nand ( n18139 , n491 , n507 );
and ( n18140 , n18138 , n18139 );
xor ( n18141 , n18136 , n18140 );
not ( n18142 , n18141 );
not ( n18143 , n18142 );
or ( n18144 , n18127 , n18143 );
buf ( n18145 , n18141 );
nand ( n18146 , n18145 , n18122 );
nand ( n18147 , n18144 , n18146 );
not ( n18148 , n18147 );
buf ( n18149 , n18031 );
not ( n18150 , n18149 );
or ( n18151 , n18148 , n18150 );
nand ( n18152 , n18126 , n18151 );
buf ( n18153 , n2026 );
not ( n18154 , n18153 );
and ( n18155 , n18138 , n18114 );
nor ( n18156 , n490 , n506 );
nor ( n18157 , n489 , n505 );
nor ( n18158 , n18156 , n18157 );
nand ( n18159 , n18155 , n18158 );
nor ( n18160 , n18128 , n18159 );
not ( n18161 , n18160 );
not ( n18162 , n18092 );
or ( n18163 , n18161 , n18162 );
not ( n18164 , n18159 );
and ( n18165 , n18110 , n18164 );
not ( n18166 , n18158 );
or ( n18167 , n18137 , n18115 );
nand ( n18168 , n18167 , n18139 );
not ( n18169 , n18168 );
or ( n18170 , n18166 , n18169 );
nand ( n18171 , n490 , n506 );
not ( n18172 , n18171 );
not ( n18173 , n18157 );
and ( n18174 , n18172 , n18173 );
and ( n18175 , n489 , n505 );
nor ( n18176 , n18174 , n18175 );
nand ( n18177 , n18170 , n18176 );
nor ( n18178 , n18165 , n18177 );
nand ( n18179 , n18163 , n18178 );
not ( n18180 , n18179 );
xor ( n18181 , n18154 , n18180 );
not ( n18182 , n18181 );
buf ( n18183 , n2014 );
xnor ( n18184 , n18183 , n18153 );
not ( n18185 , n18183 );
buf ( n18186 , n2353 );
not ( n18187 , n18186 );
not ( n18188 , n18187 );
or ( n18189 , n18185 , n18188 );
not ( n18190 , n18183 );
nand ( n18191 , n18190 , n18186 );
nand ( n18192 , n18189 , n18191 );
nor ( n18193 , n18184 , n18192 );
buf ( n18194 , n18193 );
not ( n18195 , n18194 );
or ( n18196 , n18182 , n18195 );
not ( n18197 , n18192 );
not ( n18198 , n18153 );
or ( n18199 , n18197 , n18198 );
nand ( n18200 , n18196 , n18199 );
not ( n18201 , n18200 );
xor ( n18202 , n18152 , n18201 );
not ( n18203 , n18149 );
not ( n18204 , n18124 );
or ( n18205 , n18203 , n18204 );
not ( n18206 , n18041 );
not ( n18207 , n18044 );
and ( n18208 , n18048 , n18207 );
not ( n18209 , n18208 );
nand ( n18210 , n18066 , n18058 );
nand ( n18211 , n18091 , n18210 );
not ( n18212 , n18211 );
or ( n18213 , n18209 , n18212 );
and ( n18214 , n18099 , n18207 );
not ( n18215 , n18104 );
nor ( n18216 , n18214 , n18215 );
nand ( n18217 , n18213 , n18216 );
not ( n18218 , n18107 );
nor ( n18219 , n18218 , n18043 );
xor ( n18220 , n18217 , n18219 );
not ( n18221 , n18220 );
not ( n18222 , n18221 );
or ( n18223 , n18206 , n18222 );
not ( n18224 , n18221 );
nand ( n18225 , n18224 , n18122 );
nand ( n18226 , n18223 , n18225 );
nand ( n18227 , n18226 , n18039 );
nand ( n18228 , n18205 , n18227 );
not ( n18229 , n6223 );
not ( n18230 , n18229 );
not ( n18231 , n6303 );
or ( n18232 , n18230 , n18231 );
buf ( n18233 , n2175 );
not ( n18234 , n18233 );
and ( n18235 , n18234 , n6304 );
not ( n18236 , n2301 );
and ( n18237 , n18229 , n18236 );
and ( n18238 , n18234 , n2301 );
nor ( n18239 , n18237 , n18238 );
nor ( n18240 , n18235 , n18239 );
nand ( n18241 , n18232 , n18240 );
not ( n18242 , n18241 );
not ( n18243 , n18242 );
not ( n18244 , n2301 );
not ( n18245 , n18244 );
not ( n18246 , n18047 );
not ( n18247 , n18246 );
not ( n18248 , n18092 );
or ( n18249 , n18247 , n18248 );
nand ( n18250 , n18249 , n18096 );
not ( n18251 , n18046 );
nand ( n18252 , n18251 , n18098 );
not ( n18253 , n18252 );
and ( n18254 , n18250 , n18253 );
not ( n18255 , n18250 );
and ( n18256 , n18255 , n18252 );
nor ( n18257 , n18254 , n18256 );
not ( n18258 , n18257 );
not ( n18259 , n18258 );
xor ( n18260 , n18245 , n18259 );
not ( n18261 , n18260 );
or ( n18262 , n18243 , n18261 );
not ( n18263 , n18048 );
not ( n18264 , n18211 );
or ( n18265 , n18263 , n18264 );
not ( n18266 , n18099 );
nand ( n18267 , n18265 , n18266 );
not ( n18268 , n18104 );
nor ( n18269 , n18268 , n18044 );
buf ( n18270 , n18269 );
and ( n18271 , n18267 , n18270 );
not ( n18272 , n18267 );
not ( n18273 , n18269 );
and ( n18274 , n18272 , n18273 );
nor ( n18275 , n18271 , n18274 );
not ( n18276 , n18275 );
not ( n18277 , n18276 );
xor ( n18278 , n18245 , n18277 );
and ( n18279 , n456 , n2070 );
not ( n18280 , n456 );
and ( n18281 , n18280 , n2073 );
nor ( n18282 , n18279 , n18281 );
not ( n18283 , n18282 );
not ( n18284 , n6223 );
or ( n18285 , n18283 , n18284 );
not ( n18286 , n18282 );
nand ( n18287 , n18286 , n18229 );
nand ( n18288 , n18285 , n18287 );
not ( n18289 , n18288 );
not ( n18290 , n18289 );
nand ( n18291 , n18278 , n18290 );
nand ( n18292 , n18262 , n18291 );
xor ( n18293 , n18228 , n18292 );
not ( n18294 , n18153 );
not ( n18295 , n3177 );
or ( n18296 , n18294 , n18295 );
or ( n18297 , n3177 , n18153 );
nand ( n18298 , n18296 , n18297 );
not ( n18299 , n18298 );
buf ( n18300 , n18299 );
not ( n18301 , n18300 );
buf ( n18302 , n18030 );
not ( n18303 , n18155 );
nor ( n18304 , n18303 , n18128 );
not ( n18305 , n18304 );
not ( n18306 , n18092 );
or ( n18307 , n18305 , n18306 );
and ( n18308 , n18110 , n18155 );
nor ( n18309 , n18308 , n18168 );
nand ( n18310 , n18307 , n18309 );
not ( n18311 , n18156 );
nand ( n18312 , n18311 , n18171 );
not ( n18313 , n18312 );
and ( n18314 , n18310 , n18313 );
not ( n18315 , n18310 );
and ( n18316 , n18315 , n18312 );
nor ( n18317 , n18314 , n18316 );
buf ( n18318 , n18317 );
and ( n18319 , n18302 , n18318 );
not ( n18320 , n18302 );
not ( n18321 , n18317 );
and ( n18322 , n18320 , n18321 );
nor ( n18323 , n18319 , n18322 );
not ( n18324 , n18323 );
or ( n18325 , n18301 , n18324 );
not ( n18326 , n18302 );
and ( n18327 , n18326 , n18142 );
not ( n18328 , n18326 );
and ( n18329 , n18328 , n18145 );
nor ( n18330 , n18327 , n18329 );
not ( n18331 , n18330 );
not ( n18332 , n2458 );
not ( n18333 , n18030 );
or ( n18334 , n18332 , n18333 );
or ( n18335 , n18030 , n2458 );
nand ( n18336 , n18334 , n18335 );
nand ( n18337 , n18336 , n18298 );
not ( n18338 , n18337 );
not ( n18339 , n18338 );
or ( n18340 , n18331 , n18339 );
nand ( n18341 , n18325 , n18340 );
and ( n18342 , n18293 , n18341 );
and ( n18343 , n18228 , n18292 );
or ( n18344 , n18342 , n18343 );
xor ( n18345 , n18202 , n18344 );
not ( n18346 , n2259 );
buf ( n18347 , n2387 );
not ( n18348 , n18347 );
or ( n18349 , n18346 , n18348 );
nand ( n18350 , n18348 , n18346 );
nand ( n18351 , n18349 , n18350 );
not ( n18352 , n2353 );
and ( n18353 , n2259 , n18352 );
not ( n18354 , n2259 );
and ( n18355 , n18354 , n2353 );
or ( n18356 , n18353 , n18355 );
nand ( n18357 , n18351 , n18356 );
not ( n18358 , n18357 );
buf ( n18359 , n18358 );
not ( n18360 , n18348 );
not ( n18361 , n18346 );
and ( n18362 , n18360 , n18361 );
and ( n18363 , n18348 , n18346 );
nor ( n18364 , n18362 , n18363 );
buf ( n18365 , n18364 );
or ( n18366 , n18359 , n18365 );
not ( n18367 , n18186 );
buf ( n18368 , n18367 );
buf ( n18369 , n18368 );
not ( n18370 , n18369 );
buf ( n18371 , n18370 );
not ( n18372 , n18371 );
not ( n18373 , n18372 );
nand ( n18374 , n18366 , n18373 );
not ( n18375 , n18096 );
nor ( n18376 , n18375 , n18047 );
xor ( n18377 , n18376 , n18092 );
and ( n18378 , n18245 , n18377 );
xor ( n18379 , n18374 , n18378 );
not ( n18380 , n18194 );
not ( n18381 , n18198 );
not ( n18382 , n18381 );
nor ( n18383 , n18137 , n18113 );
nand ( n18384 , n18383 , n18311 );
nor ( n18385 , n18128 , n18384 );
not ( n18386 , n18385 );
not ( n18387 , n18092 );
or ( n18388 , n18386 , n18387 );
not ( n18389 , n18384 );
and ( n18390 , n18110 , n18389 );
not ( n18391 , n18311 );
not ( n18392 , n18168 );
or ( n18393 , n18391 , n18392 );
nand ( n18394 , n18393 , n18171 );
nor ( n18395 , n18390 , n18394 );
nand ( n18396 , n18388 , n18395 );
nor ( n18397 , n18157 , n18175 );
xor ( n18398 , n18396 , n18397 );
not ( n18399 , n18398 );
not ( n18400 , n18399 );
or ( n18401 , n18382 , n18400 );
not ( n18402 , n18399 );
nand ( n18403 , n18198 , n18402 );
nand ( n18404 , n18401 , n18403 );
not ( n18405 , n18404 );
or ( n18406 , n18380 , n18405 );
not ( n18407 , n18197 );
nand ( n18408 , n18181 , n18407 );
nand ( n18409 , n18406 , n18408 );
and ( n18410 , n18379 , n18409 );
and ( n18411 , n18374 , n18378 );
or ( n18412 , n18410 , n18411 );
not ( n18413 , n18338 );
not ( n18414 , n18323 );
or ( n18415 , n18413 , n18414 );
not ( n18416 , n18302 );
not ( n18417 , n18402 );
not ( n18418 , n18417 );
or ( n18419 , n18416 , n18418 );
nand ( n18420 , n18402 , n18326 );
nand ( n18421 , n18419 , n18420 );
nand ( n18422 , n18421 , n18300 );
nand ( n18423 , n18415 , n18422 );
xor ( n18424 , n18245 , n18224 );
not ( n18425 , n18424 );
not ( n18426 , n18290 );
or ( n18427 , n18425 , n18426 );
nand ( n18428 , n18278 , n18242 );
nand ( n18429 , n18427 , n18428 );
xor ( n18430 , n18423 , n18429 );
and ( n18431 , n18245 , n18259 );
xor ( n18432 , n18430 , n18431 );
xor ( n18433 , n18412 , n18432 );
not ( n18434 , n18369 );
not ( n18435 , n18434 );
and ( n18436 , n18435 , n18180 );
not ( n18437 , n18435 );
not ( n18438 , n18180 );
and ( n18439 , n18437 , n18438 );
nor ( n18440 , n18436 , n18439 );
not ( n18441 , n18440 );
not ( n18442 , n18359 );
or ( n18443 , n18441 , n18442 );
not ( n18444 , n18365 );
not ( n18445 , n18373 );
or ( n18446 , n18444 , n18445 );
nand ( n18447 , n18443 , n18446 );
buf ( n18448 , n2301 );
not ( n18449 , n18052 );
nor ( n18450 , n18089 , n18449 );
not ( n18451 , n18450 );
nor ( n18452 , n501 , n517 );
nor ( n18453 , n502 , n518 );
nor ( n18454 , n18452 , n18453 );
not ( n18455 , n18454 );
and ( n18456 , n504 , n520 );
not ( n18457 , n18456 );
not ( n18458 , n18079 );
or ( n18459 , n18457 , n18458 );
nand ( n18460 , n503 , n519 );
nand ( n18461 , n18459 , n18460 );
not ( n18462 , n18461 );
or ( n18463 , n18455 , n18462 );
or ( n18464 , n18452 , n18070 );
nand ( n18465 , n18464 , n18069 );
not ( n18466 , n18465 );
nand ( n18467 , n18463 , n18466 );
not ( n18468 , n18467 );
or ( n18469 , n18451 , n18468 );
not ( n18470 , n18063 );
not ( n18471 , n18052 );
not ( n18472 , n18061 );
not ( n18473 , n18060 );
and ( n18474 , n18472 , n18473 );
not ( n18475 , n18064 );
nor ( n18476 , n18474 , n18475 );
nor ( n18477 , n18471 , n18476 );
nor ( n18478 , n18470 , n18477 );
nand ( n18479 , n18469 , n18478 );
and ( n18480 , n18054 , n18057 );
xor ( n18481 , n18479 , n18480 );
buf ( n18482 , n18481 );
and ( n18483 , n18448 , n18482 );
not ( n18484 , n18407 );
not ( n18485 , n18404 );
or ( n18486 , n18484 , n18485 );
not ( n18487 , n18381 );
not ( n18488 , n18321 );
or ( n18489 , n18487 , n18488 );
nand ( n18490 , n18318 , n18198 );
nand ( n18491 , n18489 , n18490 );
nand ( n18492 , n18491 , n18194 );
nand ( n18493 , n18486 , n18492 );
xor ( n18494 , n18483 , n18493 );
not ( n18495 , n18039 );
not ( n18496 , n6304 );
not ( n18497 , n18276 );
or ( n18498 , n18496 , n18497 );
nand ( n18499 , n18277 , n18122 );
nand ( n18500 , n18498 , n18499 );
not ( n18501 , n18500 );
or ( n18502 , n18495 , n18501 );
nand ( n18503 , n18226 , n18149 );
nand ( n18504 , n18502 , n18503 );
and ( n18505 , n18494 , n18504 );
and ( n18506 , n18483 , n18493 );
or ( n18507 , n18505 , n18506 );
xor ( n18508 , n18447 , n18507 );
xor ( n18509 , n18374 , n18378 );
xor ( n18510 , n18509 , n18409 );
and ( n18511 , n18508 , n18510 );
and ( n18512 , n18447 , n18507 );
or ( n18513 , n18511 , n18512 );
xor ( n18514 , n18433 , n18513 );
xor ( n18515 , n18345 , n18514 );
not ( n18516 , n18290 );
not ( n18517 , n18260 );
or ( n18518 , n18516 , n18517 );
xor ( n18519 , n18245 , n18377 );
nand ( n18520 , n18519 , n18242 );
nand ( n18521 , n18518 , n18520 );
not ( n18522 , n18338 );
and ( n18523 , n18302 , n18118 );
not ( n18524 , n18302 );
and ( n18525 , n18524 , n18119 );
nor ( n18526 , n18523 , n18525 );
not ( n18527 , n18526 );
or ( n18528 , n18522 , n18527 );
nand ( n18529 , n18330 , n18300 );
nand ( n18530 , n18528 , n18529 );
xor ( n18531 , n18521 , n18530 );
not ( n18532 , n18447 );
and ( n18533 , n18531 , n18532 );
and ( n18534 , n18521 , n18530 );
or ( n18535 , n18533 , n18534 );
xor ( n18536 , n18228 , n18292 );
xor ( n18537 , n18536 , n18341 );
xor ( n18538 , n18535 , n18537 );
xor ( n18539 , n18447 , n18507 );
xor ( n18540 , n18539 , n18510 );
and ( n18541 , n18538 , n18540 );
and ( n18542 , n18535 , n18537 );
or ( n18543 , n18541 , n18542 );
and ( n18544 , n18515 , n18543 );
and ( n18545 , n18345 , n18514 );
or ( n18546 , n18544 , n18545 );
xor ( n18547 , n18152 , n18201 );
and ( n18548 , n18547 , n18344 );
and ( n18549 , n18152 , n18201 );
or ( n18550 , n18548 , n18549 );
xor ( n18551 , n18423 , n18429 );
and ( n18552 , n18551 , n18431 );
and ( n18553 , n18423 , n18429 );
or ( n18554 , n18552 , n18553 );
not ( n18555 , n18197 );
not ( n18556 , n18195 );
or ( n18557 , n18555 , n18556 );
nand ( n18558 , n18557 , n18381 );
not ( n18559 , n18421 );
or ( n18560 , n18559 , n18339 );
not ( n18561 , n18030 );
and ( n18562 , n18561 , n18438 );
not ( n18563 , n18561 );
and ( n18564 , n18563 , n18180 );
nor ( n18565 , n18562 , n18564 );
not ( n18566 , n18300 );
or ( n18567 , n18565 , n18566 );
nand ( n18568 , n18560 , n18567 );
xor ( n18569 , n18558 , n18568 );
not ( n18570 , n18290 );
xor ( n18571 , n18245 , n18118 );
not ( n18572 , n18571 );
or ( n18573 , n18570 , n18572 );
not ( n18574 , n18424 );
or ( n18575 , n18574 , n18241 );
nand ( n18576 , n18573 , n18575 );
xor ( n18577 , n18569 , n18576 );
xor ( n18578 , n18554 , n18577 );
and ( n18579 , n18245 , n18277 );
not ( n18580 , n18149 );
not ( n18581 , n18041 );
not ( n18582 , n18321 );
or ( n18583 , n18581 , n18582 );
nand ( n18584 , n18318 , n18122 );
nand ( n18585 , n18583 , n18584 );
not ( n18586 , n18585 );
or ( n18587 , n18580 , n18586 );
nand ( n18588 , n18147 , n18039 );
nand ( n18589 , n18587 , n18588 );
xor ( n18590 , n18579 , n18589 );
xor ( n18591 , n18590 , n18200 );
xor ( n18592 , n18578 , n18591 );
xor ( n18593 , n18550 , n18592 );
xor ( n18594 , n18412 , n18432 );
and ( n18595 , n18594 , n18513 );
and ( n18596 , n18412 , n18432 );
or ( n18597 , n18595 , n18596 );
xor ( n18598 , n18593 , n18597 );
or ( n18599 , n18546 , n18598 );
not ( n18600 , n18599 );
xor ( n18601 , n18550 , n18592 );
and ( n18602 , n18601 , n18597 );
and ( n18603 , n18550 , n18592 );
or ( n18604 , n18602 , n18603 );
and ( n18605 , n18245 , n18224 );
not ( n18606 , n18039 );
not ( n18607 , n18585 );
or ( n18608 , n18606 , n18607 );
not ( n18609 , n18041 );
not ( n18610 , n18417 );
or ( n18611 , n18609 , n18610 );
nand ( n18612 , n18402 , n18122 );
nand ( n18613 , n18611 , n18612 );
nand ( n18614 , n18613 , n18149 );
nand ( n18615 , n18608 , n18614 );
xor ( n18616 , n18605 , n18615 );
not ( n18617 , n18242 );
not ( n18618 , n18571 );
or ( n18619 , n18617 , n18618 );
xor ( n18620 , n18245 , n18145 );
nand ( n18621 , n18620 , n18290 );
nand ( n18622 , n18619 , n18621 );
xor ( n18623 , n18616 , n18622 );
or ( n18624 , n18565 , n18339 );
or ( n18625 , n18566 , n18326 );
nand ( n18626 , n18624 , n18625 );
not ( n18627 , n18626 );
xor ( n18628 , n18558 , n18568 );
and ( n18629 , n18628 , n18576 );
and ( n18630 , n18558 , n18568 );
or ( n18631 , n18629 , n18630 );
xor ( n18632 , n18627 , n18631 );
xor ( n18633 , n18579 , n18589 );
and ( n18634 , n18633 , n18200 );
and ( n18635 , n18579 , n18589 );
or ( n18636 , n18634 , n18635 );
xor ( n18637 , n18632 , n18636 );
xor ( n18638 , n18623 , n18637 );
xor ( n18639 , n18554 , n18577 );
and ( n18640 , n18639 , n18591 );
and ( n18641 , n18554 , n18577 );
or ( n18642 , n18640 , n18641 );
xor ( n18643 , n18638 , n18642 );
nor ( n18644 , n18604 , n18643 );
nor ( n18645 , n18600 , n18644 );
not ( n18646 , n18645 );
not ( n18647 , n18039 );
not ( n18648 , n18041 );
not ( n18649 , n18482 );
not ( n18650 , n18649 );
or ( n18651 , n18648 , n18650 );
nand ( n18652 , n18482 , n18122 );
nand ( n18653 , n18651 , n18652 );
not ( n18654 , n18653 );
or ( n18655 , n18647 , n18654 );
not ( n18656 , n18377 );
and ( n18657 , n18656 , n18041 );
not ( n18658 , n18656 );
and ( n18659 , n18658 , n18122 );
or ( n18660 , n18657 , n18659 );
nand ( n18661 , n18660 , n18149 );
nand ( n18662 , n18655 , n18661 );
not ( n18663 , n18242 );
not ( n18664 , n18061 );
nand ( n18665 , n18664 , n18064 );
not ( n18666 , n18665 );
not ( n18667 , n18666 );
not ( n18668 , n18071 );
not ( n18669 , n18461 );
not ( n18670 , n18669 );
or ( n18671 , n18668 , n18670 );
and ( n18672 , n18071 , n18453 );
not ( n18673 , n18452 );
or ( n18674 , n500 , n516 );
nand ( n18675 , n18673 , n18674 );
nor ( n18676 , n18672 , n18675 );
nand ( n18677 , n18671 , n18676 );
nand ( n18678 , n18677 , n18060 );
not ( n18679 , n18678 );
not ( n18680 , n18679 );
or ( n18681 , n18667 , n18680 );
nand ( n18682 , n18678 , n18665 );
nand ( n18683 , n18681 , n18682 );
not ( n18684 , n18683 );
not ( n18685 , n18684 );
xor ( n18686 , n18245 , n18685 );
not ( n18687 , n18686 );
or ( n18688 , n18663 , n18687 );
not ( n18689 , n18245 );
not ( n18690 , n18089 );
not ( n18691 , n18690 );
not ( n18692 , n18467 );
or ( n18693 , n18691 , n18692 );
nand ( n18694 , n18693 , n18476 );
not ( n18695 , n18063 );
nor ( n18696 , n18695 , n18449 );
xor ( n18697 , n18694 , n18696 );
not ( n18698 , n18697 );
not ( n18699 , n18698 );
or ( n18700 , n18689 , n18699 );
not ( n18701 , n18448 );
nand ( n18702 , n18701 , n18697 );
nand ( n18703 , n18700 , n18702 );
nand ( n18704 , n18703 , n18290 );
nand ( n18705 , n18688 , n18704 );
xor ( n18706 , n18662 , n18705 );
not ( n18707 , n18117 );
and ( n18708 , n18154 , n18707 );
not ( n18709 , n18154 );
and ( n18710 , n18709 , n18118 );
nor ( n18711 , n18708 , n18710 );
nand ( n18712 , n18711 , n18407 );
not ( n18713 , n18220 );
xor ( n18714 , n18198 , n18713 );
nand ( n18715 , n18714 , n18194 );
nand ( n18716 , n18712 , n18715 );
and ( n18717 , n18706 , n18716 );
and ( n18718 , n18662 , n18705 );
or ( n18719 , n18717 , n18718 );
not ( n18720 , n18290 );
xor ( n18721 , n18448 , n18482 );
not ( n18722 , n18721 );
or ( n18723 , n18720 , n18722 );
nand ( n18724 , n18703 , n18242 );
nand ( n18725 , n18723 , n18724 );
and ( n18726 , n18245 , n18685 );
xor ( n18727 , n18725 , n18726 );
not ( n18728 , n18365 );
and ( n18729 , n18371 , n18402 );
not ( n18730 , n18371 );
and ( n18731 , n18730 , n18399 );
nor ( n18732 , n18729 , n18731 );
not ( n18733 , n18732 );
or ( n18734 , n18728 , n18733 );
not ( n18735 , n18434 );
not ( n18736 , n18321 );
or ( n18737 , n18735 , n18736 );
not ( n18738 , n18434 );
nand ( n18739 , n18318 , n18738 );
nand ( n18740 , n18737 , n18739 );
nand ( n18741 , n18740 , n18359 );
nand ( n18742 , n18734 , n18741 );
xor ( n18743 , n18727 , n18742 );
xor ( n18744 , n18719 , n18743 );
not ( n18745 , n18338 );
and ( n18746 , n18276 , n18030 );
not ( n18747 , n18276 );
and ( n18748 , n18747 , n18561 );
or ( n18749 , n18746 , n18748 );
not ( n18750 , n18749 );
or ( n18751 , n18745 , n18750 );
not ( n18752 , n18030 );
not ( n18753 , n18221 );
or ( n18754 , n18752 , n18753 );
nand ( n18755 , n18224 , n18561 );
nand ( n18756 , n18754 , n18755 );
nand ( n18757 , n18756 , n18300 );
nand ( n18758 , n18751 , n18757 );
or ( n18759 , n2638 , n456 );
not ( n18760 , n17397 );
nand ( n18761 , n18760 , n456 );
and ( n18762 , n456 , n469 );
not ( n18763 , n456 );
and ( n18764 , n18763 , n485 );
nor ( n18765 , n18762 , n18764 );
not ( n18766 , n18765 );
nand ( n18767 , n18759 , n18761 , n18766 );
not ( n18768 , n18767 );
nand ( n18769 , n18759 , n18761 );
buf ( n18770 , n18769 );
or ( n18771 , n18768 , n18770 );
buf ( n18772 , n18765 );
not ( n18773 , n18772 );
buf ( n18774 , n18773 );
nand ( n18775 , n18771 , n18774 );
not ( n18776 , n18775 );
and ( n18777 , n18674 , n18060 );
xor ( n18778 , n18777 , n18467 );
buf ( n18779 , n18778 );
not ( n18780 , n18779 );
not ( n18781 , n18780 );
nand ( n18782 , n18781 , n18245 );
nand ( n18783 , n18776 , n18782 );
xor ( n18784 , n18758 , n18783 );
not ( n18785 , n18149 );
not ( n18786 , n18041 );
not ( n18787 , n18258 );
or ( n18788 , n18786 , n18787 );
nand ( n18789 , n18259 , n18122 );
nand ( n18790 , n18788 , n18789 );
not ( n18791 , n18790 );
or ( n18792 , n18785 , n18791 );
nand ( n18793 , n18660 , n18039 );
nand ( n18794 , n18792 , n18793 );
xor ( n18795 , n18784 , n18794 );
xor ( n18796 , n18744 , n18795 );
not ( n18797 , n18775 );
not ( n18798 , n18782 );
not ( n18799 , n18798 );
or ( n18800 , n18797 , n18799 );
nand ( n18801 , n18800 , n18783 );
nand ( n18802 , n18082 , n18070 );
not ( n18803 , n18069 );
nor ( n18804 , n18803 , n18452 );
and ( n18805 , n18802 , n18804 );
not ( n18806 , n18802 );
nand ( n18807 , n18085 , n18069 );
and ( n18808 , n18806 , n18807 );
nor ( n18809 , n18805 , n18808 );
buf ( n18810 , n18809 );
and ( n18811 , n18810 , n18245 );
not ( n18812 , n18768 );
not ( n18813 , n18774 );
not ( n18814 , n18813 );
not ( n18815 , n18438 );
or ( n18816 , n18814 , n18815 );
nand ( n18817 , n18180 , n18774 );
nand ( n18818 , n18816 , n18817 );
not ( n18819 , n18818 );
or ( n18820 , n18812 , n18819 );
nand ( n18821 , n18774 , n18770 );
nand ( n18822 , n18820 , n18821 );
and ( n18823 , n18811 , n18822 );
xor ( n18824 , n18801 , n18823 );
and ( n18825 , n18780 , n18245 );
not ( n18826 , n18780 );
and ( n18827 , n18826 , n18244 );
or ( n18828 , n18825 , n18827 );
and ( n18829 , n18828 , n18288 );
not ( n18830 , n18810 );
not ( n18831 , n18244 );
and ( n18832 , n18830 , n18831 );
and ( n18833 , n18810 , n18244 );
nor ( n18834 , n18832 , n18833 );
nor ( n18835 , n18834 , n18241 );
nor ( n18836 , n18829 , n18835 );
not ( n18837 , n18453 );
nand ( n18838 , n18837 , n18070 );
and ( n18839 , n18838 , n18669 );
not ( n18840 , n18838 );
not ( n18841 , n18669 );
and ( n18842 , n18840 , n18841 );
nor ( n18843 , n18839 , n18842 );
buf ( n18844 , n18843 );
not ( n18845 , n18844 );
or ( n18846 , n18845 , n18244 );
nor ( n18847 , n18836 , n18846 );
not ( n18848 , n18149 );
not ( n18849 , n18653 );
or ( n18850 , n18848 , n18849 );
not ( n18851 , n18041 );
not ( n18852 , n18698 );
or ( n18853 , n18851 , n18852 );
nand ( n18854 , n18697 , n18122 );
nand ( n18855 , n18853 , n18854 );
nand ( n18856 , n18855 , n18039 );
nand ( n18857 , n18850 , n18856 );
xor ( n18858 , n18847 , n18857 );
not ( n18859 , n18290 );
not ( n18860 , n18686 );
or ( n18861 , n18859 , n18860 );
nand ( n18862 , n18828 , n18242 );
nand ( n18863 , n18861 , n18862 );
and ( n18864 , n18858 , n18863 );
and ( n18865 , n18847 , n18857 );
or ( n18866 , n18864 , n18865 );
and ( n18867 , n18824 , n18866 );
and ( n18868 , n18801 , n18823 );
or ( n18869 , n18867 , n18868 );
not ( n18870 , n18407 );
not ( n18871 , n18381 );
not ( n18872 , n18142 );
or ( n18873 , n18871 , n18872 );
nand ( n18874 , n18145 , n18154 );
nand ( n18875 , n18873 , n18874 );
not ( n18876 , n18875 );
or ( n18877 , n18870 , n18876 );
nand ( n18878 , n18711 , n18194 );
nand ( n18879 , n18877 , n18878 );
not ( n18880 , n18347 );
not ( n18881 , n18880 );
and ( n18882 , n18881 , n18179 );
not ( n18883 , n18881 );
and ( n18884 , n18883 , n18180 );
nor ( n18885 , n18882 , n18884 );
not ( n18886 , n2851 );
and ( n18887 , n18347 , n18886 );
not ( n18888 , n18347 );
not ( n18889 , n18886 );
and ( n18890 , n18888 , n18889 );
nor ( n18891 , n18887 , n18890 );
not ( n18892 , n18886 );
not ( n18893 , n3316 );
or ( n18894 , n18892 , n18893 );
or ( n18895 , n3316 , n18886 );
nand ( n18896 , n18894 , n18895 );
nand ( n18897 , n18891 , n18896 );
not ( n18898 , n18897 );
and ( n18899 , n18885 , n18898 );
not ( n18900 , n18896 );
and ( n18901 , n18900 , n18881 );
nor ( n18902 , n18899 , n18901 );
xor ( n18903 , n18879 , n18902 );
not ( n18904 , n18898 );
not ( n18905 , n18348 );
xor ( n18906 , n18905 , n18398 );
not ( n18907 , n18906 );
or ( n18908 , n18904 , n18907 );
nand ( n18909 , n18885 , n18900 );
nand ( n18910 , n18908 , n18909 );
not ( n18911 , n18300 );
not ( n18912 , n18749 );
or ( n18913 , n18911 , n18912 );
not ( n18914 , n18030 );
not ( n18915 , n18258 );
or ( n18916 , n18914 , n18915 );
nand ( n18917 , n18257 , n18561 );
nand ( n18918 , n18916 , n18917 );
nand ( n18919 , n18918 , n18338 );
nand ( n18920 , n18913 , n18919 );
xor ( n18921 , n18910 , n18920 );
not ( n18922 , n18365 );
not ( n18923 , n18740 );
or ( n18924 , n18922 , n18923 );
not ( n18925 , n18368 );
buf ( n18926 , n18925 );
not ( n18927 , n18926 );
not ( n18928 , n18927 );
not ( n18929 , n18928 );
not ( n18930 , n18142 );
or ( n18931 , n18929 , n18930 );
nand ( n18932 , n18145 , n18372 );
nand ( n18933 , n18931 , n18932 );
nand ( n18934 , n18933 , n18359 );
nand ( n18935 , n18924 , n18934 );
and ( n18936 , n18921 , n18935 );
and ( n18937 , n18910 , n18920 );
or ( n18938 , n18936 , n18937 );
xor ( n18939 , n18903 , n18938 );
xor ( n18940 , n18869 , n18939 );
not ( n18941 , n18194 );
not ( n18942 , n18381 );
and ( n18943 , n18267 , n18270 );
not ( n18944 , n18267 );
and ( n18945 , n18944 , n18273 );
nor ( n18946 , n18943 , n18945 );
not ( n18947 , n18946 );
not ( n18948 , n18947 );
or ( n18949 , n18942 , n18948 );
not ( n18950 , n18946 );
or ( n18951 , n18950 , n18153 );
nand ( n18952 , n18949 , n18951 );
not ( n18953 , n18952 );
or ( n18954 , n18941 , n18953 );
nand ( n18955 , n18714 , n18407 );
nand ( n18956 , n18954 , n18955 );
not ( n18957 , n18900 );
not ( n18958 , n18906 );
or ( n18959 , n18957 , n18958 );
not ( n18960 , n18880 );
not ( n18961 , n18317 );
or ( n18962 , n18960 , n18961 );
not ( n18963 , n18881 );
or ( n18964 , n18317 , n18963 );
nand ( n18965 , n18962 , n18964 );
nand ( n18966 , n18965 , n18898 );
nand ( n18967 , n18959 , n18966 );
xor ( n18968 , n18956 , n18967 );
not ( n18969 , n18338 );
not ( n18970 , n18030 );
not ( n18971 , n18656 );
or ( n18972 , n18970 , n18971 );
nand ( n18973 , n18377 , n18561 );
nand ( n18974 , n18972 , n18973 );
not ( n18975 , n18974 );
or ( n18976 , n18969 , n18975 );
nand ( n18977 , n18918 , n18300 );
nand ( n18978 , n18976 , n18977 );
and ( n18979 , n18968 , n18978 );
and ( n18980 , n18956 , n18967 );
or ( n18981 , n18979 , n18980 );
xor ( n18982 , n18662 , n18705 );
xor ( n18983 , n18982 , n18716 );
xor ( n18984 , n18981 , n18983 );
xor ( n18985 , n18910 , n18920 );
xor ( n18986 , n18985 , n18935 );
and ( n18987 , n18984 , n18986 );
and ( n18988 , n18981 , n18983 );
or ( n18989 , n18987 , n18988 );
xor ( n18990 , n18940 , n18989 );
xor ( n18991 , n18796 , n18990 );
not ( n18992 , n18359 );
not ( n18993 , n18373 );
not ( n18994 , n18119 );
or ( n18995 , n18993 , n18994 );
nand ( n18996 , n18118 , n18372 );
nand ( n18997 , n18995 , n18996 );
not ( n18998 , n18997 );
or ( n18999 , n18992 , n18998 );
nand ( n19000 , n18933 , n18365 );
nand ( n19001 , n18999 , n19000 );
xor ( n19002 , n18811 , n18822 );
xor ( n19003 , n19001 , n19002 );
xor ( n19004 , n18836 , n18846 );
not ( n19005 , n18338 );
not ( n19006 , n18030 );
not ( n19007 , n18649 );
or ( n19008 , n19006 , n19007 );
nand ( n19009 , n18482 , n18561 );
nand ( n19010 , n19008 , n19009 );
not ( n19011 , n19010 );
or ( n19012 , n19005 , n19011 );
nand ( n19013 , n18974 , n18300 );
nand ( n19014 , n19012 , n19013 );
and ( n19015 , n19004 , n19014 );
and ( n19016 , n19003 , n19015 );
and ( n19017 , n19001 , n19002 );
or ( n19018 , n19016 , n19017 );
xor ( n19019 , n18801 , n18823 );
xor ( n19020 , n19019 , n18866 );
xor ( n19021 , n19018 , n19020 );
not ( n19022 , n18039 );
and ( n19023 , n18685 , n18122 );
not ( n19024 , n18685 );
and ( n19025 , n19024 , n18041 );
or ( n19026 , n19023 , n19025 );
not ( n19027 , n19026 );
or ( n19028 , n19022 , n19027 );
nand ( n19029 , n18855 , n18149 );
nand ( n19030 , n19028 , n19029 );
and ( n19031 , n18257 , n18381 );
not ( n19032 , n18257 );
and ( n19033 , n19032 , n18154 );
nor ( n19034 , n19031 , n19033 );
not ( n19035 , n19034 );
or ( n19036 , n19035 , n18195 );
not ( n19037 , n18952 );
or ( n19038 , n19037 , n18197 );
nand ( n19039 , n19036 , n19038 );
xor ( n19040 , n19030 , n19039 );
not ( n19041 , n18818 );
not ( n19042 , n18770 );
or ( n19043 , n19041 , n19042 );
and ( n19044 , n18398 , n18774 );
not ( n19045 , n18398 );
and ( n19046 , n19045 , n18813 );
or ( n19047 , n19044 , n19046 );
or ( n19048 , n19047 , n18767 );
nand ( n19049 , n19043 , n19048 );
and ( n19050 , n19040 , n19049 );
and ( n19051 , n19030 , n19039 );
or ( n19052 , n19050 , n19051 );
xor ( n19053 , n18847 , n18857 );
xor ( n19054 , n19053 , n18863 );
xor ( n19055 , n19052 , n19054 );
xor ( n19056 , n18956 , n18967 );
xor ( n19057 , n19056 , n18978 );
and ( n19058 , n19055 , n19057 );
and ( n19059 , n19052 , n19054 );
or ( n19060 , n19058 , n19059 );
and ( n19061 , n19021 , n19060 );
and ( n19062 , n19018 , n19020 );
or ( n19063 , n19061 , n19062 );
xor ( n19064 , n18991 , n19063 );
xor ( n19065 , n18981 , n18983 );
xor ( n19066 , n19065 , n18986 );
xor ( n19067 , n19001 , n19002 );
xor ( n19068 , n19067 , n19015 );
not ( n19069 , n18898 );
not ( n19070 , n18881 );
not ( n19071 , n18142 );
or ( n19072 , n19070 , n19071 );
not ( n19073 , n18905 );
nand ( n19074 , n18141 , n19073 );
nand ( n19075 , n19072 , n19074 );
not ( n19076 , n19075 );
or ( n19077 , n19069 , n19076 );
nand ( n19078 , n18965 , n18900 );
nand ( n19079 , n19077 , n19078 );
not ( n19080 , n18359 );
not ( n19081 , n18927 );
and ( n19082 , n19081 , n18224 );
not ( n19083 , n19081 );
and ( n19084 , n19083 , n18221 );
nor ( n19085 , n19082 , n19084 );
not ( n19086 , n19085 );
or ( n19087 , n19080 , n19086 );
nand ( n19088 , n18997 , n18365 );
nand ( n19089 , n19087 , n19088 );
xor ( n19090 , n19079 , n19089 );
not ( n19091 , n18288 );
not ( n19092 , n18834 );
not ( n19093 , n19092 );
or ( n19094 , n19091 , n19093 );
not ( n19095 , n18448 );
not ( n19096 , n18844 );
not ( n19097 , n19096 );
or ( n19098 , n19095 , n19097 );
nand ( n19099 , n18844 , n18244 );
nand ( n19100 , n19098 , n19099 );
nand ( n19101 , n19100 , n18242 );
nand ( n19102 , n19094 , n19101 );
nand ( n19103 , n504 , n520 );
not ( n19104 , n19103 );
nand ( n19105 , n18079 , n18460 );
not ( n19106 , n19105 );
not ( n19107 , n19106 );
or ( n19108 , n19104 , n19107 );
not ( n19109 , n19103 );
nand ( n19110 , n19109 , n19105 );
nand ( n19111 , n19108 , n19110 );
buf ( n19112 , n19111 );
and ( n19113 , n18448 , n19112 );
xor ( n19114 , n19102 , n19113 );
not ( n19115 , n18149 );
not ( n19116 , n19026 );
or ( n19117 , n19115 , n19116 );
not ( n19118 , n18041 );
not ( n19119 , n18780 );
or ( n19120 , n19118 , n19119 );
nand ( n19121 , n18779 , n18122 );
nand ( n19122 , n19120 , n19121 );
nand ( n19123 , n19122 , n18039 );
nand ( n19124 , n19117 , n19123 );
and ( n19125 , n19114 , n19124 );
and ( n19126 , n19102 , n19113 );
or ( n19127 , n19125 , n19126 );
and ( n19128 , n19090 , n19127 );
and ( n19129 , n19079 , n19089 );
or ( n19130 , n19128 , n19129 );
xor ( n19131 , n19068 , n19130 );
xor ( n19132 , n19004 , n19014 );
not ( n19133 , n18300 );
not ( n19134 , n19010 );
or ( n19135 , n19133 , n19134 );
not ( n19136 , n18030 );
not ( n19137 , n18698 );
or ( n19138 , n19136 , n19137 );
nand ( n19139 , n18697 , n18561 );
nand ( n19140 , n19138 , n19139 );
nand ( n19141 , n19140 , n18338 );
nand ( n19142 , n19135 , n19141 );
not ( n19143 , n18407 );
not ( n19144 , n19034 );
or ( n19145 , n19143 , n19144 );
and ( n19146 , n18656 , n18381 );
not ( n19147 , n18656 );
and ( n19148 , n19147 , n18198 );
or ( n19149 , n19146 , n19148 );
nand ( n19150 , n19149 , n18194 );
nand ( n19151 , n19145 , n19150 );
xor ( n19152 , n19142 , n19151 );
not ( n19153 , n18317 );
not ( n19154 , n18813 );
and ( n19155 , n19153 , n19154 );
and ( n19156 , n18318 , n18813 );
nor ( n19157 , n19155 , n19156 );
or ( n19158 , n19157 , n18767 );
not ( n19159 , n18770 );
or ( n19160 , n19047 , n19159 );
nand ( n19161 , n19158 , n19160 );
and ( n19162 , n19152 , n19161 );
and ( n19163 , n19142 , n19151 );
or ( n19164 , n19162 , n19163 );
xor ( n19165 , n19132 , n19164 );
not ( n19166 , n18900 );
not ( n19167 , n19075 );
or ( n19168 , n19166 , n19167 );
not ( n19169 , n18880 );
not ( n19170 , n18117 );
or ( n19171 , n19169 , n19170 );
or ( n19172 , n18117 , n18963 );
nand ( n19173 , n19171 , n19172 );
nand ( n19174 , n19173 , n18898 );
nand ( n19175 , n19168 , n19174 );
xor ( n19176 , n504 , n520 );
not ( n19177 , n19176 );
not ( n19178 , n19177 );
and ( n19179 , n19178 , n18448 );
not ( n19180 , n18242 );
xor ( n19181 , n18448 , n19112 );
not ( n19182 , n19181 );
or ( n19183 , n19180 , n19182 );
nand ( n19184 , n19100 , n18288 );
nand ( n19185 , n19183 , n19184 );
xor ( n19186 , n19179 , n19185 );
not ( n19187 , n18241 );
and ( n19188 , n18448 , n19177 );
not ( n19189 , n18448 );
buf ( n19190 , n19176 );
and ( n19191 , n19189 , n19190 );
nor ( n19192 , n19188 , n19191 );
not ( n19193 , n19192 );
and ( n19194 , n19187 , n19193 );
and ( n19195 , n18288 , n19181 );
nor ( n19196 , n19194 , n19195 );
and ( n19197 , n6304 , n18229 );
nor ( n19198 , n19197 , n18236 );
not ( n19199 , n18234 );
not ( n19200 , n6303 );
or ( n19201 , n19199 , n19200 );
nand ( n19202 , n19201 , n19178 );
nand ( n19203 , n19198 , n19202 );
nor ( n19204 , n19196 , n19203 );
and ( n19205 , n19186 , n19204 );
and ( n19206 , n19179 , n19185 );
or ( n19207 , n19205 , n19206 );
xor ( n19208 , n19175 , n19207 );
not ( n19209 , n18359 );
not ( n19210 , n18371 );
not ( n19211 , n18276 );
or ( n19212 , n19210 , n19211 );
nand ( n19213 , n18277 , n18927 );
nand ( n19214 , n19212 , n19213 );
not ( n19215 , n19214 );
or ( n19216 , n19209 , n19215 );
nand ( n19217 , n19085 , n18365 );
nand ( n19218 , n19216 , n19217 );
and ( n19219 , n19208 , n19218 );
and ( n19220 , n19175 , n19207 );
or ( n19221 , n19219 , n19220 );
and ( n19222 , n19165 , n19221 );
and ( n19223 , n19132 , n19164 );
or ( n19224 , n19222 , n19223 );
and ( n19225 , n19131 , n19224 );
and ( n19226 , n19068 , n19130 );
or ( n19227 , n19225 , n19226 );
xor ( n19228 , n19066 , n19227 );
xor ( n19229 , n19018 , n19020 );
xor ( n19230 , n19229 , n19060 );
and ( n19231 , n19228 , n19230 );
and ( n19232 , n19066 , n19227 );
or ( n19233 , n19231 , n19232 );
nor ( n19234 , n19064 , n19233 );
xor ( n19235 , n19052 , n19054 );
xor ( n19236 , n19235 , n19057 );
xor ( n19237 , n19068 , n19130 );
xor ( n19238 , n19237 , n19224 );
xor ( n19239 , n19236 , n19238 );
xor ( n19240 , n19030 , n19039 );
xor ( n19241 , n19240 , n19049 );
xor ( n19242 , n19079 , n19089 );
xor ( n19243 , n19242 , n19127 );
xor ( n19244 , n19241 , n19243 );
not ( n19245 , n18031 );
not ( n19246 , n19122 );
or ( n19247 , n19245 , n19246 );
and ( n19248 , n18810 , n18122 );
not ( n19249 , n18810 );
and ( n19250 , n19249 , n18041 );
or ( n19251 , n19248 , n19250 );
nand ( n19252 , n19251 , n18039 );
nand ( n19253 , n19247 , n19252 );
not ( n19254 , n18338 );
not ( n19255 , n18684 );
and ( n19256 , n18030 , n19255 );
not ( n19257 , n18030 );
and ( n19258 , n19257 , n18684 );
nor ( n19259 , n19256 , n19258 );
not ( n19260 , n19259 );
or ( n19261 , n19254 , n19260 );
nand ( n19262 , n19140 , n18300 );
nand ( n19263 , n19261 , n19262 );
xor ( n19264 , n19253 , n19263 );
not ( n19265 , n18194 );
not ( n19266 , n18381 );
not ( n19267 , n18649 );
or ( n19268 , n19266 , n19267 );
nand ( n19269 , n18482 , n18198 );
nand ( n19270 , n19268 , n19269 );
not ( n19271 , n19270 );
or ( n19272 , n19265 , n19271 );
nand ( n19273 , n19149 , n18407 );
nand ( n19274 , n19272 , n19273 );
and ( n19275 , n19264 , n19274 );
and ( n19276 , n19253 , n19263 );
or ( n19277 , n19275 , n19276 );
xor ( n19278 , n19102 , n19113 );
xor ( n19279 , n19278 , n19124 );
xor ( n19280 , n19277 , n19279 );
xor ( n19281 , n19179 , n19185 );
xor ( n19282 , n19281 , n19204 );
not ( n19283 , n18898 );
and ( n19284 , n18880 , n18221 );
not ( n19285 , n18880 );
and ( n19286 , n19285 , n18224 );
nor ( n19287 , n19284 , n19286 );
not ( n19288 , n19287 );
or ( n19289 , n19283 , n19288 );
nand ( n19290 , n19173 , n18900 );
nand ( n19291 , n19289 , n19290 );
xor ( n19292 , n19282 , n19291 );
not ( n19293 , n18813 );
not ( n19294 , n18141 );
or ( n19295 , n19293 , n19294 );
or ( n19296 , n18145 , n18813 );
nand ( n19297 , n19295 , n19296 );
not ( n19298 , n19297 );
not ( n19299 , n18768 );
or ( n19300 , n19298 , n19299 );
or ( n19301 , n19157 , n19159 );
nand ( n19302 , n19300 , n19301 );
and ( n19303 , n19292 , n19302 );
and ( n19304 , n19282 , n19291 );
or ( n19305 , n19303 , n19304 );
and ( n19306 , n19280 , n19305 );
and ( n19307 , n19277 , n19279 );
or ( n19308 , n19306 , n19307 );
and ( n19309 , n19244 , n19308 );
and ( n19310 , n19241 , n19243 );
or ( n19311 , n19309 , n19310 );
and ( n19312 , n19239 , n19311 );
and ( n19313 , n19236 , n19238 );
or ( n19314 , n19312 , n19313 );
xor ( n19315 , n19066 , n19227 );
xor ( n19316 , n19315 , n19230 );
nor ( n19317 , n19314 , n19316 );
nor ( n19318 , n19234 , n19317 );
xor ( n19319 , n18719 , n18743 );
and ( n19320 , n19319 , n18795 );
and ( n19321 , n18719 , n18743 );
or ( n19322 , n19320 , n19321 );
not ( n19323 , n18407 );
not ( n19324 , n18491 );
or ( n19325 , n19323 , n19324 );
nand ( n19326 , n18875 , n18194 );
nand ( n19327 , n19325 , n19326 );
not ( n19328 , n18902 );
xor ( n19329 , n19327 , n19328 );
xor ( n19330 , n18725 , n18726 );
and ( n19331 , n19330 , n18742 );
and ( n19332 , n18725 , n18726 );
or ( n19333 , n19331 , n19332 );
xor ( n19334 , n19329 , n19333 );
xor ( n19335 , n18879 , n18902 );
and ( n19336 , n19335 , n18938 );
and ( n19337 , n18879 , n18902 );
or ( n19338 , n19336 , n19337 );
xor ( n19339 , n19334 , n19338 );
xor ( n19340 , n18758 , n18783 );
and ( n19341 , n19340 , n18794 );
and ( n19342 , n18758 , n18783 );
or ( n19343 , n19341 , n19342 );
not ( n19344 , n18896 );
not ( n19345 , n18897 );
or ( n19346 , n19344 , n19345 );
nand ( n19347 , n19346 , n18881 );
not ( n19348 , n18242 );
not ( n19349 , n18721 );
or ( n19350 , n19348 , n19349 );
nand ( n19351 , n18519 , n18290 );
nand ( n19352 , n19350 , n19351 );
xor ( n19353 , n19347 , n19352 );
not ( n19354 , n18245 );
nor ( n19355 , n19354 , n18698 );
xor ( n19356 , n19353 , n19355 );
xor ( n19357 , n19343 , n19356 );
not ( n19358 , n18359 );
not ( n19359 , n18732 );
or ( n19360 , n19358 , n19359 );
nand ( n19361 , n18440 , n18365 );
nand ( n19362 , n19360 , n19361 );
not ( n19363 , n18300 );
not ( n19364 , n18526 );
or ( n19365 , n19363 , n19364 );
nand ( n19366 , n18756 , n18338 );
nand ( n19367 , n19365 , n19366 );
xor ( n19368 , n19362 , n19367 );
not ( n19369 , n18149 );
not ( n19370 , n18500 );
or ( n19371 , n19369 , n19370 );
nand ( n19372 , n18790 , n18039 );
nand ( n19373 , n19371 , n19372 );
xor ( n19374 , n19368 , n19373 );
xor ( n19375 , n19357 , n19374 );
xor ( n19376 , n19339 , n19375 );
xor ( n19377 , n19322 , n19376 );
xor ( n19378 , n18869 , n18939 );
and ( n19379 , n19378 , n18989 );
and ( n19380 , n18869 , n18939 );
or ( n19381 , n19379 , n19380 );
and ( n19382 , n19377 , n19381 );
and ( n19383 , n19322 , n19376 );
or ( n19384 , n19382 , n19383 );
not ( n19385 , n19384 );
xor ( n19386 , n19347 , n19352 );
and ( n19387 , n19386 , n19355 );
and ( n19388 , n19347 , n19352 );
or ( n19389 , n19387 , n19388 );
xor ( n19390 , n19362 , n19367 );
and ( n19391 , n19390 , n19373 );
and ( n19392 , n19362 , n19367 );
or ( n19393 , n19391 , n19392 );
xor ( n19394 , n19389 , n19393 );
xor ( n19395 , n18521 , n18530 );
xor ( n19396 , n19395 , n18532 );
xor ( n19397 , n19394 , n19396 );
xor ( n19398 , n18483 , n18493 );
xor ( n19399 , n19398 , n18504 );
xor ( n19400 , n19327 , n19328 );
and ( n19401 , n19400 , n19333 );
and ( n19402 , n19327 , n19328 );
or ( n19403 , n19401 , n19402 );
xor ( n19404 , n19399 , n19403 );
xor ( n19405 , n19343 , n19356 );
and ( n19406 , n19405 , n19374 );
and ( n19407 , n19343 , n19356 );
or ( n19408 , n19406 , n19407 );
xor ( n19409 , n19404 , n19408 );
xor ( n19410 , n19397 , n19409 );
xor ( n19411 , n19334 , n19338 );
and ( n19412 , n19411 , n19375 );
and ( n19413 , n19334 , n19338 );
or ( n19414 , n19412 , n19413 );
xor ( n19415 , n19410 , n19414 );
not ( n19416 , n19415 );
nand ( n19417 , n19385 , n19416 );
xor ( n19418 , n19322 , n19376 );
xor ( n19419 , n19418 , n19381 );
not ( n19420 , n19419 );
xor ( n19421 , n18796 , n18990 );
and ( n19422 , n19421 , n19063 );
and ( n19423 , n18796 , n18990 );
or ( n19424 , n19422 , n19423 );
not ( n19425 , n19424 );
nand ( n19426 , n19420 , n19425 );
and ( n19427 , n19318 , n19417 , n19426 );
not ( n19428 , n19427 );
xor ( n19429 , n19132 , n19164 );
xor ( n19430 , n19429 , n19221 );
xor ( n19431 , n19241 , n19243 );
xor ( n19432 , n19431 , n19308 );
xor ( n19433 , n19430 , n19432 );
xor ( n19434 , n19175 , n19207 );
xor ( n19435 , n19434 , n19218 );
xor ( n19436 , n19142 , n19151 );
xor ( n19437 , n19436 , n19161 );
xor ( n19438 , n19435 , n19437 );
xor ( n19439 , n19277 , n19279 );
xor ( n19440 , n19439 , n19305 );
and ( n19441 , n19438 , n19440 );
and ( n19442 , n19435 , n19437 );
or ( n19443 , n19441 , n19442 );
xor ( n19444 , n19433 , n19443 );
not ( n19445 , n19444 );
not ( n19446 , n18365 );
not ( n19447 , n19214 );
or ( n19448 , n19446 , n19447 );
not ( n19449 , n18928 );
not ( n19450 , n18258 );
or ( n19451 , n19449 , n19450 );
nand ( n19452 , n18259 , n18738 );
nand ( n19453 , n19451 , n19452 );
nand ( n19454 , n19453 , n18359 );
nand ( n19455 , n19448 , n19454 );
not ( n19456 , n18149 );
not ( n19457 , n19251 );
or ( n19458 , n19456 , n19457 );
not ( n19459 , n6304 );
not ( n19460 , n18845 );
or ( n19461 , n19459 , n19460 );
nand ( n19462 , n18844 , n18122 );
nand ( n19463 , n19461 , n19462 );
nand ( n19464 , n19463 , n18039 );
nand ( n19465 , n19458 , n19464 );
xor ( n19466 , n19196 , n19203 );
xor ( n19467 , n19465 , n19466 );
not ( n19468 , n18300 );
not ( n19469 , n19259 );
or ( n19470 , n19468 , n19469 );
not ( n19471 , n18030 );
not ( n19472 , n18780 );
or ( n19473 , n19471 , n19472 );
nand ( n19474 , n18779 , n18561 );
nand ( n19475 , n19473 , n19474 );
nand ( n19476 , n19475 , n18338 );
nand ( n19477 , n19470 , n19476 );
and ( n19478 , n19467 , n19477 );
and ( n19479 , n19465 , n19466 );
or ( n19480 , n19478 , n19479 );
xor ( n19481 , n19455 , n19480 );
xor ( n19482 , n19253 , n19263 );
xor ( n19483 , n19482 , n19274 );
and ( n19484 , n19481 , n19483 );
and ( n19485 , n19455 , n19480 );
or ( n19486 , n19484 , n19485 );
not ( n19487 , n18407 );
not ( n19488 , n19270 );
or ( n19489 , n19487 , n19488 );
not ( n19490 , n18381 );
not ( n19491 , n18698 );
or ( n19492 , n19490 , n19491 );
nand ( n19493 , n18697 , n18198 );
nand ( n19494 , n19492 , n19493 );
nand ( n19495 , n19494 , n18194 );
nand ( n19496 , n19489 , n19495 );
not ( n19497 , n18900 );
not ( n19498 , n19287 );
or ( n19499 , n19497 , n19498 );
not ( n19500 , n18276 );
not ( n19501 , n18881 );
or ( n19502 , n19500 , n19501 );
nand ( n19503 , n18946 , n18880 );
nand ( n19504 , n19502 , n19503 );
nand ( n19505 , n19504 , n18898 );
nand ( n19506 , n19499 , n19505 );
xor ( n19507 , n19496 , n19506 );
and ( n19508 , n18288 , n19178 );
not ( n19509 , n18031 );
not ( n19510 , n19463 );
or ( n19511 , n19509 , n19510 );
not ( n19512 , n6304 );
not ( n19513 , n19112 );
not ( n19514 , n19513 );
or ( n19515 , n19512 , n19514 );
nand ( n19516 , n19112 , n6303 );
nand ( n19517 , n19515 , n19516 );
nand ( n19518 , n19517 , n18037 );
nand ( n19519 , n19511 , n19518 );
xor ( n19520 , n19508 , n19519 );
nand ( n19521 , n18561 , n6206 );
and ( n19522 , n19521 , n19178 );
not ( n19523 , n2270 );
not ( n19524 , n18030 );
or ( n19525 , n19523 , n19524 );
nand ( n19526 , n19525 , n6304 );
nor ( n19527 , n19522 , n19526 );
not ( n19528 , n18031 );
not ( n19529 , n19517 );
or ( n19530 , n19528 , n19529 );
not ( n19531 , n6304 );
not ( n19532 , n19177 );
or ( n19533 , n19531 , n19532 );
nand ( n19534 , n6303 , n19178 );
nand ( n19535 , n19533 , n19534 );
nand ( n19536 , n18037 , n19535 );
nand ( n19537 , n19530 , n19536 );
and ( n19538 , n19527 , n19537 );
and ( n19539 , n19520 , n19538 );
and ( n19540 , n19508 , n19519 );
or ( n19541 , n19539 , n19540 );
and ( n19542 , n19507 , n19541 );
and ( n19543 , n19496 , n19506 );
or ( n19544 , n19542 , n19543 );
xor ( n19545 , n19282 , n19291 );
xor ( n19546 , n19545 , n19302 );
xor ( n19547 , n19544 , n19546 );
not ( n19548 , n18768 );
not ( n19549 , n18772 );
and ( n19550 , n19549 , n18118 );
not ( n19551 , n19549 );
and ( n19552 , n19551 , n18707 );
nor ( n19553 , n19550 , n19552 );
not ( n19554 , n19553 );
or ( n19555 , n19548 , n19554 );
nand ( n19556 , n19297 , n18770 );
nand ( n19557 , n19555 , n19556 );
not ( n19558 , n18365 );
not ( n19559 , n19453 );
or ( n19560 , n19558 , n19559 );
and ( n19561 , n18926 , n18377 );
not ( n19562 , n18926 );
and ( n19563 , n19562 , n18656 );
nor ( n19564 , n19561 , n19563 );
nand ( n19565 , n19564 , n18359 );
nand ( n19566 , n19560 , n19565 );
xor ( n19567 , n19557 , n19566 );
xor ( n19568 , n19465 , n19466 );
xor ( n19569 , n19568 , n19477 );
and ( n19570 , n19567 , n19569 );
and ( n19571 , n19557 , n19566 );
or ( n19572 , n19570 , n19571 );
and ( n19573 , n19547 , n19572 );
and ( n19574 , n19544 , n19546 );
or ( n19575 , n19573 , n19574 );
xor ( n19576 , n19486 , n19575 );
xor ( n19577 , n19435 , n19437 );
xor ( n19578 , n19577 , n19440 );
and ( n19579 , n19576 , n19578 );
and ( n19580 , n19486 , n19575 );
or ( n19581 , n19579 , n19580 );
not ( n19582 , n19581 );
and ( n19583 , n19445 , n19582 );
xor ( n19584 , n19236 , n19238 );
xor ( n19585 , n19584 , n19311 );
xor ( n19586 , n19430 , n19432 );
and ( n19587 , n19586 , n19443 );
and ( n19588 , n19430 , n19432 );
or ( n19589 , n19587 , n19588 );
nor ( n19590 , n19585 , n19589 );
nor ( n19591 , n19583 , n19590 );
not ( n19592 , n19591 );
xor ( n19593 , n19486 , n19575 );
xor ( n19594 , n19593 , n19578 );
not ( n19595 , n19594 );
xor ( n19596 , n19455 , n19480 );
xor ( n19597 , n19596 , n19483 );
not ( n19598 , n18300 );
not ( n19599 , n19475 );
or ( n19600 , n19598 , n19599 );
not ( n19601 , n18030 );
not ( n19602 , n18810 );
not ( n19603 , n19602 );
or ( n19604 , n19601 , n19603 );
nand ( n19605 , n18810 , n18561 );
nand ( n19606 , n19604 , n19605 );
nand ( n19607 , n19606 , n18338 );
nand ( n19608 , n19600 , n19607 );
not ( n19609 , n18359 );
and ( n19610 , n18482 , n18434 );
not ( n19611 , n18482 );
and ( n19612 , n19611 , n18927 );
nor ( n19613 , n19610 , n19612 );
not ( n19614 , n19613 );
or ( n19615 , n19609 , n19614 );
nand ( n19616 , n19564 , n18365 );
nand ( n19617 , n19615 , n19616 );
xor ( n19618 , n19608 , n19617 );
not ( n19619 , n18407 );
not ( n19620 , n19494 );
or ( n19621 , n19619 , n19620 );
not ( n19622 , n18153 );
not ( n19623 , n18684 );
or ( n19624 , n19622 , n19623 );
nand ( n19625 , n18683 , n18198 );
nand ( n19626 , n19624 , n19625 );
nand ( n19627 , n19626 , n18194 );
nand ( n19628 , n19621 , n19627 );
and ( n19629 , n19618 , n19628 );
and ( n19630 , n19608 , n19617 );
or ( n19631 , n19629 , n19630 );
not ( n19632 , n18898 );
and ( n19633 , n18257 , n18880 );
not ( n19634 , n18257 );
and ( n19635 , n19634 , n18881 );
or ( n19636 , n19633 , n19635 );
not ( n19637 , n19636 );
or ( n19638 , n19632 , n19637 );
nand ( n19639 , n19504 , n18900 );
nand ( n19640 , n19638 , n19639 );
xor ( n19641 , n19508 , n19519 );
xor ( n19642 , n19641 , n19538 );
xor ( n19643 , n19640 , n19642 );
not ( n19644 , n18768 );
not ( n19645 , n18774 );
not ( n19646 , n18221 );
or ( n19647 , n19645 , n19646 );
nand ( n19648 , n18224 , n18813 );
nand ( n19649 , n19647 , n19648 );
not ( n19650 , n19649 );
or ( n19651 , n19644 , n19650 );
nand ( n19652 , n19553 , n18770 );
nand ( n19653 , n19651 , n19652 );
and ( n19654 , n19643 , n19653 );
and ( n19655 , n19640 , n19642 );
or ( n19656 , n19654 , n19655 );
xor ( n19657 , n19631 , n19656 );
xor ( n19658 , n19496 , n19506 );
xor ( n19659 , n19658 , n19541 );
and ( n19660 , n19657 , n19659 );
and ( n19661 , n19631 , n19656 );
or ( n19662 , n19660 , n19661 );
xor ( n19663 , n19597 , n19662 );
xor ( n19664 , n19544 , n19546 );
xor ( n19665 , n19664 , n19572 );
and ( n19666 , n19663 , n19665 );
and ( n19667 , n19597 , n19662 );
or ( n19668 , n19666 , n19667 );
not ( n19669 , n19668 );
and ( n19670 , n19595 , n19669 );
xor ( n19671 , n19597 , n19662 );
xor ( n19672 , n19671 , n19665 );
xor ( n19673 , n19557 , n19566 );
xor ( n19674 , n19673 , n19569 );
not ( n19675 , n18299 );
not ( n19676 , n19606 );
or ( n19677 , n19675 , n19676 );
not ( n19678 , n18030 );
not ( n19679 , n18845 );
or ( n19680 , n19678 , n19679 );
nand ( n19681 , n18844 , n18561 );
nand ( n19682 , n19680 , n19681 );
nand ( n19683 , n19682 , n18338 );
nand ( n19684 , n19677 , n19683 );
xor ( n19685 , n19527 , n19537 );
xor ( n19686 , n19684 , n19685 );
not ( n19687 , n18192 );
not ( n19688 , n19626 );
or ( n19689 , n19687 , n19688 );
not ( n19690 , n18153 );
not ( n19691 , n18780 );
or ( n19692 , n19690 , n19691 );
nand ( n19693 , n18779 , n18198 );
nand ( n19694 , n19692 , n19693 );
nand ( n19695 , n19694 , n18194 );
nand ( n19696 , n19689 , n19695 );
and ( n19697 , n19686 , n19696 );
and ( n19698 , n19684 , n19685 );
or ( n19699 , n19697 , n19698 );
xor ( n19700 , n19608 , n19617 );
xor ( n19701 , n19700 , n19628 );
xor ( n19702 , n19699 , n19701 );
not ( n19703 , n18359 );
not ( n19704 , n18369 );
not ( n19705 , n19704 );
not ( n19706 , n18698 );
or ( n19707 , n19705 , n19706 );
not ( n19708 , n19704 );
nand ( n19709 , n18697 , n19708 );
nand ( n19710 , n19707 , n19709 );
not ( n19711 , n19710 );
or ( n19712 , n19703 , n19711 );
nand ( n19713 , n19613 , n18365 );
nand ( n19714 , n19712 , n19713 );
and ( n19715 , n18031 , n19178 );
not ( n19716 , n18299 );
not ( n19717 , n19682 );
or ( n19718 , n19716 , n19717 );
not ( n19719 , n18030 );
not ( n19720 , n19513 );
or ( n19721 , n19719 , n19720 );
nand ( n19722 , n19112 , n18561 );
nand ( n19723 , n19721 , n19722 );
nand ( n19724 , n19723 , n18338 );
nand ( n19725 , n19718 , n19724 );
xor ( n19726 , n19715 , n19725 );
not ( n19727 , n18407 );
not ( n19728 , n19694 );
or ( n19729 , n19727 , n19728 );
not ( n19730 , n18153 );
not ( n19731 , n19602 );
or ( n19732 , n19730 , n19731 );
nand ( n19733 , n18810 , n18154 );
nand ( n19734 , n19732 , n19733 );
nand ( n19735 , n19734 , n18193 );
nand ( n19736 , n19729 , n19735 );
and ( n19737 , n19726 , n19736 );
and ( n19738 , n19715 , n19725 );
or ( n19739 , n19737 , n19738 );
xor ( n19740 , n19714 , n19739 );
not ( n19741 , n18900 );
not ( n19742 , n19636 );
or ( n19743 , n19741 , n19742 );
and ( n19744 , n18377 , n18963 );
not ( n19745 , n18377 );
and ( n19746 , n19745 , n18881 );
or ( n19747 , n19744 , n19746 );
nand ( n19748 , n19747 , n18898 );
nand ( n19749 , n19743 , n19748 );
and ( n19750 , n19740 , n19749 );
and ( n19751 , n19714 , n19739 );
or ( n19752 , n19750 , n19751 );
and ( n19753 , n19702 , n19752 );
and ( n19754 , n19699 , n19701 );
or ( n19755 , n19753 , n19754 );
xor ( n19756 , n19674 , n19755 );
xor ( n19757 , n19631 , n19656 );
xor ( n19758 , n19757 , n19659 );
and ( n19759 , n19756 , n19758 );
and ( n19760 , n19674 , n19755 );
or ( n19761 , n19759 , n19760 );
nor ( n19762 , n19672 , n19761 );
nor ( n19763 , n19670 , n19762 );
not ( n19764 , n19763 );
xor ( n19765 , n19674 , n19755 );
xor ( n19766 , n19765 , n19758 );
xor ( n19767 , n19640 , n19642 );
xor ( n19768 , n19767 , n19653 );
not ( n19769 , n18770 );
not ( n19770 , n19649 );
or ( n19771 , n19769 , n19770 );
not ( n19772 , n19549 );
not ( n19773 , n18276 );
or ( n19774 , n19772 , n19773 );
not ( n19775 , n18774 );
nand ( n19776 , n19775 , n18275 );
nand ( n19777 , n19774 , n19776 );
nand ( n19778 , n19777 , n18768 );
nand ( n19779 , n19771 , n19778 );
xor ( n19780 , n19684 , n19685 );
xor ( n19781 , n19780 , n19696 );
xor ( n19782 , n19779 , n19781 );
nand ( n19783 , n18198 , n2458 );
and ( n19784 , n19783 , n19178 );
not ( n19785 , n3177 );
not ( n19786 , n18153 );
or ( n19787 , n19785 , n19786 );
nand ( n19788 , n19787 , n18030 );
nor ( n19789 , n19784 , n19788 );
not ( n19790 , n18299 );
not ( n19791 , n19723 );
or ( n19792 , n19790 , n19791 );
not ( n19793 , n18337 );
not ( n19794 , n18030 );
not ( n19795 , n19177 );
or ( n19796 , n19794 , n19795 );
nand ( n19797 , n18561 , n19178 );
nand ( n19798 , n19796 , n19797 );
nand ( n19799 , n19793 , n19798 );
nand ( n19800 , n19792 , n19799 );
and ( n19801 , n19789 , n19800 );
not ( n19802 , n19747 );
not ( n19803 , n18900 );
or ( n19804 , n19802 , n19803 );
not ( n19805 , n18905 );
not ( n19806 , n18649 );
or ( n19807 , n19805 , n19806 );
nand ( n19808 , n18482 , n18963 );
nand ( n19809 , n19807 , n19808 );
nand ( n19810 , n19809 , n18898 );
nand ( n19811 , n19804 , n19810 );
xor ( n19812 , n19801 , n19811 );
not ( n19813 , n18359 );
not ( n19814 , n18370 );
not ( n19815 , n18684 );
or ( n19816 , n19814 , n19815 );
nand ( n19817 , n19255 , n19708 );
nand ( n19818 , n19816 , n19817 );
not ( n19819 , n19818 );
or ( n19820 , n19813 , n19819 );
nand ( n19821 , n19710 , n18365 );
nand ( n19822 , n19820 , n19821 );
and ( n19823 , n19812 , n19822 );
and ( n19824 , n19801 , n19811 );
or ( n19825 , n19823 , n19824 );
and ( n19826 , n19782 , n19825 );
and ( n19827 , n19779 , n19781 );
or ( n19828 , n19826 , n19827 );
xor ( n19829 , n19768 , n19828 );
xor ( n19830 , n19699 , n19701 );
xor ( n19831 , n19830 , n19752 );
and ( n19832 , n19829 , n19831 );
and ( n19833 , n19768 , n19828 );
or ( n19834 , n19832 , n19833 );
nor ( n19835 , n19766 , n19834 );
xor ( n19836 , n19768 , n19828 );
xor ( n19837 , n19836 , n19831 );
xor ( n19838 , n19714 , n19739 );
xor ( n19839 , n19838 , n19749 );
xor ( n19840 , n19715 , n19725 );
xor ( n19841 , n19840 , n19736 );
not ( n19842 , n18768 );
not ( n19843 , n18774 );
not ( n19844 , n18258 );
or ( n19845 , n19843 , n19844 );
nand ( n19846 , n18257 , n18813 );
nand ( n19847 , n19845 , n19846 );
not ( n19848 , n19847 );
or ( n19849 , n19842 , n19848 );
nand ( n19850 , n19777 , n18770 );
nand ( n19851 , n19849 , n19850 );
xor ( n19852 , n19841 , n19851 );
not ( n19853 , n18407 );
not ( n19854 , n19734 );
or ( n19855 , n19853 , n19854 );
not ( n19856 , n18153 );
not ( n19857 , n18845 );
or ( n19858 , n19856 , n19857 );
nand ( n19859 , n18844 , n18154 );
nand ( n19860 , n19858 , n19859 );
nand ( n19861 , n19860 , n18193 );
nand ( n19862 , n19855 , n19861 );
xor ( n19863 , n19789 , n19800 );
xor ( n19864 , n19862 , n19863 );
not ( n19865 , n18900 );
not ( n19866 , n19809 );
or ( n19867 , n19865 , n19866 );
not ( n19868 , n18881 );
not ( n19869 , n18698 );
or ( n19870 , n19868 , n19869 );
not ( n19871 , n18905 );
nand ( n19872 , n19871 , n18697 );
nand ( n19873 , n19870 , n19872 );
nand ( n19874 , n19873 , n18898 );
nand ( n19875 , n19867 , n19874 );
and ( n19876 , n19864 , n19875 );
and ( n19877 , n19862 , n19863 );
or ( n19878 , n19876 , n19877 );
and ( n19879 , n19852 , n19878 );
and ( n19880 , n19841 , n19851 );
or ( n19881 , n19879 , n19880 );
xor ( n19882 , n19839 , n19881 );
xor ( n19883 , n19779 , n19781 );
xor ( n19884 , n19883 , n19825 );
and ( n19885 , n19882 , n19884 );
and ( n19886 , n19839 , n19881 );
or ( n19887 , n19885 , n19886 );
nor ( n19888 , n19837 , n19887 );
nor ( n19889 , n19835 , n19888 );
not ( n19890 , n19889 );
xor ( n19891 , n19839 , n19881 );
xor ( n19892 , n19891 , n19884 );
not ( n19893 , n19892 );
xor ( n19894 , n19801 , n19811 );
xor ( n19895 , n19894 , n19822 );
not ( n19896 , n18365 );
not ( n19897 , n19818 );
or ( n19898 , n19896 , n19897 );
not ( n19899 , n18925 );
not ( n19900 , n18780 );
or ( n19901 , n19899 , n19900 );
buf ( n19902 , n18367 );
nand ( n19903 , n18779 , n19902 );
nand ( n19904 , n19901 , n19903 );
nand ( n19905 , n19904 , n18359 );
nand ( n19906 , n19898 , n19905 );
and ( n19907 , n18299 , n19178 );
not ( n19908 , n18407 );
not ( n19909 , n19860 );
or ( n19910 , n19908 , n19909 );
not ( n19911 , n19111 );
and ( n19912 , n18153 , n19911 );
not ( n19913 , n18153 );
and ( n19914 , n19913 , n19112 );
or ( n19915 , n19912 , n19914 );
nand ( n19916 , n19915 , n18193 );
nand ( n19917 , n19910 , n19916 );
xor ( n19918 , n19907 , n19917 );
not ( n19919 , n18364 );
not ( n19920 , n19904 );
or ( n19921 , n19919 , n19920 );
and ( n19922 , n18810 , n18368 );
not ( n19923 , n18810 );
not ( n19924 , n19902 );
and ( n19925 , n19923 , n19924 );
or ( n19926 , n19922 , n19925 );
nand ( n19927 , n19926 , n18359 );
nand ( n19928 , n19921 , n19927 );
and ( n19929 , n19918 , n19928 );
and ( n19930 , n19907 , n19917 );
or ( n19931 , n19929 , n19930 );
xor ( n19932 , n19906 , n19931 );
not ( n19933 , n18770 );
not ( n19934 , n19847 );
or ( n19935 , n19933 , n19934 );
not ( n19936 , n18774 );
not ( n19937 , n18656 );
or ( n19938 , n19936 , n19937 );
not ( n19939 , n19549 );
nand ( n19940 , n19939 , n18377 );
nand ( n19941 , n19938 , n19940 );
nand ( n19942 , n19941 , n18768 );
nand ( n19943 , n19935 , n19942 );
and ( n19944 , n19932 , n19943 );
and ( n19945 , n19906 , n19931 );
or ( n19946 , n19944 , n19945 );
xor ( n19947 , n19895 , n19946 );
xor ( n19948 , n19841 , n19851 );
xor ( n19949 , n19948 , n19878 );
and ( n19950 , n19947 , n19949 );
and ( n19951 , n19895 , n19946 );
or ( n19952 , n19950 , n19951 );
not ( n19953 , n19952 );
and ( n19954 , n19893 , n19953 );
xor ( n19955 , n19895 , n19946 );
xor ( n19956 , n19955 , n19949 );
nand ( n19957 , n19902 , n18190 );
and ( n19958 , n19957 , n19178 );
not ( n19959 , n18183 );
not ( n19960 , n18367 );
not ( n19961 , n19960 );
or ( n19962 , n19959 , n19961 );
nand ( n19963 , n19962 , n18153 );
nor ( n19964 , n19958 , n19963 );
not ( n19965 , n18192 );
not ( n19966 , n19915 );
or ( n19967 , n19965 , n19966 );
nor ( n19968 , n18184 , n18192 );
not ( n19969 , n19178 );
not ( n19970 , n18198 );
or ( n19971 , n19969 , n19970 );
nand ( n19972 , n19177 , n18153 );
nand ( n19973 , n19971 , n19972 );
nand ( n19974 , n19968 , n19973 );
nand ( n19975 , n19967 , n19974 );
and ( n19976 , n19964 , n19975 );
not ( n19977 , n18898 );
and ( n19978 , n18905 , n18684 );
not ( n19979 , n18905 );
and ( n19980 , n19979 , n18683 );
or ( n19981 , n19978 , n19980 );
not ( n19982 , n19981 );
or ( n19983 , n19977 , n19982 );
nand ( n19984 , n19873 , n18900 );
nand ( n19985 , n19983 , n19984 );
xor ( n19986 , n19976 , n19985 );
not ( n19987 , n18770 );
not ( n19988 , n19941 );
or ( n19989 , n19987 , n19988 );
not ( n19990 , n18774 );
not ( n19991 , n18649 );
or ( n19992 , n19990 , n19991 );
not ( n19993 , n19549 );
nand ( n19994 , n19993 , n18482 );
nand ( n19995 , n19992 , n19994 );
nand ( n19996 , n19995 , n18768 );
nand ( n19997 , n19989 , n19996 );
and ( n19998 , n19986 , n19997 );
and ( n19999 , n19976 , n19985 );
or ( n20000 , n19998 , n19999 );
xor ( n20001 , n19862 , n19863 );
xor ( n20002 , n20001 , n19875 );
xor ( n20003 , n20000 , n20002 );
xor ( n20004 , n19906 , n19931 );
xor ( n20005 , n20004 , n19943 );
and ( n20006 , n20003 , n20005 );
and ( n20007 , n20000 , n20002 );
or ( n20008 , n20006 , n20007 );
nor ( n20009 , n19956 , n20008 );
nor ( n20010 , n19954 , n20009 );
not ( n20011 , n20010 );
xor ( n20012 , n19907 , n19917 );
xor ( n20013 , n20012 , n19928 );
not ( n20014 , n18364 );
not ( n20015 , n19926 );
or ( n20016 , n20014 , n20015 );
not ( n20017 , n18368 );
not ( n20018 , n20017 );
not ( n20019 , n19096 );
or ( n20020 , n20018 , n20019 );
nand ( n20021 , n18844 , n19902 );
nand ( n20022 , n20020 , n20021 );
nand ( n20023 , n20022 , n18358 );
nand ( n20024 , n20016 , n20023 );
xor ( n20025 , n19964 , n19975 );
xor ( n20026 , n20024 , n20025 );
not ( n20027 , n18900 );
not ( n20028 , n19981 );
or ( n20029 , n20027 , n20028 );
not ( n20030 , n18905 );
not ( n20031 , n18780 );
or ( n20032 , n20030 , n20031 );
nand ( n20033 , n18779 , n19073 );
nand ( n20034 , n20032 , n20033 );
nand ( n20035 , n20034 , n18898 );
nand ( n20036 , n20029 , n20035 );
and ( n20037 , n20026 , n20036 );
and ( n20038 , n20024 , n20025 );
or ( n20039 , n20037 , n20038 );
xor ( n20040 , n20013 , n20039 );
xor ( n20041 , n19976 , n19985 );
xor ( n20042 , n20041 , n19997 );
and ( n20043 , n20040 , n20042 );
and ( n20044 , n20013 , n20039 );
or ( n20045 , n20043 , n20044 );
not ( n20046 , n20045 );
xor ( n20047 , n20000 , n20002 );
xor ( n20048 , n20047 , n20005 );
not ( n20049 , n20048 );
nand ( n20050 , n20046 , n20049 );
not ( n20051 , n20050 );
xor ( n20052 , n20013 , n20039 );
xor ( n20053 , n20052 , n20042 );
not ( n20054 , n20053 );
not ( n20055 , n18770 );
not ( n20056 , n19995 );
or ( n20057 , n20055 , n20056 );
xor ( n20058 , n19549 , n18697 );
nand ( n20059 , n20058 , n18768 );
nand ( n20060 , n20057 , n20059 );
nor ( n20061 , n18197 , n19177 );
not ( n20062 , n18364 );
not ( n20063 , n20022 );
or ( n20064 , n20062 , n20063 );
not ( n20065 , n18367 );
not ( n20066 , n20065 );
not ( n20067 , n19911 );
or ( n20068 , n20066 , n20067 );
nand ( n20069 , n19111 , n18367 );
nand ( n20070 , n20068 , n20069 );
nand ( n20071 , n18358 , n20070 );
nand ( n20072 , n20064 , n20071 );
xor ( n20073 , n20061 , n20072 );
not ( n20074 , n2259 );
nand ( n20075 , n20074 , n18880 );
and ( n20076 , n20075 , n19190 );
not ( n20077 , n2259 );
not ( n20078 , n18905 );
or ( n20079 , n20077 , n20078 );
nand ( n20080 , n20079 , n19960 );
nor ( n20081 , n20076 , n20080 );
not ( n20082 , n18364 );
not ( n20083 , n20070 );
or ( n20084 , n20082 , n20083 );
not ( n20085 , n18357 );
not ( n20086 , n19178 );
not ( n20087 , n18367 );
or ( n20088 , n20086 , n20087 );
not ( n20089 , n19190 );
not ( n20090 , n18367 );
nand ( n20091 , n20089 , n20090 );
nand ( n20092 , n20088 , n20091 );
nand ( n20093 , n20085 , n20092 );
nand ( n20094 , n20084 , n20093 );
and ( n20095 , n20081 , n20094 );
and ( n20096 , n20073 , n20095 );
and ( n20097 , n20061 , n20072 );
or ( n20098 , n20096 , n20097 );
xor ( n20099 , n20060 , n20098 );
xor ( n20100 , n20024 , n20025 );
xor ( n20101 , n20100 , n20036 );
and ( n20102 , n20099 , n20101 );
and ( n20103 , n20060 , n20098 );
or ( n20104 , n20102 , n20103 );
not ( n20105 , n20104 );
nand ( n20106 , n20054 , n20105 );
not ( n20107 , n20106 );
nor ( n20108 , n18351 , n19177 );
not ( n20109 , n18900 );
and ( n20110 , n18844 , n18347 );
not ( n20111 , n18844 );
and ( n20112 , n20111 , n18348 );
nor ( n20113 , n20110 , n20112 );
not ( n20114 , n20113 );
or ( n20115 , n20109 , n20114 );
not ( n20116 , n18347 );
not ( n20117 , n19911 );
or ( n20118 , n20116 , n20117 );
nand ( n20119 , n19111 , n18348 );
nand ( n20120 , n20118 , n20119 );
nand ( n20121 , n20120 , n18898 );
nand ( n20122 , n20115 , n20121 );
xor ( n20123 , n20108 , n20122 );
not ( n20124 , n18897 );
and ( n20125 , n19176 , n18348 );
not ( n20126 , n19176 );
and ( n20127 , n20126 , n18905 );
nor ( n20128 , n20125 , n20127 );
not ( n20129 , n20128 );
and ( n20130 , n20124 , n20129 );
and ( n20131 , n18900 , n20120 );
nor ( n20132 , n20130 , n20131 );
not ( n20133 , n18889 );
and ( n20134 , n18773 , n20133 );
nor ( n20135 , n20134 , n18348 );
or ( n20136 , n19549 , n20133 );
nand ( n20137 , n20136 , n19190 );
nand ( n20138 , n20135 , n20137 );
nor ( n20139 , n20132 , n20138 );
xor ( n20140 , n20123 , n20139 );
not ( n20141 , n18770 );
not ( n20142 , n19549 );
not ( n20143 , n18780 );
or ( n20144 , n20142 , n20143 );
nand ( n20145 , n18779 , n18772 );
nand ( n20146 , n20144 , n20145 );
not ( n20147 , n20146 );
or ( n20148 , n20141 , n20147 );
not ( n20149 , n18772 );
not ( n20150 , n18810 );
not ( n20151 , n20150 );
or ( n20152 , n20149 , n20151 );
or ( n20153 , n20150 , n18772 );
nand ( n20154 , n20152 , n20153 );
not ( n20155 , n20154 );
nand ( n20156 , n20155 , n18768 );
nand ( n20157 , n20148 , n20156 );
or ( n20158 , n20140 , n20157 );
and ( n20159 , n18844 , n18773 );
not ( n20160 , n18844 );
and ( n20161 , n20160 , n18772 );
nor ( n20162 , n20159 , n20161 );
not ( n20163 , n20162 );
not ( n20164 , n18768 );
or ( n20165 , n20163 , n20164 );
or ( n20166 , n20154 , n19159 );
nand ( n20167 , n20165 , n20166 );
xor ( n20168 , n20138 , n20132 );
xor ( n20169 , n20167 , n20168 );
nor ( n20170 , n18896 , n19177 );
not ( n20171 , n18770 );
not ( n20172 , n20162 );
or ( n20173 , n20171 , n20172 );
not ( n20174 , n18773 );
not ( n20175 , n19911 );
or ( n20176 , n20174 , n20175 );
nand ( n20177 , n19111 , n18772 );
nand ( n20178 , n20176 , n20177 );
nand ( n20179 , n20178 , n18768 );
nand ( n20180 , n20173 , n20179 );
xor ( n20181 , n20170 , n20180 );
and ( n20182 , n20178 , n18770 );
nand ( n20183 , n19549 , n19177 );
nand ( n20184 , n18772 , n19190 );
and ( n20185 , n20183 , n20184 );
nor ( n20186 , n20185 , n18767 );
nor ( n20187 , n20182 , n20186 );
nand ( n20188 , n19178 , n18770 );
nand ( n20189 , n20188 , n18773 );
nor ( n20190 , n20187 , n20189 );
and ( n20191 , n20181 , n20190 );
and ( n20192 , n20170 , n20180 );
or ( n20193 , n20191 , n20192 );
and ( n20194 , n20169 , n20193 );
and ( n20195 , n20167 , n20168 );
or ( n20196 , n20194 , n20195 );
and ( n20197 , n20158 , n20196 );
nand ( n20198 , n20140 , n20157 );
not ( n20199 , n20198 );
nor ( n20200 , n20197 , n20199 );
not ( n20201 , n18900 );
not ( n20202 , n18905 );
not ( n20203 , n19602 );
or ( n20204 , n20202 , n20203 );
not ( n20205 , n18347 );
nand ( n20206 , n20205 , n18810 );
nand ( n20207 , n20204 , n20206 );
not ( n20208 , n20207 );
or ( n20209 , n20201 , n20208 );
nand ( n20210 , n20113 , n18898 );
nand ( n20211 , n20209 , n20210 );
xor ( n20212 , n20081 , n20094 );
xor ( n20213 , n20211 , n20212 );
not ( n20214 , n18770 );
not ( n20215 , n18684 );
xor ( n20216 , n18773 , n20215 );
not ( n20217 , n20216 );
or ( n20218 , n20214 , n20217 );
nand ( n20219 , n20146 , n18768 );
nand ( n20220 , n20218 , n20219 );
xor ( n20221 , n20213 , n20220 );
xor ( n20222 , n20108 , n20122 );
and ( n20223 , n20222 , n20139 );
and ( n20224 , n20108 , n20122 );
or ( n20225 , n20223 , n20224 );
nor ( n20226 , n20221 , n20225 );
or ( n20227 , n20200 , n20226 );
nand ( n20228 , n20221 , n20225 );
nand ( n20229 , n20227 , n20228 );
not ( n20230 , n18900 );
not ( n20231 , n20034 );
or ( n20232 , n20230 , n20231 );
nand ( n20233 , n20207 , n18898 );
nand ( n20234 , n20232 , n20233 );
not ( n20235 , n18768 );
not ( n20236 , n20216 );
or ( n20237 , n20235 , n20236 );
nand ( n20238 , n20058 , n18770 );
nand ( n20239 , n20237 , n20238 );
xor ( n20240 , n20234 , n20239 );
xor ( n20241 , n20061 , n20072 );
xor ( n20242 , n20241 , n20095 );
xor ( n20243 , n20240 , n20242 );
not ( n20244 , n20243 );
xor ( n20245 , n20211 , n20212 );
and ( n20246 , n20245 , n20220 );
and ( n20247 , n20211 , n20212 );
or ( n20248 , n20246 , n20247 );
not ( n20249 , n20248 );
nand ( n20250 , n20244 , n20249 );
and ( n20251 , n20229 , n20250 );
and ( n20252 , n20243 , n20248 );
nor ( n20253 , n20251 , n20252 );
xor ( n20254 , n20060 , n20098 );
xor ( n20255 , n20254 , n20101 );
xor ( n20256 , n20234 , n20239 );
and ( n20257 , n20256 , n20242 );
and ( n20258 , n20234 , n20239 );
or ( n20259 , n20257 , n20258 );
nor ( n20260 , n20255 , n20259 );
or ( n20261 , n20253 , n20260 );
nand ( n20262 , n20255 , n20259 );
nand ( n20263 , n20261 , n20262 );
not ( n20264 , n20263 );
or ( n20265 , n20107 , n20264 );
nand ( n20266 , n20053 , n20104 );
nand ( n20267 , n20265 , n20266 );
not ( n20268 , n20267 );
or ( n20269 , n20051 , n20268 );
not ( n20270 , n20049 );
nand ( n20271 , n20270 , n20045 );
nand ( n20272 , n20269 , n20271 );
not ( n20273 , n20272 );
or ( n20274 , n20011 , n20273 );
not ( n20275 , n19892 );
not ( n20276 , n19952 );
nand ( n20277 , n20275 , n20276 );
and ( n20278 , n19956 , n20008 );
and ( n20279 , n20277 , n20278 );
nor ( n20280 , n20275 , n20276 );
nor ( n20281 , n20279 , n20280 );
nand ( n20282 , n20274 , n20281 );
not ( n20283 , n20282 );
or ( n20284 , n19890 , n20283 );
nor ( n20285 , n19766 , n19834 );
not ( n20286 , n20285 );
nand ( n20287 , n19837 , n19887 );
not ( n20288 , n20287 );
and ( n20289 , n20286 , n20288 );
and ( n20290 , n19766 , n19834 );
nor ( n20291 , n20289 , n20290 );
nand ( n20292 , n20284 , n20291 );
not ( n20293 , n20292 );
or ( n20294 , n19764 , n20293 );
not ( n20295 , n19594 );
not ( n20296 , n19668 );
nand ( n20297 , n20295 , n20296 );
not ( n20298 , n19672 );
not ( n20299 , n19761 );
nor ( n20300 , n20298 , n20299 );
and ( n20301 , n20297 , n20300 );
and ( n20302 , n19594 , n19668 );
nor ( n20303 , n20301 , n20302 );
nand ( n20304 , n20294 , n20303 );
not ( n20305 , n20304 );
or ( n20306 , n19592 , n20305 );
not ( n20307 , n19590 );
nand ( n20308 , n19444 , n19581 );
not ( n20309 , n20308 );
and ( n20310 , n20307 , n20309 );
and ( n20311 , n19585 , n19589 );
nor ( n20312 , n20310 , n20311 );
nand ( n20313 , n20306 , n20312 );
not ( n20314 , n20313 );
or ( n20315 , n19428 , n20314 );
not ( n20316 , n19426 );
nand ( n20317 , n19314 , n19316 );
or ( n20318 , n19234 , n20317 );
nand ( n20319 , n19064 , n19233 );
nand ( n20320 , n20318 , n20319 );
not ( n20321 , n20320 );
or ( n20322 , n20316 , n20321 );
not ( n20323 , n19420 );
nand ( n20324 , n20323 , n19424 );
nand ( n20325 , n20322 , n20324 );
not ( n20326 , n19384 );
nand ( n20327 , n19416 , n20326 );
and ( n20328 , n20325 , n20327 );
nor ( n20329 , n19416 , n20326 );
nor ( n20330 , n20328 , n20329 );
nand ( n20331 , n20315 , n20330 );
not ( n20332 , n20331 );
xor ( n20333 , n19397 , n19409 );
and ( n20334 , n20333 , n19414 );
and ( n20335 , n19397 , n19409 );
or ( n20336 , n20334 , n20335 );
xor ( n20337 , n19389 , n19393 );
and ( n20338 , n20337 , n19396 );
and ( n20339 , n19389 , n19393 );
or ( n20340 , n20338 , n20339 );
xor ( n20341 , n18535 , n18537 );
xor ( n20342 , n20341 , n18540 );
xor ( n20343 , n20340 , n20342 );
xor ( n20344 , n19399 , n19403 );
and ( n20345 , n20344 , n19408 );
and ( n20346 , n19399 , n19403 );
or ( n20347 , n20345 , n20346 );
xor ( n20348 , n20343 , n20347 );
or ( n20349 , n20336 , n20348 );
xor ( n20350 , n18345 , n18514 );
xor ( n20351 , n20350 , n18543 );
xor ( n20352 , n20340 , n20342 );
and ( n20353 , n20352 , n20347 );
and ( n20354 , n20340 , n20342 );
or ( n20355 , n20353 , n20354 );
nor ( n20356 , n20351 , n20355 );
not ( n20357 , n20356 );
nand ( n20358 , n20349 , n20357 );
not ( n20359 , n20358 );
not ( n20360 , n20359 );
or ( n20361 , n20332 , n20360 );
nand ( n20362 , n20336 , n20348 );
not ( n20363 , n20362 );
not ( n20364 , n20356 );
and ( n20365 , n20363 , n20364 );
and ( n20366 , n20351 , n20355 );
nor ( n20367 , n20365 , n20366 );
nand ( n20368 , n20361 , n20367 );
not ( n20369 , n20368 );
or ( n20370 , n18646 , n20369 );
nand ( n20371 , n18546 , n18598 );
or ( n20372 , n18644 , n20371 );
nand ( n20373 , n18604 , n18643 );
nand ( n20374 , n20372 , n20373 );
not ( n20375 , n20374 );
nand ( n20376 , n20370 , n20375 );
or ( n20377 , n18338 , n18300 );
nand ( n20378 , n20377 , n18302 );
not ( n20379 , n18149 );
or ( n20380 , n18438 , n18122 );
or ( n20381 , n18180 , n18041 );
nand ( n20382 , n20380 , n20381 );
not ( n20383 , n20382 );
or ( n20384 , n20379 , n20383 );
nand ( n20385 , n18613 , n18039 );
nand ( n20386 , n20384 , n20385 );
xor ( n20387 , n20378 , n20386 );
and ( n20388 , n18245 , n18118 );
xor ( n20389 , n20387 , n20388 );
not ( n20390 , n18242 );
not ( n20391 , n18620 );
or ( n20392 , n20390 , n20391 );
and ( n20393 , n18244 , n18318 );
not ( n20394 , n18244 );
and ( n20395 , n20394 , n18321 );
nor ( n20396 , n20393 , n20395 );
or ( n20397 , n20396 , n18289 );
nand ( n20398 , n20392 , n20397 );
xor ( n20399 , n20398 , n18626 );
xor ( n20400 , n18605 , n18615 );
and ( n20401 , n20400 , n18622 );
and ( n20402 , n18605 , n18615 );
or ( n20403 , n20401 , n20402 );
xor ( n20404 , n20399 , n20403 );
xor ( n20405 , n20389 , n20404 );
xor ( n20406 , n18627 , n18631 );
and ( n20407 , n20406 , n18636 );
and ( n20408 , n18627 , n18631 );
or ( n20409 , n20407 , n20408 );
xor ( n20410 , n20405 , n20409 );
xor ( n20411 , n18623 , n18637 );
and ( n20412 , n20411 , n18642 );
and ( n20413 , n18623 , n18637 );
or ( n20414 , n20412 , n20413 );
or ( n20415 , n20410 , n20414 );
nand ( n20416 , n20414 , n20410 );
nand ( n20417 , n20415 , n20416 );
not ( n20418 , n20417 );
and ( n20419 , n20376 , n20418 );
not ( n20420 , n20376 );
and ( n20421 , n20420 , n20417 );
nor ( n20422 , n20419 , n20421 );
and ( n20423 , n18029 , n20422 );
not ( n20424 , n18029 );
not ( n20425 , n20422 );
and ( n20426 , n20424 , n20425 );
nor ( n20427 , n20423 , n20426 );
not ( n20428 , n20427 );
or ( n20429 , n18026 , n20428 );
and ( n20430 , n18645 , n20415 );
not ( n20431 , n20430 );
not ( n20432 , n20368 );
or ( n20433 , n20431 , n20432 );
and ( n20434 , n20374 , n20415 );
not ( n20435 , n20416 );
nor ( n20436 , n20434 , n20435 );
nand ( n20437 , n20433 , n20436 );
xor ( n20438 , n20389 , n20404 );
and ( n20439 , n20438 , n20409 );
and ( n20440 , n20389 , n20404 );
or ( n20441 , n20439 , n20440 );
xor ( n20442 , n20378 , n20386 );
and ( n20443 , n20442 , n20388 );
and ( n20444 , n20378 , n20386 );
or ( n20445 , n20443 , n20444 );
or ( n20446 , n20396 , n18241 );
not ( n20447 , n18402 );
not ( n20448 , n18244 );
and ( n20449 , n20447 , n20448 );
and ( n20450 , n18402 , n18244 );
nor ( n20451 , n20449 , n20450 );
or ( n20452 , n20451 , n18289 );
nand ( n20453 , n20446 , n20452 );
and ( n20454 , n18245 , n18145 );
xor ( n20455 , n20453 , n20454 );
and ( n20456 , n20382 , n18039 );
and ( n20457 , n18149 , n18041 );
nor ( n20458 , n20456 , n20457 );
xor ( n20459 , n20455 , n20458 );
xor ( n20460 , n20445 , n20459 );
xor ( n20461 , n20398 , n18626 );
and ( n20462 , n20461 , n20403 );
and ( n20463 , n20398 , n18626 );
or ( n20464 , n20462 , n20463 );
xor ( n20465 , n20460 , n20464 );
or ( n20466 , n20441 , n20465 );
nand ( n20467 , n20441 , n20465 );
nand ( n20468 , n20466 , n20467 );
and ( n20469 , n20437 , n20468 );
not ( n20470 , n20437 );
not ( n20471 , n20468 );
and ( n20472 , n20470 , n20471 );
nor ( n20473 , n20469 , n20472 );
not ( n20474 , n20473 );
and ( n20475 , n18029 , n20474 );
not ( n20476 , n18029 );
not ( n20477 , n20474 );
and ( n20478 , n20476 , n20477 );
nor ( n20479 , n20475 , n20478 );
nand ( n20480 , n20479 , n18012 );
nand ( n20481 , n20429 , n20480 );
nor ( n20482 , n524 , n540 );
not ( n20483 , n20482 );
nand ( n20484 , n524 , n540 );
and ( n20485 , n20483 , n20484 );
nand ( n20486 , n536 , n552 );
not ( n20487 , n20486 );
not ( n20488 , n18015 );
or ( n20489 , n20487 , n20488 );
nor ( n20490 , n534 , n550 );
nor ( n20491 , n18017 , n20490 );
nand ( n20492 , n20489 , n20491 );
nand ( n20493 , n533 , n549 );
nand ( n20494 , n534 , n550 );
nand ( n20495 , n20492 , n20493 , n20494 );
not ( n20496 , n20495 );
nor ( n20497 , n529 , n545 );
nor ( n20498 , n533 , n549 );
nor ( n20499 , n530 , n546 );
nor ( n20500 , n20497 , n20498 , n20499 );
nor ( n20501 , n531 , n547 );
nor ( n20502 , n532 , n548 );
nor ( n20503 , n20501 , n20502 );
and ( n20504 , n20500 , n20503 );
not ( n20505 , n20504 );
or ( n20506 , n20496 , n20505 );
nand ( n20507 , n530 , n546 );
nand ( n20508 , n529 , n545 );
nand ( n20509 , n531 , n547 );
and ( n20510 , n20507 , n20508 , n20509 );
not ( n20511 , n20510 );
not ( n20512 , n20501 );
nand ( n20513 , n532 , n548 );
not ( n20514 , n20513 );
nand ( n20515 , n20512 , n20514 );
not ( n20516 , n20515 );
or ( n20517 , n20511 , n20516 );
not ( n20518 , n20499 );
not ( n20519 , n20518 );
not ( n20520 , n20497 );
not ( n20521 , n20520 );
or ( n20522 , n20519 , n20521 );
nand ( n20523 , n20522 , n20508 );
nand ( n20524 , n20517 , n20523 );
nand ( n20525 , n20506 , n20524 );
not ( n20526 , n20525 );
nor ( n20527 , n525 , n541 );
nor ( n20528 , n526 , n542 );
nor ( n20529 , n20527 , n20528 );
nor ( n20530 , n527 , n543 );
nor ( n20531 , n528 , n544 );
nor ( n20532 , n20530 , n20531 );
nand ( n20533 , n20529 , n20532 );
not ( n20534 , n20533 );
not ( n20535 , n20534 );
or ( n20536 , n20526 , n20535 );
nand ( n20537 , n528 , n544 );
or ( n20538 , n20530 , n20537 );
nand ( n20539 , n527 , n543 );
nand ( n20540 , n20538 , n20539 );
not ( n20541 , n20540 );
not ( n20542 , n20529 );
or ( n20543 , n20541 , n20542 );
not ( n20544 , n20527 );
nand ( n20545 , n526 , n542 );
not ( n20546 , n20545 );
and ( n20547 , n20544 , n20546 );
and ( n20548 , n525 , n541 );
nor ( n20549 , n20547 , n20548 );
nand ( n20550 , n20543 , n20549 );
not ( n20551 , n20550 );
nand ( n20552 , n20536 , n20551 );
xor ( n20553 , n20485 , n20552 );
not ( n20554 , n20553 );
not ( n20555 , n20554 );
nor ( n20556 , n20527 , n20548 );
not ( n20557 , n20528 );
and ( n20558 , n20532 , n20557 );
not ( n20559 , n20558 );
not ( n20560 , n20525 );
or ( n20561 , n20559 , n20560 );
and ( n20562 , n20540 , n20557 );
not ( n20563 , n20545 );
nor ( n20564 , n20562 , n20563 );
nand ( n20565 , n20561 , n20564 );
xor ( n20566 , n20556 , n20565 );
not ( n20567 , n20566 );
or ( n20568 , n20555 , n20567 );
not ( n20569 , n20566 );
nand ( n20570 , n20569 , n20553 );
nand ( n20571 , n20568 , n20570 );
not ( n20572 , n20571 );
not ( n20573 , n20554 );
nor ( n20574 , n20533 , n20482 );
not ( n20575 , n20574 );
not ( n20576 , n20495 );
not ( n20577 , n20504 );
or ( n20578 , n20576 , n20577 );
nand ( n20579 , n20578 , n20524 );
not ( n20580 , n20579 );
or ( n20581 , n20575 , n20580 );
not ( n20582 , n20483 );
not ( n20583 , n20550 );
or ( n20584 , n20582 , n20583 );
nand ( n20585 , n20584 , n20484 );
not ( n20586 , n20585 );
nand ( n20587 , n20581 , n20586 );
nor ( n20588 , n523 , n539 );
not ( n20589 , n20588 );
nand ( n20590 , n523 , n539 );
nand ( n20591 , n20589 , n20590 );
not ( n20592 , n20591 );
and ( n20593 , n20587 , n20592 );
not ( n20594 , n20587 );
and ( n20595 , n20594 , n20591 );
nor ( n20596 , n20593 , n20595 );
not ( n20597 , n20596 );
or ( n20598 , n20573 , n20597 );
or ( n20599 , n20596 , n20554 );
nand ( n20600 , n20598 , n20599 );
nand ( n20601 , n20572 , n20600 );
not ( n20602 , n20601 );
not ( n20603 , n20602 );
not ( n20604 , n20592 );
not ( n20605 , n20587 );
not ( n20606 , n20605 );
or ( n20607 , n20604 , n20606 );
nand ( n20608 , n20587 , n20591 );
nand ( n20609 , n20607 , n20608 );
not ( n20610 , n19888 );
and ( n20611 , n20282 , n20610 );
not ( n20612 , n20287 );
nor ( n20613 , n20611 , n20612 );
xor ( n20614 , n19766 , n19834 );
and ( n20615 , n20613 , n20614 );
not ( n20616 , n20613 );
or ( n20617 , n19835 , n20290 );
and ( n20618 , n20616 , n20617 );
nor ( n20619 , n20615 , n20618 );
not ( n20620 , n20619 );
and ( n20621 , n20609 , n20620 );
not ( n20622 , n20609 );
not ( n20623 , n20620 );
and ( n20624 , n20622 , n20623 );
nor ( n20625 , n20621 , n20624 );
not ( n20626 , n20625 );
or ( n20627 , n20603 , n20626 );
buf ( n20628 , n20609 );
not ( n20629 , n20628 );
nand ( n20630 , n19672 , n19761 );
not ( n20631 , n19672 );
nand ( n20632 , n20631 , n20299 );
nand ( n20633 , n20630 , n20632 );
not ( n20634 , n20633 );
not ( n20635 , n20634 );
not ( n20636 , n20292 );
not ( n20637 , n20636 );
or ( n20638 , n20635 , n20637 );
nand ( n20639 , n20292 , n20633 );
nand ( n20640 , n20638 , n20639 );
not ( n20641 , n20640 );
not ( n20642 , n20641 );
or ( n20643 , n20629 , n20642 );
not ( n20644 , n20609 );
nand ( n20645 , n20640 , n20644 );
nand ( n20646 , n20643 , n20645 );
buf ( n20647 , n20571 );
nand ( n20648 , n20646 , n20647 );
nand ( n20649 , n20627 , n20648 );
nor ( n20650 , n20588 , n20482 );
nor ( n20651 , n522 , n538 );
nor ( n20652 , n521 , n537 );
nor ( n20653 , n20651 , n20652 );
and ( n20654 , n20650 , n20653 );
not ( n20655 , n20654 );
nor ( n20656 , n20655 , n20533 );
not ( n20657 , n20656 );
not ( n20658 , n20579 );
or ( n20659 , n20657 , n20658 );
and ( n20660 , n20654 , n20550 );
not ( n20661 , n20653 );
not ( n20662 , n20484 );
not ( n20663 , n20662 );
not ( n20664 , n20589 );
or ( n20665 , n20663 , n20664 );
nand ( n20666 , n20665 , n20590 );
not ( n20667 , n20666 );
or ( n20668 , n20661 , n20667 );
nand ( n20669 , n522 , n538 );
nor ( n20670 , n20669 , n20652 );
and ( n20671 , n521 , n537 );
nor ( n20672 , n20670 , n20671 );
nand ( n20673 , n20668 , n20672 );
nor ( n20674 , n20660 , n20673 );
nand ( n20675 , n20659 , n20674 );
nor ( n20676 , n20671 , n20652 );
not ( n20677 , n20651 );
and ( n20678 , n20650 , n20677 );
not ( n20679 , n20678 );
nor ( n20680 , n20679 , n20533 );
not ( n20681 , n20680 );
not ( n20682 , n20525 );
or ( n20683 , n20681 , n20682 );
and ( n20684 , n20678 , n20550 );
not ( n20685 , n20677 );
not ( n20686 , n20666 );
or ( n20687 , n20685 , n20686 );
nand ( n20688 , n20687 , n20669 );
nor ( n20689 , n20684 , n20688 );
nand ( n20690 , n20683 , n20689 );
xor ( n20691 , n20676 , n20690 );
xnor ( n20692 , n20675 , n20691 );
not ( n20693 , n20692 );
not ( n20694 , n20693 );
buf ( n20695 , n20267 );
xor ( n20696 , n20045 , n20048 );
not ( n20697 , n20696 );
and ( n20698 , n20695 , n20697 );
not ( n20699 , n20695 );
and ( n20700 , n20699 , n20696 );
nor ( n20701 , n20698 , n20700 );
buf ( n20702 , n20701 );
not ( n20703 , n20702 );
not ( n20704 , n20703 );
or ( n20705 , n20694 , n20704 );
and ( n20706 , n20266 , n20106 );
buf ( n20707 , n20263 );
xor ( n20708 , n20706 , n20707 );
not ( n20709 , n20708 );
nand ( n20710 , n20692 , n20675 );
or ( n20711 , n20709 , n20710 );
nand ( n20712 , n20705 , n20711 );
not ( n20713 , n20609 );
not ( n20714 , n20650 );
nor ( n20715 , n20714 , n20533 );
not ( n20716 , n20715 );
not ( n20717 , n20579 );
or ( n20718 , n20716 , n20717 );
and ( n20719 , n20650 , n20550 );
nor ( n20720 , n20719 , n20666 );
nand ( n20721 , n20718 , n20720 );
nand ( n20722 , n20677 , n20669 );
xnor ( n20723 , n20721 , n20722 );
not ( n20724 , n20723 );
or ( n20725 , n20713 , n20724 );
or ( n20726 , n20596 , n20723 );
nand ( n20727 , n20725 , n20726 );
not ( n20728 , n20727 );
not ( n20729 , n20728 );
buf ( n20730 , n20691 );
not ( n20731 , n20730 );
not ( n20732 , n20277 );
nor ( n20733 , n20732 , n20280 );
or ( n20734 , n19956 , n20008 );
not ( n20735 , n20734 );
not ( n20736 , n20272 );
or ( n20737 , n20735 , n20736 );
not ( n20738 , n20278 );
nand ( n20739 , n20737 , n20738 );
xor ( n20740 , n20733 , n20739 );
buf ( n20741 , n20740 );
not ( n20742 , n20741 );
not ( n20743 , n20742 );
or ( n20744 , n20731 , n20743 );
not ( n20745 , n20730 );
nand ( n20746 , n20741 , n20745 );
nand ( n20747 , n20744 , n20746 );
not ( n20748 , n20747 );
or ( n20749 , n20729 , n20748 );
nand ( n20750 , n20738 , n20734 );
xnor ( n20751 , n20272 , n20750 );
not ( n20752 , n20751 );
not ( n20753 , n20752 );
and ( n20754 , n20730 , n20753 );
not ( n20755 , n20730 );
and ( n20756 , n20755 , n20752 );
nor ( n20757 , n20754 , n20756 );
and ( n20758 , n20723 , n20691 );
not ( n20759 , n20723 );
not ( n20760 , n20691 );
and ( n20761 , n20759 , n20760 );
nor ( n20762 , n20758 , n20761 );
and ( n20763 , n20762 , n20727 );
not ( n20764 , n20763 );
not ( n20765 , n20764 );
nand ( n20766 , n20757 , n20765 );
nand ( n20767 , n20749 , n20766 );
and ( n20768 , n20712 , n20767 );
xor ( n20769 , n20649 , n20768 );
not ( n20770 , n20693 );
not ( n20771 , n20753 );
or ( n20772 , n20770 , n20771 );
or ( n20773 , n20702 , n20710 );
nand ( n20774 , n20772 , n20773 );
not ( n20775 , n20765 );
not ( n20776 , n20747 );
or ( n20777 , n20775 , n20776 );
not ( n20778 , n20730 );
nand ( n20779 , n20610 , n20287 );
not ( n20780 , n20779 );
buf ( n20781 , n20282 );
not ( n20782 , n20781 );
not ( n20783 , n20782 );
or ( n20784 , n20780 , n20783 );
not ( n20785 , n20779 );
nand ( n20786 , n20785 , n20781 );
nand ( n20787 , n20784 , n20786 );
not ( n20788 , n20787 );
or ( n20789 , n20778 , n20788 );
not ( n20790 , n20779 );
not ( n20791 , n20782 );
or ( n20792 , n20790 , n20791 );
nand ( n20793 , n20792 , n20786 );
not ( n20794 , n20793 );
nand ( n20795 , n20794 , n20745 );
nand ( n20796 , n20789 , n20795 );
nand ( n20797 , n20796 , n20728 );
nand ( n20798 , n20777 , n20797 );
xor ( n20799 , n20774 , n20798 );
xor ( n20800 , n20769 , n20799 );
not ( n20801 , n20503 );
nor ( n20802 , n20801 , n20499 );
not ( n20803 , n20802 );
nor ( n20804 , n20490 , n20498 );
not ( n20805 , n20804 );
or ( n20806 , n18017 , n20486 );
nand ( n20807 , n20806 , n18015 );
not ( n20808 , n20807 );
or ( n20809 , n20805 , n20808 );
nor ( n20810 , n533 , n549 );
or ( n20811 , n20810 , n20494 );
nand ( n20812 , n20811 , n20493 );
not ( n20813 , n20812 );
nand ( n20814 , n20809 , n20813 );
not ( n20815 , n20814 );
or ( n20816 , n20803 , n20815 );
nand ( n20817 , n20515 , n20509 );
and ( n20818 , n20817 , n20518 );
not ( n20819 , n20507 );
nor ( n20820 , n20818 , n20819 );
nand ( n20821 , n20816 , n20820 );
nand ( n20822 , n20520 , n20508 );
not ( n20823 , n20822 );
and ( n20824 , n20821 , n20823 );
not ( n20825 , n20821 );
and ( n20826 , n20825 , n20822 );
nor ( n20827 , n20824 , n20826 );
buf ( n20828 , n20827 );
nand ( n20829 , n20518 , n20507 );
not ( n20830 , n20503 );
not ( n20831 , n20814 );
or ( n20832 , n20830 , n20831 );
not ( n20833 , n20817 );
nand ( n20834 , n20832 , n20833 );
xnor ( n20835 , n20829 , n20834 );
and ( n20836 , n20828 , n20835 );
not ( n20837 , n20828 );
not ( n20838 , n20835 );
and ( n20839 , n20837 , n20838 );
nor ( n20840 , n20836 , n20839 );
not ( n20841 , n20840 );
not ( n20842 , n20838 );
not ( n20843 , n20502 );
not ( n20844 , n20843 );
not ( n20845 , n20814 );
or ( n20846 , n20844 , n20845 );
nand ( n20847 , n20846 , n20513 );
nand ( n20848 , n20512 , n20509 );
not ( n20849 , n20848 );
and ( n20850 , n20847 , n20849 );
not ( n20851 , n20847 );
and ( n20852 , n20851 , n20848 );
nor ( n20853 , n20850 , n20852 );
not ( n20854 , n20853 );
or ( n20855 , n20842 , n20854 );
not ( n20856 , n20853 );
nand ( n20857 , n20835 , n20856 );
nand ( n20858 , n20855 , n20857 );
nor ( n20859 , n20841 , n20858 );
buf ( n20860 , n20859 );
not ( n20861 , n20860 );
not ( n20862 , n20827 );
not ( n20863 , n20862 );
not ( n20864 , n20863 );
not ( n20865 , n19317 );
not ( n20866 , n20865 );
not ( n20867 , n20313 );
or ( n20868 , n20866 , n20867 );
nand ( n20869 , n20868 , n20317 );
not ( n20870 , n19234 );
nand ( n20871 , n20870 , n20319 );
nor ( n20872 , n20869 , n20871 );
and ( n20873 , n20869 , n20871 );
or ( n20874 , n20872 , n20873 );
not ( n20875 , n20874 );
not ( n20876 , n20875 );
or ( n20877 , n20864 , n20876 );
buf ( n20878 , n20874 );
nand ( n20879 , n20878 , n20862 );
nand ( n20880 , n20877 , n20879 );
not ( n20881 , n20880 );
or ( n20882 , n20861 , n20881 );
not ( n20883 , n20863 );
and ( n20884 , n19425 , n19419 );
not ( n20885 , n19425 );
and ( n20886 , n20885 , n19420 );
nor ( n20887 , n20884 , n20886 );
not ( n20888 , n20887 );
not ( n20889 , n20888 );
not ( n20890 , n20313 );
not ( n20891 , n19318 );
or ( n20892 , n20890 , n20891 );
not ( n20893 , n20320 );
nand ( n20894 , n20892 , n20893 );
not ( n20895 , n20894 );
not ( n20896 , n20895 );
or ( n20897 , n20889 , n20896 );
nand ( n20898 , n20894 , n20887 );
nand ( n20899 , n20897 , n20898 );
not ( n20900 , n20899 );
not ( n20901 , n20900 );
or ( n20902 , n20883 , n20901 );
nand ( n20903 , n20899 , n20862 );
nand ( n20904 , n20902 , n20903 );
buf ( n20905 , n20858 );
nand ( n20906 , n20904 , n20905 );
nand ( n20907 , n20882 , n20906 );
xor ( n20908 , n20800 , n20907 );
not ( n20909 , n20532 );
not ( n20910 , n20579 );
or ( n20911 , n20909 , n20910 );
not ( n20912 , n20540 );
nand ( n20913 , n20911 , n20912 );
nand ( n20914 , n20557 , n20545 );
xor ( n20915 , n20913 , n20914 );
not ( n20916 , n20531 );
not ( n20917 , n20916 );
not ( n20918 , n20525 );
or ( n20919 , n20917 , n20918 );
nand ( n20920 , n20919 , n20537 );
not ( n20921 , n20530 );
nand ( n20922 , n20921 , n20539 );
and ( n20923 , n20920 , n20922 );
not ( n20924 , n20920 );
not ( n20925 , n20922 );
and ( n20926 , n20924 , n20925 );
nor ( n20927 , n20923 , n20926 );
and ( n20928 , n20915 , n20927 );
not ( n20929 , n20915 );
not ( n20930 , n20927 );
and ( n20931 , n20929 , n20930 );
or ( n20932 , n20928 , n20931 );
not ( n20933 , n20932 );
not ( n20934 , n20933 );
buf ( n20935 , n20566 );
not ( n20936 , n20935 );
or ( n20937 , n19444 , n19581 );
nand ( n20938 , n20937 , n20308 );
not ( n20939 , n20938 );
not ( n20940 , n20939 );
not ( n20941 , n20304 );
not ( n20942 , n20941 );
or ( n20943 , n20940 , n20942 );
nand ( n20944 , n20304 , n20938 );
nand ( n20945 , n20943 , n20944 );
not ( n20946 , n20945 );
not ( n20947 , n20946 );
or ( n20948 , n20936 , n20947 );
not ( n20949 , n20939 );
not ( n20950 , n20941 );
or ( n20951 , n20949 , n20950 );
nand ( n20952 , n20951 , n20944 );
not ( n20953 , n20935 );
nand ( n20954 , n20952 , n20953 );
nand ( n20955 , n20948 , n20954 );
not ( n20956 , n20955 );
or ( n20957 , n20934 , n20956 );
not ( n20958 , n20302 );
nand ( n20959 , n20958 , n20297 );
not ( n20960 , n20632 );
not ( n20961 , n20292 );
or ( n20962 , n20960 , n20961 );
nand ( n20963 , n20962 , n20630 );
and ( n20964 , n20959 , n20963 );
not ( n20965 , n20959 );
not ( n20966 , n20963 );
and ( n20967 , n20965 , n20966 );
nor ( n20968 , n20964 , n20967 );
not ( n20969 , n20968 );
and ( n20970 , n20935 , n20969 );
not ( n20971 , n20935 );
buf ( n20972 , n20968 );
and ( n20973 , n20971 , n20972 );
nor ( n20974 , n20970 , n20973 );
and ( n20975 , n20915 , n20569 );
not ( n20976 , n20915 );
and ( n20977 , n20976 , n20566 );
nor ( n20978 , n20975 , n20977 );
and ( n20979 , n20978 , n20932 );
buf ( n20980 , n20979 );
nand ( n20981 , n20974 , n20980 );
nand ( n20982 , n20957 , n20981 );
buf ( n20983 , n20930 );
nor ( n20984 , n19590 , n20311 );
and ( n20985 , n20304 , n20937 );
not ( n20986 , n20308 );
nor ( n20987 , n20985 , n20986 );
and ( n20988 , n20984 , n20987 );
not ( n20989 , n20984 );
not ( n20990 , n20987 );
and ( n20991 , n20989 , n20990 );
or ( n20992 , n20988 , n20991 );
and ( n20993 , n20983 , n20992 );
not ( n20994 , n20983 );
not ( n20995 , n20992 );
and ( n20996 , n20994 , n20995 );
nor ( n20997 , n20993 , n20996 );
not ( n20998 , n20997 );
and ( n20999 , n20916 , n20537 );
xor ( n21000 , n20999 , n20579 );
xor ( n21001 , n21000 , n20930 );
xnor ( n21002 , n21000 , n20827 );
and ( n21003 , n21001 , n21002 );
not ( n21004 , n21003 );
or ( n21005 , n20998 , n21004 );
nand ( n21006 , n20865 , n20317 );
not ( n21007 , n20313 );
not ( n21008 , n21007 );
and ( n21009 , n21006 , n21008 );
not ( n21010 , n21006 );
and ( n21011 , n21010 , n21007 );
or ( n21012 , n21009 , n21011 );
buf ( n21013 , n21012 );
and ( n21014 , n20983 , n21013 );
not ( n21015 , n20983 );
not ( n21016 , n21012 );
and ( n21017 , n21015 , n21016 );
nor ( n21018 , n21014 , n21017 );
not ( n21019 , n21002 );
buf ( n21020 , n21019 );
nand ( n21021 , n21018 , n21020 );
nand ( n21022 , n21005 , n21021 );
xor ( n21023 , n20982 , n21022 );
not ( n21024 , n20728 );
not ( n21025 , n20757 );
or ( n21026 , n21024 , n21025 );
and ( n21027 , n20730 , n20702 );
not ( n21028 , n20730 );
and ( n21029 , n21028 , n20703 );
nor ( n21030 , n21027 , n21029 );
or ( n21031 , n21030 , n20764 );
nand ( n21032 , n21026 , n21031 );
not ( n21033 , n21032 );
not ( n21034 , n20253 );
not ( n21035 , n21034 );
or ( n21036 , n20255 , n20259 );
nand ( n21037 , n21036 , n20262 );
not ( n21038 , n21037 );
or ( n21039 , n21035 , n21038 );
not ( n21040 , n21037 );
not ( n21041 , n21034 );
nand ( n21042 , n21040 , n21041 );
nand ( n21043 , n21039 , n21042 );
buf ( n21044 , n21043 );
not ( n21045 , n20710 );
and ( n21046 , n21044 , n21045 );
not ( n21047 , n20709 );
and ( n21048 , n21047 , n20693 );
nor ( n21049 , n21046 , n21048 );
nor ( n21050 , n21033 , n21049 );
not ( n21051 , n20647 );
not ( n21052 , n20625 );
or ( n21053 , n21051 , n21052 );
and ( n21054 , n20628 , n20794 );
not ( n21055 , n20628 );
and ( n21056 , n21055 , n20787 );
nor ( n21057 , n21054 , n21056 );
nand ( n21058 , n21057 , n20602 );
nand ( n21059 , n21053 , n21058 );
xor ( n21060 , n21050 , n21059 );
xor ( n21061 , n20712 , n20767 );
and ( n21062 , n21060 , n21061 );
and ( n21063 , n21050 , n21059 );
or ( n21064 , n21062 , n21063 );
xor ( n21065 , n21023 , n21064 );
and ( n21066 , n20908 , n21065 );
and ( n21067 , n20800 , n20907 );
or ( n21068 , n21066 , n21067 );
xor ( n21069 , n20481 , n21068 );
not ( n21070 , n21049 );
not ( n21071 , n21032 );
or ( n21072 , n21070 , n21071 );
or ( n21073 , n21032 , n21049 );
nand ( n21074 , n21072 , n21073 );
not ( n21075 , n20647 );
not ( n21076 , n21057 );
or ( n21077 , n21075 , n21076 );
and ( n21078 , n20609 , n20741 );
not ( n21079 , n20609 );
and ( n21080 , n21079 , n20742 );
nor ( n21081 , n21078 , n21080 );
nand ( n21082 , n21081 , n20602 );
nand ( n21083 , n21077 , n21082 );
and ( n21084 , n21074 , n21083 );
not ( n21085 , n20933 );
not ( n21086 , n20974 );
or ( n21087 , n21085 , n21086 );
buf ( n21088 , n20640 );
and ( n21089 , n20935 , n21088 );
not ( n21090 , n20935 );
and ( n21091 , n21090 , n20641 );
nor ( n21092 , n21089 , n21091 );
nand ( n21093 , n21092 , n20980 );
nand ( n21094 , n21087 , n21093 );
xor ( n21095 , n21084 , n21094 );
xor ( n21096 , n21050 , n21059 );
xor ( n21097 , n21096 , n21061 );
and ( n21098 , n21095 , n21097 );
and ( n21099 , n21084 , n21094 );
or ( n21100 , n21098 , n21099 );
not ( n21101 , n20494 );
nor ( n21102 , n21101 , n20490 );
xor ( n21103 , n21102 , n20807 );
xor ( n21104 , n21103 , n18023 );
buf ( n21105 , n21104 );
not ( n21106 , n21105 );
and ( n21107 , n20492 , n20494 );
not ( n21108 , n20810 );
nand ( n21109 , n21108 , n20493 );
xor ( n21110 , n21107 , n21109 );
buf ( n21111 , n21110 );
not ( n21112 , n21111 );
nand ( n21113 , n18599 , n20371 );
not ( n21114 , n21113 );
and ( n21115 , n20368 , n21114 );
not ( n21116 , n20368 );
and ( n21117 , n21116 , n21113 );
nor ( n21118 , n21115 , n21117 );
not ( n21119 , n21118 );
not ( n21120 , n21119 );
or ( n21121 , n21112 , n21120 );
not ( n21122 , n21110 );
not ( n21123 , n21122 );
not ( n21124 , n21123 );
nand ( n21125 , n21118 , n21124 );
nand ( n21126 , n21121 , n21125 );
not ( n21127 , n21126 );
or ( n21128 , n21106 , n21127 );
not ( n21129 , n21111 );
not ( n21130 , n20349 );
not ( n21131 , n20331 );
or ( n21132 , n21130 , n21131 );
buf ( n21133 , n20362 );
nand ( n21134 , n21132 , n21133 );
not ( n21135 , n20357 );
nor ( n21136 , n21135 , n20366 );
xor ( n21137 , n21134 , n21136 );
not ( n21138 , n21137 );
not ( n21139 , n21138 );
or ( n21140 , n21129 , n21139 );
nand ( n21141 , n21137 , n21124 );
nand ( n21142 , n21140 , n21141 );
not ( n21143 , n21104 );
and ( n21144 , n21111 , n21103 );
nor ( n21145 , n21111 , n21103 );
nor ( n21146 , n21144 , n21145 );
and ( n21147 , n21143 , n21146 );
buf ( n21148 , n21147 );
nand ( n21149 , n21142 , n21148 );
nand ( n21150 , n21128 , n21149 );
xor ( n21151 , n21100 , n21150 );
nor ( n21152 , n20514 , n20502 );
xor ( n21153 , n21152 , n20814 );
xor ( n21154 , n21153 , n20853 );
not ( n21155 , n21110 );
not ( n21156 , n21155 );
not ( n21157 , n21153 );
not ( n21158 , n21157 );
or ( n21159 , n21156 , n21158 );
nand ( n21160 , n21153 , n21110 );
nand ( n21161 , n21159 , n21160 );
and ( n21162 , n21154 , n21161 );
buf ( n21163 , n21162 );
not ( n21164 , n21163 );
not ( n21165 , n20856 );
not ( n21166 , n21165 );
not ( n21167 , n21166 );
buf ( n21168 , n19426 );
nand ( n21169 , n20894 , n21168 );
and ( n21170 , n21169 , n20324 );
not ( n21171 , n20327 );
nor ( n21172 , n21171 , n20329 );
nor ( n21173 , n21170 , n21172 );
and ( n21174 , n21168 , n20894 );
nand ( n21175 , n21172 , n20324 );
nor ( n21176 , n21174 , n21175 );
nor ( n21177 , n21173 , n21176 );
not ( n21178 , n21177 );
and ( n21179 , n21167 , n21178 );
not ( n21180 , n21167 );
not ( n21181 , n21178 );
and ( n21182 , n21180 , n21181 );
nor ( n21183 , n21179 , n21182 );
not ( n21184 , n21183 );
or ( n21185 , n21164 , n21184 );
and ( n21186 , n21133 , n20349 );
buf ( n21187 , n20331 );
not ( n21188 , n21187 );
and ( n21189 , n21186 , n21188 );
not ( n21190 , n21186 );
and ( n21191 , n21190 , n21187 );
or ( n21192 , n21189 , n21191 );
buf ( n21193 , n21192 );
and ( n21194 , n21167 , n21193 );
not ( n21195 , n21167 );
not ( n21196 , n21192 );
and ( n21197 , n21195 , n21196 );
nor ( n21198 , n21194 , n21197 );
not ( n21199 , n21161 );
nand ( n21200 , n21198 , n21199 );
nand ( n21201 , n21185 , n21200 );
and ( n21202 , n21151 , n21201 );
and ( n21203 , n21100 , n21150 );
or ( n21204 , n21202 , n21203 );
xor ( n21205 , n21069 , n21204 );
xor ( n21206 , n20800 , n20907 );
xor ( n21207 , n21206 , n21065 );
xor ( n21208 , n21100 , n21150 );
xor ( n21209 , n21208 , n21201 );
xor ( n21210 , n21207 , n21209 );
xor ( n21211 , n21083 , n21074 );
not ( n21212 , n20905 );
not ( n21213 , n20862 );
and ( n21214 , n21213 , n21013 );
not ( n21215 , n21213 );
and ( n21216 , n21215 , n21016 );
nor ( n21217 , n21214 , n21216 );
not ( n21218 , n21217 );
or ( n21219 , n21212 , n21218 );
not ( n21220 , n20863 );
not ( n21221 , n20995 );
or ( n21222 , n21220 , n21221 );
nand ( n21223 , n20992 , n20862 );
nand ( n21224 , n21222 , n21223 );
nand ( n21225 , n21224 , n20860 );
nand ( n21226 , n21219 , n21225 );
xor ( n21227 , n21211 , n21226 );
not ( n21228 , n20765 );
not ( n21229 , n20730 );
not ( n21230 , n21044 );
or ( n21231 , n21229 , n21230 );
or ( n21232 , n21044 , n20730 );
nand ( n21233 , n21231 , n21232 );
not ( n21234 , n21233 );
not ( n21235 , n21234 );
or ( n21236 , n21228 , n21235 );
and ( n21237 , n20745 , n21047 );
not ( n21238 , n20745 );
and ( n21239 , n21238 , n20709 );
nor ( n21240 , n21237 , n21239 );
not ( n21241 , n21240 );
nand ( n21242 , n21241 , n20728 );
nand ( n21243 , n21236 , n21242 );
not ( n21244 , n20693 );
not ( n21245 , n20252 );
nand ( n21246 , n21245 , n20250 );
not ( n21247 , n20200 );
not ( n21248 , n20226 );
and ( n21249 , n21247 , n21248 );
not ( n21250 , n20228 );
nor ( n21251 , n21249 , n21250 );
and ( n21252 , n21246 , n21251 );
not ( n21253 , n21246 );
and ( n21254 , n21253 , n20229 );
nor ( n21255 , n21252 , n21254 );
not ( n21256 , n21255 );
not ( n21257 , n21256 );
not ( n21258 , n21257 );
or ( n21259 , n21244 , n21258 );
not ( n21260 , n20226 );
nand ( n21261 , n21260 , n20228 );
not ( n21262 , n21261 );
not ( n21263 , n21262 );
not ( n21264 , n20200 );
or ( n21265 , n21263 , n21264 );
not ( n21266 , n20200 );
nand ( n21267 , n21261 , n21266 );
nand ( n21268 , n21265 , n21267 );
not ( n21269 , n21268 );
or ( n21270 , n21269 , n20710 );
nand ( n21271 , n21259 , n21270 );
xor ( n21272 , n21243 , n21271 );
not ( n21273 , n20647 );
not ( n21274 , n20609 );
not ( n21275 , n20752 );
or ( n21276 , n21274 , n21275 );
nand ( n21277 , n20753 , n20644 );
nand ( n21278 , n21276 , n21277 );
not ( n21279 , n21278 );
or ( n21280 , n21273 , n21279 );
not ( n21281 , n20609 );
not ( n21282 , n20702 );
or ( n21283 , n21281 , n21282 );
nand ( n21284 , n20703 , n20644 );
nand ( n21285 , n21283 , n21284 );
nand ( n21286 , n21285 , n20602 );
nand ( n21287 , n21280 , n21286 );
and ( n21288 , n21272 , n21287 );
and ( n21289 , n21243 , n21271 );
or ( n21290 , n21288 , n21289 );
not ( n21291 , n21290 );
not ( n21292 , n20933 );
and ( n21293 , n20935 , n20620 );
not ( n21294 , n20935 );
and ( n21295 , n21294 , n20623 );
nor ( n21296 , n21293 , n21295 );
not ( n21297 , n21296 );
or ( n21298 , n21292 , n21297 );
and ( n21299 , n20935 , n20794 );
not ( n21300 , n20935 );
and ( n21301 , n21300 , n20787 );
nor ( n21302 , n21299 , n21301 );
nand ( n21303 , n21302 , n20979 );
nand ( n21304 , n21298 , n21303 );
not ( n21305 , n21304 );
or ( n21306 , n21291 , n21305 );
not ( n21307 , n21290 );
not ( n21308 , n21307 );
not ( n21309 , n21304 );
not ( n21310 , n21309 );
or ( n21311 , n21308 , n21310 );
buf ( n21312 , n21256 );
or ( n21313 , n21312 , n20710 );
not ( n21314 , n21043 );
or ( n21315 , n21314 , n20692 );
nand ( n21316 , n21313 , n21315 );
or ( n21317 , n21240 , n20764 );
not ( n21318 , n20728 );
or ( n21319 , n21030 , n21318 );
nand ( n21320 , n21317 , n21319 );
xor ( n21321 , n21316 , n21320 );
not ( n21322 , n20647 );
not ( n21323 , n21081 );
or ( n21324 , n21322 , n21323 );
nand ( n21325 , n21278 , n20602 );
nand ( n21326 , n21324 , n21325 );
xor ( n21327 , n21321 , n21326 );
nand ( n21328 , n21311 , n21327 );
nand ( n21329 , n21306 , n21328 );
and ( n21330 , n21227 , n21329 );
and ( n21331 , n21211 , n21226 );
or ( n21332 , n21330 , n21331 );
not ( n21333 , n21020 );
not ( n21334 , n21333 );
not ( n21335 , n21334 );
not ( n21336 , n20997 );
or ( n21337 , n21335 , n21336 );
and ( n21338 , n20983 , n20952 );
not ( n21339 , n20983 );
and ( n21340 , n21339 , n20946 );
nor ( n21341 , n21338 , n21340 );
nand ( n21342 , n21341 , n21003 );
nand ( n21343 , n21337 , n21342 );
not ( n21344 , n20979 );
not ( n21345 , n21296 );
or ( n21346 , n21344 , n21345 );
nand ( n21347 , n21092 , n20933 );
nand ( n21348 , n21346 , n21347 );
not ( n21349 , n21348 );
not ( n21350 , n21349 );
not ( n21351 , n21003 );
and ( n21352 , n20983 , n20969 );
not ( n21353 , n20983 );
and ( n21354 , n21353 , n20972 );
nor ( n21355 , n21352 , n21354 );
not ( n21356 , n21355 );
or ( n21357 , n21351 , n21356 );
nand ( n21358 , n21341 , n21020 );
nand ( n21359 , n21357 , n21358 );
not ( n21360 , n21359 );
not ( n21361 , n21360 );
or ( n21362 , n21350 , n21361 );
xor ( n21363 , n21316 , n21320 );
and ( n21364 , n21363 , n21326 );
and ( n21365 , n21316 , n21320 );
or ( n21366 , n21364 , n21365 );
nand ( n21367 , n21362 , n21366 );
not ( n21368 , n21349 );
nand ( n21369 , n21368 , n21359 );
nand ( n21370 , n21367 , n21369 );
xor ( n21371 , n21343 , n21370 );
not ( n21372 , n20905 );
not ( n21373 , n20880 );
or ( n21374 , n21372 , n21373 );
nand ( n21375 , n21217 , n20860 );
nand ( n21376 , n21374 , n21375 );
xor ( n21377 , n21371 , n21376 );
xor ( n21378 , n21332 , n21377 );
not ( n21379 , n18012 );
not ( n21380 , n18029 );
not ( n21381 , n18599 );
not ( n21382 , n20368 );
or ( n21383 , n21381 , n21382 );
nand ( n21384 , n21383 , n20371 );
not ( n21385 , n18644 );
nand ( n21386 , n21385 , n20373 );
and ( n21387 , n21384 , n21386 );
not ( n21388 , n21384 );
not ( n21389 , n21386 );
and ( n21390 , n21388 , n21389 );
nor ( n21391 , n21387 , n21390 );
not ( n21392 , n21391 );
or ( n21393 , n21380 , n21392 );
not ( n21394 , n21391 );
nand ( n21395 , n21394 , n18028 );
nand ( n21396 , n21393 , n21395 );
not ( n21397 , n21396 );
or ( n21398 , n21379 , n21397 );
and ( n21399 , n18028 , n21119 );
not ( n21400 , n18028 );
and ( n21401 , n21400 , n21118 );
nor ( n21402 , n21399 , n21401 );
nand ( n21403 , n21402 , n18025 );
nand ( n21404 , n21398 , n21403 );
and ( n21405 , n21378 , n21404 );
and ( n21406 , n21332 , n21377 );
or ( n21407 , n21405 , n21406 );
and ( n21408 , n21210 , n21407 );
and ( n21409 , n21207 , n21209 );
or ( n21410 , n21408 , n21409 );
xor ( n21411 , n21205 , n21410 );
and ( n21412 , n20774 , n20798 );
not ( n21413 , n20628 );
not ( n21414 , n20972 );
or ( n21415 , n21413 , n21414 );
nand ( n21416 , n20969 , n20644 );
nand ( n21417 , n21415 , n21416 );
not ( n21418 , n21417 );
or ( n21419 , n21418 , n20572 );
nand ( n21420 , n20646 , n20602 );
nand ( n21421 , n21419 , n21420 );
xor ( n21422 , n21412 , n21421 );
not ( n21423 , n20763 );
not ( n21424 , n20796 );
or ( n21425 , n21423 , n21424 );
not ( n21426 , n21318 );
not ( n21427 , n20730 );
not ( n21428 , n20623 );
or ( n21429 , n21427 , n21428 );
nand ( n21430 , n20620 , n20745 );
nand ( n21431 , n21429 , n21430 );
nand ( n21432 , n21426 , n21431 );
nand ( n21433 , n21425 , n21432 );
not ( n21434 , n20752 );
not ( n21435 , n20710 );
and ( n21436 , n21434 , n21435 );
and ( n21437 , n20741 , n20693 );
nor ( n21438 , n21436 , n21437 );
xnor ( n21439 , n21433 , n21438 );
xor ( n21440 , n21422 , n21439 );
not ( n21441 , n21163 );
not ( n21442 , n21198 );
or ( n21443 , n21441 , n21442 );
not ( n21444 , n21167 );
not ( n21445 , n21138 );
or ( n21446 , n21444 , n21445 );
nand ( n21447 , n21137 , n21166 );
nand ( n21448 , n21446 , n21447 );
nand ( n21449 , n21448 , n21199 );
nand ( n21450 , n21443 , n21449 );
xor ( n21451 , n21440 , n21450 );
not ( n21452 , n20905 );
and ( n21453 , n21213 , n21178 );
not ( n21454 , n21213 );
and ( n21455 , n21454 , n21181 );
nor ( n21456 , n21453 , n21455 );
not ( n21457 , n21456 );
or ( n21458 , n21452 , n21457 );
nand ( n21459 , n20904 , n20860 );
nand ( n21460 , n21458 , n21459 );
xor ( n21461 , n21451 , n21460 );
xor ( n21462 , n20982 , n21022 );
and ( n21463 , n21462 , n21064 );
and ( n21464 , n20982 , n21022 );
or ( n21465 , n21463 , n21464 );
xor ( n21466 , n20649 , n20768 );
and ( n21467 , n21466 , n20799 );
and ( n21468 , n20649 , n20768 );
or ( n21469 , n21467 , n21468 );
not ( n21470 , n20933 );
not ( n21471 , n20935 );
not ( n21472 , n20995 );
or ( n21473 , n21471 , n21472 );
nand ( n21474 , n20992 , n20953 );
nand ( n21475 , n21473 , n21474 );
not ( n21476 , n21475 );
or ( n21477 , n21470 , n21476 );
nand ( n21478 , n20955 , n20980 );
nand ( n21479 , n21477 , n21478 );
xor ( n21480 , n21469 , n21479 );
not ( n21481 , n21003 );
not ( n21482 , n21018 );
or ( n21483 , n21481 , n21482 );
not ( n21484 , n20983 );
not ( n21485 , n20875 );
or ( n21486 , n21484 , n21485 );
not ( n21487 , n20983 );
nand ( n21488 , n20878 , n21487 );
nand ( n21489 , n21486 , n21488 );
nand ( n21490 , n21489 , n21334 );
nand ( n21491 , n21483 , n21490 );
xor ( n21492 , n21480 , n21491 );
xor ( n21493 , n21465 , n21492 );
not ( n21494 , n21148 );
not ( n21495 , n21126 );
or ( n21496 , n21494 , n21495 );
not ( n21497 , n21111 );
not ( n21498 , n21391 );
or ( n21499 , n21497 , n21498 );
nand ( n21500 , n21394 , n21124 );
nand ( n21501 , n21499 , n21500 );
nand ( n21502 , n21501 , n21105 );
nand ( n21503 , n21496 , n21502 );
xor ( n21504 , n21493 , n21503 );
xor ( n21505 , n21461 , n21504 );
xor ( n21506 , n21343 , n21370 );
and ( n21507 , n21506 , n21376 );
and ( n21508 , n21343 , n21370 );
or ( n21509 , n21507 , n21508 );
not ( n21510 , n21509 );
not ( n21511 , n18025 );
not ( n21512 , n21396 );
or ( n21513 , n21511 , n21512 );
nand ( n21514 , n20427 , n18012 );
nand ( n21515 , n21513 , n21514 );
not ( n21516 , n21515 );
or ( n21517 , n21510 , n21516 );
not ( n21518 , n21509 );
not ( n21519 , n21518 );
not ( n21520 , n21515 );
not ( n21521 , n21520 );
or ( n21522 , n21519 , n21521 );
not ( n21523 , n21105 );
not ( n21524 , n21142 );
or ( n21525 , n21523 , n21524 );
not ( n21526 , n21111 );
not ( n21527 , n21196 );
or ( n21528 , n21526 , n21527 );
nand ( n21529 , n21193 , n21122 );
nand ( n21530 , n21528 , n21529 );
nand ( n21531 , n21530 , n21148 );
nand ( n21532 , n21525 , n21531 );
xor ( n21533 , n21084 , n21094 );
xor ( n21534 , n21533 , n21097 );
xor ( n21535 , n21532 , n21534 );
not ( n21536 , n21163 );
not ( n21537 , n21167 );
not ( n21538 , n20900 );
or ( n21539 , n21537 , n21538 );
nand ( n21540 , n20899 , n21166 );
nand ( n21541 , n21539 , n21540 );
not ( n21542 , n21541 );
or ( n21543 , n21536 , n21542 );
nand ( n21544 , n21183 , n21199 );
nand ( n21545 , n21543 , n21544 );
and ( n21546 , n21535 , n21545 );
and ( n21547 , n21532 , n21534 );
or ( n21548 , n21546 , n21547 );
nand ( n21549 , n21522 , n21548 );
nand ( n21550 , n21517 , n21549 );
xor ( n21551 , n21505 , n21550 );
xnor ( n21552 , n21411 , n21551 );
not ( n21553 , n21509 );
not ( n21554 , n21520 );
or ( n21555 , n21553 , n21554 );
nand ( n21556 , n21518 , n21515 );
nand ( n21557 , n21555 , n21556 );
xnor ( n21558 , n21557 , n21548 );
not ( n21559 , n21558 );
xor ( n21560 , n21207 , n21209 );
xor ( n21561 , n21560 , n21407 );
not ( n21562 , n21561 );
not ( n21563 , n21562 );
or ( n21564 , n21559 , n21563 );
not ( n21565 , n21163 );
not ( n21566 , n21167 );
not ( n21567 , n20875 );
or ( n21568 , n21566 , n21567 );
nand ( n21569 , n20878 , n21166 );
nand ( n21570 , n21568 , n21569 );
not ( n21571 , n21570 );
or ( n21572 , n21565 , n21571 );
nand ( n21573 , n21541 , n21199 );
nand ( n21574 , n21572 , n21573 );
nand ( n21575 , n21360 , n21366 , n21349 );
not ( n21576 , n21366 );
buf ( n21577 , n21348 );
nand ( n21578 , n21576 , n21360 , n21577 );
nand ( n21579 , n21359 , n21366 , n21577 );
nor ( n21580 , n21366 , n21577 );
nand ( n21581 , n21359 , n21580 );
nand ( n21582 , n21575 , n21578 , n21579 , n21581 );
xor ( n21583 , n21574 , n21582 );
not ( n21584 , n21148 );
not ( n21585 , n21111 );
not ( n21586 , n21181 );
or ( n21587 , n21585 , n21586 );
nand ( n21588 , n21178 , n21122 );
nand ( n21589 , n21587 , n21588 );
not ( n21590 , n21589 );
or ( n21591 , n21584 , n21590 );
nand ( n21592 , n21530 , n21105 );
nand ( n21593 , n21591 , n21592 );
and ( n21594 , n21583 , n21593 );
and ( n21595 , n21574 , n21582 );
or ( n21596 , n21594 , n21595 );
xor ( n21597 , n21532 , n21534 );
xor ( n21598 , n21597 , n21545 );
xor ( n21599 , n21596 , n21598 );
and ( n21600 , n20983 , n21088 );
not ( n21601 , n20983 );
and ( n21602 , n21601 , n20641 );
nor ( n21603 , n21600 , n21602 );
not ( n21604 , n21603 );
not ( n21605 , n21003 );
or ( n21606 , n21604 , n21605 );
not ( n21607 , n21355 );
or ( n21608 , n21607 , n21333 );
nand ( n21609 , n21606 , n21608 );
not ( n21610 , n20693 );
not ( n21611 , n21268 );
or ( n21612 , n21610 , n21611 );
and ( n21613 , n20158 , n20198 );
not ( n21614 , n21613 );
buf ( n21615 , n20196 );
nand ( n21616 , n21614 , n21615 );
not ( n21617 , n21615 );
nand ( n21618 , n21613 , n21617 );
nand ( n21619 , n21616 , n21618 );
not ( n21620 , n21619 );
not ( n21621 , n21620 );
not ( n21622 , n21621 );
or ( n21623 , n21622 , n20710 );
nand ( n21624 , n21612 , n21623 );
or ( n21625 , n21233 , n20727 );
and ( n21626 , n20730 , n21312 );
not ( n21627 , n20730 );
and ( n21628 , n21627 , n21257 );
nor ( n21629 , n21626 , n21628 );
or ( n21630 , n21629 , n20764 );
nand ( n21631 , n21625 , n21630 );
xor ( n21632 , n21624 , n21631 );
not ( n21633 , n20647 );
not ( n21634 , n21285 );
or ( n21635 , n21633 , n21634 );
not ( n21636 , n20628 );
not ( n21637 , n20709 );
or ( n21638 , n21636 , n21637 );
nand ( n21639 , n21047 , n20644 );
nand ( n21640 , n21638 , n21639 );
nand ( n21641 , n21640 , n20602 );
nand ( n21642 , n21635 , n21641 );
and ( n21643 , n21632 , n21642 );
and ( n21644 , n21624 , n21631 );
or ( n21645 , n21643 , n21644 );
not ( n21646 , n20933 );
not ( n21647 , n21302 );
or ( n21648 , n21646 , n21647 );
and ( n21649 , n20935 , n20741 );
not ( n21650 , n20935 );
and ( n21651 , n21650 , n20742 );
nor ( n21652 , n21649 , n21651 );
nand ( n21653 , n21652 , n20980 );
nand ( n21654 , n21648 , n21653 );
xor ( n21655 , n21645 , n21654 );
xor ( n21656 , n21243 , n21271 );
xor ( n21657 , n21656 , n21287 );
and ( n21658 , n21655 , n21657 );
and ( n21659 , n21645 , n21654 );
or ( n21660 , n21658 , n21659 );
xor ( n21661 , n21609 , n21660 );
not ( n21662 , n20905 );
not ( n21663 , n21224 );
or ( n21664 , n21662 , n21663 );
and ( n21665 , n20863 , n20945 );
not ( n21666 , n20863 );
and ( n21667 , n21666 , n20946 );
nor ( n21668 , n21665 , n21667 );
nand ( n21669 , n21668 , n20860 );
nand ( n21670 , n21664 , n21669 );
and ( n21671 , n21661 , n21670 );
and ( n21672 , n21609 , n21660 );
or ( n21673 , n21671 , n21672 );
not ( n21674 , n21673 );
not ( n21675 , n18012 );
not ( n21676 , n21402 );
or ( n21677 , n21675 , n21676 );
not ( n21678 , n18029 );
not ( n21679 , n21138 );
or ( n21680 , n21678 , n21679 );
nand ( n21681 , n21137 , n18028 );
nand ( n21682 , n21680 , n21681 );
nand ( n21683 , n21682 , n18025 );
nand ( n21684 , n21677 , n21683 );
not ( n21685 , n21684 );
or ( n21686 , n21674 , n21685 );
and ( n21687 , n21165 , n21013 );
not ( n21688 , n21165 );
and ( n21689 , n21688 , n21016 );
nor ( n21690 , n21687 , n21689 );
not ( n21691 , n21690 );
not ( n21692 , n21163 );
or ( n21693 , n21691 , n21692 );
not ( n21694 , n21570 );
or ( n21695 , n21694 , n21161 );
nand ( n21696 , n21693 , n21695 );
xor ( n21697 , n21290 , n21309 );
xnor ( n21698 , n21697 , n21327 );
or ( n21699 , n21696 , n21698 );
not ( n21700 , n21020 );
not ( n21701 , n21603 );
or ( n21702 , n21700 , n21701 );
and ( n21703 , n20983 , n20620 );
not ( n21704 , n20983 );
and ( n21705 , n21704 , n20623 );
nor ( n21706 , n21703 , n21705 );
nand ( n21707 , n21706 , n21003 );
nand ( n21708 , n21702 , n21707 );
xor ( n21709 , n21624 , n21631 );
xor ( n21710 , n21709 , n21642 );
not ( n21711 , n21710 );
not ( n21712 , n20693 );
not ( n21713 , n21620 );
not ( n21714 , n21713 );
or ( n21715 , n21712 , n21714 );
xor ( n21716 , n20167 , n20168 );
xor ( n21717 , n21716 , n20193 );
not ( n21718 , n21717 );
or ( n21719 , n21718 , n20710 );
nand ( n21720 , n21715 , n21719 );
nor ( n21721 , n21629 , n21318 );
nor ( n21722 , n21261 , n21266 );
not ( n21723 , n21722 );
nand ( n21724 , n21723 , n21267 );
and ( n21725 , n20730 , n21724 );
not ( n21726 , n20730 );
and ( n21727 , n21726 , n21269 );
nor ( n21728 , n21725 , n21727 );
not ( n21729 , n21728 );
nor ( n21730 , n21729 , n20764 );
or ( n21731 , n21721 , n21730 );
xor ( n21732 , n21720 , n21731 );
not ( n21733 , n20647 );
not ( n21734 , n21640 );
or ( n21735 , n21733 , n21734 );
not ( n21736 , n20609 );
not ( n21737 , n21314 );
or ( n21738 , n21736 , n21737 );
nand ( n21739 , n21044 , n20644 );
nand ( n21740 , n21738 , n21739 );
nand ( n21741 , n21740 , n20602 );
nand ( n21742 , n21735 , n21741 );
and ( n21743 , n21732 , n21742 );
and ( n21744 , n21720 , n21731 );
or ( n21745 , n21743 , n21744 );
not ( n21746 , n21745 );
nand ( n21747 , n21711 , n21746 );
not ( n21748 , n21747 );
not ( n21749 , n20979 );
and ( n21750 , n20935 , n20753 );
not ( n21751 , n20935 );
and ( n21752 , n21751 , n20752 );
nor ( n21753 , n21750 , n21752 );
not ( n21754 , n21753 );
or ( n21755 , n21749 , n21754 );
nand ( n21756 , n21652 , n20933 );
nand ( n21757 , n21755 , n21756 );
not ( n21758 , n21757 );
or ( n21759 , n21748 , n21758 );
not ( n21760 , n21746 );
nand ( n21761 , n21760 , n21710 );
nand ( n21762 , n21759 , n21761 );
xor ( n21763 , n21708 , n21762 );
nand ( n21764 , n21668 , n20905 );
and ( n21765 , n20863 , n20969 );
not ( n21766 , n20863 );
and ( n21767 , n21766 , n20972 );
nor ( n21768 , n21765 , n21767 );
nand ( n21769 , n20860 , n21768 );
nand ( n21770 , n21764 , n21769 );
and ( n21771 , n21763 , n21770 );
and ( n21772 , n21708 , n21762 );
or ( n21773 , n21771 , n21772 );
nand ( n21774 , n21699 , n21773 );
nand ( n21775 , n21698 , n21696 );
nand ( n21776 , n21774 , n21775 );
not ( n21777 , n21673 );
not ( n21778 , n21684 );
nand ( n21779 , n21777 , n21778 );
nand ( n21780 , n21776 , n21779 );
nand ( n21781 , n21686 , n21780 );
and ( n21782 , n21599 , n21781 );
and ( n21783 , n21596 , n21598 );
or ( n21784 , n21782 , n21783 );
nand ( n21785 , n21564 , n21784 );
not ( n21786 , n21558 );
nand ( n21787 , n21786 , n21561 );
and ( n21788 , n21785 , n21787 );
nor ( n21789 , n21552 , n21788 );
not ( n21790 , n21789 );
nand ( n21791 , n21552 , n21788 );
nand ( n21792 , n21790 , n21791 );
xor ( n21793 , n21784 , n21558 );
and ( n21794 , n21793 , n21561 );
not ( n21795 , n21793 );
and ( n21796 , n21795 , n21562 );
nor ( n21797 , n21794 , n21796 );
xor ( n21798 , n21596 , n21598 );
xor ( n21799 , n21798 , n21781 );
xor ( n21800 , n21211 , n21226 );
xor ( n21801 , n21800 , n21329 );
xor ( n21802 , n21574 , n21582 );
xor ( n21803 , n21802 , n21593 );
xor ( n21804 , n21801 , n21803 );
not ( n21805 , n18025 );
not ( n21806 , n18029 );
not ( n21807 , n21196 );
or ( n21808 , n21806 , n21807 );
nand ( n21809 , n21193 , n18028 );
nand ( n21810 , n21808 , n21809 );
not ( n21811 , n21810 );
or ( n21812 , n21805 , n21811 );
nand ( n21813 , n21682 , n18012 );
nand ( n21814 , n21812 , n21813 );
xor ( n21815 , n21609 , n21660 );
xor ( n21816 , n21815 , n21670 );
xor ( n21817 , n21814 , n21816 );
not ( n21818 , n21148 );
and ( n21819 , n21111 , n20899 );
not ( n21820 , n21111 );
and ( n21821 , n21820 , n20900 );
nor ( n21822 , n21819 , n21821 );
not ( n21823 , n21822 );
or ( n21824 , n21818 , n21823 );
nand ( n21825 , n21589 , n21105 );
nand ( n21826 , n21824 , n21825 );
and ( n21827 , n21817 , n21826 );
and ( n21828 , n21814 , n21816 );
or ( n21829 , n21827 , n21828 );
and ( n21830 , n21804 , n21829 );
and ( n21831 , n21801 , n21803 );
or ( n21832 , n21830 , n21831 );
not ( n21833 , n21832 );
xor ( n21834 , n21332 , n21377 );
xor ( n21835 , n21834 , n21404 );
not ( n21836 , n21835 );
nand ( n21837 , n21833 , n21836 );
and ( n21838 , n21799 , n21837 );
and ( n21839 , n21835 , n21832 );
nor ( n21840 , n21838 , n21839 );
nand ( n21841 , n21797 , n21840 );
not ( n21842 , n21832 );
not ( n21843 , n21836 );
or ( n21844 , n21842 , n21843 );
nand ( n21845 , n21833 , n21835 );
nand ( n21846 , n21844 , n21845 );
not ( n21847 , n21799 );
and ( n21848 , n21846 , n21847 );
not ( n21849 , n21846 );
and ( n21850 , n21849 , n21799 );
nor ( n21851 , n21848 , n21850 );
xor ( n21852 , n21801 , n21803 );
xor ( n21853 , n21852 , n21829 );
not ( n21854 , n21853 );
not ( n21855 , n21854 );
not ( n21856 , n21778 );
not ( n21857 , n21673 );
and ( n21858 , n21856 , n21857 );
and ( n21859 , n21673 , n21778 );
nor ( n21860 , n21858 , n21859 );
xor ( n21861 , n21860 , n21776 );
not ( n21862 , n21861 );
and ( n21863 , n21855 , n21862 );
nand ( n21864 , n21854 , n21861 );
xor ( n21865 , n21645 , n21654 );
xor ( n21866 , n21865 , n21657 );
not ( n21867 , n21199 );
not ( n21868 , n21690 );
or ( n21869 , n21867 , n21868 );
and ( n21870 , n21165 , n20992 );
not ( n21871 , n21165 );
and ( n21872 , n21871 , n20995 );
nor ( n21873 , n21870 , n21872 );
nand ( n21874 , n21873 , n21162 );
nand ( n21875 , n21869 , n21874 );
buf ( n21876 , n21875 );
xor ( n21877 , n21866 , n21876 );
not ( n21878 , n21105 );
not ( n21879 , n21822 );
or ( n21880 , n21878 , n21879 );
not ( n21881 , n21111 );
not ( n21882 , n20875 );
or ( n21883 , n21881 , n21882 );
nand ( n21884 , n20878 , n21122 );
nand ( n21885 , n21883 , n21884 );
nand ( n21886 , n21885 , n21148 );
nand ( n21887 , n21880 , n21886 );
and ( n21888 , n21877 , n21887 );
and ( n21889 , n21866 , n21876 );
or ( n21890 , n21888 , n21889 );
not ( n21891 , n21757 );
nand ( n21892 , n21891 , n21711 , n21745 );
nand ( n21893 , n21891 , n21710 , n21746 );
nand ( n21894 , n21757 , n21711 , n21746 );
nand ( n21895 , n21757 , n21710 , n21745 );
nand ( n21896 , n21892 , n21893 , n21894 , n21895 );
not ( n21897 , n21896 );
not ( n21898 , n21199 );
not ( n21899 , n21873 );
or ( n21900 , n21898 , n21899 );
and ( n21901 , n21165 , n20952 );
not ( n21902 , n21165 );
and ( n21903 , n21902 , n20946 );
nor ( n21904 , n21901 , n21903 );
nand ( n21905 , n21904 , n21162 );
nand ( n21906 , n21900 , n21905 );
not ( n21907 , n21906 );
not ( n21908 , n20693 );
xor ( n21909 , n20170 , n20180 );
xor ( n21910 , n21909 , n20190 );
not ( n21911 , n21910 );
not ( n21912 , n21911 );
not ( n21913 , n21912 );
or ( n21914 , n21908 , n21913 );
not ( n21915 , n20190 );
nand ( n21916 , n20187 , n20189 );
nand ( n21917 , n21915 , n21916 );
not ( n21918 , n21917 );
not ( n21919 , n21918 );
or ( n21920 , n20710 , n21919 );
nand ( n21921 , n21914 , n21920 );
not ( n21922 , n20763 );
and ( n21923 , n20730 , n21717 );
not ( n21924 , n20730 );
and ( n21925 , n21924 , n21718 );
nor ( n21926 , n21923 , n21925 );
not ( n21927 , n21926 );
or ( n21928 , n21922 , n21927 );
and ( n21929 , n20760 , n21622 );
not ( n21930 , n20760 );
and ( n21931 , n21930 , n21713 );
nor ( n21932 , n21929 , n21931 );
nand ( n21933 , n21932 , n20728 );
nand ( n21934 , n21928 , n21933 );
xor ( n21935 , n21921 , n21934 );
or ( n21936 , n20710 , n20188 );
or ( n21937 , n21919 , n20692 );
nand ( n21938 , n21936 , n21937 );
not ( n21939 , n20728 );
not ( n21940 , n21926 );
or ( n21941 , n21939 , n21940 );
not ( n21942 , n20730 );
not ( n21943 , n21911 );
or ( n21944 , n21942 , n21943 );
buf ( n21945 , n21910 );
nand ( n21946 , n21945 , n20760 );
nand ( n21947 , n21944 , n21946 );
not ( n21948 , n21947 );
or ( n21949 , n21948 , n20764 );
nand ( n21950 , n21941 , n21949 );
xor ( n21951 , n21938 , n21950 );
nor ( n21952 , n20692 , n20188 );
not ( n21953 , n20728 );
not ( n21954 , n21947 );
or ( n21955 , n21953 , n21954 );
not ( n21956 , n20691 );
not ( n21957 , n21919 );
or ( n21958 , n21956 , n21957 );
nand ( n21959 , n21918 , n20760 );
nand ( n21960 , n21958 , n21959 );
nand ( n21961 , n21960 , n20763 );
nand ( n21962 , n21955 , n21961 );
xor ( n21963 , n21952 , n21962 );
not ( n21964 , n20188 );
and ( n21965 , n20723 , n21964 );
nor ( n21966 , n21965 , n20760 );
or ( n21967 , n20723 , n21964 );
nand ( n21968 , n21967 , n20609 );
and ( n21969 , n21966 , n21968 );
not ( n21970 , n20728 );
not ( n21971 , n21960 );
or ( n21972 , n21970 , n21971 );
or ( n21973 , n20691 , n20188 );
or ( n21974 , n20760 , n21964 );
nand ( n21975 , n21973 , n21974 );
nand ( n21976 , n20763 , n21975 );
nand ( n21977 , n21972 , n21976 );
and ( n21978 , n21969 , n21977 );
and ( n21979 , n21963 , n21978 );
and ( n21980 , n21952 , n21962 );
or ( n21981 , n21979 , n21980 );
and ( n21982 , n21951 , n21981 );
and ( n21983 , n21938 , n21950 );
or ( n21984 , n21982 , n21983 );
and ( n21985 , n21935 , n21984 );
and ( n21986 , n21921 , n21934 );
or ( n21987 , n21985 , n21986 );
or ( n21988 , n21911 , n20710 );
or ( n21989 , n21718 , n20692 );
nand ( n21990 , n21988 , n21989 );
not ( n21991 , n20728 );
not ( n21992 , n21728 );
or ( n21993 , n21991 , n21992 );
not ( n21994 , n21932 );
or ( n21995 , n21994 , n20764 );
nand ( n21996 , n21993 , n21995 );
xor ( n21997 , n21990 , n21996 );
not ( n21998 , n20647 );
not ( n21999 , n21740 );
or ( n22000 , n21998 , n21999 );
and ( n22001 , n21255 , n20609 );
not ( n22002 , n21255 );
and ( n22003 , n22002 , n20644 );
nor ( n22004 , n22001 , n22003 );
nand ( n22005 , n22004 , n20602 );
nand ( n22006 , n22000 , n22005 );
xor ( n22007 , n21997 , n22006 );
xor ( n22008 , n21987 , n22007 );
not ( n22009 , n20933 );
not ( n22010 , n20935 );
not ( n22011 , n20702 );
or ( n22012 , n22010 , n22011 );
nand ( n22013 , n20703 , n20953 );
nand ( n22014 , n22012 , n22013 );
not ( n22015 , n22014 );
or ( n22016 , n22009 , n22015 );
not ( n22017 , n20935 );
not ( n22018 , n20709 );
or ( n22019 , n22017 , n22018 );
nand ( n22020 , n21047 , n20953 );
nand ( n22021 , n22019 , n22020 );
nand ( n22022 , n22021 , n20979 );
nand ( n22023 , n22016 , n22022 );
and ( n22024 , n22008 , n22023 );
and ( n22025 , n21987 , n22007 );
or ( n22026 , n22024 , n22025 );
not ( n22027 , n21020 );
not ( n22028 , n20983 );
not ( n22029 , n20793 );
or ( n22030 , n22028 , n22029 );
or ( n22031 , n20793 , n20983 );
nand ( n22032 , n22030 , n22031 );
not ( n22033 , n22032 );
or ( n22034 , n22027 , n22033 );
and ( n22035 , n20983 , n20741 );
not ( n22036 , n20983 );
and ( n22037 , n22036 , n20742 );
nor ( n22038 , n22035 , n22037 );
nand ( n22039 , n22038 , n21003 );
nand ( n22040 , n22034 , n22039 );
xor ( n22041 , n22026 , n22040 );
not ( n22042 , n20860 );
and ( n22043 , n20863 , n20620 );
not ( n22044 , n20863 );
and ( n22045 , n22044 , n20623 );
nor ( n22046 , n22043 , n22045 );
not ( n22047 , n22046 );
or ( n22048 , n22042 , n22047 );
not ( n22049 , n20863 );
not ( n22050 , n20641 );
or ( n22051 , n22049 , n22050 );
nand ( n22052 , n20640 , n20862 );
nand ( n22053 , n22051 , n22052 );
nand ( n22054 , n22053 , n20905 );
nand ( n22055 , n22048 , n22054 );
and ( n22056 , n22041 , n22055 );
and ( n22057 , n22026 , n22040 );
or ( n22058 , n22056 , n22057 );
not ( n22059 , n22058 );
nand ( n22060 , n21907 , n22059 );
not ( n22061 , n22060 );
or ( n22062 , n21897 , n22061 );
and ( n22063 , n21906 , n22058 );
not ( n22064 , n22063 );
nand ( n22065 , n22062 , n22064 );
not ( n22066 , n22065 );
xor ( n22067 , n21708 , n21762 );
xor ( n22068 , n22067 , n21770 );
not ( n22069 , n22068 );
not ( n22070 , n21020 );
not ( n22071 , n21706 );
or ( n22072 , n22070 , n22071 );
nand ( n22073 , n22032 , n21003 );
nand ( n22074 , n22072 , n22073 );
xor ( n22075 , n21990 , n21996 );
and ( n22076 , n22075 , n22006 );
and ( n22077 , n21990 , n21996 );
or ( n22078 , n22076 , n22077 );
xor ( n22079 , n21720 , n21731 );
xor ( n22080 , n22079 , n21742 );
xor ( n22081 , n22078 , n22080 );
not ( n22082 , n20979 );
not ( n22083 , n22014 );
or ( n22084 , n22082 , n22083 );
nand ( n22085 , n21753 , n20933 );
nand ( n22086 , n22084 , n22085 );
and ( n22087 , n22081 , n22086 );
and ( n22088 , n22078 , n22080 );
or ( n22089 , n22087 , n22088 );
xor ( n22090 , n22074 , n22089 );
not ( n22091 , n20905 );
not ( n22092 , n21768 );
or ( n22093 , n22091 , n22092 );
nand ( n22094 , n22053 , n20860 );
nand ( n22095 , n22093 , n22094 );
and ( n22096 , n22090 , n22095 );
and ( n22097 , n22074 , n22089 );
or ( n22098 , n22096 , n22097 );
not ( n22099 , n22098 );
nand ( n22100 , n22069 , n22099 );
not ( n22101 , n22100 );
or ( n22102 , n22066 , n22101 );
nand ( n22103 , n22068 , n22098 );
nand ( n22104 , n22102 , n22103 );
xor ( n22105 , n21890 , n22104 );
xor ( n22106 , n21773 , n21698 );
xor ( n22107 , n22106 , n21696 );
and ( n22108 , n22105 , n22107 );
and ( n22109 , n21890 , n22104 );
or ( n22110 , n22108 , n22109 );
and ( n22111 , n21864 , n22110 );
nor ( n22112 , n21863 , n22111 );
nand ( n22113 , n21851 , n22112 );
and ( n22114 , n21841 , n22113 );
not ( n22115 , n22114 );
not ( n22116 , n21861 );
not ( n22117 , n22110 );
or ( n22118 , n22116 , n22117 );
or ( n22119 , n22110 , n21861 );
nand ( n22120 , n22118 , n22119 );
and ( n22121 , n22120 , n21853 );
not ( n22122 , n22120 );
and ( n22123 , n22122 , n21854 );
nor ( n22124 , n22121 , n22123 );
xor ( n22125 , n21814 , n21816 );
xor ( n22126 , n22125 , n21826 );
nand ( n22127 , n21810 , n18012 );
not ( n22128 , n18029 );
not ( n22129 , n21181 );
or ( n22130 , n22128 , n22129 );
nand ( n22131 , n21178 , n18028 );
nand ( n22132 , n22130 , n22131 );
nand ( n22133 , n22132 , n18025 );
nand ( n22134 , n22127 , n22133 );
xor ( n22135 , n21866 , n21876 );
xor ( n22136 , n22135 , n21887 );
xor ( n22137 , n22134 , n22136 );
xor ( n22138 , n22074 , n22089 );
xor ( n22139 , n22138 , n22095 );
not ( n22140 , n22139 );
not ( n22141 , n21105 );
not ( n22142 , n21885 );
or ( n22143 , n22141 , n22142 );
not ( n22144 , n21111 );
not ( n22145 , n21016 );
or ( n22146 , n22144 , n22145 );
nand ( n22147 , n21013 , n21122 );
nand ( n22148 , n22146 , n22147 );
nand ( n22149 , n22148 , n21148 );
nand ( n22150 , n22143 , n22149 );
not ( n22151 , n22150 );
or ( n22152 , n22140 , n22151 );
or ( n22153 , n22150 , n22139 );
xor ( n22154 , n22078 , n22080 );
xor ( n22155 , n22154 , n22086 );
not ( n22156 , n21199 );
not ( n22157 , n21904 );
or ( n22158 , n22156 , n22157 );
and ( n22159 , n21165 , n20969 );
not ( n22160 , n21165 );
and ( n22161 , n22160 , n20972 );
nor ( n22162 , n22159 , n22161 );
nand ( n22163 , n22162 , n21162 );
nand ( n22164 , n22158 , n22163 );
xor ( n22165 , n22155 , n22164 );
xor ( n22166 , n22026 , n22040 );
xor ( n22167 , n22166 , n22055 );
and ( n22168 , n22165 , n22167 );
and ( n22169 , n22155 , n22164 );
or ( n22170 , n22168 , n22169 );
nand ( n22171 , n22153 , n22170 );
nand ( n22172 , n22152 , n22171 );
and ( n22173 , n22137 , n22172 );
and ( n22174 , n22134 , n22136 );
or ( n22175 , n22173 , n22174 );
xor ( n22176 , n22126 , n22175 );
xor ( n22177 , n21890 , n22104 );
xor ( n22178 , n22177 , n22107 );
and ( n22179 , n22176 , n22178 );
and ( n22180 , n22126 , n22175 );
or ( n22181 , n22179 , n22180 );
nor ( n22182 , n22124 , n22181 );
xor ( n22183 , n22126 , n22175 );
xor ( n22184 , n22183 , n22178 );
not ( n22185 , n18012 );
not ( n22186 , n22132 );
or ( n22187 , n22185 , n22186 );
and ( n22188 , n18029 , n20899 );
not ( n22189 , n18029 );
and ( n22190 , n22189 , n20900 );
nor ( n22191 , n22188 , n22190 );
nand ( n22192 , n22191 , n18025 );
nand ( n22193 , n22187 , n22192 );
not ( n22194 , n21896 );
and ( n22195 , n22194 , n21906 , n22059 );
not ( n22196 , n22195 );
not ( n22197 , n22194 );
nand ( n22198 , n22197 , n22063 );
nand ( n22199 , n21907 , n21896 , n22059 );
not ( n22200 , n21906 );
nand ( n22201 , n22200 , n22194 , n22058 );
nand ( n22202 , n22196 , n22198 , n22199 , n22201 );
xor ( n22203 , n22193 , n22202 );
not ( n22204 , n20647 );
not ( n22205 , n22004 );
or ( n22206 , n22204 , n22205 );
and ( n22207 , n20609 , n21724 );
not ( n22208 , n20609 );
and ( n22209 , n22208 , n21269 );
nor ( n22210 , n22207 , n22209 );
nand ( n22211 , n22210 , n20602 );
nand ( n22212 , n22206 , n22211 );
xor ( n22213 , n21921 , n21934 );
xor ( n22214 , n22213 , n21984 );
and ( n22215 , n22212 , n22214 );
not ( n22216 , n20933 );
not ( n22217 , n22021 );
or ( n22218 , n22216 , n22217 );
and ( n22219 , n20935 , n21044 );
not ( n22220 , n20935 );
and ( n22221 , n22220 , n21314 );
nor ( n22222 , n22219 , n22221 );
nand ( n22223 , n22222 , n20979 );
nand ( n22224 , n22218 , n22223 );
xor ( n22225 , n21921 , n21934 );
xor ( n22226 , n22225 , n21984 );
and ( n22227 , n22224 , n22226 );
and ( n22228 , n22212 , n22224 );
or ( n22229 , n22215 , n22227 , n22228 );
not ( n22230 , n21020 );
not ( n22231 , n22038 );
or ( n22232 , n22230 , n22231 );
and ( n22233 , n20983 , n20753 );
not ( n22234 , n20983 );
and ( n22235 , n22234 , n20752 );
nor ( n22236 , n22233 , n22235 );
nand ( n22237 , n22236 , n21003 );
nand ( n22238 , n22232 , n22237 );
xor ( n22239 , n22229 , n22238 );
not ( n22240 , n20905 );
not ( n22241 , n22046 );
or ( n22242 , n22240 , n22241 );
and ( n22243 , n20863 , n20794 );
not ( n22244 , n20863 );
not ( n22245 , n20779 );
not ( n22246 , n20782 );
or ( n22247 , n22245 , n22246 );
nand ( n22248 , n22247 , n20786 );
and ( n22249 , n22244 , n22248 );
nor ( n22250 , n22243 , n22249 );
nand ( n22251 , n22250 , n20860 );
nand ( n22252 , n22242 , n22251 );
and ( n22253 , n22239 , n22252 );
and ( n22254 , n22229 , n22238 );
or ( n22255 , n22253 , n22254 );
not ( n22256 , n22255 );
not ( n22257 , n21105 );
not ( n22258 , n22148 );
or ( n22259 , n22257 , n22258 );
not ( n22260 , n21111 );
not ( n22261 , n20995 );
or ( n22262 , n22260 , n22261 );
nand ( n22263 , n21124 , n20992 );
nand ( n22264 , n22262 , n22263 );
nand ( n22265 , n22264 , n21148 );
nand ( n22266 , n22259 , n22265 );
not ( n22267 , n22266 );
or ( n22268 , n22256 , n22267 );
or ( n22269 , n22266 , n22255 );
xor ( n22270 , n21987 , n22007 );
xor ( n22271 , n22270 , n22023 );
xor ( n22272 , n21938 , n21950 );
xor ( n22273 , n22272 , n21981 );
not ( n22274 , n20647 );
not ( n22275 , n22210 );
or ( n22276 , n22274 , n22275 );
nand ( n22277 , n21713 , n20644 );
not ( n22278 , n21621 );
nand ( n22279 , n22278 , n20609 );
nand ( n22280 , n22277 , n22279 );
nand ( n22281 , n22280 , n20602 );
nand ( n22282 , n22276 , n22281 );
xor ( n22283 , n22273 , n22282 );
xor ( n22284 , n21952 , n21962 );
xor ( n22285 , n22284 , n21978 );
not ( n22286 , n20571 );
not ( n22287 , n22280 );
or ( n22288 , n22286 , n22287 );
and ( n22289 , n20609 , n21717 );
not ( n22290 , n20609 );
and ( n22291 , n22290 , n21718 );
nor ( n22292 , n22289 , n22291 );
nand ( n22293 , n22292 , n20602 );
nand ( n22294 , n22288 , n22293 );
xor ( n22295 , n22285 , n22294 );
xor ( n22296 , n21969 , n21977 );
not ( n22297 , n20571 );
not ( n22298 , n22292 );
or ( n22299 , n22297 , n22298 );
not ( n22300 , n20609 );
not ( n22301 , n21945 );
not ( n22302 , n22301 );
or ( n22303 , n22300 , n22302 );
nand ( n22304 , n21912 , n20644 );
nand ( n22305 , n22303 , n22304 );
nand ( n22306 , n22305 , n20602 );
nand ( n22307 , n22299 , n22306 );
xor ( n22308 , n22296 , n22307 );
nor ( n22309 , n20727 , n20188 );
not ( n22310 , n20571 );
not ( n22311 , n22305 );
or ( n22312 , n22310 , n22311 );
not ( n22313 , n20609 );
not ( n22314 , n21918 );
not ( n22315 , n22314 );
or ( n22316 , n22313 , n22315 );
not ( n22317 , n22314 );
nand ( n22318 , n22317 , n20644 );
nand ( n22319 , n22316 , n22318 );
nand ( n22320 , n22319 , n20602 );
nand ( n22321 , n22312 , n22320 );
xor ( n22322 , n22309 , n22321 );
and ( n22323 , n20553 , n21964 );
and ( n22324 , n20554 , n20188 );
nor ( n22325 , n22324 , n20953 );
nor ( n22326 , n22323 , n22325 , n20644 );
not ( n22327 , n20571 );
not ( n22328 , n22319 );
or ( n22329 , n22327 , n22328 );
or ( n22330 , n20609 , n20188 );
or ( n22331 , n20644 , n21964 );
nand ( n22332 , n22330 , n22331 );
nand ( n22333 , n20602 , n22332 );
nand ( n22334 , n22329 , n22333 );
and ( n22335 , n22326 , n22334 );
and ( n22336 , n22322 , n22335 );
and ( n22337 , n22309 , n22321 );
or ( n22338 , n22336 , n22337 );
and ( n22339 , n22308 , n22338 );
and ( n22340 , n22296 , n22307 );
or ( n22341 , n22339 , n22340 );
and ( n22342 , n22295 , n22341 );
and ( n22343 , n22285 , n22294 );
or ( n22344 , n22342 , n22343 );
and ( n22345 , n22283 , n22344 );
and ( n22346 , n22273 , n22282 );
or ( n22347 , n22345 , n22346 );
not ( n22348 , n21020 );
not ( n22349 , n22236 );
or ( n22350 , n22348 , n22349 );
and ( n22351 , n20703 , n20983 );
not ( n22352 , n20703 );
and ( n22353 , n22352 , n21487 );
nor ( n22354 , n22351 , n22353 );
nand ( n22355 , n22354 , n21003 );
nand ( n22356 , n22350 , n22355 );
xor ( n22357 , n22347 , n22356 );
xor ( n22358 , n21921 , n21934 );
xor ( n22359 , n22358 , n21984 );
xor ( n22360 , n22212 , n22224 );
xor ( n22361 , n22359 , n22360 );
and ( n22362 , n22357 , n22361 );
and ( n22363 , n22347 , n22356 );
or ( n22364 , n22362 , n22363 );
xor ( n22365 , n22271 , n22364 );
not ( n22366 , n21199 );
not ( n22367 , n22162 );
or ( n22368 , n22366 , n22367 );
and ( n22369 , n21165 , n21088 );
not ( n22370 , n21165 );
and ( n22371 , n22370 , n20641 );
nor ( n22372 , n22369 , n22371 );
nand ( n22373 , n22372 , n21162 );
nand ( n22374 , n22368 , n22373 );
and ( n22375 , n22365 , n22374 );
and ( n22376 , n22271 , n22364 );
or ( n22377 , n22375 , n22376 );
nand ( n22378 , n22269 , n22377 );
nand ( n22379 , n22268 , n22378 );
and ( n22380 , n22203 , n22379 );
and ( n22381 , n22193 , n22202 );
or ( n22382 , n22380 , n22381 );
xor ( n22383 , n22099 , n22068 );
xnor ( n22384 , n22383 , n22065 );
xor ( n22385 , n22382 , n22384 );
xor ( n22386 , n22134 , n22136 );
xor ( n22387 , n22386 , n22172 );
and ( n22388 , n22385 , n22387 );
and ( n22389 , n22382 , n22384 );
or ( n22390 , n22388 , n22389 );
nor ( n22391 , n22184 , n22390 );
nor ( n22392 , n22182 , n22391 );
not ( n22393 , n22392 );
xor ( n22394 , n22382 , n22384 );
xor ( n22395 , n22394 , n22387 );
xor ( n22396 , n22193 , n22202 );
xor ( n22397 , n22396 , n22379 );
xor ( n22398 , n22139 , n22150 );
xnor ( n22399 , n22398 , n22170 );
not ( n22400 , n22399 );
or ( n22401 , n22397 , n22400 );
not ( n22402 , n18025 );
not ( n22403 , n18029 );
not ( n22404 , n20875 );
or ( n22405 , n22403 , n22404 );
nand ( n22406 , n20878 , n18028 );
nand ( n22407 , n22405 , n22406 );
not ( n22408 , n22407 );
or ( n22409 , n22402 , n22408 );
nand ( n22410 , n22191 , n18012 );
nand ( n22411 , n22409 , n22410 );
not ( n22412 , n22411 );
xor ( n22413 , n22155 , n22164 );
xor ( n22414 , n22413 , n22167 );
not ( n22415 , n22414 );
or ( n22416 , n22412 , n22415 );
or ( n22417 , n22411 , n22414 );
xor ( n22418 , n22229 , n22238 );
xor ( n22419 , n22418 , n22252 );
not ( n22420 , n21105 );
not ( n22421 , n22264 );
or ( n22422 , n22420 , n22421 );
and ( n22423 , n21111 , n20945 );
not ( n22424 , n21111 );
and ( n22425 , n22424 , n20946 );
nor ( n22426 , n22423 , n22425 );
nand ( n22427 , n22426 , n21148 );
nand ( n22428 , n22422 , n22427 );
xor ( n22429 , n22419 , n22428 );
not ( n22430 , n20905 );
not ( n22431 , n22250 );
or ( n22432 , n22430 , n22431 );
and ( n22433 , n20863 , n20741 );
not ( n22434 , n20863 );
and ( n22435 , n22434 , n20742 );
nor ( n22436 , n22433 , n22435 );
nand ( n22437 , n22436 , n20860 );
nand ( n22438 , n22432 , n22437 );
not ( n22439 , n20933 );
not ( n22440 , n22222 );
or ( n22441 , n22439 , n22440 );
and ( n22442 , n20935 , n21312 );
not ( n22443 , n20935 );
and ( n22444 , n22443 , n21257 );
nor ( n22445 , n22442 , n22444 );
not ( n22446 , n22445 );
nand ( n22447 , n22446 , n20979 );
nand ( n22448 , n22441 , n22447 );
xor ( n22449 , n22273 , n22282 );
xor ( n22450 , n22449 , n22344 );
xor ( n22451 , n22448 , n22450 );
not ( n22452 , n21003 );
and ( n22453 , n20983 , n21047 );
not ( n22454 , n20983 );
and ( n22455 , n22454 , n20709 );
nor ( n22456 , n22453 , n22455 );
not ( n22457 , n22456 );
or ( n22458 , n22452 , n22457 );
nand ( n22459 , n21020 , n22354 );
nand ( n22460 , n22458 , n22459 );
and ( n22461 , n22451 , n22460 );
and ( n22462 , n22448 , n22450 );
or ( n22463 , n22461 , n22462 );
xor ( n22464 , n22438 , n22463 );
not ( n22465 , n21199 );
not ( n22466 , n22372 );
or ( n22467 , n22465 , n22466 );
not ( n22468 , n21165 );
not ( n22469 , n20623 );
or ( n22470 , n22468 , n22469 );
nand ( n22471 , n20620 , n21166 );
nand ( n22472 , n22470 , n22471 );
nand ( n22473 , n22472 , n21162 );
nand ( n22474 , n22467 , n22473 );
and ( n22475 , n22464 , n22474 );
and ( n22476 , n22438 , n22463 );
or ( n22477 , n22475 , n22476 );
and ( n22478 , n22429 , n22477 );
and ( n22479 , n22419 , n22428 );
or ( n22480 , n22478 , n22479 );
nand ( n22481 , n22417 , n22480 );
nand ( n22482 , n22416 , n22481 );
nand ( n22483 , n22401 , n22482 );
nand ( n22484 , n22397 , n22400 );
nand ( n22485 , n22483 , n22484 );
xor ( n22486 , n22395 , n22485 );
xor ( n22487 , n22266 , n22255 );
xnor ( n22488 , n22487 , n22377 );
xor ( n22489 , n22347 , n22356 );
xor ( n22490 , n22489 , n22361 );
not ( n22491 , n22490 );
not ( n22492 , n21105 );
not ( n22493 , n22426 );
or ( n22494 , n22492 , n22493 );
and ( n22495 , n20969 , n21111 );
not ( n22496 , n20969 );
and ( n22497 , n22496 , n21122 );
nor ( n22498 , n22495 , n22497 );
nand ( n22499 , n22498 , n21148 );
nand ( n22500 , n22494 , n22499 );
not ( n22501 , n22500 );
or ( n22502 , n22491 , n22501 );
not ( n22503 , n22490 );
not ( n22504 , n22503 );
not ( n22505 , n22500 );
not ( n22506 , n22505 );
or ( n22507 , n22504 , n22506 );
not ( n22508 , n20980 );
not ( n22509 , n20935 );
not ( n22510 , n21724 );
not ( n22511 , n22510 );
or ( n22512 , n22509 , n22511 );
or ( n22513 , n22510 , n20935 );
nand ( n22514 , n22512 , n22513 );
not ( n22515 , n22514 );
or ( n22516 , n22508 , n22515 );
or ( n22517 , n22445 , n20932 );
nand ( n22518 , n22516 , n22517 );
xor ( n22519 , n22285 , n22294 );
xor ( n22520 , n22519 , n22341 );
xor ( n22521 , n22518 , n22520 );
not ( n22522 , n21020 );
not ( n22523 , n22456 );
or ( n22524 , n22522 , n22523 );
and ( n22525 , n20983 , n21314 );
not ( n22526 , n20983 );
and ( n22527 , n22526 , n21044 );
nor ( n22528 , n22525 , n22527 );
not ( n22529 , n22528 );
nand ( n22530 , n22529 , n21003 );
nand ( n22531 , n22524 , n22530 );
and ( n22532 , n22521 , n22531 );
and ( n22533 , n22518 , n22520 );
or ( n22534 , n22532 , n22533 );
not ( n22535 , n20905 );
not ( n22536 , n22436 );
or ( n22537 , n22535 , n22536 );
and ( n22538 , n20863 , n20753 );
not ( n22539 , n20863 );
and ( n22540 , n22539 , n20752 );
nor ( n22541 , n22538 , n22540 );
nand ( n22542 , n22541 , n20860 );
nand ( n22543 , n22537 , n22542 );
xor ( n22544 , n22534 , n22543 );
xor ( n22545 , n22448 , n22450 );
xor ( n22546 , n22545 , n22460 );
and ( n22547 , n22544 , n22546 );
and ( n22548 , n22534 , n22543 );
or ( n22549 , n22547 , n22548 );
nand ( n22550 , n22507 , n22549 );
nand ( n22551 , n22502 , n22550 );
xor ( n22552 , n22271 , n22364 );
xor ( n22553 , n22552 , n22374 );
xor ( n22554 , n22551 , n22553 );
not ( n22555 , n18025 );
not ( n22556 , n18029 );
not ( n22557 , n21016 );
or ( n22558 , n22556 , n22557 );
nand ( n22559 , n21013 , n18028 );
nand ( n22560 , n22558 , n22559 );
not ( n22561 , n22560 );
or ( n22562 , n22555 , n22561 );
nand ( n22563 , n22407 , n18012 );
nand ( n22564 , n22562 , n22563 );
and ( n22565 , n22554 , n22564 );
and ( n22566 , n22551 , n22553 );
or ( n22567 , n22565 , n22566 );
not ( n22568 , n22567 );
xor ( n22569 , n22488 , n22568 );
xor ( n22570 , n22411 , n22414 );
xnor ( n22571 , n22570 , n22480 );
xor ( n22572 , n22569 , n22571 );
xor ( n22573 , n22419 , n22428 );
xor ( n22574 , n22573 , n22477 );
not ( n22575 , n18012 );
not ( n22576 , n22560 );
or ( n22577 , n22575 , n22576 );
not ( n22578 , n18029 );
not ( n22579 , n20995 );
or ( n22580 , n22578 , n22579 );
nand ( n22581 , n20992 , n18028 );
nand ( n22582 , n22580 , n22581 );
nand ( n22583 , n22582 , n18025 );
nand ( n22584 , n22577 , n22583 );
xor ( n22585 , n22438 , n22463 );
xor ( n22586 , n22585 , n22474 );
xor ( n22587 , n22584 , n22586 );
not ( n22588 , n21199 );
not ( n22589 , n22472 );
or ( n22590 , n22588 , n22589 );
not ( n22591 , n21165 );
not ( n22592 , n20787 );
or ( n22593 , n22591 , n22592 );
nand ( n22594 , n20794 , n21166 );
nand ( n22595 , n22593 , n22594 );
nand ( n22596 , n22595 , n21162 );
nand ( n22597 , n22590 , n22596 );
not ( n22598 , n22597 );
not ( n22599 , n21105 );
not ( n22600 , n22498 );
or ( n22601 , n22599 , n22600 );
and ( n22602 , n21111 , n21088 );
not ( n22603 , n21111 );
and ( n22604 , n22603 , n20641 );
nor ( n22605 , n22602 , n22604 );
nand ( n22606 , n22605 , n21148 );
nand ( n22607 , n22601 , n22606 );
not ( n22608 , n22607 );
or ( n22609 , n22598 , n22608 );
or ( n22610 , n22607 , n22597 );
not ( n22611 , n20905 );
not ( n22612 , n22541 );
or ( n22613 , n22611 , n22612 );
not ( n22614 , n20863 );
not ( n22615 , n20702 );
or ( n22616 , n22614 , n22615 );
nand ( n22617 , n20703 , n20862 );
nand ( n22618 , n22616 , n22617 );
nand ( n22619 , n22618 , n20860 );
nand ( n22620 , n22613 , n22619 );
xor ( n22621 , n22296 , n22307 );
xor ( n22622 , n22621 , n22338 );
not ( n22623 , n22622 );
not ( n22624 , n20933 );
not ( n22625 , n22514 );
or ( n22626 , n22624 , n22625 );
and ( n22627 , n20935 , n21713 );
not ( n22628 , n20935 );
and ( n22629 , n22628 , n22278 );
nor ( n22630 , n22627 , n22629 );
nand ( n22631 , n22630 , n20979 );
nand ( n22632 , n22626 , n22631 );
not ( n22633 , n22632 );
or ( n22634 , n22623 , n22633 );
or ( n22635 , n22632 , n22622 );
xor ( n22636 , n22309 , n22321 );
xor ( n22637 , n22636 , n22335 );
not ( n22638 , n20933 );
not ( n22639 , n22630 );
or ( n22640 , n22638 , n22639 );
and ( n22641 , n20935 , n21717 );
not ( n22642 , n20935 );
and ( n22643 , n22642 , n21718 );
nor ( n22644 , n22641 , n22643 );
nand ( n22645 , n22644 , n20979 );
nand ( n22646 , n22640 , n22645 );
xor ( n22647 , n22637 , n22646 );
xor ( n22648 , n22326 , n22334 );
not ( n22649 , n20933 );
not ( n22650 , n22644 );
or ( n22651 , n22649 , n22650 );
and ( n22652 , n20935 , n21945 );
not ( n22653 , n20935 );
and ( n22654 , n22653 , n22301 );
nor ( n22655 , n22652 , n22654 );
nand ( n22656 , n22655 , n20979 );
nand ( n22657 , n22651 , n22656 );
xor ( n22658 , n22648 , n22657 );
and ( n22659 , n20571 , n21964 );
not ( n22660 , n20933 );
and ( n22661 , n20569 , n21919 );
not ( n22662 , n20569 );
and ( n22663 , n22662 , n21918 );
nor ( n22664 , n22661 , n22663 );
not ( n22665 , n22664 );
or ( n22666 , n22660 , n22665 );
and ( n22667 , n20569 , n21964 );
and ( n22668 , n20566 , n20188 );
nor ( n22669 , n22667 , n22668 );
not ( n22670 , n22669 );
nand ( n22671 , n22670 , n20979 );
nand ( n22672 , n22666 , n22671 );
not ( n22673 , n20915 );
and ( n22674 , n22673 , n21964 );
nor ( n22675 , n22674 , n20953 );
or ( n22676 , n21964 , n22673 );
nand ( n22677 , n22676 , n20983 );
and ( n22678 , n22675 , n22677 );
and ( n22679 , n22672 , n22678 );
xor ( n22680 , n22659 , n22679 );
not ( n22681 , n20933 );
not ( n22682 , n22655 );
or ( n22683 , n22681 , n22682 );
nand ( n22684 , n22664 , n20979 );
nand ( n22685 , n22683 , n22684 );
and ( n22686 , n22680 , n22685 );
or ( n22687 , n22686 , C0 );
and ( n22688 , n22658 , n22687 );
and ( n22689 , n22648 , n22657 );
or ( n22690 , n22688 , n22689 );
and ( n22691 , n22647 , n22690 );
and ( n22692 , n22637 , n22646 );
or ( n22693 , n22691 , n22692 );
nand ( n22694 , n22635 , n22693 );
nand ( n22695 , n22634 , n22694 );
or ( n22696 , n22620 , n22695 );
xor ( n22697 , n22518 , n22520 );
xor ( n22698 , n22697 , n22531 );
and ( n22699 , n22696 , n22698 );
and ( n22700 , n22695 , n22620 );
nor ( n22701 , n22699 , n22700 );
not ( n22702 , n22701 );
nand ( n22703 , n22610 , n22702 );
nand ( n22704 , n22609 , n22703 );
and ( n22705 , n22587 , n22704 );
and ( n22706 , n22584 , n22586 );
or ( n22707 , n22705 , n22706 );
xor ( n22708 , n22574 , n22707 );
xor ( n22709 , n22551 , n22553 );
xor ( n22710 , n22709 , n22564 );
and ( n22711 , n22708 , n22710 );
and ( n22712 , n22574 , n22707 );
nor ( n22713 , n22711 , n22712 );
and ( n22714 , n22572 , n22713 );
xnor ( n22715 , n22482 , n22399 );
not ( n22716 , n22397 );
and ( n22717 , n22715 , n22716 );
not ( n22718 , n22715 );
and ( n22719 , n22718 , n22397 );
nor ( n22720 , n22717 , n22719 );
xor ( n22721 , n22488 , n22568 );
and ( n22722 , n22721 , n22571 );
and ( n22723 , n22488 , n22568 );
or ( n22724 , n22722 , n22723 );
and ( n22725 , n22720 , n22724 );
nor ( n22726 , n22714 , n22725 );
not ( n22727 , n22726 );
xor ( n22728 , n22584 , n22586 );
xor ( n22729 , n22728 , n22704 );
not ( n22730 , n22729 );
xor ( n22731 , n22534 , n22543 );
xor ( n22732 , n22731 , n22546 );
not ( n22733 , n22732 );
not ( n22734 , n22528 );
not ( n22735 , n21333 );
and ( n22736 , n22734 , n22735 );
not ( n22737 , n20983 );
not ( n22738 , n21312 );
or ( n22739 , n22737 , n22738 );
nand ( n22740 , n21257 , n21487 );
nand ( n22741 , n22739 , n22740 );
and ( n22742 , n22741 , n21003 );
nor ( n22743 , n22736 , n22742 );
not ( n22744 , n22743 );
not ( n22745 , n22744 );
xor ( n22746 , n22632 , n22622 );
xnor ( n22747 , n22746 , n22693 );
not ( n22748 , n22747 );
not ( n22749 , n22748 );
or ( n22750 , n22745 , n22749 );
and ( n22751 , n22618 , n20905 );
and ( n22752 , n20863 , n20709 );
not ( n22753 , n20863 );
and ( n22754 , n22753 , n21047 );
or ( n22755 , n22752 , n22754 );
and ( n22756 , n22755 , n20860 );
nor ( n22757 , n22751 , n22756 );
nand ( n22758 , n22750 , n22757 );
nand ( n22759 , n22747 , n22743 );
nand ( n22760 , n22758 , n22759 );
not ( n22761 , n22760 );
and ( n22762 , n21166 , n20741 );
not ( n22763 , n21166 );
and ( n22764 , n22763 , n20742 );
nor ( n22765 , n22762 , n22764 );
not ( n22766 , n22765 );
not ( n22767 , n21162 );
not ( n22768 , n22767 );
and ( n22769 , n22766 , n22768 );
and ( n22770 , n22595 , n21199 );
nor ( n22771 , n22769 , n22770 );
not ( n22772 , n22771 );
or ( n22773 , n22761 , n22772 );
xor ( n22774 , n22695 , n22620 );
xor ( n22775 , n22774 , n22698 );
nand ( n22776 , n22773 , n22775 );
not ( n22777 , n22771 );
not ( n22778 , n22760 );
nand ( n22779 , n22777 , n22778 );
and ( n22780 , n22776 , n22779 );
not ( n22781 , n22780 );
not ( n22782 , n22781 );
or ( n22783 , n22733 , n22782 );
not ( n22784 , n22732 );
not ( n22785 , n22784 );
not ( n22786 , n22780 );
or ( n22787 , n22785 , n22786 );
and ( n22788 , n18029 , n20952 );
not ( n22789 , n18029 );
and ( n22790 , n22789 , n20946 );
nor ( n22791 , n22788 , n22790 );
not ( n22792 , n22791 );
not ( n22793 , n18025 );
or ( n22794 , n22792 , n22793 );
not ( n22795 , n18012 );
not ( n22796 , n22795 );
nand ( n22797 , n22796 , n22582 );
nand ( n22798 , n22794 , n22797 );
nand ( n22799 , n22787 , n22798 );
nand ( n22800 , n22783 , n22799 );
not ( n22801 , n22800 );
and ( n22802 , n22500 , n22503 );
not ( n22803 , n22500 );
and ( n22804 , n22803 , n22490 );
or ( n22805 , n22802 , n22804 );
not ( n22806 , n22549 );
and ( n22807 , n22805 , n22806 );
not ( n22808 , n22805 );
and ( n22809 , n22808 , n22549 );
nor ( n22810 , n22807 , n22809 );
nand ( n22811 , n22801 , n22810 );
not ( n22812 , n22811 );
or ( n22813 , n22730 , n22812 );
not ( n22814 , n22810 );
nand ( n22815 , n22800 , n22814 );
nand ( n22816 , n22813 , n22815 );
xor ( n22817 , n22574 , n22707 );
xor ( n22818 , n22817 , n22710 );
xor ( n22819 , n22816 , n22818 );
not ( n22820 , n20860 );
not ( n22821 , n20862 );
and ( n22822 , n22821 , n21257 );
not ( n22823 , n22821 );
and ( n22824 , n22823 , n21312 );
nor ( n22825 , n22822 , n22824 );
not ( n22826 , n22825 );
or ( n22827 , n22820 , n22826 );
and ( n22828 , n20862 , n21044 );
not ( n22829 , n20862 );
and ( n22830 , n22829 , n21314 );
nor ( n22831 , n22828 , n22830 );
not ( n22832 , n20905 );
or ( n22833 , n22831 , n22832 );
nand ( n22834 , n22827 , n22833 );
xor ( n22835 , n22648 , n22657 );
xor ( n22836 , n22835 , n22687 );
not ( n22837 , n21020 );
and ( n22838 , n20983 , n21268 );
not ( n22839 , n20983 );
and ( n22840 , n22839 , n22510 );
nor ( n22841 , n22838 , n22840 );
not ( n22842 , n22841 );
or ( n22843 , n22837 , n22842 );
and ( n22844 , n20983 , n21713 );
not ( n22845 , n20983 );
and ( n22846 , n22845 , n21622 );
nor ( n22847 , n22844 , n22846 );
nand ( n22848 , n22847 , n21003 );
nand ( n22849 , n22843 , n22848 );
xor ( n22850 , n22836 , n22849 );
xor ( n22851 , n22659 , n22679 );
xor ( n22852 , n22851 , n22685 );
not ( n22853 , n21020 );
not ( n22854 , n22847 );
or ( n22855 , n22853 , n22854 );
and ( n22856 , n20983 , n21717 );
not ( n22857 , n20983 );
and ( n22858 , n22857 , n21718 );
nor ( n22859 , n22856 , n22858 );
nand ( n22860 , n22859 , n21003 );
nand ( n22861 , n22855 , n22860 );
xor ( n22862 , n22852 , n22861 );
xor ( n22863 , n22672 , n22678 );
not ( n22864 , n21020 );
not ( n22865 , n22859 );
or ( n22866 , n22864 , n22865 );
and ( n22867 , n20983 , n21945 );
not ( n22868 , n20983 );
and ( n22869 , n22868 , n21911 );
nor ( n22870 , n22867 , n22869 );
nand ( n22871 , n22870 , n21003 );
nand ( n22872 , n22866 , n22871 );
xor ( n22873 , n22863 , n22872 );
and ( n22874 , n20933 , n21964 );
not ( n22875 , n21020 );
not ( n22876 , n22870 );
or ( n22877 , n22875 , n22876 );
and ( n22878 , n20983 , n22317 );
not ( n22879 , n20983 );
and ( n22880 , n22879 , n22314 );
nor ( n22881 , n22878 , n22880 );
nand ( n22882 , n22881 , n21003 );
nand ( n22883 , n22877 , n22882 );
xor ( n22884 , n22874 , n22883 );
or ( n22885 , n21000 , n21964 );
nand ( n22886 , n22885 , n22821 );
nand ( n22887 , n21000 , n21964 );
and ( n22888 , n22886 , n20983 , n22887 );
not ( n22889 , n21020 );
not ( n22890 , n22881 );
or ( n22891 , n22889 , n22890 );
or ( n22892 , n20983 , n20188 );
or ( n22893 , n21487 , n21964 );
nand ( n22894 , n22892 , n22893 );
nand ( n22895 , n21003 , n22894 );
nand ( n22896 , n22891 , n22895 );
and ( n22897 , n22888 , n22896 );
and ( n22898 , n22884 , n22897 );
and ( n22899 , n22874 , n22883 );
or ( n22900 , n22898 , n22899 );
and ( n22901 , n22873 , n22900 );
and ( n22902 , n22863 , n22872 );
or ( n22903 , n22901 , n22902 );
and ( n22904 , n22862 , n22903 );
and ( n22905 , n22852 , n22861 );
or ( n22906 , n22904 , n22905 );
xor ( n22907 , n22850 , n22906 );
xor ( n22908 , n22834 , n22907 );
not ( n22909 , n21162 );
and ( n22910 , n21165 , n21047 );
not ( n22911 , n21165 );
and ( n22912 , n22911 , n20709 );
nor ( n22913 , n22910 , n22912 );
not ( n22914 , n22913 );
or ( n22915 , n22909 , n22914 );
not ( n22916 , n21165 );
not ( n22917 , n20702 );
or ( n22918 , n22916 , n22917 );
nand ( n22919 , n20703 , n21166 );
nand ( n22920 , n22918 , n22919 );
nand ( n22921 , n22920 , n21199 );
nand ( n22922 , n22915 , n22921 );
and ( n22923 , n22908 , n22922 );
and ( n22924 , n22834 , n22907 );
or ( n22925 , n22923 , n22924 );
not ( n22926 , n21105 );
not ( n22927 , n22248 );
and ( n22928 , n22927 , n21111 );
not ( n22929 , n22927 );
and ( n22930 , n22929 , n21124 );
nor ( n22931 , n22928 , n22930 );
not ( n22932 , n22931 );
or ( n22933 , n22926 , n22932 );
and ( n22934 , n20740 , n21122 );
not ( n22935 , n20740 );
and ( n22936 , n22935 , n21111 );
or ( n22937 , n22934 , n22936 );
nand ( n22938 , n22937 , n21148 );
nand ( n22939 , n22933 , n22938 );
xor ( n22940 , n22925 , n22939 );
and ( n22941 , n18028 , n20641 );
not ( n22942 , n18028 );
and ( n22943 , n22942 , n20640 );
nor ( n22944 , n22941 , n22943 );
not ( n22945 , n22944 );
not ( n22946 , n18012 );
or ( n22947 , n22945 , n22946 );
and ( n22948 , n18029 , n20620 );
not ( n22949 , n18029 );
and ( n22950 , n22949 , n20623 );
nor ( n22951 , n22948 , n22950 );
nand ( n22952 , n22951 , n18025 );
nand ( n22953 , n22947 , n22952 );
and ( n22954 , n22940 , n22953 );
and ( n22955 , n22925 , n22939 );
or ( n22956 , n22954 , n22955 );
xor ( n22957 , n22637 , n22646 );
xor ( n22958 , n22957 , n22690 );
not ( n22959 , n21020 );
not ( n22960 , n22741 );
or ( n22961 , n22959 , n22960 );
nand ( n22962 , n22841 , n21003 );
nand ( n22963 , n22961 , n22962 );
xor ( n22964 , n22958 , n22963 );
not ( n22965 , n20905 );
not ( n22966 , n22755 );
or ( n22967 , n22965 , n22966 );
not ( n22968 , n22831 );
nand ( n22969 , n22968 , n20860 );
nand ( n22970 , n22967 , n22969 );
and ( n22971 , n22964 , n22970 );
and ( n22972 , n22958 , n22963 );
or ( n22973 , n22971 , n22972 );
not ( n22974 , n21199 );
not ( n22975 , n22765 );
not ( n22976 , n22975 );
or ( n22977 , n22974 , n22976 );
and ( n22978 , n21165 , n20753 );
not ( n22979 , n21165 );
and ( n22980 , n22979 , n20752 );
or ( n22981 , n22978 , n22980 );
not ( n22982 , n22981 );
nand ( n22983 , n22982 , n21162 );
nand ( n22984 , n22977 , n22983 );
xor ( n22985 , n22973 , n22984 );
not ( n22986 , n21105 );
not ( n22987 , n21111 );
not ( n22988 , n20623 );
or ( n22989 , n22987 , n22988 );
nand ( n22990 , n20620 , n21124 );
nand ( n22991 , n22989 , n22990 );
not ( n22992 , n22991 );
or ( n22993 , n22986 , n22992 );
nand ( n22994 , n22931 , n21148 );
nand ( n22995 , n22993 , n22994 );
xor ( n22996 , n22985 , n22995 );
xor ( n22997 , n22956 , n22996 );
xor ( n22998 , n22743 , n22748 );
xnor ( n22999 , n22998 , n22757 );
xor ( n23000 , n22836 , n22849 );
and ( n23001 , n23000 , n22906 );
and ( n23002 , n22836 , n22849 );
or ( n23003 , n23001 , n23002 );
not ( n23004 , n22920 );
not ( n23005 , n21162 );
or ( n23006 , n23004 , n23005 );
or ( n23007 , n22981 , n21161 );
nand ( n23008 , n23006 , n23007 );
xor ( n23009 , n23003 , n23008 );
xor ( n23010 , n22958 , n22963 );
xor ( n23011 , n23010 , n22970 );
and ( n23012 , n23009 , n23011 );
and ( n23013 , n23003 , n23008 );
or ( n23014 , n23012 , n23013 );
xor ( n23015 , n22999 , n23014 );
xor ( n23016 , n18029 , n20959 );
xor ( n23017 , n23016 , n20966 );
not ( n23018 , n23017 );
not ( n23019 , n18012 );
or ( n23020 , n23018 , n23019 );
nand ( n23021 , n22944 , n18025 );
nand ( n23022 , n23020 , n23021 );
not ( n23023 , n23022 );
and ( n23024 , n23015 , n23023 );
not ( n23025 , n23015 );
and ( n23026 , n23025 , n23022 );
nor ( n23027 , n23024 , n23026 );
and ( n23028 , n22997 , n23027 );
and ( n23029 , n22956 , n22996 );
or ( n23030 , n23028 , n23029 );
not ( n23031 , n23030 );
xor ( n23032 , n22777 , n22778 );
xnor ( n23033 , n23032 , n22775 );
not ( n23034 , n22999 );
not ( n23035 , n23023 );
or ( n23036 , n23034 , n23035 );
nand ( n23037 , n23036 , n23014 );
not ( n23038 , n22999 );
nand ( n23039 , n23038 , n23022 );
and ( n23040 , n23037 , n23039 );
xor ( n23041 , n23033 , n23040 );
not ( n23042 , n21105 );
not ( n23043 , n22605 );
or ( n23044 , n23042 , n23043 );
nand ( n23045 , n22991 , n21148 );
nand ( n23046 , n23044 , n23045 );
not ( n23047 , n18012 );
not ( n23048 , n22791 );
or ( n23049 , n23047 , n23048 );
nand ( n23050 , n23017 , n18025 );
nand ( n23051 , n23049 , n23050 );
xor ( n23052 , n23046 , n23051 );
xor ( n23053 , n22973 , n22984 );
and ( n23054 , n23053 , n22995 );
and ( n23055 , n22973 , n22984 );
or ( n23056 , n23054 , n23055 );
xnor ( n23057 , n23052 , n23056 );
xor ( n23058 , n23041 , n23057 );
nand ( n23059 , n23031 , n23058 );
not ( n23060 , n23059 );
xor ( n23061 , n23003 , n23008 );
xor ( n23062 , n23061 , n23011 );
not ( n23063 , n23062 );
xor ( n23064 , n22925 , n22939 );
xor ( n23065 , n23064 , n22953 );
not ( n23066 , n23065 );
or ( n23067 , n23063 , n23066 );
not ( n23068 , n23062 );
not ( n23069 , n23068 );
not ( n23070 , n23065 );
not ( n23071 , n23070 );
or ( n23072 , n23069 , n23071 );
not ( n23073 , n21105 );
not ( n23074 , n22937 );
or ( n23075 , n23073 , n23074 );
not ( n23076 , n21111 );
not ( n23077 , n20752 );
or ( n23078 , n23076 , n23077 );
nand ( n23079 , n20751 , n21122 );
nand ( n23080 , n23078 , n23079 );
nand ( n23081 , n23080 , n21148 );
nand ( n23082 , n23075 , n23081 );
not ( n23083 , n20905 );
not ( n23084 , n22825 );
or ( n23085 , n23083 , n23084 );
and ( n23086 , n22821 , n21268 );
not ( n23087 , n22821 );
and ( n23088 , n23087 , n21269 );
nor ( n23089 , n23086 , n23088 );
nand ( n23090 , n23089 , n20860 );
nand ( n23091 , n23085 , n23090 );
xor ( n23092 , n22852 , n22861 );
xor ( n23093 , n23092 , n22903 );
xor ( n23094 , n23091 , n23093 );
not ( n23095 , n21199 );
not ( n23096 , n22913 );
or ( n23097 , n23095 , n23096 );
and ( n23098 , n21165 , n21044 );
not ( n23099 , n21165 );
and ( n23100 , n23099 , n21314 );
nor ( n23101 , n23098 , n23100 );
nand ( n23102 , n23101 , n21162 );
nand ( n23103 , n23097 , n23102 );
and ( n23104 , n23094 , n23103 );
and ( n23105 , n23091 , n23093 );
or ( n23106 , n23104 , n23105 );
or ( n23107 , n23082 , n23106 );
not ( n23108 , n23107 );
xor ( n23109 , n22863 , n22872 );
xor ( n23110 , n23109 , n22900 );
not ( n23111 , n20905 );
not ( n23112 , n23089 );
or ( n23113 , n23111 , n23112 );
xor ( n23114 , n22821 , n21713 );
nand ( n23115 , n23114 , n20860 );
nand ( n23116 , n23113 , n23115 );
xor ( n23117 , n23110 , n23116 );
xor ( n23118 , n22874 , n22883 );
xor ( n23119 , n23118 , n22897 );
not ( n23120 , n20905 );
not ( n23121 , n23114 );
or ( n23122 , n23120 , n23121 );
not ( n23123 , n22821 );
not ( n23124 , n21718 );
or ( n23125 , n23123 , n23124 );
nand ( n23126 , n21717 , n20862 );
nand ( n23127 , n23125 , n23126 );
nand ( n23128 , n23127 , n20860 );
nand ( n23129 , n23122 , n23128 );
xor ( n23130 , n23119 , n23129 );
xor ( n23131 , n22888 , n22896 );
not ( n23132 , n20905 );
not ( n23133 , n23127 );
or ( n23134 , n23132 , n23133 );
and ( n23135 , n21910 , n20862 );
not ( n23136 , n21910 );
and ( n23137 , n23136 , n22821 );
or ( n23138 , n23135 , n23137 );
nand ( n23139 , n23138 , n20859 );
nand ( n23140 , n23134 , n23139 );
xor ( n23141 , n23131 , n23140 );
not ( n23142 , n20905 );
not ( n23143 , n23138 );
or ( n23144 , n23142 , n23143 );
not ( n23145 , n20862 );
not ( n23146 , n23145 );
not ( n23147 , n21919 );
or ( n23148 , n23146 , n23147 );
nand ( n23149 , n21918 , n20862 );
nand ( n23150 , n23148 , n23149 );
nand ( n23151 , n23150 , n20859 );
nand ( n23152 , n23144 , n23151 );
nand ( n23153 , n21019 , n21964 );
not ( n23154 , n23153 );
or ( n23155 , n23152 , n23154 );
not ( n23156 , n20858 );
not ( n23157 , n23150 );
or ( n23158 , n23156 , n23157 );
or ( n23159 , n23145 , n20188 );
or ( n23160 , n20862 , n21964 );
nand ( n23161 , n23159 , n23160 );
nand ( n23162 , n20859 , n23161 );
nand ( n23163 , n23158 , n23162 );
or ( n23164 , n20835 , n21964 );
nand ( n23165 , n23164 , n21165 );
nand ( n23166 , n20835 , n21964 );
and ( n23167 , n23165 , n22821 , n23166 );
nand ( n23168 , n23155 , n23163 , n23167 );
nand ( n23169 , n23152 , n23154 );
nand ( n23170 , n23168 , n23169 );
and ( n23171 , n23141 , n23170 );
and ( n23172 , n23131 , n23140 );
or ( n23173 , n23171 , n23172 );
and ( n23174 , n23130 , n23173 );
and ( n23175 , n23119 , n23129 );
or ( n23176 , n23174 , n23175 );
and ( n23177 , n23117 , n23176 );
and ( n23178 , n23110 , n23116 );
or ( n23179 , n23177 , n23178 );
not ( n23180 , n23179 );
not ( n23181 , n21105 );
not ( n23182 , n23080 );
or ( n23183 , n23181 , n23182 );
and ( n23184 , n20701 , n21111 );
not ( n23185 , n20701 );
and ( n23186 , n23185 , n21122 );
or ( n23187 , n23184 , n23186 );
nand ( n23188 , n23187 , n21148 );
nand ( n23189 , n23183 , n23188 );
not ( n23190 , n23189 );
nand ( n23191 , n23180 , n23190 );
not ( n23192 , n23191 );
xor ( n23193 , n23091 , n23093 );
xor ( n23194 , n23193 , n23103 );
not ( n23195 , n23194 );
or ( n23196 , n23192 , n23195 );
nand ( n23197 , n23189 , n23179 );
nand ( n23198 , n23196 , n23197 );
not ( n23199 , n23198 );
or ( n23200 , n23108 , n23199 );
nand ( n23201 , n23082 , n23106 );
nand ( n23202 , n23200 , n23201 );
nand ( n23203 , n23072 , n23202 );
nand ( n23204 , n23067 , n23203 );
xor ( n23205 , n22956 , n22996 );
xor ( n23206 , n23205 , n23027 );
xor ( n23207 , n23204 , n23206 );
xor ( n23208 , n22834 , n22907 );
xor ( n23209 , n23208 , n22922 );
not ( n23210 , n18012 );
not ( n23211 , n22951 );
or ( n23212 , n23210 , n23211 );
not ( n23213 , n22248 );
not ( n23214 , n18029 );
or ( n23215 , n23213 , n23214 );
nand ( n23216 , n22927 , n18028 );
nand ( n23217 , n23215 , n23216 );
nand ( n23218 , n23217 , n18025 );
nand ( n23219 , n23212 , n23218 );
xor ( n23220 , n23209 , n23219 );
not ( n23221 , n23198 );
not ( n23222 , n23106 );
not ( n23223 , n23082 );
or ( n23224 , n23222 , n23223 );
or ( n23225 , n23082 , n23106 );
nand ( n23226 , n23224 , n23225 );
not ( n23227 , n23226 );
or ( n23228 , n23221 , n23227 );
or ( n23229 , n23226 , n23198 );
nand ( n23230 , n23228 , n23229 );
and ( n23231 , n23220 , n23230 );
and ( n23232 , n23209 , n23219 );
or ( n23233 , n23231 , n23232 );
xor ( n23234 , n23202 , n23068 );
xnor ( n23235 , n23234 , n23065 );
xor ( n23236 , n23233 , n23235 );
not ( n23237 , n21199 );
nand ( n23238 , n22510 , n21165 );
nand ( n23239 , n21724 , n21166 );
nand ( n23240 , n23238 , n23239 );
not ( n23241 , n23240 );
or ( n23242 , n23237 , n23241 );
or ( n23243 , n21165 , n21622 );
nand ( n23244 , n21620 , n21165 );
nand ( n23245 , n23243 , n23244 );
nand ( n23246 , n23245 , n21162 );
nand ( n23247 , n23242 , n23246 );
xor ( n23248 , n23131 , n23140 );
xor ( n23249 , n23248 , n23170 );
xor ( n23250 , n23247 , n23249 );
and ( n23251 , n23152 , n23153 );
not ( n23252 , n23152 );
and ( n23253 , n23252 , n23154 );
or ( n23254 , n23251 , n23253 );
and ( n23255 , n23167 , n23163 );
xnor ( n23256 , n23254 , n23255 );
not ( n23257 , n23256 );
not ( n23258 , n21165 );
nand ( n23259 , n23258 , n21199 );
or ( n23260 , n21622 , n23259 );
not ( n23261 , n23244 );
nand ( n23262 , n23261 , n21199 );
not ( n23263 , n21165 );
not ( n23264 , n21718 );
or ( n23265 , n23263 , n23264 );
nand ( n23266 , n21717 , n20856 );
nand ( n23267 , n23265 , n23266 );
nand ( n23268 , n23267 , n21162 );
nand ( n23269 , n23260 , n23262 , n23268 );
not ( n23270 , n23269 );
not ( n23271 , n23270 );
or ( n23272 , n23257 , n23271 );
xor ( n23273 , n23167 , n23163 );
not ( n23274 , n21199 );
not ( n23275 , n23267 );
or ( n23276 , n23274 , n23275 );
and ( n23277 , n21910 , n20856 );
not ( n23278 , n21910 );
and ( n23279 , n23278 , n21165 );
or ( n23280 , n23277 , n23279 );
nand ( n23281 , n23280 , n21162 );
nand ( n23282 , n23276 , n23281 );
xor ( n23283 , n23273 , n23282 );
nand ( n23284 , n20858 , n21964 );
not ( n23285 , n23284 );
not ( n23286 , n21199 );
not ( n23287 , n23280 );
or ( n23288 , n23286 , n23287 );
not ( n23289 , n21165 );
not ( n23290 , n22314 );
or ( n23291 , n23289 , n23290 );
nand ( n23292 , n21918 , n20856 );
nand ( n23293 , n23291 , n23292 );
nand ( n23294 , n23293 , n21162 );
nand ( n23295 , n23288 , n23294 );
not ( n23296 , n23295 );
not ( n23297 , n23296 );
or ( n23298 , n23285 , n23297 );
not ( n23299 , n21199 );
not ( n23300 , n23293 );
or ( n23301 , n23299 , n23300 );
or ( n23302 , n21165 , n20188 );
or ( n23303 , n20856 , n21964 );
nand ( n23304 , n23302 , n23303 );
nand ( n23305 , n21162 , n23304 );
nand ( n23306 , n23301 , n23305 );
or ( n23307 , n21153 , n21964 );
nand ( n23308 , n23307 , n21111 );
nand ( n23309 , n21153 , n21964 );
and ( n23310 , n21165 , n23308 , n23309 );
and ( n23311 , n23306 , n23310 );
nand ( n23312 , n23298 , n23311 );
not ( n23313 , n23284 );
nand ( n23314 , n23295 , n23313 );
nand ( n23315 , n23312 , n23314 );
and ( n23316 , n23283 , n23315 );
and ( n23317 , n23273 , n23282 );
or ( n23318 , n23316 , n23317 );
nand ( n23319 , n23272 , n23318 );
not ( n23320 , n23256 );
nand ( n23321 , n23320 , n23269 );
nand ( n23322 , n23319 , n23321 );
and ( n23323 , n23250 , n23322 );
and ( n23324 , n23247 , n23249 );
or ( n23325 , n23323 , n23324 );
not ( n23326 , n18012 );
not ( n23327 , n18029 );
not ( n23328 , n20752 );
or ( n23329 , n23327 , n23328 );
nand ( n23330 , n20751 , n18028 );
nand ( n23331 , n23329 , n23330 );
not ( n23332 , n23331 );
or ( n23333 , n23326 , n23332 );
not ( n23334 , n18029 );
not ( n23335 , n20701 );
or ( n23336 , n23334 , n23335 );
or ( n23337 , n20701 , n18029 );
nand ( n23338 , n23336 , n23337 );
nand ( n23339 , n23338 , n18025 );
nand ( n23340 , n23333 , n23339 );
xor ( n23341 , n23325 , n23340 );
not ( n23342 , n21105 );
not ( n23343 , n21111 );
not ( n23344 , n20709 );
or ( n23345 , n23343 , n23344 );
nand ( n23346 , n20708 , n21122 );
nand ( n23347 , n23345 , n23346 );
not ( n23348 , n23347 );
or ( n23349 , n23342 , n23348 );
not ( n23350 , n21111 );
not ( n23351 , n21314 );
or ( n23352 , n23350 , n23351 );
nand ( n23353 , n21044 , n21122 );
nand ( n23354 , n23352 , n23353 );
nand ( n23355 , n23354 , n21148 );
nand ( n23356 , n23349 , n23355 );
not ( n23357 , n21165 );
not ( n23358 , n21312 );
or ( n23359 , n23357 , n23358 );
nand ( n23360 , n21257 , n21166 );
nand ( n23361 , n23359 , n23360 );
and ( n23362 , n23361 , n21199 );
and ( n23363 , n23240 , n21162 );
nor ( n23364 , n23362 , n23363 );
not ( n23365 , n23364 );
xor ( n23366 , n23119 , n23129 );
xor ( n23367 , n23366 , n23173 );
not ( n23368 , n23367 );
or ( n23369 , n23365 , n23368 );
or ( n23370 , n23367 , n23364 );
nand ( n23371 , n23369 , n23370 );
xor ( n23372 , n23356 , n23371 );
and ( n23373 , n23341 , n23372 );
and ( n23374 , n23325 , n23340 );
or ( n23375 , n23373 , n23374 );
not ( n23376 , n23375 );
not ( n23377 , n18012 );
xor ( n23378 , n18029 , n20740 );
not ( n23379 , n23378 );
or ( n23380 , n23377 , n23379 );
nand ( n23381 , n23331 , n18025 );
nand ( n23382 , n23380 , n23381 );
not ( n23383 , n23356 );
not ( n23384 , n23383 );
not ( n23385 , n23364 );
and ( n23386 , n23384 , n23385 );
nand ( n23387 , n23383 , n23364 );
and ( n23388 , n23387 , n23367 );
nor ( n23389 , n23386 , n23388 );
xor ( n23390 , n23382 , n23389 );
not ( n23391 , n23390 );
and ( n23392 , n23376 , n23391 );
and ( n23393 , n23375 , n23390 );
nor ( n23394 , n23392 , n23393 );
not ( n23395 , n23394 );
not ( n23396 , n21105 );
not ( n23397 , n23187 );
or ( n23398 , n23396 , n23397 );
nand ( n23399 , n23347 , n21148 );
nand ( n23400 , n23398 , n23399 );
not ( n23401 , n23400 );
xor ( n23402 , n23110 , n23116 );
xor ( n23403 , n23402 , n23176 );
not ( n23404 , n21199 );
not ( n23405 , n23101 );
or ( n23406 , n23404 , n23405 );
nand ( n23407 , n23361 , n21162 );
nand ( n23408 , n23406 , n23407 );
xnor ( n23409 , n23403 , n23408 );
not ( n23410 , n23409 );
or ( n23411 , n23401 , n23410 );
or ( n23412 , n23409 , n23400 );
nand ( n23413 , n23411 , n23412 );
nand ( n23414 , n23395 , n23413 );
not ( n23415 , n21105 );
not ( n23416 , n23354 );
or ( n23417 , n23415 , n23416 );
xor ( n23418 , n21111 , n21255 );
nand ( n23419 , n23418 , n21148 );
nand ( n23420 , n23417 , n23419 );
xor ( n23421 , n23247 , n23249 );
xor ( n23422 , n23421 , n23322 );
xor ( n23423 , n23420 , n23422 );
not ( n23424 , n18025 );
xor ( n23425 , n18023 , n20708 );
not ( n23426 , n23425 );
or ( n23427 , n23424 , n23426 );
nand ( n23428 , n23338 , n18012 );
nand ( n23429 , n23427 , n23428 );
and ( n23430 , n23423 , n23429 );
and ( n23431 , n23420 , n23422 );
or ( n23432 , n23430 , n23431 );
xor ( n23433 , n23325 , n23340 );
xor ( n23434 , n23433 , n23372 );
xor ( n23435 , n23432 , n23434 );
not ( n23436 , n18012 );
not ( n23437 , n23425 );
or ( n23438 , n23436 , n23437 );
not ( n23439 , n18029 );
not ( n23440 , n21314 );
or ( n23441 , n23439 , n23440 );
nand ( n23442 , n21044 , n18028 );
nand ( n23443 , n23441 , n23442 );
nand ( n23444 , n23443 , n18025 );
nand ( n23445 , n23438 , n23444 );
not ( n23446 , n23445 );
not ( n23447 , n23446 );
not ( n23448 , n21105 );
not ( n23449 , n23418 );
or ( n23450 , n23448 , n23449 );
not ( n23451 , n21122 );
not ( n23452 , n21724 );
or ( n23453 , n23451 , n23452 );
or ( n23454 , n21122 , n21724 );
nand ( n23455 , n23453 , n23454 );
nand ( n23456 , n23455 , n21147 );
nand ( n23457 , n23450 , n23456 );
not ( n23458 , n23457 );
not ( n23459 , n23458 );
or ( n23460 , n23447 , n23459 );
buf ( n23461 , n23256 );
and ( n23462 , n23270 , n23461 );
not ( n23463 , n23270 );
not ( n23464 , n23256 );
and ( n23465 , n23463 , n23464 );
nor ( n23466 , n23462 , n23465 );
not ( n23467 , n23318 );
and ( n23468 , n23466 , n23467 );
not ( n23469 , n23466 );
and ( n23470 , n23469 , n23318 );
nor ( n23471 , n23468 , n23470 );
not ( n23472 , n23471 );
nand ( n23473 , n23460 , n23472 );
nand ( n23474 , n23445 , n23457 );
nand ( n23475 , n23473 , n23474 );
xor ( n23476 , n23420 , n23422 );
xor ( n23477 , n23476 , n23429 );
xor ( n23478 , n23475 , n23477 );
xor ( n23479 , n23273 , n23282 );
xor ( n23480 , n23479 , n23315 );
not ( n23481 , n21105 );
not ( n23482 , n23455 );
or ( n23483 , n23481 , n23482 );
not ( n23484 , n21111 );
not ( n23485 , n22278 );
or ( n23486 , n23484 , n23485 );
not ( n23487 , n21110 );
nand ( n23488 , n23487 , n21619 );
nand ( n23489 , n23486 , n23488 );
nand ( n23490 , n23489 , n21147 );
nand ( n23491 , n23483 , n23490 );
or ( n23492 , n23480 , n23491 );
not ( n23493 , n23492 );
not ( n23494 , n23313 );
not ( n23495 , n23296 );
or ( n23496 , n23494 , n23495 );
nand ( n23497 , n23295 , n23284 );
nand ( n23498 , n23496 , n23497 );
xnor ( n23499 , n23498 , n23311 );
not ( n23500 , n23499 );
not ( n23501 , n23500 );
not ( n23502 , n21105 );
not ( n23503 , n23489 );
or ( n23504 , n23502 , n23503 );
and ( n23505 , n21111 , n21717 );
not ( n23506 , n21111 );
and ( n23507 , n23506 , n21718 );
nor ( n23508 , n23505 , n23507 );
nand ( n23509 , n23508 , n21147 );
nand ( n23510 , n23504 , n23509 );
not ( n23511 , n23510 );
or ( n23512 , n23501 , n23511 );
or ( n23513 , n23510 , n23500 );
xor ( n23514 , n23310 , n23306 );
not ( n23515 , n21105 );
not ( n23516 , n23508 );
or ( n23517 , n23515 , n23516 );
and ( n23518 , n21111 , n21945 );
not ( n23519 , n21111 );
and ( n23520 , n23519 , n21911 );
nor ( n23521 , n23518 , n23520 );
nand ( n23522 , n23521 , n21147 );
nand ( n23523 , n23517 , n23522 );
xor ( n23524 , n23514 , n23523 );
and ( n23525 , n21199 , n21964 );
not ( n23526 , n21104 );
not ( n23527 , n23521 );
or ( n23528 , n23526 , n23527 );
not ( n23529 , n21111 );
not ( n23530 , n22314 );
or ( n23531 , n23529 , n23530 );
nand ( n23532 , n21918 , n21122 );
nand ( n23533 , n23531 , n23532 );
nand ( n23534 , n23533 , n21147 );
nand ( n23535 , n23528 , n23534 );
xor ( n23536 , n23525 , n23535 );
not ( n23537 , n21104 );
not ( n23538 , n23533 );
or ( n23539 , n23537 , n23538 );
or ( n23540 , n21111 , n20188 );
or ( n23541 , n21122 , n21964 );
nand ( n23542 , n23540 , n23541 );
nand ( n23543 , n21147 , n23542 );
nand ( n23544 , n23539 , n23543 );
not ( n23545 , n23544 );
or ( n23546 , n21964 , n21103 );
nand ( n23547 , n23546 , n18023 );
nand ( n23548 , n21964 , n21103 );
nand ( n23549 , n23547 , n21111 , n23548 );
nor ( n23550 , n23545 , n23549 );
and ( n23551 , n23536 , n23550 );
and ( n23552 , n23525 , n23535 );
or ( n23553 , n23551 , n23552 );
and ( n23554 , n23524 , n23553 );
and ( n23555 , n23514 , n23523 );
or ( n23556 , n23554 , n23555 );
nand ( n23557 , n23513 , n23556 );
nand ( n23558 , n23512 , n23557 );
not ( n23559 , n23558 );
or ( n23560 , n23493 , n23559 );
nand ( n23561 , n23491 , n23480 );
nand ( n23562 , n23560 , n23561 );
not ( n23563 , n23562 );
not ( n23564 , n23472 );
not ( n23565 , n23458 );
or ( n23566 , n23564 , n23565 );
nand ( n23567 , n23471 , n23457 );
nand ( n23568 , n23566 , n23567 );
and ( n23569 , n23568 , n23446 );
not ( n23570 , n23568 );
and ( n23571 , n23570 , n23445 );
nor ( n23572 , n23569 , n23571 );
nand ( n23573 , n23563 , n23572 );
not ( n23574 , n23573 );
not ( n23575 , n23443 );
or ( n23576 , n23575 , n22795 );
and ( n23577 , n21312 , n18029 );
not ( n23578 , n21312 );
and ( n23579 , n23578 , n18028 );
nor ( n23580 , n23577 , n23579 );
or ( n23581 , n23580 , n18024 );
nand ( n23582 , n23576 , n23581 );
not ( n23583 , n23582 );
or ( n23584 , n23480 , n23491 );
nand ( n23585 , n23480 , n23491 );
nand ( n23586 , n23584 , n23585 );
xor ( n23587 , n23586 , n23558 );
nand ( n23588 , n23583 , n23587 );
not ( n23589 , n23588 );
not ( n23590 , n18027 );
not ( n23591 , n21713 );
or ( n23592 , n23590 , n23591 );
nand ( n23593 , n21616 , n21618 , n18023 );
nand ( n23594 , n23592 , n23593 );
not ( n23595 , n23594 );
not ( n23596 , n18025 );
or ( n23597 , n23595 , n23596 );
not ( n23598 , n21724 );
not ( n23599 , n18027 );
and ( n23600 , n23598 , n23599 );
and ( n23601 , n21268 , n18027 );
nor ( n23602 , n23600 , n23601 );
or ( n23603 , n23602 , n22795 );
nand ( n23604 , n23597 , n23603 );
xor ( n23605 , n23514 , n23523 );
xor ( n23606 , n23605 , n23553 );
nor ( n23607 , n23604 , n23606 );
xor ( n23608 , n23525 , n23535 );
xor ( n23609 , n23608 , n23550 );
not ( n23610 , n18012 );
not ( n23611 , n23594 );
or ( n23612 , n23610 , n23611 );
and ( n23613 , n18027 , n21717 );
not ( n23614 , n18027 );
and ( n23615 , n23614 , n21718 );
nor ( n23616 , n23613 , n23615 );
or ( n23617 , n23616 , n18024 );
nand ( n23618 , n23612 , n23617 );
xor ( n23619 , n23609 , n23618 );
not ( n23620 , n23549 );
not ( n23621 , n23544 );
or ( n23622 , n23620 , n23621 );
or ( n23623 , n23544 , n23549 );
nand ( n23624 , n23622 , n23623 );
or ( n23625 , n23616 , n22795 );
and ( n23626 , n18023 , n21911 );
not ( n23627 , n18023 );
and ( n23628 , n23627 , n21945 );
nor ( n23629 , n23626 , n23628 );
or ( n23630 , n23629 , n18024 );
nand ( n23631 , n23625 , n23630 );
xor ( n23632 , n23624 , n23631 );
nor ( n23633 , n21143 , n20188 );
not ( n23634 , n21964 );
not ( n23635 , n18024 );
and ( n23636 , n23634 , n23635 );
not ( n23637 , n18023 );
not ( n23638 , n22314 );
or ( n23639 , n23637 , n23638 );
nand ( n23640 , n21918 , n18027 );
nand ( n23641 , n23639 , n23640 );
and ( n23642 , n23641 , n18012 );
nor ( n23643 , n23636 , n23642 );
nand ( n23644 , n21964 , n18012 );
nand ( n23645 , n23644 , n18023 );
nor ( n23646 , n23643 , n23645 );
xor ( n23647 , n23633 , n23646 );
not ( n23648 , n18025 );
not ( n23649 , n23641 );
or ( n23650 , n23648 , n23649 );
or ( n23651 , n23629 , n22795 );
nand ( n23652 , n23650 , n23651 );
and ( n23653 , n23647 , n23652 );
or ( n23654 , n23653 , C0 );
and ( n23655 , n23632 , n23654 );
and ( n23656 , n23624 , n23631 );
or ( n23657 , n23655 , n23656 );
and ( n23658 , n23619 , n23657 );
and ( n23659 , n23609 , n23618 );
or ( n23660 , n23658 , n23659 );
not ( n23661 , n23660 );
or ( n23662 , n23607 , n23661 );
nand ( n23663 , n23604 , n23606 );
nand ( n23664 , n23662 , n23663 );
not ( n23665 , n23664 );
xor ( n23666 , n23499 , n23510 );
xor ( n23667 , n23666 , n23556 );
not ( n23668 , n23580 );
not ( n23669 , n22795 );
and ( n23670 , n23668 , n23669 );
not ( n23671 , n23602 );
and ( n23672 , n23671 , n18025 );
nor ( n23673 , n23670 , n23672 );
nand ( n23674 , n23667 , n23673 );
not ( n23675 , n23674 );
or ( n23676 , n23665 , n23675 );
or ( n23677 , n23667 , n23673 );
nand ( n23678 , n23676 , n23677 );
not ( n23679 , n23678 );
or ( n23680 , n23589 , n23679 );
not ( n23681 , n23587 );
nand ( n23682 , n23681 , n23582 );
nand ( n23683 , n23680 , n23682 );
not ( n23684 , n23683 );
or ( n23685 , n23574 , n23684 );
not ( n23686 , n23572 );
nand ( n23687 , n23686 , n23562 );
nand ( n23688 , n23685 , n23687 );
and ( n23689 , n23478 , n23688 );
and ( n23690 , n23475 , n23477 );
or ( n23691 , n23689 , n23690 );
and ( n23692 , n23435 , n23691 );
and ( n23693 , n23432 , n23434 );
or ( n23694 , n23692 , n23693 );
not ( n23695 , n23413 );
nand ( n23696 , n23695 , n23394 );
nand ( n23697 , n23694 , n23696 );
nand ( n23698 , n23414 , n23697 );
and ( n23699 , n23179 , n23190 );
not ( n23700 , n23179 );
and ( n23701 , n23700 , n23189 );
or ( n23702 , n23699 , n23701 );
xnor ( n23703 , n23194 , n23702 );
not ( n23704 , n23703 );
or ( n23705 , n23400 , n23408 );
nand ( n23706 , n23705 , n23403 );
nand ( n23707 , n23400 , n23408 );
and ( n23708 , n23706 , n23707 );
and ( n23709 , n23217 , n18012 );
not ( n23710 , n23378 );
nor ( n23711 , n23710 , n18024 );
nor ( n23712 , n23709 , n23711 );
xor ( n23713 , n23708 , n23712 );
not ( n23714 , n23713 );
and ( n23715 , n23704 , n23714 );
and ( n23716 , n23703 , n23713 );
nor ( n23717 , n23715 , n23716 );
not ( n23718 , n23382 );
not ( n23719 , n23718 );
not ( n23720 , n23389 );
and ( n23721 , n23719 , n23720 );
nand ( n23722 , n23718 , n23389 );
and ( n23723 , n23375 , n23722 );
nor ( n23724 , n23721 , n23723 );
and ( n23725 , n23717 , n23724 );
not ( n23726 , n23725 );
and ( n23727 , n23698 , n23726 );
or ( n23728 , n23717 , n23724 );
not ( n23729 , n23728 );
nor ( n23730 , n23727 , n23729 );
xor ( n23731 , n23209 , n23219 );
xor ( n23732 , n23731 , n23230 );
and ( n23733 , n23708 , n23712 );
or ( n23734 , n23703 , n23733 );
or ( n23735 , n23712 , n23708 );
nand ( n23736 , n23734 , n23735 );
buf ( n23737 , n23736 );
nor ( n23738 , n23732 , n23737 );
or ( n23739 , n23730 , n23738 );
nand ( n23740 , n23732 , n23737 );
nand ( n23741 , n23739 , n23740 );
and ( n23742 , n23236 , n23741 );
and ( n23743 , n23233 , n23235 );
or ( n23744 , n23742 , n23743 );
and ( n23745 , n23207 , n23744 );
and ( n23746 , n23204 , n23206 );
or ( n23747 , n23745 , n23746 );
not ( n23748 , n23747 );
or ( n23749 , n23060 , n23748 );
not ( n23750 , n23058 );
nand ( n23751 , n23750 , n23030 );
nand ( n23752 , n23749 , n23751 );
not ( n23753 , n23752 );
not ( n23754 , n22814 );
not ( n23755 , n22801 );
or ( n23756 , n23754 , n23755 );
nand ( n23757 , n22800 , n22810 );
nand ( n23758 , n23756 , n23757 );
not ( n23759 , n22729 );
and ( n23760 , n23758 , n23759 );
not ( n23761 , n23758 );
and ( n23762 , n23761 , n22729 );
nor ( n23763 , n23760 , n23762 );
xor ( n23764 , n22597 , n22701 );
xor ( n23765 , n23764 , n22607 );
not ( n23766 , n23765 );
not ( n23767 , n23046 );
not ( n23768 , n23051 );
or ( n23769 , n23767 , n23768 );
or ( n23770 , n23051 , n23046 );
nand ( n23771 , n23770 , n23056 );
nand ( n23772 , n23769 , n23771 );
not ( n23773 , n23772 );
not ( n23774 , n23773 );
or ( n23775 , n23766 , n23774 );
xor ( n23776 , n22732 , n22780 );
xnor ( n23777 , n23776 , n22798 );
nand ( n23778 , n23775 , n23777 );
not ( n23779 , n23765 );
nand ( n23780 , n23772 , n23779 );
and ( n23781 , n23778 , n23780 );
nand ( n23782 , n23763 , n23781 );
not ( n23783 , n23779 );
not ( n23784 , n23773 );
or ( n23785 , n23783 , n23784 );
nand ( n23786 , n23772 , n23765 );
nand ( n23787 , n23785 , n23786 );
not ( n23788 , n23777 );
and ( n23789 , n23787 , n23788 );
not ( n23790 , n23787 );
buf ( n23791 , n23777 );
and ( n23792 , n23790 , n23791 );
nor ( n23793 , n23789 , n23792 );
xor ( n23794 , n23033 , n23040 );
and ( n23795 , n23794 , n23057 );
and ( n23796 , n23033 , n23040 );
or ( n23797 , n23795 , n23796 );
nand ( n23798 , n23793 , n23797 );
and ( n23799 , n23782 , n23798 );
not ( n23800 , n23799 );
or ( n23801 , n23753 , n23800 );
nor ( n23802 , n23793 , n23797 );
and ( n23803 , n23802 , n23782 );
nor ( n23804 , n23763 , n23781 );
nor ( n23805 , n23803 , n23804 );
nand ( n23806 , n23801 , n23805 );
and ( n23807 , n22819 , n23806 );
and ( n23808 , n22816 , n22818 );
or ( n23809 , n23807 , n23808 );
not ( n23810 , n23809 );
or ( n23811 , n22727 , n23810 );
nand ( n23812 , n22720 , n22724 );
nor ( n23813 , n22572 , n22713 );
and ( n23814 , n23812 , n23813 );
nor ( n23815 , n22720 , n22724 );
nor ( n23816 , n23814 , n23815 );
nand ( n23817 , n23811 , n23816 );
and ( n23818 , n22486 , n23817 );
and ( n23819 , n22395 , n22485 );
or ( n23820 , n23818 , n23819 );
not ( n23821 , n23820 );
or ( n23822 , n22393 , n23821 );
not ( n23823 , n22182 );
and ( n23824 , n22184 , n22390 );
and ( n23825 , n23823 , n23824 );
and ( n23826 , n22181 , n22124 );
nor ( n23827 , n23825 , n23826 );
nand ( n23828 , n23822 , n23827 );
not ( n23829 , n23828 );
or ( n23830 , n22115 , n23829 );
nor ( n23831 , n21851 , n22112 );
and ( n23832 , n21841 , n23831 );
nor ( n23833 , n21797 , n21840 );
nor ( n23834 , n23832 , n23833 );
nand ( n23835 , n23830 , n23834 );
xor ( n23836 , n21792 , n23835 );
not ( n23837 , n18007 );
or ( n23838 , n23836 , n23837 );
nand ( n23839 , n18008 , n23838 );
and ( n23840 , n17228 , n472 );
and ( n23841 , n17247 , n471 );
nor ( n23842 , n23840 , n23841 );
nor ( n23843 , n17306 , n23842 );
buf ( n23844 , n18007 );
not ( n23845 , n23844 );
and ( n23846 , n23843 , n23845 );
and ( n23847 , n23643 , n23645 );
nor ( n23848 , n23847 , n23646 );
and ( n23849 , n23848 , n23844 );
nor ( n23850 , n23846 , n23849 );
or ( n23851 , n17648 , n17680 );
not ( n23852 , n23851 );
not ( n23853 , n23852 );
buf ( n23854 , n17662 );
not ( n23855 , n23854 );
not ( n23856 , n23855 );
not ( n23857 , n17669 );
not ( n23858 , n23857 );
not ( n23859 , n17627 );
or ( n23860 , n23858 , n23859 );
buf ( n23861 , n17674 );
nand ( n23862 , n23860 , n23861 );
not ( n23863 , n23862 );
or ( n23864 , n23856 , n23863 );
buf ( n23865 , n17676 );
nand ( n23866 , n23864 , n23865 );
not ( n23867 , n23866 );
or ( n23868 , n23853 , n23867 );
not ( n23869 , n23851 );
or ( n23870 , n23866 , n23869 );
nand ( n23871 , n23868 , n23870 );
or ( n23872 , n23871 , n18007 );
not ( n23873 , n23826 );
nand ( n23874 , n23873 , n23823 );
not ( n23875 , n22391 );
not ( n23876 , n23875 );
not ( n23877 , n23820 );
or ( n23878 , n23876 , n23877 );
not ( n23879 , n23824 );
nand ( n23880 , n23878 , n23879 );
xor ( n23881 , n23874 , n23880 );
or ( n23882 , n23881 , n23837 );
nand ( n23883 , n23872 , n23882 );
nand ( n23884 , n23855 , n23865 );
and ( n23885 , n23862 , n23884 );
not ( n23886 , n23862 );
not ( n23887 , n23884 );
and ( n23888 , n23886 , n23887 );
nor ( n23889 , n23885 , n23888 );
or ( n23890 , n23889 , n18007 );
nand ( n23891 , n23879 , n23875 );
xor ( n23892 , n23891 , n23820 );
or ( n23893 , n23892 , n23837 );
nand ( n23894 , n23890 , n23893 );
nand ( n23895 , n23857 , n23861 );
not ( n23896 , n23895 );
and ( n23897 , n17627 , n23896 );
not ( n23898 , n17627 );
and ( n23899 , n23898 , n23895 );
or ( n23900 , n23897 , n23899 );
or ( n23901 , n23900 , n18007 );
xor ( n23902 , n22395 , n22485 );
xor ( n23903 , n23902 , n23817 );
not ( n23904 , n23903 );
or ( n23905 , n23904 , n23837 );
nand ( n23906 , n23901 , n23905 );
not ( n23907 , n17600 );
not ( n23908 , n17534 );
not ( n23909 , n16951 );
not ( n23910 , n17357 );
or ( n23911 , n23909 , n23910 );
not ( n23912 , n17605 );
nand ( n23913 , n23911 , n23912 );
not ( n23914 , n23913 );
or ( n23915 , n23908 , n23914 );
nand ( n23916 , n23915 , n17616 );
not ( n23917 , n23916 );
or ( n23918 , n23907 , n23917 );
nand ( n23919 , n23918 , n17624 );
not ( n23920 , n23919 );
not ( n23921 , n17591 );
and ( n23922 , n23921 , n17595 );
not ( n23923 , n23922 );
or ( n23924 , n23920 , n23923 );
or ( n23925 , n23922 , n23919 );
nand ( n23926 , n23924 , n23925 );
or ( n23927 , n23926 , n18007 );
not ( n23928 , n23813 );
nand ( n23929 , n22572 , n22713 );
nand ( n23930 , n23928 , n23929 );
xor ( n23931 , n23930 , n23809 );
or ( n23932 , n23931 , n23837 );
nand ( n23933 , n23927 , n23932 );
not ( n23934 , n17621 );
nand ( n23935 , n23934 , n17586 );
xor ( n23936 , n23916 , n23935 );
or ( n23937 , n23936 , n23844 );
not ( n23938 , n23804 );
nand ( n23939 , n23938 , n23782 );
and ( n23940 , n23747 , n23059 );
not ( n23941 , n23751 );
nor ( n23942 , n23940 , n23941 );
not ( n23943 , n23798 );
or ( n23944 , n23942 , n23943 );
not ( n23945 , n23802 );
nand ( n23946 , n23944 , n23945 );
xor ( n23947 , n23939 , n23946 );
not ( n23948 , n23844 );
or ( n23949 , n23947 , n23948 );
nand ( n23950 , n23937 , n23949 );
not ( n23951 , n10190 );
or ( n23952 , n12789 , n12743 );
nand ( n23953 , n23952 , n499 );
not ( n23954 , n12882 );
xor ( n23955 , n489 , n13133 );
not ( n23956 , n23955 );
or ( n23957 , n23954 , n23956 );
xor ( n23958 , n489 , n13450 );
nand ( n23959 , n23958 , n12635 );
nand ( n23960 , n23957 , n23959 );
xor ( n23961 , n23953 , n23960 );
and ( n23962 , n12922 , n489 );
and ( n23963 , n23961 , n23962 );
and ( n23964 , n23953 , n23960 );
or ( n23965 , n23963 , n23964 );
not ( n23966 , n12845 );
not ( n23967 , n493 );
not ( n23968 , n15576 );
or ( n23969 , n23967 , n23968 );
nand ( n23970 , n15575 , n12862 );
nand ( n23971 , n23969 , n23970 );
not ( n23972 , n23971 );
or ( n23973 , n23966 , n23972 );
not ( n23974 , n493 );
not ( n23975 , n13336 );
or ( n23976 , n23974 , n23975 );
nand ( n23977 , n13339 , n12862 );
nand ( n23978 , n23976 , n23977 );
nand ( n23979 , n23978 , n15386 );
nand ( n23980 , n23973 , n23979 );
and ( n23981 , n12764 , n489 );
xor ( n23982 , n23980 , n23981 );
not ( n23983 , n12731 );
not ( n23984 , n491 );
not ( n23985 , n12512 );
or ( n23986 , n23984 , n23985 );
nand ( n23987 , n12515 , n12703 );
nand ( n23988 , n23986 , n23987 );
not ( n23989 , n23988 );
or ( n23990 , n23983 , n23989 );
not ( n23991 , n491 );
not ( n23992 , n12546 );
or ( n23993 , n23991 , n23992 );
nand ( n23994 , n12549 , n12703 );
nand ( n23995 , n23993 , n23994 );
nand ( n23996 , n23995 , n12688 );
nand ( n23997 , n23990 , n23996 );
and ( n23998 , n23982 , n23997 );
and ( n23999 , n23980 , n23981 );
or ( n24000 , n23998 , n23999 );
xor ( n24001 , n23965 , n24000 );
and ( n24002 , n489 , n13450 );
not ( n24003 , n12845 );
not ( n24004 , n15727 );
and ( n24005 , n24004 , n12862 );
not ( n24006 , n24004 );
and ( n24007 , n24006 , n493 );
or ( n24008 , n24005 , n24007 );
not ( n24009 , n24008 );
or ( n24010 , n24003 , n24009 );
nand ( n24011 , n23971 , n15386 );
nand ( n24012 , n24010 , n24011 );
xor ( n24013 , n24002 , n24012 );
not ( n24014 , n12688 );
not ( n24015 , n23988 );
or ( n24016 , n24014 , n24015 );
not ( n24017 , n491 );
not ( n24018 , n13336 );
or ( n24019 , n24017 , n24018 );
nand ( n24020 , n17764 , n12703 );
nand ( n24021 , n24019 , n24020 );
nand ( n24022 , n24021 , n12731 );
nand ( n24023 , n24016 , n24022 );
xor ( n24024 , n24013 , n24023 );
xor ( n24025 , n24001 , n24024 );
not ( n24026 , n13119 );
not ( n24027 , n16336 );
and ( n24028 , n495 , n24027 );
not ( n24029 , n495 );
and ( n24030 , n24029 , n16336 );
or ( n24031 , n24028 , n24030 );
not ( n24032 , n24031 );
or ( n24033 , n24026 , n24032 );
not ( n24034 , n15952 );
and ( n24035 , n495 , n24034 );
not ( n24036 , n495 );
not ( n24037 , n24034 );
and ( n24038 , n24036 , n24037 );
or ( n24039 , n24035 , n24038 );
nand ( n24040 , n24039 , n13056 );
nand ( n24041 , n24033 , n24040 );
not ( n24042 , n12610 );
buf ( n24043 , n16648 );
and ( n24044 , n497 , n24043 );
not ( n24045 , n497 );
not ( n24046 , n24043 );
and ( n24047 , n24045 , n24046 );
nor ( n24048 , n24044 , n24047 );
not ( n24049 , n24048 );
or ( n24050 , n24042 , n24049 );
nand ( n24051 , n24050 , n16583 );
xor ( n24052 , n24041 , n24051 );
not ( n24053 , n12635 );
not ( n24054 , n23955 );
or ( n24055 , n24053 , n24054 );
xor ( n24056 , n489 , n15602 );
nand ( n24057 , n24056 , n12673 );
nand ( n24058 , n24055 , n24057 );
not ( n24059 , n24058 );
xor ( n24060 , n24052 , n24059 );
not ( n24061 , n13056 );
not ( n24062 , n15727 );
xor ( n24063 , n495 , n24062 );
not ( n24064 , n24063 );
or ( n24065 , n24061 , n24064 );
nand ( n24066 , n24039 , n13119 );
nand ( n24067 , n24065 , n24066 );
not ( n24068 , n12563 );
not ( n24069 , n24048 );
or ( n24070 , n24068 , n24069 );
and ( n24071 , n497 , n16336 );
not ( n24072 , n497 );
and ( n24073 , n24072 , n24027 );
nor ( n24074 , n24071 , n24073 );
nand ( n24075 , n24074 , n12610 );
nand ( n24076 , n24070 , n24075 );
xor ( n24077 , n24067 , n24076 );
not ( n24078 , n12688 );
not ( n24079 , n491 );
not ( n24080 , n15883 );
or ( n24081 , n24079 , n24080 );
nand ( n24082 , n13133 , n12703 );
nand ( n24083 , n24081 , n24082 );
not ( n24084 , n24083 );
or ( n24085 , n24078 , n24084 );
nand ( n24086 , n23995 , n12731 );
nand ( n24087 , n24085 , n24086 );
not ( n24088 , n12673 );
not ( n24089 , n23958 );
or ( n24090 , n24088 , n24089 );
not ( n24091 , n489 );
not ( n24092 , n12923 );
or ( n24093 , n24091 , n24092 );
nand ( n24094 , n12922 , n12653 );
nand ( n24095 , n24093 , n24094 );
nand ( n24096 , n24095 , n12635 );
nand ( n24097 , n24090 , n24096 );
xor ( n24098 , n24087 , n24097 );
not ( n24099 , n13056 );
and ( n24100 , n495 , n15575 );
not ( n24101 , n495 );
and ( n24102 , n24101 , n15579 );
nor ( n24103 , n24100 , n24102 );
not ( n24104 , n24103 );
or ( n24105 , n24099 , n24104 );
nand ( n24106 , n24063 , n13119 );
nand ( n24107 , n24105 , n24106 );
and ( n24108 , n24098 , n24107 );
and ( n24109 , n24087 , n24097 );
or ( n24110 , n24108 , n24109 );
and ( n24111 , n24077 , n24110 );
and ( n24112 , n24067 , n24076 );
or ( n24113 , n24111 , n24112 );
xor ( n24114 , n24060 , n24113 );
xor ( n24115 , n23953 , n23960 );
xor ( n24116 , n24115 , n23962 );
xor ( n24117 , n23980 , n23981 );
xor ( n24118 , n24117 , n23997 );
xor ( n24119 , n24116 , n24118 );
not ( n24120 , n12845 );
not ( n24121 , n23978 );
or ( n24122 , n24120 , n24121 );
not ( n24123 , n493 );
not ( n24124 , n12512 );
or ( n24125 , n24123 , n24124 );
nand ( n24126 , n12862 , n12511 );
nand ( n24127 , n24125 , n24126 );
nand ( n24128 , n24127 , n15386 );
nand ( n24129 , n24122 , n24128 );
not ( n24130 , n23981 );
xor ( n24131 , n24129 , n24130 );
not ( n24132 , n12610 );
xnor ( n24133 , n497 , n15955 );
not ( n24134 , n24133 );
or ( n24135 , n24132 , n24134 );
nand ( n24136 , n24074 , n12563 );
nand ( n24137 , n24135 , n24136 );
and ( n24138 , n24131 , n24137 );
and ( n24139 , n24129 , n24130 );
or ( n24140 , n24138 , n24139 );
and ( n24141 , n24119 , n24140 );
and ( n24142 , n24116 , n24118 );
or ( n24143 , n24141 , n24142 );
xor ( n24144 , n24114 , n24143 );
xor ( n24145 , n24025 , n24144 );
or ( n24146 , n12909 , n12930 );
nand ( n24147 , n24146 , n501 );
and ( n24148 , n13558 , n489 );
xor ( n24149 , n24147 , n24148 );
nand ( n24150 , n13774 , n489 );
not ( n24151 , n24150 );
and ( n24152 , n24149 , n24151 );
and ( n24153 , n24147 , n24148 );
or ( n24154 , n24152 , n24153 );
not ( n24155 , n12789 );
and ( n24156 , n499 , n16649 );
not ( n24157 , n499 );
and ( n24158 , n24157 , n16648 );
or ( n24159 , n24156 , n24158 );
not ( n24160 , n24159 );
or ( n24161 , n24155 , n24160 );
nand ( n24162 , n24161 , n13645 );
xor ( n24163 , n24154 , n24162 );
not ( n24164 , n12731 );
not ( n24165 , n24083 );
or ( n24166 , n24164 , n24165 );
not ( n24167 , n491 );
not ( n24168 , n13451 );
or ( n24169 , n24167 , n24168 );
nand ( n24170 , n12703 , n13450 );
nand ( n24171 , n24169 , n24170 );
nand ( n24172 , n24171 , n12688 );
nand ( n24173 , n24166 , n24172 );
not ( n24174 , n12673 );
not ( n24175 , n24095 );
or ( n24176 , n24174 , n24175 );
and ( n24177 , n489 , n12764 );
not ( n24178 , n489 );
and ( n24179 , n24178 , n13438 );
nor ( n24180 , n24177 , n24179 );
nand ( n24181 , n24180 , n12635 );
nand ( n24182 , n24176 , n24181 );
xor ( n24183 , n24173 , n24182 );
not ( n24184 , n13119 );
not ( n24185 , n24103 );
or ( n24186 , n24184 , n24185 );
not ( n24187 , n495 );
not ( n24188 , n13336 );
or ( n24189 , n24187 , n24188 );
not ( n24190 , n495 );
nand ( n24191 , n24190 , n13339 );
nand ( n24192 , n24189 , n24191 );
nand ( n24193 , n24192 , n13056 );
nand ( n24194 , n24186 , n24193 );
and ( n24195 , n24183 , n24194 );
and ( n24196 , n24173 , n24182 );
or ( n24197 , n24195 , n24196 );
and ( n24198 , n24163 , n24197 );
and ( n24199 , n24154 , n24162 );
or ( n24200 , n24198 , n24199 );
xor ( n24201 , n24067 , n24076 );
xor ( n24202 , n24201 , n24110 );
xor ( n24203 , n24200 , n24202 );
xor ( n24204 , n24087 , n24097 );
xor ( n24205 , n24204 , n24107 );
not ( n24206 , n12845 );
not ( n24207 , n24127 );
or ( n24208 , n24206 , n24207 );
not ( n24209 , n493 );
not ( n24210 , n15599 );
or ( n24211 , n24209 , n24210 );
nand ( n24212 , n15602 , n12862 );
nand ( n24213 , n24211 , n24212 );
nand ( n24214 , n24213 , n15386 );
nand ( n24215 , n24208 , n24214 );
not ( n24216 , n12563 );
not ( n24217 , n24133 );
or ( n24218 , n24216 , n24217 );
xor ( n24219 , n497 , n16271 );
nand ( n24220 , n24219 , n12610 );
nand ( n24221 , n24218 , n24220 );
xor ( n24222 , n24215 , n24221 );
not ( n24223 , n12743 );
not ( n24224 , n24159 );
or ( n24225 , n24223 , n24224 );
not ( n24226 , n499 );
not ( n24227 , n16333 );
or ( n24228 , n24226 , n24227 );
nand ( n24229 , n12560 , n16336 );
nand ( n24230 , n24228 , n24229 );
nand ( n24231 , n24230 , n12789 );
nand ( n24232 , n24225 , n24231 );
and ( n24233 , n24222 , n24232 );
and ( n24234 , n24215 , n24221 );
or ( n24235 , n24233 , n24234 );
xor ( n24236 , n24205 , n24235 );
xor ( n24237 , n24129 , n24130 );
xor ( n24238 , n24237 , n24137 );
and ( n24239 , n24236 , n24238 );
and ( n24240 , n24205 , n24235 );
or ( n24241 , n24239 , n24240 );
and ( n24242 , n24203 , n24241 );
and ( n24243 , n24200 , n24202 );
or ( n24244 , n24242 , n24243 );
xor ( n24245 , n24145 , n24244 );
not ( n24246 , n24245 );
xor ( n24247 , n24116 , n24118 );
xor ( n24248 , n24247 , n24140 );
xor ( n24249 , n24200 , n24202 );
xor ( n24250 , n24249 , n24241 );
xor ( n24251 , n24248 , n24250 );
not ( n24252 , n12635 );
not ( n24253 , n489 );
not ( n24254 , n12781 );
or ( n24255 , n24253 , n24254 );
not ( n24256 , n489 );
nand ( n24257 , n24256 , n12780 );
nand ( n24258 , n24255 , n24257 );
not ( n24259 , n24258 );
or ( n24260 , n24252 , n24259 );
nand ( n24261 , n24180 , n12673 );
nand ( n24262 , n24260 , n24261 );
xor ( n24263 , n24262 , n24150 );
nand ( n24264 , n12602 , n489 );
not ( n24265 , n12555 );
nand ( n24266 , n24265 , n699 );
nand ( n24267 , n24264 , n24266 );
and ( n24268 , n24263 , n24267 );
and ( n24269 , n24262 , n24150 );
or ( n24270 , n24268 , n24269 );
xor ( n24271 , n24147 , n24148 );
xor ( n24272 , n24271 , n24151 );
xor ( n24273 , n24270 , n24272 );
not ( n24274 , n24213 );
not ( n24275 , n12845 );
or ( n24276 , n24274 , n24275 );
not ( n24277 , n12972 );
not ( n24278 , n12862 );
or ( n24279 , n24277 , n24278 );
nand ( n24280 , n12973 , n493 );
nand ( n24281 , n24279 , n24280 );
nand ( n24282 , n24281 , n15386 );
nand ( n24283 , n24276 , n24282 );
not ( n24284 , n12731 );
not ( n24285 , n24171 );
or ( n24286 , n24284 , n24285 );
not ( n24287 , n12911 );
not ( n24288 , n12916 );
or ( n24289 , n24287 , n24288 );
nand ( n24290 , n24289 , n12921 );
and ( n24291 , n24290 , n12703 );
not ( n24292 , n24290 );
and ( n24293 , n24292 , n491 );
or ( n24294 , n24291 , n24293 );
nand ( n24295 , n24294 , n12688 );
nand ( n24296 , n24286 , n24295 );
xor ( n24297 , n24283 , n24296 );
not ( n24298 , n12563 );
not ( n24299 , n24219 );
or ( n24300 , n24298 , n24299 );
and ( n24301 , n15574 , n497 );
not ( n24302 , n15574 );
and ( n24303 , n24302 , n864 );
nor ( n24304 , n24301 , n24303 );
nand ( n24305 , n24304 , n12610 );
nand ( n24306 , n24300 , n24305 );
and ( n24307 , n24297 , n24306 );
and ( n24308 , n24283 , n24296 );
or ( n24309 , n24307 , n24308 );
and ( n24310 , n24273 , n24309 );
and ( n24311 , n24270 , n24272 );
or ( n24312 , n24310 , n24311 );
xor ( n24313 , n24154 , n24162 );
xor ( n24314 , n24313 , n24197 );
xor ( n24315 , n24312 , n24314 );
xor ( n24316 , n24173 , n24182 );
xor ( n24317 , n24316 , n24194 );
xor ( n24318 , n24215 , n24221 );
xor ( n24319 , n24318 , n24232 );
xor ( n24320 , n24317 , n24319 );
not ( n24321 , n13119 );
not ( n24322 , n24192 );
or ( n24323 , n24321 , n24322 );
not ( n24324 , n3583 );
not ( n24325 , n12511 );
or ( n24326 , n24324 , n24325 );
nand ( n24327 , n495 , n15474 );
nand ( n24328 , n24326 , n24327 );
nand ( n24329 , n24328 , n13056 );
nand ( n24330 , n24323 , n24329 );
not ( n24331 , n12743 );
not ( n24332 , n24230 );
or ( n24333 , n24331 , n24332 );
not ( n24334 , n499 );
not ( n24335 , n24034 );
or ( n24336 , n24334 , n24335 );
nand ( n24337 , n15952 , n12560 );
nand ( n24338 , n24336 , n24337 );
nand ( n24339 , n24338 , n12789 );
nand ( n24340 , n24333 , n24339 );
xor ( n24341 , n24330 , n24340 );
not ( n24342 , n12909 );
not ( n24343 , n501 );
not ( n24344 , n16649 );
or ( n24345 , n24343 , n24344 );
nand ( n24346 , n1845 , n16648 );
nand ( n24347 , n24345 , n24346 );
not ( n24348 , n24347 );
or ( n24349 , n24342 , n24348 );
nand ( n24350 , n24349 , n16272 );
and ( n24351 , n24341 , n24350 );
and ( n24352 , n24330 , n24340 );
or ( n24353 , n24351 , n24352 );
and ( n24354 , n24320 , n24353 );
and ( n24355 , n24317 , n24319 );
or ( n24356 , n24354 , n24355 );
and ( n24357 , n24315 , n24356 );
and ( n24358 , n24312 , n24314 );
or ( n24359 , n24357 , n24358 );
and ( n24360 , n24251 , n24359 );
and ( n24361 , n24248 , n24250 );
or ( n24362 , n24360 , n24361 );
not ( n24363 , n24362 );
nand ( n24364 , n24246 , n24363 );
not ( n24365 , n24364 );
xor ( n24366 , n24205 , n24235 );
xor ( n24367 , n24366 , n24238 );
xor ( n24368 , n24312 , n24314 );
xor ( n24369 , n24368 , n24356 );
xor ( n24370 , n24367 , n24369 );
xor ( n24371 , n24270 , n24272 );
xor ( n24372 , n24371 , n24309 );
not ( n24373 , n12673 );
not ( n24374 , n24258 );
or ( n24375 , n24373 , n24374 );
nand ( n24376 , n17806 , n12635 );
nand ( n24377 , n24375 , n24376 );
not ( n24378 , n17799 );
and ( n24379 , n17810 , n24378 );
xor ( n24380 , n24377 , n24379 );
or ( n24381 , n24264 , n24266 );
nand ( n24382 , n24381 , n24267 );
and ( n24383 , n24380 , n24382 );
and ( n24384 , n24377 , n24379 );
or ( n24385 , n24383 , n24384 );
xor ( n24386 , n24262 , n24150 );
xor ( n24387 , n24386 , n24267 );
xor ( n24388 , n24385 , n24387 );
xor ( n24389 , n24283 , n24296 );
xor ( n24390 , n24389 , n24306 );
and ( n24391 , n24388 , n24390 );
and ( n24392 , n24385 , n24387 );
or ( n24393 , n24391 , n24392 );
xor ( n24394 , n24372 , n24393 );
not ( n24395 , n12845 );
not ( n24396 , n24281 );
or ( n24397 , n24395 , n24396 );
nand ( n24398 , n17728 , n15386 );
nand ( n24399 , n24397 , n24398 );
not ( n24400 , n12731 );
not ( n24401 , n24294 );
or ( n24402 , n24400 , n24401 );
nand ( n24403 , n12688 , n17794 );
nand ( n24404 , n24402 , n24403 );
xor ( n24405 , n24399 , n24404 );
not ( n24406 , n12563 );
not ( n24407 , n24304 );
or ( n24408 , n24406 , n24407 );
not ( n24409 , n497 );
not ( n24410 , n13336 );
or ( n24411 , n24409 , n24410 );
nand ( n24412 , n13339 , n12579 );
nand ( n24413 , n24411 , n24412 );
nand ( n24414 , n24413 , n12610 );
nand ( n24415 , n24408 , n24414 );
and ( n24416 , n24405 , n24415 );
and ( n24417 , n24399 , n24404 );
or ( n24418 , n24416 , n24417 );
not ( n24419 , n13119 );
not ( n24420 , n24328 );
or ( n24421 , n24419 , n24420 );
nand ( n24422 , n17718 , n13056 );
nand ( n24423 , n24421 , n24422 );
not ( n24424 , n12789 );
not ( n24425 , n17739 );
or ( n24426 , n24424 , n24425 );
nand ( n24427 , n24338 , n12743 );
nand ( n24428 , n24426 , n24427 );
xor ( n24429 , n24423 , n24428 );
not ( n24430 , n12930 );
not ( n24431 , n24347 );
or ( n24432 , n24430 , n24431 );
not ( n24433 , n501 );
not ( n24434 , n16333 );
or ( n24435 , n24433 , n24434 );
nand ( n24436 , n16336 , n12943 );
nand ( n24437 , n24435 , n24436 );
nand ( n24438 , n24437 , n12909 );
nand ( n24439 , n24432 , n24438 );
and ( n24440 , n24429 , n24439 );
and ( n24441 , n24423 , n24428 );
or ( n24442 , n24440 , n24441 );
xor ( n24443 , n24418 , n24442 );
xor ( n24444 , n24330 , n24340 );
xor ( n24445 , n24444 , n24350 );
and ( n24446 , n24443 , n24445 );
and ( n24447 , n24418 , n24442 );
or ( n24448 , n24446 , n24447 );
and ( n24449 , n24394 , n24448 );
and ( n24450 , n24372 , n24393 );
or ( n24451 , n24449 , n24450 );
xor ( n24452 , n24370 , n24451 );
xor ( n24453 , n24317 , n24319 );
xor ( n24454 , n24453 , n24353 );
xor ( n24455 , n17796 , n17797 );
and ( n24456 , n24455 , n17814 );
and ( n24457 , n17796 , n17797 );
or ( n24458 , n24456 , n24457 );
xor ( n24459 , n24377 , n24379 );
xor ( n24460 , n24459 , n24382 );
xor ( n24461 , n24458 , n24460 );
xor ( n24462 , n17720 , n17730 );
and ( n24463 , n24462 , n17741 );
and ( n24464 , n17720 , n17730 );
or ( n24465 , n24463 , n24464 );
and ( n24466 , n24461 , n24465 );
and ( n24467 , n24458 , n24460 );
or ( n24468 , n24466 , n24467 );
xor ( n24469 , n24385 , n24387 );
xor ( n24470 , n24469 , n24390 );
xor ( n24471 , n24468 , n24470 );
xor ( n24472 , n24399 , n24404 );
xor ( n24473 , n24472 , n24415 );
xor ( n24474 , n17767 , n17776 );
and ( n24475 , n24474 , n17781 );
and ( n24476 , n17767 , n17776 );
or ( n24477 , n24475 , n24476 );
xor ( n24478 , n24473 , n24477 );
xor ( n24479 , n24423 , n24428 );
xor ( n24480 , n24479 , n24439 );
and ( n24481 , n24478 , n24480 );
and ( n24482 , n24473 , n24477 );
or ( n24483 , n24481 , n24482 );
and ( n24484 , n24471 , n24483 );
and ( n24485 , n24468 , n24470 );
or ( n24486 , n24484 , n24485 );
xor ( n24487 , n24454 , n24486 );
xor ( n24488 , n24372 , n24393 );
xor ( n24489 , n24488 , n24448 );
and ( n24490 , n24487 , n24489 );
and ( n24491 , n24454 , n24486 );
or ( n24492 , n24490 , n24491 );
nor ( n24493 , n24452 , n24492 );
xor ( n24494 , n24248 , n24250 );
xor ( n24495 , n24494 , n24359 );
xor ( n24496 , n24367 , n24369 );
and ( n24497 , n24496 , n24451 );
and ( n24498 , n24367 , n24369 );
or ( n24499 , n24497 , n24498 );
nor ( n24500 , n24495 , n24499 );
nor ( n24501 , n24493 , n24500 );
not ( n24502 , n24501 );
xor ( n24503 , n17752 , n17827 );
and ( n24504 , n24503 , n17832 );
and ( n24505 , n17752 , n17827 );
or ( n24506 , n24504 , n24505 );
xor ( n24507 , n17742 , n17746 );
and ( n24508 , n24507 , n17751 );
and ( n24509 , n17742 , n17746 );
or ( n24510 , n24508 , n24509 );
xor ( n24511 , n17782 , n17821 );
and ( n24512 , n24511 , n17826 );
and ( n24513 , n17782 , n17821 );
or ( n24514 , n24512 , n24513 );
xor ( n24515 , n24510 , n24514 );
xor ( n24516 , n17786 , n17815 );
and ( n24517 , n24516 , n17820 );
and ( n24518 , n17786 , n17815 );
or ( n24519 , n24517 , n24518 );
xor ( n24520 , n24458 , n24460 );
xor ( n24521 , n24520 , n24465 );
xor ( n24522 , n24519 , n24521 );
xor ( n24523 , n24473 , n24477 );
xor ( n24524 , n24523 , n24480 );
xor ( n24525 , n24522 , n24524 );
xor ( n24526 , n24515 , n24525 );
nor ( n24527 , n24506 , n24526 );
not ( n24528 , n24527 );
xor ( n24529 , n24418 , n24442 );
xor ( n24530 , n24529 , n24445 );
xor ( n24531 , n24468 , n24470 );
xor ( n24532 , n24531 , n24483 );
xor ( n24533 , n24530 , n24532 );
xor ( n24534 , n24519 , n24521 );
and ( n24535 , n24534 , n24524 );
and ( n24536 , n24519 , n24521 );
or ( n24537 , n24535 , n24536 );
xor ( n24538 , n24533 , n24537 );
xor ( n24539 , n24510 , n24514 );
and ( n24540 , n24539 , n24525 );
and ( n24541 , n24510 , n24514 );
or ( n24542 , n24540 , n24541 );
nor ( n24543 , n24538 , n24542 );
not ( n24544 , n24543 );
xor ( n24545 , n24530 , n24532 );
and ( n24546 , n24545 , n24537 );
and ( n24547 , n24530 , n24532 );
or ( n24548 , n24546 , n24547 );
not ( n24549 , n24548 );
xor ( n24550 , n24454 , n24486 );
xor ( n24551 , n24550 , n24489 );
not ( n24552 , n24551 );
nand ( n24553 , n24549 , n24552 );
nand ( n24554 , n24528 , n17843 , n24544 , n24553 );
nor ( n24555 , n17709 , n24554 );
not ( n24556 , n24526 );
not ( n24557 , n24506 );
or ( n24558 , n24556 , n24557 );
nand ( n24559 , n24551 , n24548 );
nand ( n24560 , n24558 , n24559 );
and ( n24561 , n24538 , n24542 );
nor ( n24562 , n24560 , n24561 );
not ( n24563 , n24527 );
nand ( n24564 , n24563 , n17840 );
and ( n24565 , n24562 , n24564 );
not ( n24566 , n24538 );
not ( n24567 , n24542 );
nand ( n24568 , n24566 , n24567 );
nand ( n24569 , n24553 , n24568 );
nand ( n24570 , n24548 , n24551 );
and ( n24571 , n24569 , n24570 );
nor ( n24572 , n24565 , n24571 );
nor ( n24573 , n24555 , n24572 );
not ( n24574 , n15807 );
not ( n24575 , n15801 );
or ( n24576 , n24574 , n24575 );
nor ( n24577 , n24554 , n17704 );
nand ( n24578 , n24576 , n24577 );
nand ( n24579 , n24573 , n24578 );
not ( n24580 , n24579 );
or ( n24581 , n24502 , n24580 );
nor ( n24582 , n24495 , n24499 );
nand ( n24583 , n24452 , n24492 );
or ( n24584 , n24582 , n24583 );
nand ( n24585 , n24495 , n24499 );
nand ( n24586 , n24584 , n24585 );
not ( n24587 , n24586 );
nand ( n24588 , n24581 , n24587 );
not ( n24589 , n24588 );
or ( n24590 , n24365 , n24589 );
nand ( n24591 , n24245 , n24362 );
nand ( n24592 , n24590 , n24591 );
xor ( n24593 , n24025 , n24144 );
and ( n24594 , n24593 , n24244 );
and ( n24595 , n24025 , n24144 );
or ( n24596 , n24594 , n24595 );
xor ( n24597 , n23965 , n24000 );
and ( n24598 , n24597 , n24024 );
and ( n24599 , n23965 , n24000 );
or ( n24600 , n24598 , n24599 );
xor ( n24601 , n24041 , n24051 );
and ( n24602 , n24601 , n24059 );
and ( n24603 , n24041 , n24051 );
or ( n24604 , n24602 , n24603 );
not ( n24605 , n12673 );
not ( n24606 , n489 );
not ( n24607 , n12512 );
or ( n24608 , n24606 , n24607 );
nand ( n24609 , n12515 , n12653 );
nand ( n24610 , n24608 , n24609 );
not ( n24611 , n24610 );
or ( n24612 , n24605 , n24611 );
nand ( n24613 , n24056 , n12635 );
nand ( n24614 , n24612 , n24613 );
not ( n24615 , n15386 );
not ( n24616 , n24008 );
or ( n24617 , n24615 , n24616 );
not ( n24618 , n493 );
not ( n24619 , n24034 );
or ( n24620 , n24618 , n24619 );
nand ( n24621 , n24037 , n12862 );
nand ( n24622 , n24620 , n24621 );
nand ( n24623 , n24622 , n12845 );
nand ( n24624 , n24617 , n24623 );
xor ( n24625 , n24614 , n24624 );
not ( n24626 , n13119 );
and ( n24627 , n495 , n24046 );
not ( n24628 , n495 );
and ( n24629 , n24628 , n24043 );
or ( n24630 , n24627 , n24629 );
not ( n24631 , n24630 );
or ( n24632 , n24626 , n24631 );
nand ( n24633 , n24031 , n13056 );
nand ( n24634 , n24632 , n24633 );
xor ( n24635 , n24625 , n24634 );
xor ( n24636 , n24604 , n24635 );
xor ( n24637 , n24002 , n24012 );
and ( n24638 , n24637 , n24023 );
and ( n24639 , n24002 , n24012 );
or ( n24640 , n24638 , n24639 );
xor ( n24641 , n24058 , n24640 );
or ( n24642 , n12610 , n12563 );
nand ( n24643 , n24642 , n497 );
and ( n24644 , n489 , n13133 );
xor ( n24645 , n24643 , n24644 );
not ( n24646 , n12731 );
not ( n24647 , n491 );
not ( n24648 , n15579 );
or ( n24649 , n24647 , n24648 );
nand ( n24650 , n15580 , n12703 );
nand ( n24651 , n24649 , n24650 );
not ( n24652 , n24651 );
or ( n24653 , n24646 , n24652 );
nand ( n24654 , n24021 , n12688 );
nand ( n24655 , n24653 , n24654 );
xor ( n24656 , n24645 , n24655 );
xor ( n24657 , n24641 , n24656 );
xor ( n24658 , n24636 , n24657 );
xor ( n24659 , n24600 , n24658 );
xor ( n24660 , n24060 , n24113 );
and ( n24661 , n24660 , n24143 );
and ( n24662 , n24060 , n24113 );
or ( n24663 , n24661 , n24662 );
xor ( n24664 , n24659 , n24663 );
or ( n24665 , n24596 , n24664 );
nand ( n24666 , n24664 , n24596 );
nand ( n24667 , n24665 , n24666 );
not ( n24668 , n24667 );
and ( n24669 , n24592 , n24668 );
not ( n24670 , n24592 );
xnor ( n24671 , n24596 , n24664 );
and ( n24672 , n24670 , n24671 );
nor ( n24673 , n24669 , n24672 );
not ( n24674 , n24673 );
or ( n24675 , n23951 , n24674 );
nand ( n24676 , n16517 , n16414 );
and ( n24677 , n16408 , n24676 );
not ( n24678 , n17974 );
not ( n24679 , n16513 );
not ( n24680 , n16414 );
nand ( n24681 , n24679 , n24680 );
nand ( n24682 , n24678 , n24681 );
nor ( n24683 , n24677 , n24682 );
not ( n24684 , n17977 );
nor ( n24685 , n24683 , n24684 );
not ( n24686 , n16403 );
not ( n24687 , n17974 );
nand ( n24688 , n24687 , n24681 );
nor ( n24689 , n24686 , n24688 );
nand ( n24690 , n24689 , n10051 );
nand ( n24691 , n24685 , n24690 );
or ( n24692 , n7127 , n6983 );
nand ( n24693 , n24692 , n547 );
not ( n24694 , n537 );
nor ( n24695 , n24694 , n7544 );
xor ( n24696 , n24693 , n24695 );
nor ( n24697 , n7057 , n5325 );
and ( n24698 , n24696 , n24697 );
and ( n24699 , n24693 , n24695 );
or ( n24700 , n24698 , n24699 );
not ( n24701 , n5341 );
and ( n24702 , n9688 , n4666 );
not ( n24703 , n9688 );
and ( n24704 , n24703 , n545 );
or ( n24705 , n24702 , n24704 );
not ( n24706 , n24705 );
or ( n24707 , n24701 , n24706 );
not ( n24708 , n793 );
not ( n24709 , n9974 );
or ( n24710 , n24708 , n24709 );
nand ( n24711 , n9923 , n455 );
nand ( n24712 , n24710 , n24711 );
and ( n24713 , n24712 , n545 );
not ( n24714 , n24712 );
and ( n24715 , n24714 , n5470 );
nor ( n24716 , n24713 , n24715 );
nand ( n24717 , n24716 , n5595 );
nand ( n24718 , n24707 , n24717 );
not ( n24719 , n5786 );
not ( n24720 , n541 );
not ( n24721 , n9867 );
or ( n24722 , n24720 , n24721 );
nand ( n24723 , n9866 , n5734 );
nand ( n24724 , n24722 , n24723 );
not ( n24725 , n24724 );
or ( n24726 , n24719 , n24725 );
not ( n24727 , n541 );
not ( n24728 , n10074 );
or ( n24729 , n24727 , n24728 );
nand ( n24730 , n6967 , n5734 );
nand ( n24731 , n24729 , n24730 );
nand ( n24732 , n24731 , n10067 );
nand ( n24733 , n24726 , n24732 );
xor ( n24734 , n24718 , n24733 );
not ( n24735 , n4660 );
not ( n24736 , n539 );
not ( n24737 , n7039 );
or ( n24738 , n24736 , n24737 );
not ( n24739 , n7039 );
nand ( n24740 , n24739 , n4477 );
nand ( n24741 , n24738 , n24740 );
not ( n24742 , n24741 );
or ( n24743 , n24735 , n24742 );
not ( n24744 , n4477 );
not ( n24745 , n7341 );
not ( n24746 , n24745 );
or ( n24747 , n24744 , n24746 );
nand ( n24748 , n7341 , n539 );
nand ( n24749 , n24747 , n24748 );
nand ( n24750 , n24749 , n4450 );
nand ( n24751 , n24743 , n24750 );
and ( n24752 , n24734 , n24751 );
and ( n24753 , n24718 , n24733 );
or ( n24754 , n24752 , n24753 );
xor ( n24755 , n24700 , n24754 );
not ( n24756 , n5786 );
not ( n24757 , n541 );
not ( n24758 , n9517 );
or ( n24759 , n24757 , n24758 );
nand ( n24760 , n7326 , n5734 );
nand ( n24761 , n24759 , n24760 );
not ( n24762 , n24761 );
or ( n24763 , n24756 , n24762 );
nand ( n24764 , n24724 , n10067 );
nand ( n24765 , n24763 , n24764 );
nand ( n24766 , n7470 , n537 );
xor ( n24767 , n24765 , n24766 );
not ( n24768 , n5341 );
and ( n24769 , n24712 , n545 );
not ( n24770 , n24712 );
and ( n24771 , n24770 , n4666 );
nor ( n24772 , n24769 , n24771 );
not ( n24773 , n24772 );
or ( n24774 , n24768 , n24773 );
nand ( n24775 , n5595 , n545 );
nand ( n24776 , n24774 , n24775 );
xor ( n24777 , n24767 , n24776 );
and ( n24778 , n24755 , n24777 );
and ( n24779 , n24700 , n24754 );
or ( n24780 , n24778 , n24779 );
not ( n24781 , n5697 );
not ( n24782 , n537 );
not ( n24783 , n7039 );
or ( n24784 , n24782 , n24783 );
nand ( n24785 , n24739 , n5605 );
nand ( n24786 , n24784 , n24785 );
not ( n24787 , n24786 );
or ( n24788 , n24781 , n24787 );
not ( n24789 , n537 );
not ( n24790 , n7341 );
or ( n24791 , n24789 , n24790 );
nand ( n24792 , n24745 , n5605 );
nand ( n24793 , n24791 , n24792 );
nand ( n24794 , n24793 , n16173 );
nand ( n24795 , n24788 , n24794 );
not ( n24796 , n5786 );
not ( n24797 , n541 );
not ( n24798 , n9692 );
or ( n24799 , n24797 , n24798 );
not ( n24800 , n9692 );
nand ( n24801 , n24800 , n5734 );
nand ( n24802 , n24799 , n24801 );
not ( n24803 , n24802 );
or ( n24804 , n24796 , n24803 );
nand ( n24805 , n24761 , n10067 );
nand ( n24806 , n24804 , n24805 );
xor ( n24807 , n24795 , n24806 );
and ( n24808 , n537 , n7020 );
xor ( n24809 , n24807 , n24808 );
or ( n24810 , n5341 , n5595 );
nand ( n24811 , n24810 , n545 );
not ( n24812 , n4671 );
not ( n24813 , n543 );
not ( n24814 , n9689 );
or ( n24815 , n24813 , n24814 );
nand ( n24816 , n9886 , n5146 );
nand ( n24817 , n24815 , n24816 );
not ( n24818 , n24817 );
or ( n24819 , n24812 , n24818 );
not ( n24820 , n543 );
not ( n24821 , n9977 );
or ( n24822 , n24820 , n24821 );
buf ( n24823 , n9976 );
nand ( n24824 , n24823 , n5146 );
nand ( n24825 , n24822 , n24824 );
nand ( n24826 , n24825 , n9730 );
nand ( n24827 , n24819 , n24826 );
xor ( n24828 , n24811 , n24827 );
not ( n24829 , n4660 );
not ( n24830 , n539 );
not ( n24831 , n9867 );
or ( n24832 , n24830 , n24831 );
not ( n24833 , n9867 );
nand ( n24834 , n24833 , n4477 );
nand ( n24835 , n24832 , n24834 );
not ( n24836 , n24835 );
or ( n24837 , n24829 , n24836 );
not ( n24838 , n539 );
buf ( n24839 , n6967 );
not ( n24840 , n24839 );
not ( n24841 , n24840 );
or ( n24842 , n24838 , n24841 );
nand ( n24843 , n24839 , n4477 );
nand ( n24844 , n24842 , n24843 );
nand ( n24845 , n4450 , n24844 );
nand ( n24846 , n24837 , n24845 );
xor ( n24847 , n24828 , n24846 );
xor ( n24848 , n24809 , n24847 );
not ( n24849 , n24766 );
not ( n24850 , n4671 );
not ( n24851 , n543 );
not ( n24852 , n9692 );
or ( n24853 , n24851 , n24852 );
nand ( n24854 , n24800 , n5146 );
nand ( n24855 , n24853 , n24854 );
not ( n24856 , n24855 );
or ( n24857 , n24850 , n24856 );
nand ( n24858 , n24817 , n9730 );
nand ( n24859 , n24857 , n24858 );
not ( n24860 , n4659 );
not ( n24861 , n24844 );
or ( n24862 , n24860 , n24861 );
nand ( n24863 , n24741 , n4450 );
nand ( n24864 , n24862 , n24863 );
xor ( n24865 , n24859 , n24864 );
not ( n24866 , n24793 );
not ( n24867 , n5697 );
or ( n24868 , n24866 , n24867 );
xor ( n24869 , n537 , n7020 );
not ( n24870 , n24869 );
not ( n24871 , n16173 );
or ( n24872 , n24870 , n24871 );
nand ( n24873 , n24868 , n24872 );
and ( n24874 , n24865 , n24873 );
and ( n24875 , n24859 , n24864 );
or ( n24876 , n24874 , n24875 );
xor ( n24877 , n24849 , n24876 );
xor ( n24878 , n24765 , n24766 );
and ( n24879 , n24878 , n24776 );
and ( n24880 , n24765 , n24766 );
or ( n24881 , n24879 , n24880 );
xor ( n24882 , n24877 , n24881 );
xor ( n24883 , n24848 , n24882 );
xor ( n24884 , n24780 , n24883 );
xor ( n24885 , n24859 , n24864 );
xor ( n24886 , n24885 , n24873 );
not ( n24887 , n5697 );
not ( n24888 , n24869 );
or ( n24889 , n24887 , n24888 );
not ( n24890 , n537 );
not ( n24891 , n7469 );
or ( n24892 , n24890 , n24891 );
nand ( n24893 , n5588 , n5605 );
nand ( n24894 , n24892 , n24893 );
nand ( n24895 , n24894 , n16173 );
nand ( n24896 , n24889 , n24895 );
not ( n24897 , n9730 );
not ( n24898 , n24855 );
or ( n24899 , n24897 , n24898 );
not ( n24900 , n543 );
not ( n24901 , n9517 );
or ( n24902 , n24900 , n24901 );
not ( n24903 , n9517 );
nand ( n24904 , n24903 , n5146 );
nand ( n24905 , n24902 , n24904 );
nand ( n24906 , n24905 , n4671 );
nand ( n24907 , n24899 , n24906 );
xor ( n24908 , n24896 , n24907 );
xor ( n24909 , n24693 , n24695 );
xor ( n24910 , n24909 , n24697 );
and ( n24911 , n24908 , n24910 );
and ( n24912 , n24896 , n24907 );
or ( n24913 , n24911 , n24912 );
xor ( n24914 , n24886 , n24913 );
not ( n24915 , n5697 );
not ( n24916 , n24894 );
or ( n24917 , n24915 , n24916 );
nand ( n24918 , n17910 , n16173 );
nand ( n24919 , n24917 , n24918 );
not ( n24920 , n24697 );
xor ( n24921 , n24919 , n24920 );
not ( n24922 , n17898 );
or ( n24923 , n24922 , n5340 );
not ( n24924 , n24705 );
or ( n24925 , n24924 , n7809 );
nand ( n24926 , n24923 , n24925 );
and ( n24927 , n24921 , n24926 );
and ( n24928 , n24919 , n24920 );
or ( n24929 , n24927 , n24928 );
not ( n24930 , n5786 );
not ( n24931 , n24731 );
or ( n24932 , n24930 , n24931 );
nand ( n24933 , n17874 , n10067 );
nand ( n24934 , n24932 , n24933 );
xor ( n24935 , n17939 , n17940 );
and ( n24936 , n24935 , n17942 );
and ( n24937 , n17939 , n17940 );
or ( n24938 , n24936 , n24937 );
xor ( n24939 , n24934 , n24938 );
not ( n24940 , n24749 );
or ( n24941 , n24940 , n5970 );
not ( n24942 , n17883 );
or ( n24943 , n24942 , n5961 );
nand ( n24944 , n24941 , n24943 );
and ( n24945 , n24939 , n24944 );
and ( n24946 , n24934 , n24938 );
or ( n24947 , n24945 , n24946 );
xor ( n24948 , n24929 , n24947 );
xor ( n24949 , n24718 , n24733 );
xor ( n24950 , n24949 , n24751 );
and ( n24951 , n24948 , n24950 );
and ( n24952 , n24929 , n24947 );
or ( n24953 , n24951 , n24952 );
and ( n24954 , n24914 , n24953 );
and ( n24955 , n24886 , n24913 );
or ( n24956 , n24954 , n24955 );
xor ( n24957 , n24884 , n24956 );
not ( n24958 , n24957 );
xor ( n24959 , n24700 , n24754 );
xor ( n24960 , n24959 , n24777 );
xor ( n24961 , n24886 , n24913 );
xor ( n24962 , n24961 , n24953 );
xor ( n24963 , n24960 , n24962 );
xor ( n24964 , n24896 , n24907 );
xor ( n24965 , n24964 , n24910 );
not ( n24966 , n7026 );
not ( n24967 , n17931 );
or ( n24968 , n24966 , n24967 );
nand ( n24969 , n24968 , n7797 );
not ( n24970 , n4671 );
not ( n24971 , n17920 );
or ( n24972 , n24970 , n24971 );
nand ( n24973 , n24905 , n9730 );
nand ( n24974 , n24972 , n24973 );
xor ( n24975 , n24969 , n24974 );
xor ( n24976 , n17878 , n17891 );
and ( n24977 , n24976 , n17902 );
and ( n24978 , n17878 , n17891 );
or ( n24979 , n24977 , n24978 );
and ( n24980 , n24975 , n24979 );
and ( n24981 , n24969 , n24974 );
or ( n24982 , n24980 , n24981 );
xor ( n24983 , n24965 , n24982 );
xor ( n24984 , n24929 , n24947 );
xor ( n24985 , n24984 , n24950 );
and ( n24986 , n24983 , n24985 );
and ( n24987 , n24965 , n24982 );
or ( n24988 , n24986 , n24987 );
and ( n24989 , n24963 , n24988 );
and ( n24990 , n24960 , n24962 );
or ( n24991 , n24989 , n24990 );
not ( n24992 , n24991 );
nand ( n24993 , n24958 , n24992 );
xor ( n24994 , n17914 , n17924 );
and ( n24995 , n24994 , n17935 );
and ( n24996 , n17914 , n17924 );
or ( n24997 , n24995 , n24996 );
xor ( n24998 , n24919 , n24920 );
xor ( n24999 , n24998 , n24926 );
xor ( n25000 , n24997 , n24999 );
xor ( n25001 , n24934 , n24938 );
xor ( n25002 , n25001 , n24944 );
and ( n25003 , n25000 , n25002 );
and ( n25004 , n24997 , n24999 );
or ( n25005 , n25003 , n25004 );
xor ( n25006 , n24965 , n24982 );
xor ( n25007 , n25006 , n24985 );
xor ( n25008 , n25005 , n25007 );
xor ( n25009 , n24969 , n24974 );
xor ( n25010 , n25009 , n24979 );
xor ( n25011 , n17943 , n17947 );
and ( n25012 , n25011 , n17952 );
and ( n25013 , n17943 , n17947 );
or ( n25014 , n25012 , n25013 );
xor ( n25015 , n25010 , n25014 );
xor ( n25016 , n17868 , n17903 );
and ( n25017 , n25016 , n17936 );
and ( n25018 , n17868 , n17903 );
or ( n25019 , n25017 , n25018 );
and ( n25020 , n25015 , n25019 );
and ( n25021 , n25010 , n25014 );
or ( n25022 , n25020 , n25021 );
xor ( n25023 , n25008 , n25022 );
xor ( n25024 , n24997 , n24999 );
xor ( n25025 , n25024 , n25002 );
xor ( n25026 , n25010 , n25014 );
xor ( n25027 , n25026 , n25019 );
xor ( n25028 , n25025 , n25027 );
xor ( n25029 , n17953 , n17957 );
and ( n25030 , n25029 , n17962 );
and ( n25031 , n17953 , n17957 );
or ( n25032 , n25030 , n25031 );
and ( n25033 , n25028 , n25032 );
and ( n25034 , n25025 , n25027 );
or ( n25035 , n25033 , n25034 );
nor ( n25036 , n25023 , n25035 );
xor ( n25037 , n24960 , n24962 );
xor ( n25038 , n25037 , n24988 );
xor ( n25039 , n25005 , n25007 );
and ( n25040 , n25039 , n25022 );
and ( n25041 , n25005 , n25007 );
or ( n25042 , n25040 , n25041 );
nor ( n25043 , n25038 , n25042 );
xor ( n25044 , n25025 , n25027 );
xor ( n25045 , n25044 , n25032 );
xor ( n25046 , n17937 , n17963 );
and ( n25047 , n25046 , n17968 );
and ( n25048 , n17937 , n17963 );
or ( n25049 , n25047 , n25048 );
nor ( n25050 , n25045 , n25049 );
nor ( n25051 , n25036 , n25043 , n25050 );
nand ( n25052 , n24993 , n25051 );
xor ( n25053 , n24780 , n24883 );
and ( n25054 , n25053 , n24956 );
and ( n25055 , n24780 , n24883 );
or ( n25056 , n25054 , n25055 );
not ( n25057 , n25056 );
xor ( n25058 , n24849 , n24876 );
and ( n25059 , n25058 , n24881 );
and ( n25060 , n24849 , n24876 );
or ( n25061 , n25059 , n25060 );
xor ( n25062 , n24811 , n24827 );
and ( n25063 , n25062 , n24846 );
and ( n25064 , n24811 , n24827 );
or ( n25065 , n25063 , n25064 );
not ( n25066 , n5697 );
not ( n25067 , n537 );
not ( n25068 , n24840 );
or ( n25069 , n25067 , n25068 );
nand ( n25070 , n24839 , n5605 );
nand ( n25071 , n25069 , n25070 );
not ( n25072 , n25071 );
or ( n25073 , n25066 , n25072 );
nand ( n25074 , n24786 , n16173 );
nand ( n25075 , n25073 , n25074 );
not ( n25076 , n24745 );
nor ( n25077 , n25076 , n5605 );
xor ( n25078 , n25075 , n25077 );
not ( n25079 , n4671 );
not ( n25080 , n24825 );
or ( n25081 , n25079 , n25080 );
nand ( n25082 , n25081 , n7610 );
xor ( n25083 , n25078 , n25082 );
xor ( n25084 , n25065 , n25083 );
not ( n25085 , n4660 );
and ( n25086 , n24903 , n4477 );
not ( n25087 , n24903 );
and ( n25088 , n25087 , n539 );
or ( n25089 , n25086 , n25088 );
not ( n25090 , n25089 );
or ( n25091 , n25085 , n25090 );
nand ( n25092 , n24835 , n4450 );
nand ( n25093 , n25091 , n25092 );
not ( n25094 , n5786 );
nand ( n25095 , n541 , n9887 );
nand ( n25096 , n9886 , n5734 );
nand ( n25097 , n25095 , n25096 );
not ( n25098 , n25097 );
or ( n25099 , n25094 , n25098 );
nand ( n25100 , n10067 , n24802 );
nand ( n25101 , n25099 , n25100 );
not ( n25102 , n25101 );
xor ( n25103 , n25093 , n25102 );
xor ( n25104 , n24795 , n24806 );
and ( n25105 , n25104 , n24808 );
and ( n25106 , n24795 , n24806 );
or ( n25107 , n25105 , n25106 );
xor ( n25108 , n25103 , n25107 );
xor ( n25109 , n25084 , n25108 );
xor ( n25110 , n25061 , n25109 );
xor ( n25111 , n24809 , n24847 );
and ( n25112 , n25111 , n24882 );
and ( n25113 , n24809 , n24847 );
or ( n25114 , n25112 , n25113 );
xor ( n25115 , n25110 , n25114 );
not ( n25116 , n25115 );
nand ( n25117 , n25057 , n25116 );
xor ( n25118 , n25061 , n25109 );
and ( n25119 , n25118 , n25114 );
and ( n25120 , n25061 , n25109 );
or ( n25121 , n25119 , n25120 );
xor ( n25122 , n25093 , n25102 );
and ( n25123 , n25122 , n25107 );
and ( n25124 , n25093 , n25102 );
or ( n25125 , n25123 , n25124 );
xor ( n25126 , n25075 , n25077 );
and ( n25127 , n25126 , n25082 );
and ( n25128 , n25075 , n25077 );
or ( n25129 , n25127 , n25128 );
or ( n25130 , n4671 , n9730 );
nand ( n25131 , n25130 , n543 );
not ( n25132 , n10067 );
not ( n25133 , n25097 );
or ( n25134 , n25132 , n25133 );
not ( n25135 , n541 );
not ( n25136 , n9977 );
or ( n25137 , n25135 , n25136 );
nand ( n25138 , n24823 , n5734 );
nand ( n25139 , n25137 , n25138 );
nand ( n25140 , n25139 , n5786 );
nand ( n25141 , n25134 , n25140 );
xor ( n25142 , n25131 , n25141 );
not ( n25143 , n5697 );
not ( n25144 , n537 );
not ( n25145 , n9867 );
or ( n25146 , n25144 , n25145 );
nand ( n25147 , n24833 , n5605 );
nand ( n25148 , n25146 , n25147 );
not ( n25149 , n25148 );
or ( n25150 , n25143 , n25149 );
nand ( n25151 , n25071 , n16173 );
nand ( n25152 , n25150 , n25151 );
xor ( n25153 , n25142 , n25152 );
xor ( n25154 , n25129 , n25153 );
and ( n25155 , n24739 , n537 );
not ( n25156 , n4660 );
not ( n25157 , n539 );
not ( n25158 , n9692 );
or ( n25159 , n25157 , n25158 );
nand ( n25160 , n4477 , n24800 );
nand ( n25161 , n25159 , n25160 );
not ( n25162 , n25161 );
or ( n25163 , n25156 , n25162 );
nand ( n25164 , n25089 , n4450 );
nand ( n25165 , n25163 , n25164 );
xor ( n25166 , n25155 , n25165 );
xor ( n25167 , n25166 , n25101 );
xor ( n25168 , n25154 , n25167 );
xor ( n25169 , n25125 , n25168 );
xor ( n25170 , n25065 , n25083 );
and ( n25171 , n25170 , n25108 );
and ( n25172 , n25065 , n25083 );
or ( n25173 , n25171 , n25172 );
xor ( n25174 , n25169 , n25173 );
nor ( n25175 , n25121 , n25174 );
not ( n25176 , n25175 );
nand ( n25177 , n25117 , n25176 );
nor ( n25178 , n25052 , n25177 );
nand ( n25179 , n24691 , n25178 );
nand ( n25180 , n24957 , n24991 );
not ( n25181 , n25180 );
nand ( n25182 , n25042 , n25038 );
not ( n25183 , n25182 );
nand ( n25184 , n25045 , n25049 );
nor ( n25185 , n25023 , n25035 );
or ( n25186 , n25184 , n25185 );
nand ( n25187 , n25023 , n25035 );
nand ( n25188 , n25186 , n25187 );
not ( n25189 , n25042 );
not ( n25190 , n25038 );
nand ( n25191 , n25189 , n25190 );
nand ( n25192 , n25188 , n25191 );
not ( n25193 , n25192 );
or ( n25194 , n25183 , n25193 );
nand ( n25195 , n24958 , n24992 );
nand ( n25196 , n25194 , n25195 );
not ( n25197 , n25196 );
or ( n25198 , n25181 , n25197 );
not ( n25199 , n25177 );
nand ( n25200 , n25198 , n25199 );
nand ( n25201 , n25056 , n25115 );
nor ( n25202 , n25121 , n25174 );
or ( n25203 , n25201 , n25202 );
nand ( n25204 , n25121 , n25174 );
nand ( n25205 , n25203 , n25204 );
not ( n25206 , n25205 );
nand ( n25207 , n25179 , n25200 , n25206 );
xor ( n25208 , n25155 , n25165 );
and ( n25209 , n25208 , n25101 );
and ( n25210 , n25155 , n25165 );
or ( n25211 , n25209 , n25210 );
not ( n25212 , n7606 );
not ( n25213 , n5734 );
and ( n25214 , n25212 , n25213 );
and ( n25215 , n25139 , n10067 );
nor ( n25216 , n25214 , n25215 );
xor ( n25217 , n25131 , n25141 );
and ( n25218 , n25217 , n25152 );
and ( n25219 , n25131 , n25141 );
or ( n25220 , n25218 , n25219 );
xor ( n25221 , n25216 , n25220 );
and ( n25222 , n24839 , n537 );
not ( n25223 , n4660 );
not ( n25224 , n539 );
not ( n25225 , n9887 );
or ( n25226 , n25224 , n25225 );
nand ( n25227 , n4477 , n9886 );
nand ( n25228 , n25226 , n25227 );
not ( n25229 , n25228 );
or ( n25230 , n25223 , n25229 );
nand ( n25231 , n25161 , n4450 );
nand ( n25232 , n25230 , n25231 );
xor ( n25233 , n25222 , n25232 );
not ( n25234 , n16173 );
not ( n25235 , n25148 );
or ( n25236 , n25234 , n25235 );
xor ( n25237 , n537 , n24903 );
nand ( n25238 , n25237 , n5697 );
nand ( n25239 , n25236 , n25238 );
xor ( n25240 , n25233 , n25239 );
xor ( n25241 , n25221 , n25240 );
xor ( n25242 , n25211 , n25241 );
xor ( n25243 , n25129 , n25153 );
and ( n25244 , n25243 , n25167 );
and ( n25245 , n25129 , n25153 );
or ( n25246 , n25244 , n25245 );
xor ( n25247 , n25242 , n25246 );
xor ( n25248 , n25125 , n25168 );
and ( n25249 , n25248 , n25173 );
and ( n25250 , n25125 , n25168 );
or ( n25251 , n25249 , n25250 );
or ( n25252 , n25247 , n25251 );
nand ( n25253 , n25251 , n25247 );
nand ( n25254 , n25252 , n25253 );
not ( n25255 , n25254 );
and ( n25256 , n25207 , n25255 );
not ( n25257 , n25207 );
and ( n25258 , n25257 , n25254 );
nor ( n25259 , n25256 , n25258 );
nand ( n25260 , n25259 , n454 );
nand ( n25261 , n24675 , n25260 );
and ( n25262 , n25261 , n472 );
not ( n25263 , n10190 );
buf ( n25264 , n24579 );
nand ( n25265 , n24452 , n24492 );
not ( n25266 , n25265 );
nor ( n25267 , n25266 , n24493 );
and ( n25268 , n25264 , n25267 );
not ( n25269 , n25264 );
not ( n25270 , n25267 );
and ( n25271 , n25269 , n25270 );
nor ( n25272 , n25268 , n25271 );
not ( n25273 , n25272 );
or ( n25274 , n25263 , n25273 );
and ( n25275 , n25195 , n25180 );
not ( n25276 , n25275 );
buf ( n25277 , n25051 );
not ( n25278 , n25277 );
not ( n25279 , n24683 );
nand ( n25280 , n25279 , n24690 );
not ( n25281 , n25280 );
or ( n25282 , n25278 , n25281 );
nand ( n25283 , n25277 , n24684 );
buf ( n25284 , n25192 );
nand ( n25285 , n25283 , n25284 , n25182 );
not ( n25286 , n25285 );
nand ( n25287 , n25282 , n25286 );
not ( n25288 , n25287 );
or ( n25289 , n25276 , n25288 );
nand ( n25290 , n25280 , n25277 );
nor ( n25291 , n25285 , n25275 );
and ( n25292 , n25290 , n25291 );
not ( n25293 , n454 );
nor ( n25294 , n25292 , n25293 );
nand ( n25295 , n25289 , n25294 );
nand ( n25296 , n25274 , n25295 );
and ( n25297 , n25296 , n470 );
nor ( n25298 , n24683 , n24684 );
not ( n25299 , n25298 );
not ( n25300 , n24690 );
or ( n25301 , n25299 , n25300 );
buf ( n25302 , n25050 );
not ( n25303 , n25302 );
nand ( n25304 , n25301 , n25303 );
buf ( n25305 , n25185 );
or ( n25306 , n25304 , n25305 );
buf ( n25307 , n25188 );
not ( n25308 , n25307 );
and ( n25309 , n25042 , n25190 );
not ( n25310 , n25042 );
and ( n25311 , n25310 , n25038 );
nor ( n25312 , n25309 , n25311 );
not ( n25313 , n25312 );
and ( n25314 , n25308 , n25313 );
nand ( n25315 , n25306 , n25314 );
not ( n25316 , n25315 );
not ( n25317 , n25304 );
not ( n25318 , n25305 );
nand ( n25319 , n25318 , n25312 );
not ( n25320 , n25319 );
and ( n25321 , n25317 , n25320 );
nor ( n25322 , n25308 , n25313 );
nor ( n25323 , n25321 , n25322 );
not ( n25324 , n25323 );
or ( n25325 , n25316 , n25324 );
nand ( n25326 , n25325 , n454 );
not ( n25327 , n24561 );
or ( n25328 , n24506 , n24526 );
nand ( n25329 , n25328 , n17840 );
buf ( n25330 , n24506 );
nand ( n25331 , n25330 , n24526 );
and ( n25332 , n25329 , n25331 );
nand ( n25333 , n25327 , n25332 );
not ( n25334 , n25333 );
and ( n25335 , n24553 , n24570 );
not ( n25336 , n25335 );
nand ( n25337 , n17706 , n17710 );
nor ( n25338 , n25336 , n25337 );
nand ( n25339 , n25334 , n25338 );
buf ( n25340 , n24568 );
not ( n25341 , n25340 );
nor ( n25342 , n25341 , n25332 );
not ( n25343 , n25327 );
or ( n25344 , n25342 , n25343 );
nand ( n25345 , n25344 , n25336 );
not ( n25346 , n17843 );
not ( n25347 , n25328 );
nor ( n25348 , n25346 , n25347 );
nor ( n25349 , n25348 , n25333 );
not ( n25350 , n25327 );
nor ( n25351 , n25350 , n25340 );
or ( n25352 , n25349 , n25351 );
nand ( n25353 , n25352 , n25335 );
nand ( n25354 , n25339 , n25345 , n25353 );
nand ( n25355 , n17706 , n17710 );
and ( n25356 , n25336 , n25355 , n25348 , n25340 );
or ( n25357 , n25354 , n25356 );
nand ( n25358 , n25357 , n10190 );
and ( n25359 , n25326 , n25358 );
nor ( n25360 , n25359 , n16080 );
xor ( n25361 , n25297 , n25360 );
not ( n25362 , n10190 );
nand ( n25363 , n24364 , n24591 );
xnor ( n25364 , n24588 , n25363 );
not ( n25365 , n25364 );
or ( n25366 , n25362 , n25365 );
not ( n25367 , n25298 );
not ( n25368 , n24690 );
or ( n25369 , n25367 , n25368 );
not ( n25370 , n25056 );
nand ( n25371 , n25370 , n25116 );
buf ( n25372 , n25371 );
not ( n25373 , n25372 );
nor ( n25374 , n25373 , n25052 );
nand ( n25375 , n25369 , n25374 );
xnor ( n25376 , n25121 , n25174 );
and ( n25377 , n25376 , n454 );
or ( n25378 , n25375 , n25377 );
not ( n25379 , n25180 );
not ( n25380 , n25196 );
or ( n25381 , n25379 , n25380 );
nand ( n25382 , n25381 , n25372 );
not ( n25383 , n25382 );
not ( n25384 , n25377 );
and ( n25385 , n25383 , n25384 );
not ( n25386 , n25377 );
not ( n25387 , n25201 );
and ( n25388 , n25386 , n25387 );
nor ( n25389 , n25385 , n25388 );
not ( n25390 , n25376 );
and ( n25391 , n25390 , n454 );
nor ( n25392 , n25391 , n25387 );
nand ( n25393 , n25375 , n25382 , n25392 );
nand ( n25394 , n25378 , n25389 , n25393 );
nand ( n25395 , n25366 , n25394 );
and ( n25396 , n25395 , n472 );
and ( n25397 , n25361 , n25396 );
and ( n25398 , n25297 , n25360 );
or ( n25399 , n25397 , n25398 );
xor ( n25400 , n25262 , n25399 );
not ( n25401 , n10190 );
not ( n25402 , n25272 );
or ( n25403 , n25401 , n25402 );
nand ( n25404 , n25403 , n25295 );
and ( n25405 , n25404 , n469 );
and ( n25406 , n25395 , n471 );
xor ( n25407 , n25405 , n25406 );
not ( n25408 , n454 );
not ( n25409 , n25052 );
not ( n25410 , n25409 );
not ( n25411 , n24691 );
or ( n25412 , n25410 , n25411 );
and ( n25413 , n25196 , n25180 );
nand ( n25414 , n25412 , n25413 );
nand ( n25415 , n25372 , n25201 );
not ( n25416 , n25415 );
and ( n25417 , n25414 , n25416 );
not ( n25418 , n25414 );
and ( n25419 , n25418 , n25415 );
nor ( n25420 , n25417 , n25419 );
not ( n25421 , n25420 );
or ( n25422 , n25408 , n25421 );
not ( n25423 , n24493 );
not ( n25424 , n25423 );
not ( n25425 , n25264 );
or ( n25426 , n25424 , n25425 );
nand ( n25427 , n25426 , n25265 );
not ( n25428 , n24500 );
nand ( n25429 , n25428 , n24585 );
not ( n25430 , n25429 );
and ( n25431 , n25427 , n25430 );
not ( n25432 , n25427 );
and ( n25433 , n25432 , n25429 );
nor ( n25434 , n25431 , n25433 );
nand ( n25435 , n25434 , n10190 );
nand ( n25436 , n25422 , n25435 );
and ( n25437 , n25436 , n470 );
xor ( n25438 , n25407 , n25437 );
xor ( n25439 , n25400 , n25438 );
not ( n25440 , n25439 );
buf ( n25441 , n25436 );
and ( n25442 , n25441 , n471 );
and ( n25443 , n25404 , n471 );
not ( n25444 , n10190 );
not ( n25445 , n25348 );
not ( n25446 , n25355 );
or ( n25447 , n25445 , n25446 );
buf ( n25448 , n25332 );
nand ( n25449 , n25447 , n25448 );
and ( n25450 , n25340 , n25327 );
xor ( n25451 , n25449 , n25450 );
not ( n25452 , n25451 );
or ( n25453 , n25444 , n25452 );
buf ( n25454 , n25184 );
and ( n25455 , n25304 , n25454 );
not ( n25456 , n25305 );
buf ( n25457 , n25187 );
nand ( n25458 , n25456 , n25457 );
and ( n25459 , n25458 , n454 );
or ( n25460 , n25455 , n25459 );
not ( n25461 , n25458 );
nand ( n25462 , n25461 , n454 );
nand ( n25463 , n25462 , n25304 , n25454 );
nand ( n25464 , n25460 , n25463 );
nand ( n25465 , n25453 , n25464 );
not ( n25466 , n25465 );
nor ( n25467 , n25466 , n16080 );
xor ( n25468 , n25443 , n25467 );
nand ( n25469 , n25358 , n25326 );
not ( n25470 , n25469 );
nor ( n25471 , n25470 , n2635 );
and ( n25472 , n25468 , n25471 );
and ( n25473 , n25443 , n25467 );
or ( n25474 , n25472 , n25473 );
xor ( n25475 , n25442 , n25474 );
xor ( n25476 , n25297 , n25360 );
xor ( n25477 , n25476 , n25396 );
and ( n25478 , n25475 , n25477 );
and ( n25479 , n25442 , n25474 );
or ( n25480 , n25478 , n25479 );
not ( n25481 , n25480 );
and ( n25482 , n25440 , n25481 );
and ( n25483 , n25441 , n472 );
and ( n25484 , n25296 , n472 );
not ( n25485 , n10190 );
not ( n25486 , n17844 );
not ( n25487 , n25355 );
or ( n25488 , n25486 , n25487 );
nand ( n25489 , n25488 , n17841 );
not ( n25490 , n25331 );
nor ( n25491 , n25490 , n25347 );
xor ( n25492 , n25489 , n25491 );
not ( n25493 , n25492 );
or ( n25494 , n25485 , n25493 );
nand ( n25495 , n25303 , n25184 );
xnor ( n25496 , n24691 , n25495 );
nand ( n25497 , n25496 , n454 );
nand ( n25498 , n25494 , n25497 );
and ( n25499 , n25498 , n469 );
xor ( n25500 , n25484 , n25499 );
and ( n25501 , n25465 , n470 );
and ( n25502 , n25500 , n25501 );
and ( n25503 , n25484 , n25499 );
or ( n25504 , n25502 , n25503 );
xor ( n25505 , n25483 , n25504 );
xor ( n25506 , n25443 , n25467 );
xor ( n25507 , n25506 , n25471 );
and ( n25508 , n25505 , n25507 );
and ( n25509 , n25483 , n25504 );
or ( n25510 , n25508 , n25509 );
not ( n25511 , n25510 );
xor ( n25512 , n25442 , n25474 );
xor ( n25513 , n25512 , n25477 );
not ( n25514 , n25513 );
and ( n25515 , n25511 , n25514 );
nor ( n25516 , n25482 , n25515 );
buf ( n25517 , n25516 );
not ( n25518 , n25517 );
xor ( n25519 , n25483 , n25504 );
xor ( n25520 , n25519 , n25507 );
not ( n25521 , n25520 );
not ( n25522 , n25470 );
and ( n25523 , n25522 , n471 );
not ( n25524 , n454 );
not ( n25525 , n17983 );
or ( n25526 , n25524 , n25525 );
and ( n25527 , n25337 , n17846 );
not ( n25528 , n25337 );
and ( n25529 , n25528 , n17845 );
nor ( n25530 , n25527 , n25529 );
nand ( n25531 , n25530 , n10190 );
nand ( n25532 , n25526 , n25531 );
and ( n25533 , n25532 , n469 );
nor ( n25534 , n25466 , n17257 );
xor ( n25535 , n25533 , n25534 );
and ( n25536 , n25498 , n470 );
and ( n25537 , n25535 , n25536 );
and ( n25538 , n25533 , n25534 );
or ( n25539 , n25537 , n25538 );
xor ( n25540 , n25523 , n25539 );
xor ( n25541 , n25484 , n25499 );
xor ( n25542 , n25541 , n25501 );
and ( n25543 , n25540 , n25542 );
and ( n25544 , n25523 , n25539 );
or ( n25545 , n25543 , n25544 );
not ( n25546 , n25545 );
nand ( n25547 , n25521 , n25546 );
not ( n25548 , n25547 );
xor ( n25549 , n25523 , n25539 );
xor ( n25550 , n25549 , n25542 );
and ( n25551 , n25522 , n472 );
and ( n25552 , n25532 , n470 );
and ( n25553 , n16710 , n469 );
xor ( n25554 , n25552 , n25553 );
and ( n25555 , n25465 , n472 );
and ( n25556 , n25554 , n25555 );
and ( n25557 , n25552 , n25553 );
or ( n25558 , n25556 , n25557 );
xor ( n25559 , n25551 , n25558 );
xor ( n25560 , n25533 , n25534 );
xor ( n25561 , n25560 , n25536 );
and ( n25562 , n25559 , n25561 );
and ( n25563 , n25551 , n25558 );
or ( n25564 , n25562 , n25563 );
nor ( n25565 , n25550 , n25564 );
xor ( n25566 , n25551 , n25558 );
xor ( n25567 , n25566 , n25561 );
and ( n25568 , n25498 , n471 );
and ( n25569 , n17984 , n17851 );
not ( n25570 , n471 );
nor ( n25571 , n25569 , n25570 );
and ( n25572 , n16393 , n469 );
xor ( n25573 , n25571 , n25572 );
and ( n25574 , n16710 , n470 );
and ( n25575 , n25573 , n25574 );
and ( n25576 , n25571 , n25572 );
or ( n25577 , n25575 , n25576 );
xor ( n25578 , n25568 , n25577 );
xor ( n25579 , n25552 , n25553 );
xor ( n25580 , n25579 , n25555 );
and ( n25581 , n25578 , n25580 );
and ( n25582 , n25568 , n25577 );
or ( n25583 , n25581 , n25582 );
nand ( n25584 , n25567 , n25583 );
or ( n25585 , n25565 , n25584 );
nand ( n25586 , n25550 , n25564 );
nand ( n25587 , n25585 , n25586 );
not ( n25588 , n25587 );
or ( n25589 , n25548 , n25588 );
buf ( n25590 , n25520 );
nand ( n25591 , n25590 , n25545 );
nand ( n25592 , n25589 , n25591 );
not ( n25593 , n25592 );
not ( n25594 , n17691 );
not ( n25595 , n17681 );
nand ( n25596 , n17478 , n17495 );
nand ( n25597 , n17625 , n17590 , n25596 );
nand ( n25598 , n17589 , n25597 , n17592 , n17594 );
nand ( n25599 , n25598 , n17670 , n17647 );
not ( n25600 , n25599 );
or ( n25601 , n25595 , n25600 );
nand ( n25602 , n25601 , n16772 );
not ( n25603 , n25602 );
or ( n25604 , n25594 , n25603 );
and ( n25605 , n25498 , n472 );
xor ( n25606 , n17986 , n17987 );
and ( n25607 , n25606 , n17989 );
and ( n25608 , n17986 , n17987 );
or ( n25609 , n25607 , n25608 );
xor ( n25610 , n25605 , n25609 );
xor ( n25611 , n25571 , n25572 );
xor ( n25612 , n25611 , n25574 );
and ( n25613 , n25610 , n25612 );
and ( n25614 , n25605 , n25609 );
or ( n25615 , n25613 , n25614 );
not ( n25616 , n25615 );
not ( n25617 , n25616 );
xor ( n25618 , n25568 , n25577 );
xor ( n25619 , n25618 , n25580 );
not ( n25620 , n25619 );
not ( n25621 , n25620 );
or ( n25622 , n25617 , n25621 );
xor ( n25623 , n25605 , n25609 );
xor ( n25624 , n25623 , n25612 );
not ( n25625 , n25624 );
xor ( n25626 , n17693 , n17697 );
and ( n25627 , n25626 , n17990 );
and ( n25628 , n17693 , n17697 );
or ( n25629 , n25627 , n25628 );
not ( n25630 , n25629 );
and ( n25631 , n25625 , n25630 );
nor ( n25632 , n25631 , n17996 );
nand ( n25633 , n25622 , n25632 );
not ( n25634 , n25633 );
nand ( n25635 , n25604 , n25634 );
not ( n25636 , n25635 );
nor ( n25637 , n25624 , n25629 );
or ( n25638 , n25637 , n17999 );
nand ( n25639 , n25624 , n25629 );
nand ( n25640 , n25638 , n25639 );
nand ( n25641 , n25616 , n25620 );
and ( n25642 , n25640 , n25641 );
nand ( n25643 , n25619 , n25615 );
not ( n25644 , n25643 );
nor ( n25645 , n25642 , n25644 );
not ( n25646 , n25645 );
or ( n25647 , n25636 , n25646 );
not ( n25648 , n25550 );
not ( n25649 , n25564 );
nand ( n25650 , n25648 , n25649 );
not ( n25651 , n25567 );
not ( n25652 , n25583 );
nand ( n25653 , n25651 , n25652 );
and ( n25654 , n25650 , n25653 , n25547 );
nand ( n25655 , n25647 , n25654 );
nand ( n25656 , n25593 , n25655 );
not ( n25657 , n25656 );
or ( n25658 , n25518 , n25657 );
not ( n25659 , n25439 );
nand ( n25660 , n25659 , n25481 );
not ( n25661 , n25660 );
nand ( n25662 , n25510 , n25513 );
not ( n25663 , n25662 );
not ( n25664 , n25663 );
or ( n25665 , n25661 , n25664 );
nand ( n25666 , n25439 , n25480 );
nand ( n25667 , n25665 , n25666 );
buf ( n25668 , n25667 );
not ( n25669 , n25668 );
nand ( n25670 , n25658 , n25669 );
and ( n25671 , n25261 , n471 );
xor ( n25672 , n25405 , n25406 );
and ( n25673 , n25672 , n25437 );
and ( n25674 , n25405 , n25406 );
or ( n25675 , n25673 , n25674 );
xor ( n25676 , n25671 , n25675 );
nand ( n25677 , n24246 , n24363 );
and ( n25678 , n24501 , n25677 , n24665 );
not ( n25679 , n25678 );
not ( n25680 , n24579 );
or ( n25681 , n25679 , n25680 );
not ( n25682 , n24665 );
not ( n25683 , n25677 );
not ( n25684 , n24586 );
or ( n25685 , n25683 , n25684 );
nand ( n25686 , n25685 , n24591 );
not ( n25687 , n25686 );
or ( n25688 , n25682 , n25687 );
nand ( n25689 , n25688 , n24666 );
not ( n25690 , n25689 );
nand ( n25691 , n25681 , n25690 );
and ( n25692 , n489 , n15602 );
not ( n25693 , n25692 );
not ( n25694 , n13056 );
not ( n25695 , n24630 );
or ( n25696 , n25694 , n25695 );
nand ( n25697 , n13119 , n495 );
nand ( n25698 , n25696 , n25697 );
xor ( n25699 , n25693 , n25698 );
xor ( n25700 , n24643 , n24644 );
and ( n25701 , n25700 , n24655 );
and ( n25702 , n24643 , n24644 );
or ( n25703 , n25701 , n25702 );
xor ( n25704 , n25699 , n25703 );
xor ( n25705 , n24614 , n24624 );
and ( n25706 , n25705 , n24634 );
and ( n25707 , n24614 , n24624 );
or ( n25708 , n25706 , n25707 );
not ( n25709 , n12731 );
and ( n25710 , n15726 , n12703 );
not ( n25711 , n15726 );
and ( n25712 , n25711 , n491 );
or ( n25713 , n25710 , n25712 );
not ( n25714 , n25713 );
or ( n25715 , n25709 , n25714 );
nand ( n25716 , n12688 , n24651 );
nand ( n25717 , n25715 , n25716 );
not ( n25718 , n12635 );
not ( n25719 , n24610 );
or ( n25720 , n25718 , n25719 );
xor ( n25721 , n489 , n17764 );
nand ( n25722 , n25721 , n12882 );
nand ( n25723 , n25720 , n25722 );
xor ( n25724 , n25717 , n25723 );
not ( n25725 , n12845 );
not ( n25726 , n493 );
not ( n25727 , n16336 );
not ( n25728 , n25727 );
or ( n25729 , n25726 , n25728 );
nand ( n25730 , n16336 , n12862 );
nand ( n25731 , n25729 , n25730 );
not ( n25732 , n25731 );
or ( n25733 , n25725 , n25732 );
nand ( n25734 , n24622 , n15386 );
nand ( n25735 , n25733 , n25734 );
xor ( n25736 , n25724 , n25735 );
xor ( n25737 , n25708 , n25736 );
xor ( n25738 , n24058 , n24640 );
and ( n25739 , n25738 , n24656 );
and ( n25740 , n24058 , n24640 );
or ( n25741 , n25739 , n25740 );
xor ( n25742 , n25737 , n25741 );
xor ( n25743 , n25704 , n25742 );
xor ( n25744 , n24604 , n24635 );
and ( n25745 , n25744 , n24657 );
and ( n25746 , n24604 , n24635 );
or ( n25747 , n25745 , n25746 );
xor ( n25748 , n25743 , n25747 );
not ( n25749 , n25748 );
xor ( n25750 , n24600 , n24658 );
and ( n25751 , n25750 , n24663 );
and ( n25752 , n24600 , n24658 );
or ( n25753 , n25751 , n25752 );
not ( n25754 , n25753 );
nand ( n25755 , n25749 , n25754 );
buf ( n25756 , n25755 );
and ( n25757 , n25753 , n25748 );
not ( n25758 , n25757 );
nand ( n25759 , n25756 , n25758 );
not ( n25760 , n25759 );
and ( n25761 , n25691 , n25760 );
not ( n25762 , n25691 );
and ( n25763 , n25762 , n25759 );
nor ( n25764 , n25761 , n25763 );
nand ( n25765 , n25764 , n10190 );
not ( n25766 , n25765 );
not ( n25767 , n25252 );
not ( n25768 , n25205 );
or ( n25769 , n25767 , n25768 );
nand ( n25770 , n25769 , n25253 );
not ( n25771 , n25770 );
not ( n25772 , n25771 );
or ( n25773 , n25280 , n24684 );
or ( n25774 , n25247 , n25251 );
nand ( n25775 , n25371 , n25176 , n25774 );
nor ( n25776 , n25775 , n25052 );
nand ( n25777 , n25773 , n25776 );
not ( n25778 , n25777 );
or ( n25779 , n25772 , n25778 );
or ( n25780 , n10067 , n5786 );
nand ( n25781 , n25780 , n541 );
not ( n25782 , n4450 );
not ( n25783 , n25228 );
or ( n25784 , n25782 , n25783 );
not ( n25785 , n539 );
not ( n25786 , n9977 );
or ( n25787 , n25785 , n25786 );
not ( n25788 , n9977 );
nand ( n25789 , n25788 , n4477 );
nand ( n25790 , n25787 , n25789 );
nand ( n25791 , n25790 , n4660 );
nand ( n25792 , n25784 , n25791 );
xor ( n25793 , n25781 , n25792 );
nor ( n25794 , n9867 , n5605 );
xor ( n25795 , n25793 , n25794 );
not ( n25796 , n5697 );
xor ( n25797 , n24800 , n537 );
not ( n25798 , n25797 );
or ( n25799 , n25796 , n25798 );
nand ( n25800 , n25237 , n16173 );
nand ( n25801 , n25799 , n25800 );
not ( n25802 , n25216 );
xor ( n25803 , n25801 , n25802 );
xor ( n25804 , n25222 , n25232 );
and ( n25805 , n25804 , n25239 );
and ( n25806 , n25222 , n25232 );
or ( n25807 , n25805 , n25806 );
xor ( n25808 , n25803 , n25807 );
xor ( n25809 , n25795 , n25808 );
xor ( n25810 , n25216 , n25220 );
and ( n25811 , n25810 , n25240 );
and ( n25812 , n25216 , n25220 );
or ( n25813 , n25811 , n25812 );
xor ( n25814 , n25809 , n25813 );
xor ( n25815 , n25211 , n25241 );
and ( n25816 , n25815 , n25246 );
and ( n25817 , n25211 , n25241 );
or ( n25818 , n25816 , n25817 );
and ( n25819 , n25814 , n25818 );
not ( n25820 , n25819 );
nor ( n25821 , n25818 , n25814 );
not ( n25822 , n25821 );
and ( n25823 , n25820 , n25822 );
nand ( n25824 , n25779 , n25823 );
not ( n25825 , n25180 );
not ( n25826 , n25196 );
or ( n25827 , n25825 , n25826 );
not ( n25828 , n25775 );
nand ( n25829 , n25827 , n25828 );
not ( n25830 , n25823 );
or ( n25831 , n25829 , n25830 );
nand ( n25832 , n25831 , n454 );
not ( n25833 , n25832 );
nor ( n25834 , n25770 , n25823 );
nand ( n25835 , n25777 , n25829 , n25834 );
nand ( n25836 , n25824 , n25833 , n25835 );
not ( n25837 , n25836 );
or ( n25838 , n25766 , n25837 );
nand ( n25839 , n25838 , n472 );
not ( n25840 , n25839 );
and ( n25841 , n25436 , n469 );
xor ( n25842 , n25840 , n25841 );
and ( n25843 , n25395 , n470 );
xor ( n25844 , n25842 , n25843 );
xor ( n25845 , n25676 , n25844 );
xor ( n25846 , n25262 , n25399 );
and ( n25847 , n25846 , n25438 );
and ( n25848 , n25262 , n25399 );
or ( n25849 , n25847 , n25848 );
or ( n25850 , n25845 , n25849 );
nand ( n25851 , n25845 , n25849 );
nand ( n25852 , n25850 , n25851 );
and ( n25853 , n25670 , n25852 );
nand ( n25854 , n25656 , n25517 );
nor ( n25855 , n25852 , n25668 );
and ( n25856 , n25854 , n25855 );
nor ( n25857 , n25853 , n25856 );
or ( n25858 , n25857 , n18007 );
not ( n25859 , n20693 );
not ( n25860 , n20878 );
or ( n25861 , n25859 , n25860 );
nand ( n25862 , n21013 , n21045 );
nand ( n25863 , n25861 , n25862 );
not ( n25864 , n25863 );
not ( n25865 , n20647 );
not ( n25866 , n20628 );
not ( n25867 , n21138 );
or ( n25868 , n25866 , n25867 );
nand ( n25869 , n21137 , n20644 );
nand ( n25870 , n25868 , n25869 );
not ( n25871 , n25870 );
or ( n25872 , n25865 , n25871 );
not ( n25873 , n20628 );
not ( n25874 , n21196 );
or ( n25875 , n25873 , n25874 );
nand ( n25876 , n21193 , n20644 );
nand ( n25877 , n25875 , n25876 );
nand ( n25878 , n25877 , n20602 );
nand ( n25879 , n25872 , n25878 );
xor ( n25880 , n25864 , n25879 );
not ( n25881 , n20728 );
not ( n25882 , n20730 );
not ( n25883 , n21181 );
or ( n25884 , n25882 , n25883 );
nand ( n25885 , n21178 , n20745 );
nand ( n25886 , n25884 , n25885 );
not ( n25887 , n25886 );
or ( n25888 , n25881 , n25887 );
not ( n25889 , n20730 );
not ( n25890 , n20900 );
or ( n25891 , n25889 , n25890 );
nand ( n25892 , n20899 , n20745 );
nand ( n25893 , n25891 , n25892 );
nand ( n25894 , n25893 , n20765 );
nand ( n25895 , n25888 , n25894 );
xor ( n25896 , n25880 , n25895 );
not ( n25897 , n21163 );
not ( n25898 , n21167 );
not ( n25899 , n20458 );
or ( n25900 , n18039 , n18149 );
nand ( n25901 , n25900 , n18041 );
or ( n25902 , n20451 , n18241 );
and ( n25903 , n18180 , n18245 );
and ( n25904 , n18438 , n18244 );
nor ( n25905 , n25903 , n25904 );
or ( n25906 , n25905 , n18289 );
nand ( n25907 , n25902 , n25906 );
xor ( n25908 , n25901 , n25907 );
nor ( n25909 , n18321 , n18244 );
xor ( n25910 , n25908 , n25909 );
xor ( n25911 , n25899 , n25910 );
xor ( n25912 , n20453 , n20454 );
and ( n25913 , n25912 , n20458 );
and ( n25914 , n20453 , n20454 );
or ( n25915 , n25913 , n25914 );
and ( n25916 , n25911 , n25915 );
and ( n25917 , n25899 , n25910 );
or ( n25918 , n25916 , n25917 );
nor ( n25919 , n18417 , n18244 );
not ( n25920 , n25905 );
and ( n25921 , n25920 , n18242 );
and ( n25922 , n18290 , n18245 );
nor ( n25923 , n25921 , n25922 );
xor ( n25924 , n25919 , n25923 );
xor ( n25925 , n25901 , n25907 );
and ( n25926 , n25925 , n25909 );
and ( n25927 , n25901 , n25907 );
or ( n25928 , n25926 , n25927 );
xor ( n25929 , n25924 , n25928 );
or ( n25930 , n25918 , n25929 );
nand ( n25931 , n25918 , n25929 );
nand ( n25932 , n25930 , n25931 );
not ( n25933 , n25932 );
not ( n25934 , n25933 );
nand ( n25935 , n20466 , n20415 );
nor ( n25936 , n18644 , n25935 );
nand ( n25937 , n18599 , n25936 );
nor ( n25938 , n20358 , n25937 );
not ( n25939 , n25938 );
not ( n25940 , n20331 );
or ( n25941 , n25939 , n25940 );
or ( n25942 , n20367 , n18600 );
nand ( n25943 , n25942 , n20371 );
buf ( n25944 , n25936 );
and ( n25945 , n25943 , n25944 );
not ( n25946 , n20466 );
not ( n25947 , n20415 );
or ( n25948 , n20373 , n25947 );
nand ( n25949 , n25948 , n20416 );
not ( n25950 , n25949 );
or ( n25951 , n25946 , n25950 );
nand ( n25952 , n25951 , n20467 );
nor ( n25953 , n25945 , n25952 );
nand ( n25954 , n25941 , n25953 );
xor ( n25955 , n20445 , n20459 );
and ( n25956 , n25955 , n20464 );
and ( n25957 , n20445 , n20459 );
or ( n25958 , n25956 , n25957 );
xor ( n25959 , n25899 , n25910 );
xor ( n25960 , n25959 , n25915 );
or ( n25961 , n25958 , n25960 );
and ( n25962 , n25954 , n25961 );
and ( n25963 , n25958 , n25960 );
nor ( n25964 , n25962 , n25963 );
not ( n25965 , n25964 );
or ( n25966 , n25934 , n25965 );
not ( n25967 , n25964 );
nand ( n25968 , n25967 , n25932 );
nand ( n25969 , n25966 , n25968 );
not ( n25970 , n25969 );
not ( n25971 , n25970 );
or ( n25972 , n25898 , n25971 );
not ( n25973 , n25933 );
not ( n25974 , n25964 );
or ( n25975 , n25973 , n25974 );
nand ( n25976 , n25975 , n25968 );
nand ( n25977 , n25976 , n21166 );
nand ( n25978 , n25972 , n25977 );
not ( n25979 , n25978 );
or ( n25980 , n25897 , n25979 );
and ( n25981 , n25961 , n25930 );
not ( n25982 , n25981 );
not ( n25983 , n25954 );
or ( n25984 , n25982 , n25983 );
and ( n25985 , n25930 , n25963 );
not ( n25986 , n25931 );
nor ( n25987 , n25985 , n25986 );
nand ( n25988 , n25984 , n25987 );
xor ( n25989 , n25919 , n25923 );
and ( n25990 , n25989 , n25928 );
and ( n25991 , n25919 , n25923 );
or ( n25992 , n25990 , n25991 );
or ( n25993 , n18242 , n18290 );
nand ( n25994 , n25993 , n18245 );
nor ( n25995 , n18180 , n18244 );
xor ( n25996 , n25994 , n25995 );
not ( n25997 , n25923 );
xor ( n25998 , n25996 , n25997 );
xor ( n25999 , n25992 , n25998 );
xor ( n26000 , n25988 , n25999 );
buf ( n26001 , n26000 );
and ( n26002 , n21167 , n26001 );
not ( n26003 , n21167 );
not ( n26004 , n26000 );
and ( n26005 , n26003 , n26004 );
nor ( n26006 , n26002 , n26005 );
nand ( n26007 , n26006 , n21199 );
nand ( n26008 , n25980 , n26007 );
not ( n26009 , n21003 );
and ( n26010 , n20983 , n21394 );
not ( n26011 , n20983 );
and ( n26012 , n26011 , n21391 );
nor ( n26013 , n26010 , n26012 );
not ( n26014 , n26013 );
or ( n26015 , n26009 , n26014 );
and ( n26016 , n20983 , n20422 );
not ( n26017 , n20983 );
and ( n26018 , n26017 , n20425 );
nor ( n26019 , n26016 , n26018 );
nand ( n26020 , n26019 , n21334 );
nand ( n26021 , n26015 , n26020 );
xor ( n26022 , n26008 , n26021 );
not ( n26023 , n20905 );
not ( n26024 , n20863 );
not ( n26025 , n25963 );
nand ( n26026 , n26025 , n25961 );
and ( n26027 , n25954 , n26026 );
not ( n26028 , n25954 );
not ( n26029 , n26026 );
and ( n26030 , n26028 , n26029 );
or ( n26031 , n26027 , n26030 );
not ( n26032 , n26031 );
not ( n26033 , n26032 );
or ( n26034 , n26024 , n26033 );
nand ( n26035 , n26031 , n20862 );
nand ( n26036 , n26034 , n26035 );
not ( n26037 , n26036 );
or ( n26038 , n26023 , n26037 );
and ( n26039 , n21213 , n20474 );
not ( n26040 , n21213 );
and ( n26041 , n26040 , n20477 );
nor ( n26042 , n26039 , n26041 );
nand ( n26043 , n26042 , n20860 );
nand ( n26044 , n26038 , n26043 );
and ( n26045 , n26022 , n26044 );
and ( n26046 , n26008 , n26021 );
or ( n26047 , n26045 , n26046 );
xor ( n26048 , n25896 , n26047 );
not ( n26049 , n21167 );
not ( n26050 , n21199 );
or ( n26051 , n26049 , n26050 );
nand ( n26052 , n26006 , n21163 );
nand ( n26053 , n26051 , n26052 );
not ( n26054 , n21045 );
not ( n26055 , n20992 );
or ( n26056 , n26054 , n26055 );
nand ( n26057 , n21013 , n20693 );
nand ( n26058 , n26056 , n26057 );
or ( n26059 , n21148 , n21105 );
nand ( n26060 , n26059 , n21111 );
or ( n26061 , n26058 , n26060 );
not ( n26062 , n26061 );
not ( n26063 , n20728 );
not ( n26064 , n25893 );
or ( n26065 , n26063 , n26064 );
not ( n26066 , n20730 );
not ( n26067 , n20875 );
or ( n26068 , n26066 , n26067 );
nand ( n26069 , n20878 , n20745 );
nand ( n26070 , n26068 , n26069 );
nand ( n26071 , n26070 , n20765 );
nand ( n26072 , n26065 , n26071 );
not ( n26073 , n26072 );
or ( n26074 , n26062 , n26073 );
nand ( n26075 , n26058 , n26060 );
nand ( n26076 , n26074 , n26075 );
xor ( n26077 , n26053 , n26076 );
not ( n26078 , n20980 );
not ( n26079 , n20935 );
not ( n26080 , n21119 );
or ( n26081 , n26079 , n26080 );
nand ( n26082 , n21118 , n20953 );
nand ( n26083 , n26081 , n26082 );
not ( n26084 , n26083 );
or ( n26085 , n26078 , n26084 );
and ( n26086 , n20935 , n21394 );
not ( n26087 , n20935 );
and ( n26088 , n26087 , n21391 );
nor ( n26089 , n26086 , n26088 );
nand ( n26090 , n26089 , n20933 );
nand ( n26091 , n26085 , n26090 );
xor ( n26092 , n26077 , n26091 );
xor ( n26093 , n26048 , n26092 );
not ( n26094 , n21334 );
and ( n26095 , n20983 , n20474 );
not ( n26096 , n20983 );
and ( n26097 , n26096 , n20477 );
nor ( n26098 , n26095 , n26097 );
not ( n26099 , n26098 );
or ( n26100 , n26094 , n26099 );
nand ( n26101 , n26019 , n21003 );
nand ( n26102 , n26100 , n26101 );
not ( n26103 , n20905 );
and ( n26104 , n21213 , n25969 );
not ( n26105 , n21213 );
and ( n26106 , n26105 , n25970 );
nor ( n26107 , n26104 , n26106 );
not ( n26108 , n26107 );
or ( n26109 , n26103 , n26108 );
nand ( n26110 , n26036 , n20860 );
nand ( n26111 , n26109 , n26110 );
xor ( n26112 , n26102 , n26111 );
and ( n26113 , n20992 , n20693 );
and ( n26114 , n20945 , n21045 );
nor ( n26115 , n26113 , n26114 );
not ( n26116 , n26115 );
not ( n26117 , n20933 );
not ( n26118 , n26083 );
or ( n26119 , n26117 , n26118 );
not ( n26120 , n20935 );
not ( n26121 , n21138 );
or ( n26122 , n26120 , n26121 );
nand ( n26123 , n21137 , n20953 );
nand ( n26124 , n26122 , n26123 );
nand ( n26125 , n26124 , n20979 );
nand ( n26126 , n26119 , n26125 );
xor ( n26127 , n26116 , n26126 );
not ( n26128 , n20647 );
not ( n26129 , n25877 );
or ( n26130 , n26128 , n26129 );
not ( n26131 , n20628 );
not ( n26132 , n21181 );
or ( n26133 , n26131 , n26132 );
nand ( n26134 , n21178 , n20644 );
nand ( n26135 , n26133 , n26134 );
nand ( n26136 , n26135 , n20602 );
nand ( n26137 , n26130 , n26136 );
and ( n26138 , n26127 , n26137 );
and ( n26139 , n26116 , n26126 );
or ( n26140 , n26138 , n26139 );
xor ( n26141 , n26112 , n26140 );
and ( n26142 , n20945 , n20693 );
and ( n26143 , n20969 , n21045 );
nor ( n26144 , n26142 , n26143 );
and ( n26145 , n18024 , n22795 );
nor ( n26146 , n26145 , n18028 );
nand ( n26147 , n26144 , n26146 );
xor ( n26148 , n26147 , n26115 );
not ( n26149 , n20728 );
not ( n26150 , n26070 );
or ( n26151 , n26149 , n26150 );
not ( n26152 , n21006 );
not ( n26153 , n20745 );
and ( n26154 , n26152 , n26153 );
not ( n26155 , n26152 );
not ( n26156 , n20730 );
and ( n26157 , n26155 , n26156 );
or ( n26158 , n26154 , n26157 );
and ( n26159 , n21008 , n26158 );
not ( n26160 , n21008 );
not ( n26161 , n20745 );
and ( n26162 , n21006 , n26161 );
not ( n26163 , n21006 );
not ( n26164 , n20730 );
and ( n26165 , n26163 , n26164 );
or ( n26166 , n26162 , n26165 );
and ( n26167 , n26160 , n26166 );
or ( n26168 , n26159 , n26167 );
nand ( n26169 , n26168 , n20765 );
nand ( n26170 , n26151 , n26169 );
and ( n26171 , n26148 , n26170 );
and ( n26172 , n26147 , n26115 );
or ( n26173 , n26171 , n26172 );
xor ( n26174 , n26058 , n26060 );
xor ( n26175 , n26072 , n26174 );
xor ( n26176 , n26173 , n26175 );
xor ( n26177 , n26116 , n26126 );
xor ( n26178 , n26177 , n26137 );
and ( n26179 , n26176 , n26178 );
and ( n26180 , n26173 , n26175 );
or ( n26181 , n26179 , n26180 );
xor ( n26182 , n26141 , n26181 );
not ( n26183 , n20933 );
not ( n26184 , n26124 );
or ( n26185 , n26183 , n26184 );
and ( n26186 , n21192 , n20935 );
not ( n26187 , n21192 );
and ( n26188 , n26187 , n20953 );
nor ( n26189 , n26186 , n26188 );
nand ( n26190 , n26189 , n20980 );
nand ( n26191 , n26185 , n26190 );
not ( n26192 , n20647 );
not ( n26193 , n26135 );
or ( n26194 , n26192 , n26193 );
not ( n26195 , n20628 );
not ( n26196 , n20900 );
or ( n26197 , n26195 , n26196 );
nand ( n26198 , n20899 , n20644 );
nand ( n26199 , n26197 , n26198 );
nand ( n26200 , n26199 , n20602 );
nand ( n26201 , n26194 , n26200 );
xor ( n26202 , n26191 , n26201 );
not ( n26203 , n21003 );
not ( n26204 , n20983 );
not ( n26205 , n21119 );
or ( n26206 , n26204 , n26205 );
nand ( n26207 , n21118 , n21487 );
nand ( n26208 , n26206 , n26207 );
not ( n26209 , n26208 );
or ( n26210 , n26203 , n26209 );
nand ( n26211 , n26013 , n21334 );
nand ( n26212 , n26210 , n26211 );
and ( n26213 , n26202 , n26212 );
and ( n26214 , n26191 , n26201 );
or ( n26215 , n26213 , n26214 );
or ( n26216 , n26144 , n26146 );
nand ( n26217 , n26216 , n26147 );
not ( n26218 , n20765 );
not ( n26219 , n20730 );
not ( n26220 , n20995 );
or ( n26221 , n26219 , n26220 );
nand ( n26222 , n20992 , n20745 );
nand ( n26223 , n26221 , n26222 );
not ( n26224 , n26223 );
or ( n26225 , n26218 , n26224 );
nand ( n26226 , n26168 , n20728 );
nand ( n26227 , n26225 , n26226 );
xor ( n26228 , n26217 , n26227 );
not ( n26229 , n20602 );
not ( n26230 , n20609 );
not ( n26231 , n20875 );
or ( n26232 , n26230 , n26231 );
or ( n26233 , n20875 , n20609 );
nand ( n26234 , n26232 , n26233 );
not ( n26235 , n26234 );
or ( n26236 , n26229 , n26235 );
nand ( n26237 , n26199 , n20647 );
nand ( n26238 , n26236 , n26237 );
and ( n26239 , n26228 , n26238 );
and ( n26240 , n26217 , n26227 );
or ( n26241 , n26239 , n26240 );
not ( n26242 , n21148 );
not ( n26243 , n21111 );
not ( n26244 , n26004 );
or ( n26245 , n26243 , n26244 );
nand ( n26246 , n26001 , n21124 );
nand ( n26247 , n26245 , n26246 );
not ( n26248 , n26247 );
or ( n26249 , n26242 , n26248 );
nand ( n26250 , n21105 , n21111 );
nand ( n26251 , n26249 , n26250 );
xor ( n26252 , n26241 , n26251 );
and ( n26253 , n21167 , n26031 );
not ( n26254 , n21167 );
and ( n26255 , n26254 , n26032 );
nor ( n26256 , n26253 , n26255 );
not ( n26257 , n26256 );
not ( n26258 , n21163 );
or ( n26259 , n26257 , n26258 );
not ( n26260 , n25978 );
or ( n26261 , n26260 , n21161 );
nand ( n26262 , n26259 , n26261 );
and ( n26263 , n26252 , n26262 );
and ( n26264 , n26241 , n26251 );
or ( n26265 , n26263 , n26264 );
xor ( n26266 , n26215 , n26265 );
xor ( n26267 , n26008 , n26021 );
xor ( n26268 , n26267 , n26044 );
and ( n26269 , n26266 , n26268 );
and ( n26270 , n26215 , n26265 );
or ( n26271 , n26269 , n26270 );
xor ( n26272 , n26182 , n26271 );
xor ( n26273 , n26093 , n26272 );
xor ( n26274 , n26173 , n26175 );
xor ( n26275 , n26274 , n26178 );
not ( n26276 , n20905 );
not ( n26277 , n26042 );
or ( n26278 , n26276 , n26277 );
and ( n26279 , n21213 , n20422 );
not ( n26280 , n21213 );
and ( n26281 , n26280 , n20425 );
nor ( n26282 , n26279 , n26281 );
nand ( n26283 , n26282 , n20860 );
nand ( n26284 , n26278 , n26283 );
not ( n26285 , n26284 );
not ( n26286 , n20693 );
not ( n26287 , n20969 );
or ( n26288 , n26286 , n26287 );
or ( n26289 , n20641 , n20710 );
nand ( n26290 , n26288 , n26289 );
not ( n26291 , n20728 );
not ( n26292 , n26223 );
or ( n26293 , n26291 , n26292 );
not ( n26294 , n20730 );
not ( n26295 , n20946 );
or ( n26296 , n26294 , n26295 );
nand ( n26297 , n20952 , n20745 );
nand ( n26298 , n26296 , n26297 );
nand ( n26299 , n26298 , n20765 );
nand ( n26300 , n26293 , n26299 );
and ( n26301 , n26290 , n26300 );
not ( n26302 , n20979 );
not ( n26303 , n20935 );
not ( n26304 , n21181 );
or ( n26305 , n26303 , n26304 );
nand ( n26306 , n21178 , n20953 );
nand ( n26307 , n26305 , n26306 );
not ( n26308 , n26307 );
or ( n26309 , n26302 , n26308 );
nand ( n26310 , n26189 , n20933 );
nand ( n26311 , n26309 , n26310 );
xor ( n26312 , n26301 , n26311 );
not ( n26313 , n21334 );
not ( n26314 , n26208 );
or ( n26315 , n26313 , n26314 );
not ( n26316 , n20983 );
not ( n26317 , n21138 );
or ( n26318 , n26316 , n26317 );
nand ( n26319 , n21137 , n21487 );
nand ( n26320 , n26318 , n26319 );
nand ( n26321 , n26320 , n21003 );
nand ( n26322 , n26315 , n26321 );
and ( n26323 , n26312 , n26322 );
and ( n26324 , n26301 , n26311 );
or ( n26325 , n26323 , n26324 );
not ( n26326 , n26325 );
or ( n26327 , n26285 , n26326 );
or ( n26328 , n26325 , n26284 );
xor ( n26329 , n26147 , n26115 );
xor ( n26330 , n26329 , n26170 );
nand ( n26331 , n26328 , n26330 );
nand ( n26332 , n26327 , n26331 );
xor ( n26333 , n26275 , n26332 );
xor ( n26334 , n26215 , n26265 );
xor ( n26335 , n26334 , n26268 );
and ( n26336 , n26333 , n26335 );
and ( n26337 , n26275 , n26332 );
or ( n26338 , n26336 , n26337 );
xor ( n26339 , n26273 , n26338 );
xor ( n26340 , n26275 , n26332 );
xor ( n26341 , n26340 , n26335 );
xor ( n26342 , n26191 , n26201 );
xor ( n26343 , n26342 , n26212 );
not ( n26344 , n21148 );
not ( n26345 , n21111 );
not ( n26346 , n25970 );
or ( n26347 , n26345 , n26346 );
nand ( n26348 , n25976 , n21124 );
nand ( n26349 , n26347 , n26348 );
not ( n26350 , n26349 );
or ( n26351 , n26344 , n26350 );
nand ( n26352 , n26247 , n21105 );
nand ( n26353 , n26351 , n26352 );
not ( n26354 , n21199 );
not ( n26355 , n26256 );
or ( n26356 , n26354 , n26355 );
not ( n26357 , n21167 );
not ( n26358 , n20477 );
or ( n26359 , n26357 , n26358 );
nand ( n26360 , n20474 , n21166 );
nand ( n26361 , n26359 , n26360 );
nand ( n26362 , n26361 , n21163 );
nand ( n26363 , n26356 , n26362 );
xor ( n26364 , n26353 , n26363 );
not ( n26365 , n20860 );
and ( n26366 , n21213 , n21394 );
not ( n26367 , n21213 );
and ( n26368 , n26367 , n21391 );
nor ( n26369 , n26366 , n26368 );
not ( n26370 , n26369 );
or ( n26371 , n26365 , n26370 );
nand ( n26372 , n26282 , n20905 );
nand ( n26373 , n26371 , n26372 );
and ( n26374 , n26364 , n26373 );
and ( n26375 , n26353 , n26363 );
or ( n26376 , n26374 , n26375 );
xor ( n26377 , n26343 , n26376 );
xor ( n26378 , n26241 , n26251 );
xor ( n26379 , n26378 , n26262 );
and ( n26380 , n26377 , n26379 );
and ( n26381 , n26343 , n26376 );
or ( n26382 , n26380 , n26381 );
or ( n26383 , n26341 , n26382 );
and ( n26384 , n26284 , n26330 );
not ( n26385 , n26284 );
not ( n26386 , n26330 );
and ( n26387 , n26385 , n26386 );
or ( n26388 , n26384 , n26387 );
xor ( n26389 , n26325 , n26388 );
not ( n26390 , n26389 );
not ( n26391 , n26390 );
xor ( n26392 , n26343 , n26376 );
xor ( n26393 , n26392 , n26379 );
not ( n26394 , n26393 );
or ( n26395 , n26391 , n26394 );
or ( n26396 , n26393 , n26390 );
xor ( n26397 , n26217 , n26227 );
xor ( n26398 , n26397 , n26238 );
xor ( n26399 , n26290 , n26300 );
buf ( n26400 , n26399 );
not ( n26401 , n26400 );
not ( n26402 , n20693 );
not ( n26403 , n21088 );
or ( n26404 , n26402 , n26403 );
or ( n26405 , n20623 , n20710 );
nand ( n26406 , n26404 , n26405 );
not ( n26407 , n20728 );
not ( n26408 , n26298 );
or ( n26409 , n26407 , n26408 );
and ( n26410 , n20730 , n20969 );
not ( n26411 , n20730 );
and ( n26412 , n26411 , n20972 );
nor ( n26413 , n26410 , n26412 );
nand ( n26414 , n26413 , n20765 );
nand ( n26415 , n26409 , n26414 );
and ( n26416 , n26406 , n26415 );
buf ( n26417 , n26416 );
not ( n26418 , n26417 );
or ( n26419 , n26401 , n26418 );
not ( n26420 , n26417 );
not ( n26421 , n26420 );
not ( n26422 , n26400 );
not ( n26423 , n26422 );
or ( n26424 , n26421 , n26423 );
and ( n26425 , n20628 , n21013 );
not ( n26426 , n20628 );
and ( n26427 , n26426 , n21016 );
nor ( n26428 , n26425 , n26427 );
and ( n26429 , n26428 , n20602 );
and ( n26430 , n26234 , n20571 );
nor ( n26431 , n26429 , n26430 );
not ( n26432 , n26431 );
nand ( n26433 , n26424 , n26432 );
nand ( n26434 , n26419 , n26433 );
xor ( n26435 , n26398 , n26434 );
not ( n26436 , n21003 );
and ( n26437 , n20983 , n21193 );
not ( n26438 , n20983 );
and ( n26439 , n26438 , n21196 );
nor ( n26440 , n26437 , n26439 );
not ( n26441 , n26440 );
or ( n26442 , n26436 , n26441 );
nand ( n26443 , n26320 , n21334 );
nand ( n26444 , n26442 , n26443 );
not ( n26445 , n26307 );
or ( n26446 , n26445 , n20932 );
not ( n26447 , n20935 );
not ( n26448 , n20900 );
or ( n26449 , n26447 , n26448 );
nand ( n26450 , n20899 , n20953 );
nand ( n26451 , n26449 , n26450 );
nand ( n26452 , n26451 , n20979 );
nand ( n26453 , n26446 , n26452 );
xor ( n26454 , n26444 , n26453 );
xor ( n26455 , n26406 , n26415 );
not ( n26456 , n20693 );
not ( n26457 , n20620 );
or ( n26458 , n26456 , n26457 );
or ( n26459 , n20787 , n20710 );
nand ( n26460 , n26458 , n26459 );
not ( n26461 , n20728 );
not ( n26462 , n26413 );
or ( n26463 , n26461 , n26462 );
not ( n26464 , n20730 );
not ( n26465 , n20641 );
or ( n26466 , n26464 , n26465 );
nand ( n26467 , n21088 , n20745 );
nand ( n26468 , n26466 , n26467 );
nand ( n26469 , n26468 , n20765 );
nand ( n26470 , n26463 , n26469 );
and ( n26471 , n26460 , n26470 );
xor ( n26472 , n26455 , n26471 );
not ( n26473 , n20602 );
not ( n26474 , n20628 );
not ( n26475 , n20995 );
or ( n26476 , n26474 , n26475 );
nand ( n26477 , n20992 , n20644 );
nand ( n26478 , n26476 , n26477 );
not ( n26479 , n26478 );
or ( n26480 , n26473 , n26479 );
nand ( n26481 , n26428 , n20647 );
nand ( n26482 , n26480 , n26481 );
and ( n26483 , n26472 , n26482 );
and ( n26484 , n26455 , n26471 );
or ( n26485 , n26483 , n26484 );
and ( n26486 , n26454 , n26485 );
and ( n26487 , n26444 , n26453 );
or ( n26488 , n26486 , n26487 );
and ( n26489 , n26435 , n26488 );
and ( n26490 , n26398 , n26434 );
or ( n26491 , n26489 , n26490 );
nand ( n26492 , n26396 , n26491 );
nand ( n26493 , n26395 , n26492 );
nand ( n26494 , n26383 , n26493 );
nand ( n26495 , n26341 , n26382 );
nand ( n26496 , n26494 , n26495 );
or ( n26497 , n26339 , n26496 );
nand ( n26498 , n26339 , n26496 );
nand ( n26499 , n26497 , n26498 );
not ( n26500 , n20905 );
not ( n26501 , n20863 );
not ( n26502 , n21119 );
or ( n26503 , n26501 , n26502 );
nand ( n26504 , n21118 , n20862 );
nand ( n26505 , n26503 , n26504 );
not ( n26506 , n26505 );
or ( n26507 , n26500 , n26506 );
not ( n26508 , n20863 );
not ( n26509 , n21138 );
or ( n26510 , n26508 , n26509 );
nand ( n26511 , n21137 , n20862 );
nand ( n26512 , n26510 , n26511 );
nand ( n26513 , n26512 , n20860 );
nand ( n26514 , n26507 , n26513 );
not ( n26515 , n18012 );
not ( n26516 , n18029 );
not ( n26517 , n26004 );
or ( n26518 , n26516 , n26517 );
nand ( n26519 , n26001 , n18028 );
nand ( n26520 , n26518 , n26519 );
not ( n26521 , n26520 );
or ( n26522 , n26515 , n26521 );
not ( n26523 , n18029 );
not ( n26524 , n25970 );
or ( n26525 , n26523 , n26524 );
nand ( n26526 , n25976 , n18028 );
nand ( n26527 , n26525 , n26526 );
nand ( n26528 , n26527 , n18025 );
nand ( n26529 , n26522 , n26528 );
xor ( n26530 , n26514 , n26529 );
not ( n26531 , n21148 );
and ( n26532 , n21124 , n20477 );
not ( n26533 , n21124 );
and ( n26534 , n26533 , n20474 );
or ( n26535 , n26532 , n26534 );
not ( n26536 , n26535 );
not ( n26537 , n26536 );
or ( n26538 , n26531 , n26537 );
not ( n26539 , n21111 );
not ( n26540 , n26032 );
or ( n26541 , n26539 , n26540 );
nand ( n26542 , n26031 , n21124 );
nand ( n26543 , n26541 , n26542 );
nand ( n26544 , n26543 , n21105 );
nand ( n26545 , n26538 , n26544 );
and ( n26546 , n26530 , n26545 );
and ( n26547 , n26514 , n26529 );
or ( n26548 , n26546 , n26547 );
xor ( n26549 , n26444 , n26453 );
xor ( n26550 , n26549 , n26485 );
xor ( n26551 , n26548 , n26550 );
not ( n26552 , n20905 );
not ( n26553 , n26369 );
or ( n26554 , n26552 , n26553 );
nand ( n26555 , n26505 , n20860 );
nand ( n26556 , n26554 , n26555 );
not ( n26557 , n21148 );
not ( n26558 , n26543 );
or ( n26559 , n26557 , n26558 );
nand ( n26560 , n26349 , n21105 );
nand ( n26561 , n26559 , n26560 );
xor ( n26562 , n26556 , n26561 );
not ( n26563 , n18029 );
not ( n26564 , n18012 );
or ( n26565 , n26563 , n26564 );
not ( n26566 , n26520 );
or ( n26567 , n26566 , n18024 );
nand ( n26568 , n26565 , n26567 );
xor ( n26569 , n26562 , n26568 );
xor ( n26570 , n26551 , n26569 );
xor ( n26571 , n26455 , n26471 );
xor ( n26572 , n26571 , n26482 );
not ( n26573 , n21163 );
not ( n26574 , n21167 );
not ( n26575 , n21391 );
or ( n26576 , n26574 , n26575 );
nand ( n26577 , n21394 , n21166 );
nand ( n26578 , n26576 , n26577 );
not ( n26579 , n26578 );
or ( n26580 , n26573 , n26579 );
not ( n26581 , n21167 );
not ( n26582 , n20425 );
or ( n26583 , n26581 , n26582 );
nand ( n26584 , n20422 , n21166 );
nand ( n26585 , n26583 , n26584 );
nand ( n26586 , n26585 , n21199 );
nand ( n26587 , n26580 , n26586 );
xor ( n26588 , n26572 , n26587 );
not ( n26589 , n21433 );
nor ( n26590 , n26589 , n21438 );
not ( n26591 , n20647 );
not ( n26592 , n20644 );
not ( n26593 , n20945 );
or ( n26594 , n26592 , n26593 );
nand ( n26595 , n20946 , n20628 );
nand ( n26596 , n26594 , n26595 );
not ( n26597 , n26596 );
or ( n26598 , n26591 , n26597 );
nand ( n26599 , n21417 , n20602 );
nand ( n26600 , n26598 , n26599 );
xor ( n26601 , n26590 , n26600 );
not ( n26602 , n20693 );
not ( n26603 , n20794 );
or ( n26604 , n26602 , n26603 );
nand ( n26605 , n20741 , n21045 );
nand ( n26606 , n26604 , n26605 );
not ( n26607 , n20765 );
not ( n26608 , n21431 );
or ( n26609 , n26607 , n26608 );
nand ( n26610 , n26468 , n20728 );
nand ( n26611 , n26609 , n26610 );
xor ( n26612 , n26606 , n26611 );
and ( n26613 , n26601 , n26612 );
and ( n26614 , n26590 , n26600 );
or ( n26615 , n26613 , n26614 );
not ( n26616 , n20935 );
not ( n26617 , n20875 );
or ( n26618 , n26616 , n26617 );
nand ( n26619 , n20878 , n20953 );
nand ( n26620 , n26618 , n26619 );
not ( n26621 , n26620 );
or ( n26622 , n26621 , n20932 );
not ( n26623 , n20935 );
not ( n26624 , n21016 );
or ( n26625 , n26623 , n26624 );
nand ( n26626 , n21013 , n20953 );
nand ( n26627 , n26625 , n26626 );
nand ( n26628 , n26627 , n20980 );
nand ( n26629 , n26622 , n26628 );
xor ( n26630 , n26615 , n26629 );
not ( n26631 , n21003 );
not ( n26632 , n20983 );
not ( n26633 , n20900 );
or ( n26634 , n26632 , n26633 );
nand ( n26635 , n20899 , n21487 );
nand ( n26636 , n26634 , n26635 );
not ( n26637 , n26636 );
or ( n26638 , n26631 , n26637 );
and ( n26639 , n20983 , n21178 );
not ( n26640 , n20983 );
and ( n26641 , n26640 , n21181 );
nor ( n26642 , n26639 , n26641 );
nand ( n26643 , n26642 , n21334 );
nand ( n26644 , n26638 , n26643 );
and ( n26645 , n26630 , n26644 );
and ( n26646 , n26615 , n26629 );
or ( n26647 , n26645 , n26646 );
and ( n26648 , n26588 , n26647 );
and ( n26649 , n26572 , n26587 );
or ( n26650 , n26648 , n26649 );
not ( n26651 , n21163 );
not ( n26652 , n26585 );
or ( n26653 , n26651 , n26652 );
nand ( n26654 , n26361 , n21199 );
nand ( n26655 , n26653 , n26654 );
xor ( n26656 , n26431 , n26417 );
and ( n26657 , n26656 , n26422 );
not ( n26658 , n26656 );
and ( n26659 , n26658 , n26400 );
nor ( n26660 , n26657 , n26659 );
xor ( n26661 , n26655 , n26660 );
not ( n26662 , n20979 );
not ( n26663 , n26620 );
or ( n26664 , n26662 , n26663 );
nand ( n26665 , n26451 , n20933 );
nand ( n26666 , n26664 , n26665 );
not ( n26667 , n21334 );
not ( n26668 , n26440 );
or ( n26669 , n26667 , n26668 );
nand ( n26670 , n26642 , n21003 );
nand ( n26671 , n26669 , n26670 );
xor ( n26672 , n26666 , n26671 );
and ( n26673 , n26606 , n26611 );
not ( n26674 , n20647 );
not ( n26675 , n26478 );
or ( n26676 , n26674 , n26675 );
nand ( n26677 , n26596 , n20602 );
nand ( n26678 , n26676 , n26677 );
xor ( n26679 , n26673 , n26678 );
xor ( n26680 , n26460 , n26470 );
and ( n26681 , n26679 , n26680 );
and ( n26682 , n26673 , n26678 );
or ( n26683 , n26681 , n26682 );
and ( n26684 , n26672 , n26683 );
and ( n26685 , n26666 , n26671 );
or ( n26686 , n26684 , n26685 );
xor ( n26687 , n26661 , n26686 );
xor ( n26688 , n26650 , n26687 );
xor ( n26689 , n26666 , n26671 );
xor ( n26690 , n26689 , n26683 );
not ( n26691 , n20905 );
not ( n26692 , n26512 );
or ( n26693 , n26691 , n26692 );
not ( n26694 , n21213 );
not ( n26695 , n21196 );
or ( n26696 , n26694 , n26695 );
nand ( n26697 , n21193 , n20862 );
nand ( n26698 , n26696 , n26697 );
nand ( n26699 , n26698 , n20860 );
nand ( n26700 , n26693 , n26699 );
not ( n26701 , n18012 );
not ( n26702 , n26527 );
or ( n26703 , n26701 , n26702 );
not ( n26704 , n18029 );
not ( n26705 , n26032 );
or ( n26706 , n26704 , n26705 );
nand ( n26707 , n26031 , n18028 );
nand ( n26708 , n26706 , n26707 );
nand ( n26709 , n26708 , n18025 );
nand ( n26710 , n26703 , n26709 );
xor ( n26711 , n26700 , n26710 );
not ( n26712 , n21111 );
not ( n26713 , n20425 );
or ( n26714 , n26712 , n26713 );
nand ( n26715 , n21124 , n20422 );
nand ( n26716 , n26714 , n26715 );
not ( n26717 , n26716 );
not ( n26718 , n21148 );
or ( n26719 , n26717 , n26718 );
not ( n26720 , n21105 );
or ( n26721 , n26535 , n26720 );
nand ( n26722 , n26719 , n26721 );
and ( n26723 , n26711 , n26722 );
and ( n26724 , n26700 , n26710 );
or ( n26725 , n26723 , n26724 );
xor ( n26726 , n26690 , n26725 );
xor ( n26727 , n26673 , n26678 );
xor ( n26728 , n26727 , n26680 );
not ( n26729 , n20933 );
not ( n26730 , n26627 );
or ( n26731 , n26729 , n26730 );
nand ( n26732 , n21475 , n20979 );
nand ( n26733 , n26731 , n26732 );
not ( n26734 , n21334 );
not ( n26735 , n26636 );
or ( n26736 , n26734 , n26735 );
nand ( n26737 , n21489 , n21003 );
nand ( n26738 , n26736 , n26737 );
xor ( n26739 , n26733 , n26738 );
xor ( n26740 , n21412 , n21421 );
and ( n26741 , n26740 , n21439 );
and ( n26742 , n21412 , n21421 );
or ( n26743 , n26741 , n26742 );
and ( n26744 , n26739 , n26743 );
and ( n26745 , n26733 , n26738 );
or ( n26746 , n26744 , n26745 );
xor ( n26747 , n26728 , n26746 );
not ( n26748 , n26578 );
or ( n26749 , n26748 , n21161 );
not ( n26750 , n21167 );
not ( n26751 , n21119 );
or ( n26752 , n26750 , n26751 );
nand ( n26753 , n21118 , n21166 );
nand ( n26754 , n26752 , n26753 );
nand ( n26755 , n26754 , n21163 );
nand ( n26756 , n26749 , n26755 );
and ( n26757 , n26747 , n26756 );
and ( n26758 , n26728 , n26746 );
or ( n26759 , n26757 , n26758 );
and ( n26760 , n26726 , n26759 );
and ( n26761 , n26690 , n26725 );
or ( n26762 , n26760 , n26761 );
xor ( n26763 , n26688 , n26762 );
xor ( n26764 , n26570 , n26763 );
xor ( n26765 , n26514 , n26529 );
xor ( n26766 , n26765 , n26545 );
xor ( n26767 , n26572 , n26587 );
xor ( n26768 , n26767 , n26647 );
xor ( n26769 , n26766 , n26768 );
xor ( n26770 , n26615 , n26629 );
xor ( n26771 , n26770 , n26644 );
not ( n26772 , n26771 );
not ( n26773 , n21148 );
not ( n26774 , n21501 );
or ( n26775 , n26773 , n26774 );
nand ( n26776 , n26716 , n21105 );
nand ( n26777 , n26775 , n26776 );
not ( n26778 , n18025 );
not ( n26779 , n20479 );
or ( n26780 , n26778 , n26779 );
nand ( n26781 , n26708 , n18012 );
nand ( n26782 , n26780 , n26781 );
xor ( n26783 , n26777 , n26782 );
xor ( n26784 , n21469 , n21479 );
and ( n26785 , n26784 , n21491 );
and ( n26786 , n21469 , n21479 );
or ( n26787 , n26785 , n26786 );
and ( n26788 , n26783 , n26787 );
and ( n26789 , n26777 , n26782 );
or ( n26790 , n26788 , n26789 );
not ( n26791 , n26790 );
or ( n26792 , n26772 , n26791 );
or ( n26793 , n26790 , n26771 );
xor ( n26794 , n26590 , n26600 );
xor ( n26795 , n26794 , n26612 );
not ( n26796 , n20860 );
not ( n26797 , n21456 );
or ( n26798 , n26796 , n26797 );
nand ( n26799 , n26698 , n20905 );
nand ( n26800 , n26798 , n26799 );
xor ( n26801 , n26795 , n26800 );
not ( n26802 , n21199 );
not ( n26803 , n26754 );
or ( n26804 , n26802 , n26803 );
nand ( n26805 , n21448 , n21163 );
nand ( n26806 , n26804 , n26805 );
and ( n26807 , n26801 , n26806 );
and ( n26808 , n26795 , n26800 );
or ( n26809 , n26807 , n26808 );
nand ( n26810 , n26793 , n26809 );
nand ( n26811 , n26792 , n26810 );
and ( n26812 , n26769 , n26811 );
and ( n26813 , n26766 , n26768 );
or ( n26814 , n26812 , n26813 );
xor ( n26815 , n26764 , n26814 );
xor ( n26816 , n26690 , n26725 );
xor ( n26817 , n26816 , n26759 );
buf ( n26818 , n26817 );
not ( n26819 , n26818 );
xor ( n26820 , n26766 , n26768 );
xor ( n26821 , n26820 , n26811 );
not ( n26822 , n26821 );
or ( n26823 , n26819 , n26822 );
or ( n26824 , n26821 , n26818 );
xor ( n26825 , n26700 , n26710 );
xor ( n26826 , n26825 , n26722 );
xor ( n26827 , n26728 , n26746 );
xor ( n26828 , n26827 , n26756 );
xor ( n26829 , n26826 , n26828 );
xor ( n26830 , n26733 , n26738 );
xor ( n26831 , n26830 , n26743 );
xor ( n26832 , n21440 , n21450 );
and ( n26833 , n26832 , n21460 );
and ( n26834 , n21440 , n21450 );
or ( n26835 , n26833 , n26834 );
xor ( n26836 , n26831 , n26835 );
xor ( n26837 , n21465 , n21492 );
and ( n26838 , n26837 , n21503 );
and ( n26839 , n21465 , n21492 );
or ( n26840 , n26838 , n26839 );
and ( n26841 , n26836 , n26840 );
and ( n26842 , n26831 , n26835 );
or ( n26843 , n26841 , n26842 );
and ( n26844 , n26829 , n26843 );
and ( n26845 , n26826 , n26828 );
or ( n26846 , n26844 , n26845 );
nand ( n26847 , n26824 , n26846 );
nand ( n26848 , n26823 , n26847 );
nor ( n26849 , n26815 , n26848 );
xor ( n26850 , n26655 , n26660 );
and ( n26851 , n26850 , n26686 );
and ( n26852 , n26655 , n26660 );
or ( n26853 , n26851 , n26852 );
xor ( n26854 , n26398 , n26434 );
xor ( n26855 , n26854 , n26488 );
xor ( n26856 , n26853 , n26855 );
xor ( n26857 , n26301 , n26311 );
xor ( n26858 , n26857 , n26322 );
xor ( n26859 , n26556 , n26561 );
and ( n26860 , n26859 , n26568 );
and ( n26861 , n26556 , n26561 );
or ( n26862 , n26860 , n26861 );
xor ( n26863 , n26858 , n26862 );
xor ( n26864 , n26353 , n26363 );
xor ( n26865 , n26864 , n26373 );
xor ( n26866 , n26863 , n26865 );
xor ( n26867 , n26856 , n26866 );
not ( n26868 , n26867 );
xor ( n26869 , n26650 , n26687 );
and ( n26870 , n26869 , n26762 );
and ( n26871 , n26650 , n26687 );
or ( n26872 , n26870 , n26871 );
not ( n26873 , n26872 );
xor ( n26874 , n26548 , n26550 );
and ( n26875 , n26874 , n26569 );
and ( n26876 , n26548 , n26550 );
or ( n26877 , n26875 , n26876 );
not ( n26878 , n26877 );
not ( n26879 , n26878 );
and ( n26880 , n26873 , n26879 );
and ( n26881 , n26872 , n26878 );
nor ( n26882 , n26880 , n26881 );
not ( n26883 , n26882 );
or ( n26884 , n26868 , n26883 );
or ( n26885 , n26867 , n26882 );
nand ( n26886 , n26884 , n26885 );
xor ( n26887 , n26570 , n26763 );
and ( n26888 , n26887 , n26814 );
and ( n26889 , n26570 , n26763 );
or ( n26890 , n26888 , n26889 );
nor ( n26891 , n26886 , n26890 );
nor ( n26892 , n26849 , n26891 );
xor ( n26893 , n26858 , n26862 );
and ( n26894 , n26893 , n26865 );
and ( n26895 , n26858 , n26862 );
or ( n26896 , n26894 , n26895 );
not ( n26897 , n26896 );
not ( n26898 , n26897 );
not ( n26899 , n26393 );
xor ( n26900 , n26491 , n26389 );
not ( n26901 , n26900 );
and ( n26902 , n26899 , n26901 );
and ( n26903 , n26393 , n26900 );
nor ( n26904 , n26902 , n26903 );
not ( n26905 , n26904 );
not ( n26906 , n26905 );
or ( n26907 , n26898 , n26906 );
nand ( n26908 , n26904 , n26896 );
nand ( n26909 , n26907 , n26908 );
xor ( n26910 , n26853 , n26855 );
and ( n26911 , n26910 , n26866 );
and ( n26912 , n26853 , n26855 );
or ( n26913 , n26911 , n26912 );
not ( n26914 , n26913 );
and ( n26915 , n26909 , n26914 );
not ( n26916 , n26909 );
and ( n26917 , n26916 , n26913 );
nor ( n26918 , n26915 , n26917 );
not ( n26919 , n26872 );
not ( n26920 , n26919 );
not ( n26921 , n26878 );
and ( n26922 , n26920 , n26921 );
nand ( n26923 , n26919 , n26878 );
and ( n26924 , n26867 , n26923 );
nor ( n26925 , n26922 , n26924 );
nand ( n26926 , n26918 , n26925 );
not ( n26927 , n26897 );
not ( n26928 , n26904 );
or ( n26929 , n26927 , n26928 );
nand ( n26930 , n26929 , n26913 );
nand ( n26931 , n26905 , n26896 );
and ( n26932 , n26930 , n26931 );
xor ( n26933 , n26382 , n26341 );
xnor ( n26934 , n26933 , n26493 );
nand ( n26935 , n26932 , n26934 );
and ( n26936 , n26892 , n26926 , n26935 );
not ( n26937 , n26936 );
xor ( n26938 , n26817 , n26846 );
xnor ( n26939 , n26938 , n26821 );
xor ( n26940 , n26826 , n26828 );
xor ( n26941 , n26940 , n26843 );
xor ( n26942 , n26771 , n26809 );
xnor ( n26943 , n26942 , n26790 );
not ( n26944 , n26943 );
or ( n26945 , n26941 , n26944 );
xor ( n26946 , n26795 , n26800 );
xor ( n26947 , n26946 , n26806 );
xor ( n26948 , n26777 , n26782 );
xor ( n26949 , n26948 , n26787 );
xor ( n26950 , n26947 , n26949 );
xor ( n26951 , n20481 , n21068 );
and ( n26952 , n26951 , n21204 );
and ( n26953 , n20481 , n21068 );
or ( n26954 , n26952 , n26953 );
and ( n26955 , n26950 , n26954 );
and ( n26956 , n26947 , n26949 );
or ( n26957 , n26955 , n26956 );
nand ( n26958 , n26945 , n26957 );
nand ( n26959 , n26941 , n26944 );
and ( n26960 , n26958 , n26959 );
nand ( n26961 , n26939 , n26960 );
xor ( n26962 , n26957 , n26943 );
xor ( n26963 , n26962 , n26941 );
xor ( n26964 , n26947 , n26949 );
xor ( n26965 , n26964 , n26954 );
xor ( n26966 , n26831 , n26835 );
xor ( n26967 , n26966 , n26840 );
or ( n26968 , n26965 , n26967 );
xor ( n26969 , n21461 , n21504 );
and ( n26970 , n26969 , n21550 );
and ( n26971 , n21461 , n21504 );
or ( n26972 , n26970 , n26971 );
and ( n26973 , n26968 , n26972 );
and ( n26974 , n26967 , n26965 );
nor ( n26975 , n26973 , n26974 );
nand ( n26976 , n26963 , n26975 );
and ( n26977 , n26961 , n26976 );
not ( n26978 , n26977 );
xor ( n26979 , n26967 , n26965 );
xor ( n26980 , n26979 , n26972 );
not ( n26981 , n26980 );
or ( n26982 , n21551 , n21205 );
nand ( n26983 , n26982 , n21410 );
nand ( n26984 , n21551 , n21205 );
nand ( n26985 , n26983 , n26984 );
not ( n26986 , n26985 );
nand ( n26987 , n26981 , n26986 );
and ( n26988 , n26987 , n21791 );
not ( n26989 , n26988 );
not ( n26990 , n23835 );
or ( n26991 , n26989 , n26990 );
and ( n26992 , n26987 , n21789 );
and ( n26993 , n26980 , n26985 );
nor ( n26994 , n26992 , n26993 );
nand ( n26995 , n26991 , n26994 );
not ( n26996 , n26995 );
or ( n26997 , n26978 , n26996 );
nor ( n26998 , n26963 , n26975 );
and ( n26999 , n26961 , n26998 );
nor ( n27000 , n26939 , n26960 );
nor ( n27001 , n26999 , n27000 );
nand ( n27002 , n26997 , n27001 );
not ( n27003 , n27002 );
or ( n27004 , n26937 , n27003 );
not ( n27005 , n26926 );
nand ( n27006 , n26815 , n26848 );
or ( n27007 , n27006 , n26891 );
nand ( n27008 , n26886 , n26890 );
nand ( n27009 , n27007 , n27008 );
not ( n27010 , n27009 );
or ( n27011 , n27005 , n27010 );
not ( n27012 , n26918 );
not ( n27013 , n26925 );
nand ( n27014 , n27012 , n27013 );
nand ( n27015 , n27011 , n27014 );
and ( n27016 , n27015 , n26935 );
nor ( n27017 , n26932 , n26934 );
nor ( n27018 , n27016 , n27017 );
nand ( n27019 , n27004 , n27018 );
xor ( n27020 , n26499 , n27019 );
or ( n27021 , n27020 , n23837 );
nand ( n27022 , n25858 , n27021 );
not ( n27023 , n17533 );
not ( n27024 , n27023 );
not ( n27025 , n23913 );
or ( n27026 , n27024 , n27025 );
not ( n27027 , n17612 );
nand ( n27028 , n27026 , n27027 );
not ( n27029 , n17611 );
nor ( n27030 , n27029 , n17615 );
and ( n27031 , n27028 , n27030 );
not ( n27032 , n27028 );
not ( n27033 , n27030 );
and ( n27034 , n27032 , n27033 );
or ( n27035 , n27031 , n27034 );
or ( n27036 , n27035 , n23844 );
nor ( n27037 , n23943 , n23802 );
xor ( n27038 , n27037 , n23942 );
or ( n27039 , n27038 , n23845 );
nand ( n27040 , n27036 , n27039 );
nand ( n27041 , n27023 , n27027 );
xor ( n27042 , n23913 , n27041 );
or ( n27043 , n27042 , n23844 );
nand ( n27044 , n23751 , n23059 );
xor ( n27045 , n27044 , n23747 );
or ( n27046 , n27045 , n23948 );
nand ( n27047 , n27043 , n27046 );
not ( n27048 , n17604 );
nor ( n27049 , n27048 , n16909 );
not ( n27050 , n27049 );
not ( n27051 , n16950 );
not ( n27052 , n27051 );
buf ( n27053 , n17357 );
not ( n27054 , n27053 );
or ( n27055 , n27052 , n27054 );
nand ( n27056 , n27055 , n17602 );
not ( n27057 , n27056 );
or ( n27058 , n27050 , n27057 );
or ( n27059 , n27049 , n27056 );
nand ( n27060 , n27058 , n27059 );
or ( n27061 , n27060 , n23844 );
xor ( n27062 , n23204 , n23206 );
xor ( n27063 , n27062 , n23744 );
not ( n27064 , n27063 );
or ( n27065 , n27064 , n23948 );
nand ( n27066 , n27061 , n27065 );
nor ( n27067 , n25510 , n25513 );
not ( n27068 , n27067 );
not ( n27069 , n25663 );
nand ( n27070 , n27068 , n27069 );
not ( n27071 , n25656 );
and ( n27072 , n27070 , n27071 );
not ( n27073 , n27070 );
and ( n27074 , n27073 , n25656 );
or ( n27075 , n27072 , n27074 );
or ( n27076 , n27075 , n18007 );
and ( n27077 , n27014 , n26926 );
and ( n27078 , n27002 , n26892 );
buf ( n27079 , n27009 );
nor ( n27080 , n27078 , n27079 );
xor ( n27081 , n27077 , n27080 );
or ( n27082 , n27081 , n23837 );
nand ( n27083 , n27076 , n27082 );
and ( n27084 , n27051 , n17602 );
not ( n27085 , n27084 );
not ( n27086 , n27053 );
or ( n27087 , n27085 , n27086 );
or ( n27088 , n27084 , n27053 );
nand ( n27089 , n27087 , n27088 );
or ( n27090 , n27089 , n23844 );
xor ( n27091 , n23233 , n23235 );
xor ( n27092 , n27091 , n23741 );
not ( n27093 , n27092 );
or ( n27094 , n27093 , n23948 );
nand ( n27095 , n27090 , n27094 );
nand ( n27096 , n17033 , n17352 );
xor ( n27097 , n27096 , n17348 );
or ( n27098 , n27097 , n23844 );
not ( n27099 , n23725 );
nand ( n27100 , n27099 , n23728 );
not ( n27101 , n27100 );
nand ( n27102 , n23697 , n23414 );
not ( n27103 , n27102 );
or ( n27104 , n27101 , n27103 );
or ( n27105 , n27102 , n27100 );
nand ( n27106 , n27104 , n27105 );
not ( n27107 , n27106 );
or ( n27108 , n27107 , n23948 );
nand ( n27109 , n27098 , n27108 );
not ( n27110 , n17336 );
and ( n27111 , n17138 , n17339 );
not ( n27112 , n27111 );
or ( n27113 , n27110 , n27112 );
or ( n27114 , n27111 , n17336 );
nand ( n27115 , n27113 , n27114 );
or ( n27116 , n27115 , n23844 );
xor ( n27117 , n23475 , n23477 );
xor ( n27118 , n27117 , n23688 );
not ( n27119 , n27118 );
or ( n27120 , n27119 , n23845 );
nand ( n27121 , n27116 , n27120 );
not ( n27122 , n17332 );
and ( n27123 , n17176 , n17335 );
not ( n27124 , n27123 );
or ( n27125 , n27122 , n27124 );
or ( n27126 , n27123 , n17332 );
nand ( n27127 , n27125 , n27126 );
or ( n27128 , n27127 , n23844 );
nand ( n27129 , n23687 , n23573 );
xor ( n27130 , n23683 , n27129 );
or ( n27131 , n27130 , n23948 );
nand ( n27132 , n27128 , n27131 );
not ( n27133 , n17691 );
not ( n27134 , n25602 );
or ( n27135 , n27133 , n27134 );
nand ( n27136 , n27135 , n25634 );
nand ( n27137 , n25645 , n27136 );
nand ( n27138 , n25653 , n25584 );
xor ( n27139 , n27137 , n27138 );
or ( n27140 , n27139 , n18007 );
not ( n27141 , n27000 );
nand ( n27142 , n27141 , n26961 );
not ( n27143 , n26976 );
not ( n27144 , n26995 );
or ( n27145 , n27143 , n27144 );
not ( n27146 , n26998 );
nand ( n27147 , n27145 , n27146 );
xor ( n27148 , n27142 , n27147 );
or ( n27149 , n27148 , n23837 );
nand ( n27150 , n27140 , n27149 );
and ( n27151 , n17331 , n17211 );
xnor ( n27152 , n17328 , n27151 );
or ( n27153 , n27152 , n23844 );
nand ( n27154 , n23682 , n23588 );
xor ( n27155 , n23678 , n27154 );
or ( n27156 , n27155 , n23948 );
nand ( n27157 , n27153 , n27156 );
not ( n27158 , n23837 );
not ( n27159 , n25637 );
nand ( n27160 , n27159 , n25639 );
not ( n27161 , n27160 );
nand ( n27162 , n17692 , n17998 );
nand ( n27163 , n27162 , n17999 );
not ( n27164 , n27163 );
or ( n27165 , n27161 , n27164 );
or ( n27166 , n27160 , n27163 );
nand ( n27167 , n27165 , n27166 );
not ( n27168 , n27167 );
or ( n27169 , n27158 , n27168 );
not ( n27170 , n26993 );
nand ( n27171 , n27170 , n26987 );
not ( n27172 , n27171 );
not ( n27173 , n21791 );
not ( n27174 , n23835 );
or ( n27175 , n27173 , n27174 );
nand ( n27176 , n27175 , n21790 );
not ( n27177 , n27176 );
or ( n27178 , n27172 , n27177 );
or ( n27179 , n27176 , n27171 );
nand ( n27180 , n27178 , n27179 );
nand ( n27181 , n27180 , n18007 );
nand ( n27182 , n27169 , n27181 );
and ( n27183 , n20878 , n21045 );
and ( n27184 , n20899 , n20693 );
nor ( n27185 , n27183 , n27184 );
not ( n27186 , n27185 );
or ( n27187 , n21162 , n21199 );
nand ( n27188 , n27187 , n21167 );
not ( n27189 , n27188 );
and ( n27190 , n27186 , n27189 );
and ( n27191 , n27185 , n27188 );
nor ( n27192 , n27190 , n27191 );
not ( n27193 , n27192 );
not ( n27194 , n20647 );
not ( n27195 , n20628 );
not ( n27196 , n21119 );
or ( n27197 , n27195 , n27196 );
nand ( n27198 , n21118 , n20644 );
nand ( n27199 , n27197 , n27198 );
not ( n27200 , n27199 );
or ( n27201 , n27194 , n27200 );
nand ( n27202 , n25870 , n20602 );
nand ( n27203 , n27201 , n27202 );
not ( n27204 , n27203 );
or ( n27205 , n27193 , n27204 );
or ( n27206 , n27203 , n27192 );
nand ( n27207 , n27205 , n27206 );
not ( n27208 , n20765 );
not ( n27209 , n25886 );
or ( n27210 , n27208 , n27209 );
and ( n27211 , n20730 , n21193 );
not ( n27212 , n20730 );
and ( n27213 , n27212 , n21196 );
nor ( n27214 , n27211 , n27213 );
nand ( n27215 , n27214 , n20728 );
nand ( n27216 , n27210 , n27215 );
xor ( n27217 , n25863 , n27216 );
not ( n27218 , n20933 );
not ( n27219 , n20935 );
not ( n27220 , n20425 );
or ( n27221 , n27219 , n27220 );
nand ( n27222 , n20953 , n20422 );
nand ( n27223 , n27221 , n27222 );
not ( n27224 , n27223 );
or ( n27225 , n27218 , n27224 );
nand ( n27226 , n26089 , n20979 );
nand ( n27227 , n27225 , n27226 );
xor ( n27228 , n27217 , n27227 );
xor ( n27229 , n27207 , n27228 );
xor ( n27230 , n26053 , n26076 );
and ( n27231 , n27230 , n26091 );
and ( n27232 , n26053 , n26076 );
or ( n27233 , n27231 , n27232 );
xor ( n27234 , n27229 , n27233 );
not ( n27235 , n21003 );
not ( n27236 , n26098 );
or ( n27237 , n27235 , n27236 );
not ( n27238 , n20983 );
not ( n27239 , n26032 );
or ( n27240 , n27238 , n27239 );
nand ( n27241 , n26031 , n21487 );
nand ( n27242 , n27240 , n27241 );
nand ( n27243 , n27242 , n21334 );
nand ( n27244 , n27237 , n27243 );
not ( n27245 , n20860 );
not ( n27246 , n26107 );
or ( n27247 , n27245 , n27246 );
not ( n27248 , n20863 );
not ( n27249 , n26004 );
or ( n27250 , n27248 , n27249 );
nand ( n27251 , n26001 , n20862 );
nand ( n27252 , n27250 , n27251 );
nand ( n27253 , n27252 , n20905 );
nand ( n27254 , n27247 , n27253 );
xor ( n27255 , n27244 , n27254 );
xor ( n27256 , n25864 , n25879 );
and ( n27257 , n27256 , n25895 );
and ( n27258 , n25864 , n25879 );
or ( n27259 , n27257 , n27258 );
xor ( n27260 , n27255 , n27259 );
xor ( n27261 , n26102 , n26111 );
and ( n27262 , n27261 , n26140 );
and ( n27263 , n26102 , n26111 );
or ( n27264 , n27262 , n27263 );
not ( n27265 , n27264 );
xor ( n27266 , n27260 , n27265 );
xor ( n27267 , n25896 , n26047 );
and ( n27268 , n27267 , n26092 );
and ( n27269 , n25896 , n26047 );
or ( n27270 , n27268 , n27269 );
xnor ( n27271 , n27266 , n27270 );
xor ( n27272 , n27234 , n27271 );
xor ( n27273 , n26141 , n26181 );
and ( n27274 , n27273 , n26271 );
and ( n27275 , n26141 , n26181 );
or ( n27276 , n27274 , n27275 );
xor ( n27277 , n27272 , n27276 );
xor ( n27278 , n26093 , n26272 );
and ( n27279 , n27278 , n26338 );
and ( n27280 , n26093 , n26272 );
or ( n27281 , n27279 , n27280 );
nand ( n27282 , n27277 , n27281 );
nor ( n27283 , n27277 , n27281 );
not ( n27284 , n27283 );
nand ( n27285 , n27282 , n27284 );
not ( n27286 , n27285 );
not ( n27287 , n26936 );
not ( n27288 , n27002 );
or ( n27289 , n27287 , n27288 );
nand ( n27290 , n27289 , n27018 );
nand ( n27291 , n27290 , n26497 );
nand ( n27292 , n27291 , n26498 );
not ( n27293 , n27292 );
or ( n27294 , n27286 , n27293 );
or ( n27295 , n27292 , n27285 );
nand ( n27296 , n27294 , n27295 );
nand ( n27297 , n27296 , n18007 );
not ( n27298 , n23694 );
nand ( n27299 , n23414 , n23696 );
not ( n27300 , n27299 );
or ( n27301 , n27298 , n27300 );
or ( n27302 , n27299 , n23694 );
nand ( n27303 , n27301 , n27302 );
and ( n27304 , n27303 , n23844 );
not ( n27305 , n454 );
not ( n27306 , n9233 );
or ( n27307 , n27305 , n27306 );
or ( n27308 , n15047 , n454 );
nand ( n27309 , n27307 , n27308 );
not ( n27310 , n27309 );
not ( n27311 , n23607 );
nand ( n27312 , n27311 , n23663 );
xor ( n27313 , n23661 , n27312 );
and ( n27314 , n23844 , n27313 );
not ( n27315 , n23844 );
not ( n27316 , n17321 );
not ( n27317 , n27316 );
not ( n27318 , n17288 );
nand ( n27319 , n27318 , n17323 );
not ( n27320 , n27319 );
or ( n27321 , n27317 , n27320 );
or ( n27322 , n27316 , n27319 );
nand ( n27323 , n27321 , n27322 );
and ( n27324 , n27315 , n27323 );
or ( n27325 , n27314 , n27324 );
not ( n27326 , n454 );
nand ( n27327 , n25176 , n25117 , n25774 );
xor ( n27328 , n25781 , n25792 );
and ( n27329 , n27328 , n25794 );
and ( n27330 , n25781 , n25792 );
or ( n27331 , n27329 , n27330 );
not ( n27332 , n16173 );
not ( n27333 , n25797 );
or ( n27334 , n27332 , n27333 );
and ( n27335 , n537 , n9886 );
not ( n27336 , n537 );
and ( n27337 , n27336 , n9887 );
nor ( n27338 , n27335 , n27337 );
nand ( n27339 , n27338 , n5697 );
nand ( n27340 , n27334 , n27339 );
and ( n27341 , n537 , n24903 );
xor ( n27342 , n27340 , n27341 );
and ( n27343 , n25790 , n4450 );
nor ( n27344 , n27343 , n5971 );
xor ( n27345 , n27342 , n27344 );
xor ( n27346 , n27331 , n27345 );
xor ( n27347 , n25801 , n25802 );
and ( n27348 , n27347 , n25807 );
and ( n27349 , n25801 , n25802 );
or ( n27350 , n27348 , n27349 );
xor ( n27351 , n27346 , n27350 );
not ( n27352 , n27351 );
xor ( n27353 , n25795 , n25808 );
and ( n27354 , n27353 , n25813 );
and ( n27355 , n25795 , n25808 );
or ( n27356 , n27354 , n27355 );
not ( n27357 , n27356 );
nand ( n27358 , n27352 , n27357 );
not ( n27359 , n27358 );
nor ( n27360 , n27359 , n25821 );
not ( n27361 , n27344 );
or ( n27362 , n4450 , n4659 );
nand ( n27363 , n27362 , n539 );
not ( n27364 , n16173 );
not ( n27365 , n27338 );
or ( n27366 , n27364 , n27365 );
xor ( n27367 , n537 , n25788 );
nand ( n27368 , n27367 , n5697 );
nand ( n27369 , n27366 , n27368 );
xor ( n27370 , n27363 , n27369 );
and ( n27371 , n24800 , n537 );
xor ( n27372 , n27370 , n27371 );
xor ( n27373 , n27361 , n27372 );
xor ( n27374 , n27340 , n27341 );
and ( n27375 , n27374 , n27344 );
and ( n27376 , n27340 , n27341 );
or ( n27377 , n27375 , n27376 );
xor ( n27378 , n27373 , n27377 );
xor ( n27379 , n27331 , n27345 );
and ( n27380 , n27379 , n27350 );
and ( n27381 , n27331 , n27345 );
or ( n27382 , n27380 , n27381 );
or ( n27383 , n27378 , n27382 );
nand ( n27384 , n27360 , n27383 );
nor ( n27385 , n27327 , n27384 );
not ( n27386 , n27385 );
not ( n27387 , n25414 );
or ( n27388 , n27386 , n27387 );
and ( n27389 , n25819 , n27358 );
and ( n27390 , n27356 , n27351 );
nor ( n27391 , n27389 , n27390 );
not ( n27392 , n27391 );
and ( n27393 , n27378 , n27382 );
nor ( n27394 , n27392 , n27393 );
not ( n27395 , n27394 );
not ( n27396 , n25771 );
or ( n27397 , n27395 , n27396 );
not ( n27398 , n27383 );
not ( n27399 , n27393 );
and ( n27400 , n27398 , n27399 );
nor ( n27401 , n27393 , n27360 );
and ( n27402 , n27391 , n27401 );
nor ( n27403 , n27400 , n27402 );
nand ( n27404 , n27397 , n27403 );
nand ( n27405 , n27388 , n27404 );
not ( n27406 , n27367 );
or ( n27407 , n27406 , n24871 );
or ( n27408 , n5604 , n5605 );
nand ( n27409 , n27407 , n27408 );
nand ( n27410 , n9886 , n537 );
xor ( n27411 , n27409 , n27410 );
xor ( n27412 , n27363 , n27369 );
and ( n27413 , n27412 , n27371 );
and ( n27414 , n27363 , n27369 );
or ( n27415 , n27413 , n27414 );
xor ( n27416 , n27411 , n27415 );
not ( n27417 , n27416 );
not ( n27418 , n27417 );
xor ( n27419 , n27361 , n27372 );
and ( n27420 , n27419 , n27377 );
and ( n27421 , n27361 , n27372 );
or ( n27422 , n27420 , n27421 );
not ( n27423 , n27422 );
not ( n27424 , n27423 );
or ( n27425 , n27418 , n27424 );
or ( n27426 , n27423 , n27417 );
nand ( n27427 , n27425 , n27426 );
not ( n27428 , n27427 );
and ( n27429 , n27405 , n27428 );
not ( n27430 , n27405 );
and ( n27431 , n27430 , n27427 );
nor ( n27432 , n27429 , n27431 );
not ( n27433 , n27432 );
or ( n27434 , n27326 , n27433 );
xor ( n27435 , n25704 , n25742 );
and ( n27436 , n27435 , n25747 );
and ( n27437 , n25704 , n25742 );
or ( n27438 , n27436 , n27437 );
not ( n27439 , n27438 );
xor ( n27440 , n25693 , n25698 );
and ( n27441 , n27440 , n25703 );
and ( n27442 , n25693 , n25698 );
or ( n27443 , n27441 , n27442 );
or ( n27444 , n13056 , n13119 );
nand ( n27445 , n27444 , n495 );
not ( n27446 , n12635 );
not ( n27447 , n25721 );
or ( n27448 , n27446 , n27447 );
xor ( n27449 , n489 , n15580 );
nand ( n27450 , n12882 , n27449 );
nand ( n27451 , n27448 , n27450 );
xor ( n27452 , n27445 , n27451 );
and ( n27453 , n12515 , n489 );
xor ( n27454 , n27452 , n27453 );
xor ( n27455 , n25717 , n25723 );
and ( n27456 , n27455 , n25735 );
and ( n27457 , n25717 , n25723 );
or ( n27458 , n27456 , n27457 );
xor ( n27459 , n27454 , n27458 );
not ( n27460 , n12688 );
not ( n27461 , n25713 );
or ( n27462 , n27460 , n27461 );
not ( n27463 , n491 );
not ( n27464 , n24034 );
or ( n27465 , n27463 , n27464 );
nand ( n27466 , n24037 , n12703 );
nand ( n27467 , n27465 , n27466 );
nand ( n27468 , n27467 , n12731 );
nand ( n27469 , n27462 , n27468 );
not ( n27470 , n12845 );
and ( n27471 , n493 , n24043 );
not ( n27472 , n493 );
and ( n27473 , n27472 , n24046 );
nor ( n27474 , n27471 , n27473 );
not ( n27475 , n27474 );
or ( n27476 , n27470 , n27475 );
nand ( n27477 , n25731 , n15386 );
nand ( n27478 , n27476 , n27477 );
xor ( n27479 , n27469 , n27478 );
xor ( n27480 , n27479 , n25692 );
xor ( n27481 , n27459 , n27480 );
xor ( n27482 , n27443 , n27481 );
xor ( n27483 , n25708 , n25736 );
and ( n27484 , n27483 , n25741 );
and ( n27485 , n25708 , n25736 );
or ( n27486 , n27484 , n27485 );
xor ( n27487 , n27482 , n27486 );
not ( n27488 , n27487 );
nand ( n27489 , n27439 , n27488 );
nand ( n27490 , n27489 , n25755 );
xor ( n27491 , n27443 , n27481 );
and ( n27492 , n27491 , n27486 );
and ( n27493 , n27443 , n27481 );
or ( n27494 , n27492 , n27493 );
and ( n27495 , n489 , n17764 );
not ( n27496 , n12731 );
not ( n27497 , n491 );
not ( n27498 , n25727 );
or ( n27499 , n27497 , n27498 );
not ( n27500 , n25727 );
nand ( n27501 , n27500 , n12703 );
nand ( n27502 , n27499 , n27501 );
not ( n27503 , n27502 );
or ( n27504 , n27496 , n27503 );
nand ( n27505 , n27467 , n12688 );
nand ( n27506 , n27504 , n27505 );
xor ( n27507 , n27495 , n27506 );
not ( n27508 , n15386 );
not ( n27509 , n27474 );
or ( n27510 , n27508 , n27509 );
nand ( n27511 , n12845 , n493 );
nand ( n27512 , n27510 , n27511 );
xor ( n27513 , n27507 , n27512 );
buf ( n27514 , n24004 );
and ( n27515 , n27514 , n12653 );
not ( n27516 , n27514 );
and ( n27517 , n27516 , n489 );
or ( n27518 , n27515 , n27517 );
not ( n27519 , n27518 );
nor ( n27520 , n27519 , n12632 );
not ( n27521 , n27449 );
nor ( n27522 , n27521 , n12634 );
nor ( n27523 , n27520 , n27522 );
xor ( n27524 , n27445 , n27451 );
and ( n27525 , n27524 , n27453 );
and ( n27526 , n27445 , n27451 );
or ( n27527 , n27525 , n27526 );
xor ( n27528 , n27523 , n27527 );
xor ( n27529 , n27469 , n27478 );
and ( n27530 , n27529 , n25692 );
and ( n27531 , n27469 , n27478 );
or ( n27532 , n27530 , n27531 );
xor ( n27533 , n27528 , n27532 );
xor ( n27534 , n27513 , n27533 );
xor ( n27535 , n27454 , n27458 );
and ( n27536 , n27535 , n27480 );
and ( n27537 , n27454 , n27458 );
or ( n27538 , n27536 , n27537 );
xor ( n27539 , n27534 , n27538 );
nor ( n27540 , n27494 , n27539 );
nor ( n27541 , n27490 , n27540 );
buf ( n27542 , n27541 );
not ( n27543 , n27542 );
not ( n27544 , n25691 );
or ( n27545 , n27543 , n27544 );
not ( n27546 , n27540 );
not ( n27547 , n27546 );
not ( n27548 , n27489 );
not ( n27549 , n25757 );
or ( n27550 , n27548 , n27549 );
nand ( n27551 , n27438 , n27487 );
nand ( n27552 , n27550 , n27551 );
not ( n27553 , n27552 );
or ( n27554 , n27547 , n27553 );
nand ( n27555 , n27494 , n27539 );
nand ( n27556 , n27554 , n27555 );
not ( n27557 , n27556 );
nand ( n27558 , n27545 , n27557 );
xor ( n27559 , n27513 , n27533 );
and ( n27560 , n27559 , n27538 );
and ( n27561 , n27513 , n27533 );
or ( n27562 , n27560 , n27561 );
not ( n27563 , n27562 );
xor ( n27564 , n27495 , n27506 );
and ( n27565 , n27564 , n27512 );
and ( n27566 , n27495 , n27506 );
or ( n27567 , n27565 , n27566 );
not ( n27568 , n12731 );
and ( n27569 , n491 , n24046 );
not ( n27570 , n491 );
and ( n27571 , n27570 , n24043 );
or ( n27572 , n27569 , n27571 );
not ( n27573 , n27572 );
or ( n27574 , n27568 , n27573 );
nand ( n27575 , n27502 , n12688 );
nand ( n27576 , n27574 , n27575 );
not ( n27577 , n27523 );
xor ( n27578 , n27576 , n27577 );
or ( n27579 , n15386 , n12845 );
nand ( n27580 , n27579 , n493 );
and ( n27581 , n489 , n15580 );
xor ( n27582 , n27580 , n27581 );
not ( n27583 , n12673 );
xor ( n27584 , n489 , n24037 );
not ( n27585 , n27584 );
or ( n27586 , n27583 , n27585 );
nand ( n27587 , n27518 , n12635 );
nand ( n27588 , n27586 , n27587 );
xor ( n27589 , n27582 , n27588 );
xor ( n27590 , n27578 , n27589 );
xor ( n27591 , n27567 , n27590 );
xor ( n27592 , n27523 , n27527 );
and ( n27593 , n27592 , n27532 );
and ( n27594 , n27523 , n27527 );
or ( n27595 , n27593 , n27594 );
xor ( n27596 , n27591 , n27595 );
not ( n27597 , n27596 );
nand ( n27598 , n27563 , n27597 );
buf ( n27599 , n27598 );
not ( n27600 , n27597 );
nand ( n27601 , n27600 , n27562 );
nand ( n27602 , n27599 , n27601 );
not ( n27603 , n27602 );
and ( n27604 , n27558 , n27603 );
not ( n27605 , n27558 );
and ( n27606 , n27605 , n27602 );
nor ( n27607 , n27604 , n27606 );
nand ( n27608 , n27607 , n10190 );
nand ( n27609 , n27434 , n27608 );
xor ( n27610 , n27409 , n27410 );
and ( n27611 , n27610 , n27415 );
and ( n27612 , n27409 , n27410 );
or ( n27613 , n27611 , n27612 );
or ( n27614 , n27423 , n27417 );
nand ( n27615 , n27423 , n27417 );
not ( n27616 , n9248 );
not ( n27617 , n9250 );
nand ( n27618 , n27617 , n9213 );
not ( n27619 , n27618 );
or ( n27620 , n27616 , n27619 );
or ( n27621 , n9248 , n27618 );
nand ( n27622 , n27620 , n27621 );
not ( n27623 , n9243 );
nand ( n27624 , n9222 , n9247 );
not ( n27625 , n27624 );
or ( n27626 , n27623 , n27625 );
or ( n27627 , n9243 , n27624 );
nand ( n27628 , n27626 , n27627 );
xor ( n27629 , n9224 , n9235 );
xor ( n27630 , n27629 , n9241 );
and ( n27631 , n9232 , n9234 );
nor ( n27632 , n27631 , n9235 );
or ( n27633 , n16173 , n5697 );
nand ( n27634 , n27633 , n537 );
not ( n27635 , n27410 );
and ( n27636 , n537 , n25788 );
xor ( n27637 , n27634 , n27636 );
xor ( n27638 , n27637 , n27635 );
not ( n27639 , n20730 );
not ( n27640 , n26004 );
or ( n27641 , n27639 , n27640 );
buf ( n27642 , n26000 );
nand ( n27643 , n27642 , n20745 );
nand ( n27644 , n27641 , n27643 );
not ( n27645 , n27644 );
or ( n27646 , n27645 , n20764 );
or ( n27647 , n21318 , n20745 );
nand ( n27648 , n27646 , n27647 );
not ( n27649 , n26032 );
not ( n27650 , n20710 );
and ( n27651 , n27649 , n27650 );
and ( n27652 , n25969 , n20693 );
nor ( n27653 , n27651 , n27652 );
xor ( n27654 , n27648 , n27653 );
or ( n27655 , n20602 , n20647 );
nand ( n27656 , n27655 , n20628 );
not ( n27657 , n27656 );
not ( n27658 , n21045 );
not ( n27659 , n20474 );
or ( n27660 , n27658 , n27659 );
nand ( n27661 , n26031 , n20693 );
nand ( n27662 , n27660 , n27661 );
not ( n27663 , n27662 );
or ( n27664 , n27657 , n27663 );
or ( n27665 , n27662 , n27656 );
not ( n27666 , n20728 );
not ( n27667 , n27644 );
or ( n27668 , n27666 , n27667 );
not ( n27669 , n20730 );
not ( n27670 , n25970 );
or ( n27671 , n27669 , n27670 );
nand ( n27672 , n25976 , n20745 );
nand ( n27673 , n27671 , n27672 );
nand ( n27674 , n27673 , n20765 );
nand ( n27675 , n27668 , n27674 );
nand ( n27676 , n27665 , n27675 );
nand ( n27677 , n27664 , n27676 );
and ( n27678 , n27654 , n27677 );
and ( n27679 , n27648 , n27653 );
nor ( n27680 , n27678 , n27679 );
and ( n27681 , n20764 , n21318 );
nor ( n27682 , n27681 , n20745 );
xor ( n27683 , n27653 , n27682 );
and ( n27684 , n25969 , n21045 );
and ( n27685 , n27642 , n20693 );
nor ( n27686 , n27684 , n27685 );
xor ( n27687 , n27683 , n27686 );
nand ( n27688 , n27680 , n27687 );
or ( n27689 , n27680 , n27687 );
nand ( n27690 , n27688 , n27689 );
not ( n27691 , n27690 );
not ( n27692 , n20693 );
not ( n27693 , n21394 );
or ( n27694 , n27692 , n27693 );
nand ( n27695 , n21118 , n21045 );
nand ( n27696 , n27694 , n27695 );
not ( n27697 , n20728 );
not ( n27698 , n20730 );
not ( n27699 , n20477 );
or ( n27700 , n27698 , n27699 );
nand ( n27701 , n20474 , n20745 );
nand ( n27702 , n27700 , n27701 );
not ( n27703 , n27702 );
or ( n27704 , n27697 , n27703 );
buf ( n27705 , n20422 );
and ( n27706 , n20730 , n27705 );
not ( n27707 , n20730 );
and ( n27708 , n27707 , n20425 );
nor ( n27709 , n27706 , n27708 );
nand ( n27710 , n27709 , n20765 );
nand ( n27711 , n27704 , n27710 );
xor ( n27712 , n27696 , n27711 );
not ( n27713 , n20647 );
and ( n27714 , n20628 , n25969 );
not ( n27715 , n20628 );
and ( n27716 , n27715 , n25970 );
nor ( n27717 , n27714 , n27716 );
not ( n27718 , n27717 );
or ( n27719 , n27713 , n27718 );
not ( n27720 , n20628 );
not ( n27721 , n26032 );
or ( n27722 , n27720 , n27721 );
nand ( n27723 , n26031 , n20644 );
nand ( n27724 , n27722 , n27723 );
nand ( n27725 , n27724 , n20602 );
nand ( n27726 , n27719 , n27725 );
xor ( n27727 , n27712 , n27726 );
not ( n27728 , n20932 );
not ( n27729 , n20953 );
and ( n27730 , n27728 , n27729 );
not ( n27731 , n20935 );
not ( n27732 , n26004 );
or ( n27733 , n27731 , n27732 );
nand ( n27734 , n27642 , n20953 );
nand ( n27735 , n27733 , n27734 );
and ( n27736 , n27735 , n20980 );
nor ( n27737 , n27730 , n27736 );
or ( n27738 , n21003 , n21334 );
nand ( n27739 , n27738 , n20983 );
not ( n27740 , n20693 );
not ( n27741 , n21118 );
or ( n27742 , n27740 , n27741 );
nand ( n27743 , n21137 , n21045 );
nand ( n27744 , n27742 , n27743 );
xor ( n27745 , n27739 , n27744 );
not ( n27746 , n20765 );
not ( n27747 , n20730 );
not ( n27748 , n21391 );
or ( n27749 , n27747 , n27748 );
nand ( n27750 , n21394 , n20745 );
nand ( n27751 , n27749 , n27750 );
not ( n27752 , n27751 );
or ( n27753 , n27746 , n27752 );
nand ( n27754 , n27709 , n20728 );
nand ( n27755 , n27753 , n27754 );
and ( n27756 , n27745 , n27755 );
and ( n27757 , n27739 , n27744 );
or ( n27758 , n27756 , n27757 );
xor ( n27759 , n27737 , n27758 );
not ( n27760 , n21196 );
not ( n27761 , n20710 );
and ( n27762 , n27760 , n27761 );
and ( n27763 , n21137 , n20693 );
nor ( n27764 , n27762 , n27763 );
not ( n27765 , n27764 );
not ( n27766 , n20933 );
not ( n27767 , n27735 );
or ( n27768 , n27766 , n27767 );
and ( n27769 , n20935 , n25969 );
not ( n27770 , n20935 );
and ( n27771 , n27770 , n25970 );
nor ( n27772 , n27769 , n27771 );
nand ( n27773 , n27772 , n20979 );
nand ( n27774 , n27768 , n27773 );
xor ( n27775 , n27765 , n27774 );
not ( n27776 , n20602 );
not ( n27777 , n20628 );
not ( n27778 , n20477 );
or ( n27779 , n27777 , n27778 );
nand ( n27780 , n20474 , n20644 );
nand ( n27781 , n27779 , n27780 );
not ( n27782 , n27781 );
or ( n27783 , n27776 , n27782 );
nand ( n27784 , n27724 , n20647 );
nand ( n27785 , n27783 , n27784 );
and ( n27786 , n27775 , n27785 );
and ( n27787 , n27765 , n27774 );
or ( n27788 , n27786 , n27787 );
xor ( n27789 , n27759 , n27788 );
xor ( n27790 , n27727 , n27789 );
xor ( n27791 , n27739 , n27744 );
xor ( n27792 , n27791 , n27755 );
xor ( n27793 , n27765 , n27774 );
xor ( n27794 , n27793 , n27785 );
xor ( n27795 , n27792 , n27794 );
not ( n27796 , n21003 );
not ( n27797 , n20983 );
not ( n27798 , n26004 );
or ( n27799 , n27797 , n27798 );
nand ( n27800 , n27642 , n21487 );
nand ( n27801 , n27799 , n27800 );
not ( n27802 , n27801 );
or ( n27803 , n27796 , n27802 );
nand ( n27804 , n21334 , n20983 );
nand ( n27805 , n27803 , n27804 );
not ( n27806 , n20979 );
not ( n27807 , n20935 );
not ( n27808 , n26032 );
or ( n27809 , n27807 , n27808 );
nand ( n27810 , n20953 , n26031 );
nand ( n27811 , n27809 , n27810 );
not ( n27812 , n27811 );
or ( n27813 , n27806 , n27812 );
nand ( n27814 , n27772 , n20933 );
nand ( n27815 , n27813 , n27814 );
xor ( n27816 , n27805 , n27815 );
not ( n27817 , n20728 );
not ( n27818 , n27751 );
or ( n27819 , n27817 , n27818 );
and ( n27820 , n20730 , n21118 );
not ( n27821 , n20730 );
and ( n27822 , n27821 , n21119 );
nor ( n27823 , n27820 , n27822 );
nand ( n27824 , n27823 , n20765 );
nand ( n27825 , n27819 , n27824 );
and ( n27826 , n27816 , n27825 );
and ( n27827 , n27805 , n27815 );
or ( n27828 , n27826 , n27827 );
and ( n27829 , n27795 , n27828 );
and ( n27830 , n27792 , n27794 );
or ( n27831 , n27829 , n27830 );
and ( n27832 , n27790 , n27831 );
and ( n27833 , n27727 , n27789 );
or ( n27834 , n27832 , n27833 );
or ( n27835 , n20980 , n20933 );
nand ( n27836 , n27835 , n20935 );
not ( n27837 , n21045 );
not ( n27838 , n21394 );
or ( n27839 , n27837 , n27838 );
nand ( n27840 , n27705 , n20693 );
nand ( n27841 , n27839 , n27840 );
xor ( n27842 , n27836 , n27841 );
not ( n27843 , n20647 );
and ( n27844 , n20628 , n27642 );
not ( n27845 , n20628 );
and ( n27846 , n27845 , n26004 );
nor ( n27847 , n27844 , n27846 );
not ( n27848 , n27847 );
or ( n27849 , n27843 , n27848 );
nand ( n27850 , n27717 , n20602 );
nand ( n27851 , n27849 , n27850 );
xor ( n27852 , n27842 , n27851 );
xor ( n27853 , n27737 , n27758 );
and ( n27854 , n27853 , n27788 );
and ( n27855 , n27737 , n27758 );
or ( n27856 , n27854 , n27855 );
xor ( n27857 , n27852 , n27856 );
not ( n27858 , n27737 );
and ( n27859 , n20745 , n26031 );
not ( n27860 , n20745 );
and ( n27861 , n27860 , n26032 );
nor ( n27862 , n27859 , n27861 );
nor ( n27863 , n27862 , n21318 );
not ( n27864 , n27702 );
nor ( n27865 , n27864 , n20764 );
or ( n27866 , n27863 , n27865 );
xor ( n27867 , n27858 , n27866 );
xor ( n27868 , n27696 , n27711 );
and ( n27869 , n27868 , n27726 );
and ( n27870 , n27696 , n27711 );
or ( n27871 , n27869 , n27870 );
xor ( n27872 , n27867 , n27871 );
xor ( n27873 , n27857 , n27872 );
nor ( n27874 , n27834 , n27873 );
not ( n27875 , n27874 );
not ( n27876 , n20647 );
not ( n27877 , n27781 );
or ( n27878 , n27876 , n27877 );
not ( n27879 , n20628 );
not ( n27880 , n20425 );
or ( n27881 , n27879 , n27880 );
nand ( n27882 , n27705 , n20644 );
nand ( n27883 , n27881 , n27882 );
nand ( n27884 , n27883 , n20602 );
nand ( n27885 , n27878 , n27884 );
xor ( n27886 , n27764 , n27885 );
or ( n27887 , n20860 , n20905 );
nand ( n27888 , n27887 , n21213 );
not ( n27889 , n21045 );
not ( n27890 , n21178 );
or ( n27891 , n27889 , n27890 );
nand ( n27892 , n20693 , n21193 );
nand ( n27893 , n27891 , n27892 );
xor ( n27894 , n27888 , n27893 );
not ( n27895 , n20728 );
not ( n27896 , n27823 );
or ( n27897 , n27895 , n27896 );
and ( n27898 , n20730 , n21137 );
not ( n27899 , n20730 );
and ( n27900 , n27899 , n21138 );
nor ( n27901 , n27898 , n27900 );
nand ( n27902 , n27901 , n20765 );
nand ( n27903 , n27897 , n27902 );
and ( n27904 , n27894 , n27903 );
and ( n27905 , n27888 , n27893 );
or ( n27906 , n27904 , n27905 );
and ( n27907 , n27886 , n27906 );
and ( n27908 , n27764 , n27885 );
or ( n27909 , n27907 , n27908 );
xor ( n27910 , n27792 , n27794 );
xor ( n27911 , n27910 , n27828 );
xor ( n27912 , n27909 , n27911 );
not ( n27913 , n21334 );
not ( n27914 , n27801 );
or ( n27915 , n27913 , n27914 );
not ( n27916 , n20983 );
not ( n27917 , n25970 );
or ( n27918 , n27916 , n27917 );
nand ( n27919 , n25976 , n21487 );
nand ( n27920 , n27918 , n27919 );
nand ( n27921 , n27920 , n21003 );
nand ( n27922 , n27915 , n27921 );
not ( n27923 , n20980 );
not ( n27924 , n20935 );
not ( n27925 , n20477 );
or ( n27926 , n27924 , n27925 );
nand ( n27927 , n20474 , n20953 );
nand ( n27928 , n27926 , n27927 );
not ( n27929 , n27928 );
or ( n27930 , n27923 , n27929 );
nand ( n27931 , n27811 , n20933 );
nand ( n27932 , n27930 , n27931 );
xor ( n27933 , n27922 , n27932 );
not ( n27934 , n20602 );
not ( n27935 , n20628 );
not ( n27936 , n21391 );
or ( n27937 , n27935 , n27936 );
nand ( n27938 , n21394 , n20644 );
nand ( n27939 , n27937 , n27938 );
not ( n27940 , n27939 );
or ( n27941 , n27934 , n27940 );
nand ( n27942 , n27883 , n20647 );
nand ( n27943 , n27941 , n27942 );
and ( n27944 , n27933 , n27943 );
and ( n27945 , n27922 , n27932 );
or ( n27946 , n27944 , n27945 );
xor ( n27947 , n27805 , n27815 );
xor ( n27948 , n27947 , n27825 );
xor ( n27949 , n27946 , n27948 );
xor ( n27950 , n27764 , n27885 );
xor ( n27951 , n27950 , n27906 );
and ( n27952 , n27949 , n27951 );
and ( n27953 , n27946 , n27948 );
or ( n27954 , n27952 , n27953 );
and ( n27955 , n27912 , n27954 );
and ( n27956 , n27909 , n27911 );
or ( n27957 , n27955 , n27956 );
xor ( n27958 , n27727 , n27789 );
xor ( n27959 , n27958 , n27831 );
or ( n27960 , n27957 , n27959 );
nand ( n27961 , n27875 , n27960 );
xor ( n27962 , n27836 , n27841 );
and ( n27963 , n27962 , n27851 );
and ( n27964 , n27836 , n27841 );
or ( n27965 , n27963 , n27964 );
not ( n27966 , n20765 );
not ( n27967 , n27862 );
not ( n27968 , n27967 );
or ( n27969 , n27966 , n27968 );
nand ( n27970 , n27673 , n20728 );
nand ( n27971 , n27969 , n27970 );
not ( n27972 , n27971 );
not ( n27973 , n20425 );
not ( n27974 , n20710 );
and ( n27975 , n27973 , n27974 );
and ( n27976 , n20474 , n20693 );
nor ( n27977 , n27975 , n27976 );
not ( n27978 , n27977 );
and ( n27979 , n27972 , n27978 );
and ( n27980 , n27971 , n27977 );
nor ( n27981 , n27979 , n27980 );
not ( n27982 , n27847 );
not ( n27983 , n20602 );
or ( n27984 , n27982 , n27983 );
nand ( n27985 , n20647 , n20628 );
nand ( n27986 , n27984 , n27985 );
and ( n27987 , n27981 , n27986 );
not ( n27988 , n27981 );
not ( n27989 , n27986 );
and ( n27990 , n27988 , n27989 );
nor ( n27991 , n27987 , n27990 );
xor ( n27992 , n27965 , n27991 );
xor ( n27993 , n27858 , n27866 );
and ( n27994 , n27993 , n27871 );
and ( n27995 , n27858 , n27866 );
or ( n27996 , n27994 , n27995 );
xor ( n27997 , n27992 , n27996 );
xor ( n27998 , n27852 , n27856 );
and ( n27999 , n27998 , n27872 );
and ( n28000 , n27852 , n27856 );
or ( n28001 , n27999 , n28000 );
or ( n28002 , n27997 , n28001 );
xor ( n28003 , n27656 , n27662 );
xnor ( n28004 , n28003 , n27675 );
and ( n28005 , n28004 , n27986 );
not ( n28006 , n28004 );
and ( n28007 , n28006 , n27989 );
or ( n28008 , n28005 , n28007 );
not ( n28009 , n27977 );
not ( n28010 , n27986 );
or ( n28011 , n28009 , n28010 );
nand ( n28012 , n28011 , n27971 );
not ( n28013 , n27977 );
nand ( n28014 , n28013 , n27989 );
and ( n28015 , n28012 , n28014 );
xnor ( n28016 , n28008 , n28015 );
xor ( n28017 , n27965 , n27991 );
and ( n28018 , n28017 , n27996 );
and ( n28019 , n27965 , n27991 );
or ( n28020 , n28018 , n28019 );
or ( n28021 , n28016 , n28020 );
xor ( n28022 , n27648 , n27653 );
xor ( n28023 , n28022 , n27677 );
not ( n28024 , n28023 );
not ( n28025 , n28004 );
not ( n28026 , n27989 );
and ( n28027 , n28025 , n28026 );
and ( n28028 , n28004 , n27989 );
nor ( n28029 , n28028 , n28015 );
nor ( n28030 , n28027 , n28029 );
nand ( n28031 , n28024 , n28030 );
nand ( n28032 , n28002 , n28021 , n28031 );
nor ( n28033 , n27961 , n28032 );
not ( n28034 , n28033 );
not ( n28035 , n20765 );
not ( n28036 , n27214 );
or ( n28037 , n28035 , n28036 );
nand ( n28038 , n27901 , n20728 );
nand ( n28039 , n28037 , n28038 );
xor ( n28040 , n27888 , n27893 );
xor ( n28041 , n28040 , n27903 );
xor ( n28042 , n28039 , n28041 );
not ( n28043 , n20647 );
not ( n28044 , n27939 );
or ( n28045 , n28043 , n28044 );
nand ( n28046 , n27199 , n20602 );
nand ( n28047 , n28045 , n28046 );
not ( n28048 , n20900 );
not ( n28049 , n20710 );
and ( n28050 , n28048 , n28049 );
and ( n28051 , n21178 , n20693 );
nor ( n28052 , n28050 , n28051 );
not ( n28053 , n28052 );
nor ( n28054 , n28047 , n28053 );
not ( n28055 , n20860 );
not ( n28056 , n27252 );
or ( n28057 , n28055 , n28056 );
nand ( n28058 , n20905 , n21213 );
nand ( n28059 , n28057 , n28058 );
not ( n28060 , n28059 );
or ( n28061 , n28054 , n28060 );
nand ( n28062 , n28047 , n28053 );
nand ( n28063 , n28061 , n28062 );
and ( n28064 , n28042 , n28063 );
and ( n28065 , n28039 , n28041 );
or ( n28066 , n28064 , n28065 );
xor ( n28067 , n27946 , n27948 );
xor ( n28068 , n28067 , n27951 );
xor ( n28069 , n28066 , n28068 );
xor ( n28070 , n27922 , n27932 );
xor ( n28071 , n28070 , n27943 );
not ( n28072 , n28071 );
and ( n28073 , n27920 , n21334 );
and ( n28074 , n27242 , n21003 );
nor ( n28075 , n28073 , n28074 );
xor ( n28076 , n28039 , n28075 );
and ( n28077 , n27223 , n20979 );
and ( n28078 , n27928 , n20933 );
nor ( n28079 , n28077 , n28078 );
and ( n28080 , n28076 , n28079 );
and ( n28081 , n28039 , n28075 );
or ( n28082 , n28080 , n28081 );
nand ( n28083 , n28072 , n28082 );
not ( n28084 , n28083 );
xor ( n28085 , n28039 , n28041 );
xor ( n28086 , n28085 , n28063 );
not ( n28087 , n28086 );
or ( n28088 , n28084 , n28087 );
not ( n28089 , n28082 );
nand ( n28090 , n28089 , n28071 );
nand ( n28091 , n28088 , n28090 );
xor ( n28092 , n28069 , n28091 );
xor ( n28093 , n28082 , n28071 );
xor ( n28094 , n28093 , n28086 );
not ( n28095 , n28094 );
not ( n28096 , n28095 );
not ( n28097 , n27185 );
not ( n28098 , n27203 );
not ( n28099 , n28098 );
or ( n28100 , n28097 , n28099 );
nand ( n28101 , n28100 , n27188 );
not ( n28102 , n27185 );
nand ( n28103 , n28102 , n27203 );
and ( n28104 , n28101 , n28103 );
not ( n28105 , n28104 );
not ( n28106 , n28105 );
xor ( n28107 , n28039 , n28075 );
xor ( n28108 , n28107 , n28079 );
not ( n28109 , n28108 );
not ( n28110 , n28109 );
or ( n28111 , n28106 , n28110 );
not ( n28112 , n28104 );
not ( n28113 , n28108 );
or ( n28114 , n28112 , n28113 );
xor ( n28115 , n25863 , n27216 );
and ( n28116 , n28115 , n27227 );
and ( n28117 , n25863 , n27216 );
or ( n28118 , n28116 , n28117 );
nand ( n28119 , n28114 , n28118 );
nand ( n28120 , n28111 , n28119 );
not ( n28121 , n28120 );
or ( n28122 , n28096 , n28121 );
not ( n28123 , n28120 );
not ( n28124 , n28123 );
not ( n28125 , n28094 );
or ( n28126 , n28124 , n28125 );
xor ( n28127 , n27244 , n27254 );
and ( n28128 , n28127 , n27259 );
and ( n28129 , n27244 , n27254 );
or ( n28130 , n28128 , n28129 );
not ( n28131 , n28130 );
xor ( n28132 , n28059 , n28052 );
xor ( n28133 , n28132 , n28047 );
nand ( n28134 , n28131 , n28133 );
not ( n28135 , n28134 );
xor ( n28136 , n27207 , n27228 );
and ( n28137 , n28136 , n27233 );
and ( n28138 , n27207 , n27228 );
or ( n28139 , n28137 , n28138 );
not ( n28140 , n28139 );
or ( n28141 , n28135 , n28140 );
not ( n28142 , n28133 );
nand ( n28143 , n28142 , n28130 );
nand ( n28144 , n28141 , n28143 );
nand ( n28145 , n28126 , n28144 );
nand ( n28146 , n28122 , n28145 );
or ( n28147 , n28092 , n28146 );
xor ( n28148 , n28066 , n28068 );
and ( n28149 , n28148 , n28091 );
and ( n28150 , n28066 , n28068 );
or ( n28151 , n28149 , n28150 );
xor ( n28152 , n27909 , n27911 );
xor ( n28153 , n28152 , n27954 );
nor ( n28154 , n28151 , n28153 );
not ( n28155 , n28154 );
and ( n28156 , n28147 , n28155 );
not ( n28157 , n28156 );
and ( n28158 , n28118 , n28104 );
not ( n28159 , n28118 );
and ( n28160 , n28159 , n28105 );
nor ( n28161 , n28158 , n28160 );
and ( n28162 , n28161 , n28109 );
not ( n28163 , n28161 );
and ( n28164 , n28163 , n28108 );
nor ( n28165 , n28162 , n28164 );
not ( n28166 , n28130 );
not ( n28167 , n28133 );
and ( n28168 , n28166 , n28167 );
and ( n28169 , n28130 , n28133 );
nor ( n28170 , n28168 , n28169 );
xor ( n28171 , n28139 , n28170 );
xor ( n28172 , n28165 , n28171 );
not ( n28173 , n27260 );
nand ( n28174 , n28173 , n27265 );
and ( n28175 , n27270 , n28174 );
nor ( n28176 , n28173 , n27265 );
nor ( n28177 , n28175 , n28176 );
xor ( n28178 , n28172 , n28177 );
or ( n28179 , n27234 , n27271 );
and ( n28180 , n28179 , n27276 );
and ( n28181 , n27234 , n27271 );
nor ( n28182 , n28180 , n28181 );
nand ( n28183 , n28178 , n28182 );
and ( n28184 , n28144 , n28120 );
not ( n28185 , n28144 );
and ( n28186 , n28185 , n28123 );
nor ( n28187 , n28184 , n28186 );
and ( n28188 , n28187 , n28094 );
not ( n28189 , n28187 );
and ( n28190 , n28189 , n28095 );
nor ( n28191 , n28188 , n28190 );
xor ( n28192 , n28165 , n28171 );
and ( n28193 , n28192 , n28177 );
and ( n28194 , n28165 , n28171 );
or ( n28195 , n28193 , n28194 );
nand ( n28196 , n28191 , n28195 );
nand ( n28197 , n26497 , n27284 , n28183 , n28196 );
not ( n28198 , n28197 );
not ( n28199 , n28198 );
not ( n28200 , n27290 );
or ( n28201 , n28199 , n28200 );
not ( n28202 , n28196 );
not ( n28203 , n28183 );
or ( n28204 , n26498 , n27283 );
nand ( n28205 , n28204 , n27282 );
not ( n28206 , n28205 );
or ( n28207 , n28203 , n28206 );
or ( n28208 , n28178 , n28182 );
nand ( n28209 , n28207 , n28208 );
not ( n28210 , n28209 );
or ( n28211 , n28202 , n28210 );
or ( n28212 , n28191 , n28195 );
nand ( n28213 , n28211 , n28212 );
not ( n28214 , n28213 );
nand ( n28215 , n28201 , n28214 );
not ( n28216 , n28215 );
or ( n28217 , n28157 , n28216 );
nand ( n28218 , n28092 , n28146 );
or ( n28219 , n28218 , n28154 );
nand ( n28220 , n28151 , n28153 );
nand ( n28221 , n28219 , n28220 );
not ( n28222 , n28221 );
nand ( n28223 , n28217 , n28222 );
not ( n28224 , n28223 );
or ( n28225 , n28034 , n28224 );
nand ( n28226 , n27957 , n27959 );
not ( n28227 , n28226 );
not ( n28228 , n27874 );
and ( n28229 , n28227 , n28228 );
and ( n28230 , n27834 , n27873 );
nor ( n28231 , n28229 , n28230 );
or ( n28232 , n28231 , n28032 );
nand ( n28233 , n27997 , n28001 );
nor ( n28234 , n28016 , n28020 );
or ( n28235 , n28233 , n28234 );
nand ( n28236 , n28016 , n28020 );
nand ( n28237 , n28235 , n28236 );
and ( n28238 , n28237 , n28031 );
not ( n28239 , n28023 );
nor ( n28240 , n28239 , n28030 );
nor ( n28241 , n28238 , n28240 );
nand ( n28242 , n28232 , n28241 );
not ( n28243 , n28242 );
nand ( n28244 , n28225 , n28243 );
not ( n28245 , n28244 );
or ( n28246 , n27691 , n28245 );
or ( n28247 , n28244 , n27690 );
nand ( n28248 , n28246 , n28247 );
nor ( n28249 , n27291 , n27283 );
nor ( n28250 , n28249 , n28205 );
not ( n28251 , n28250 );
nand ( n28252 , n28251 , n28183 );
nand ( n28253 , n28252 , n28208 );
not ( n28254 , n26926 );
or ( n28255 , n27080 , n28254 );
nand ( n28256 , n28255 , n27014 );
not ( n28257 , n27002 );
or ( n28258 , n28257 , n26849 );
nand ( n28259 , n28258 , n27006 );
not ( n28260 , n23833 );
nand ( n28261 , n28260 , n21841 );
not ( n28262 , n28261 );
not ( n28263 , n23828 );
not ( n28264 , n22113 );
or ( n28265 , n28263 , n28264 );
not ( n28266 , n23831 );
nand ( n28267 , n28265 , n28266 );
not ( n28268 , n28267 );
or ( n28269 , n28262 , n28268 );
or ( n28270 , n28267 , n28261 );
nand ( n28271 , n28269 , n28270 );
nor ( n28272 , n23831 , n28264 );
and ( n28273 , n28272 , n23828 );
not ( n28274 , n28272 );
and ( n28275 , n28274 , n28263 );
nor ( n28276 , n28273 , n28275 );
and ( n28277 , n23809 , n23929 );
nor ( n28278 , n28277 , n23813 );
xor ( n28279 , n22816 , n22818 );
xor ( n28280 , n28279 , n23806 );
not ( n28281 , n23812 );
nor ( n28282 , n28281 , n23815 );
not ( n28283 , n27006 );
nor ( n28284 , n28283 , n26849 );
not ( n28285 , n26891 );
nand ( n28286 , n28285 , n27008 );
nand ( n28287 , n26976 , n27146 );
xor ( n28288 , n23432 , n23434 );
xor ( n28289 , n28288 , n23691 );
not ( n28290 , n27017 );
nand ( n28291 , n28290 , n26935 );
nand ( n28292 , n28156 , n28033 , n27688 );
nor ( n28293 , n28292 , n28197 );
and ( n28294 , n28033 , n28221 );
nor ( n28295 , n28294 , n28242 );
not ( n28296 , n27688 );
or ( n28297 , n28295 , n28296 );
nand ( n28298 , n28297 , n27689 );
nand ( n28299 , n28212 , n28196 );
and ( n28300 , n28208 , n28183 );
nor ( n28301 , n28230 , n27874 );
not ( n28302 , n28226 );
not ( n28303 , n27960 );
nor ( n28304 , n28302 , n28303 );
not ( n28305 , n23664 );
nand ( n28306 , n23674 , n23677 );
not ( n28307 , n28306 );
or ( n28308 , n28305 , n28307 );
or ( n28309 , n28306 , n23664 );
nand ( n28310 , n28308 , n28309 );
nand ( n28311 , n28002 , n28233 );
nand ( n28312 , n28021 , n28236 );
xor ( n28313 , n23624 , n23631 );
xor ( n28314 , n28313 , n23654 );
nor ( n28315 , n26004 , n20710 );
not ( n28316 , n28315 );
xor ( n28317 , n27653 , n27682 );
and ( n28318 , n28317 , n27686 );
and ( n28319 , n27653 , n27682 );
or ( n28320 , n28318 , n28319 );
not ( n28321 , n28320 );
or ( n28322 , n28316 , n28321 );
or ( n28323 , n28320 , n28315 );
nand ( n28324 , n28322 , n28323 );
xor ( n28325 , n23633 , n23646 );
xor ( n28326 , n28325 , n23652 );
not ( n28327 , n28002 );
not ( n28328 , n27961 );
nand ( n28329 , n28328 , n28223 );
nand ( n28330 , n28329 , n28231 );
not ( n28331 , n28330 );
or ( n28332 , n28327 , n28331 );
nand ( n28333 , n28332 , n28233 );
xnor ( n28334 , n28333 , n28312 );
xor ( n28335 , n27580 , n27581 );
and ( n28336 , n28335 , n27588 );
and ( n28337 , n27580 , n27581 );
or ( n28338 , n28336 , n28337 );
xor ( n28339 , n27576 , n27577 );
and ( n28340 , n28339 , n27589 );
and ( n28341 , n27576 , n27577 );
or ( n28342 , n28340 , n28341 );
xor ( n28343 , n27567 , n27590 );
and ( n28344 , n28343 , n27595 );
and ( n28345 , n27567 , n27590 );
or ( n28346 , n28344 , n28345 );
not ( n28347 , n12673 );
not ( n28348 , n489 );
not ( n28349 , n25727 );
or ( n28350 , n28348 , n28349 );
nand ( n28351 , n27500 , n12653 );
nand ( n28352 , n28350 , n28351 );
not ( n28353 , n28352 );
or ( n28354 , n28347 , n28353 );
nand ( n28355 , n27584 , n12635 );
nand ( n28356 , n28354 , n28355 );
not ( n28357 , n12688 );
not ( n28358 , n27572 );
or ( n28359 , n28357 , n28358 );
nand ( n28360 , n12731 , n491 );
nand ( n28361 , n28359 , n28360 );
xor ( n28362 , n28356 , n28361 );
nand ( n28363 , n27514 , n489 );
xor ( n28364 , n28362 , n28363 );
xor ( n28365 , n28356 , n28361 );
and ( n28366 , n28365 , n28363 );
and ( n28367 , n28356 , n28361 );
or ( n28368 , n28366 , n28367 );
xor ( n28369 , n28338 , n28364 );
xor ( n28370 , n28369 , n28342 );
xor ( n28371 , n28338 , n28364 );
and ( n28372 , n28371 , n28342 );
and ( n28373 , n28338 , n28364 );
or ( n28374 , n28372 , n28373 );
or ( n28375 , n12688 , n12731 );
nand ( n28376 , n28375 , n491 );
and ( n28377 , n489 , n24037 );
xor ( n28378 , n28376 , n28377 );
not ( n28379 , n12673 );
xor ( n28380 , n489 , n24043 );
not ( n28381 , n28380 );
or ( n28382 , n28379 , n28381 );
nand ( n28383 , n28352 , n12635 );
nand ( n28384 , n28382 , n28383 );
xor ( n28385 , n28378 , n28384 );
xor ( n28386 , n28376 , n28377 );
and ( n28387 , n28386 , n28384 );
and ( n28388 , n28376 , n28377 );
or ( n28389 , n28387 , n28388 );
not ( n28390 , n28363 );
xor ( n28391 , n28390 , n28385 );
xor ( n28392 , n28391 , n28368 );
xor ( n28393 , n28390 , n28385 );
and ( n28394 , n28393 , n28368 );
and ( n28395 , n28390 , n28385 );
or ( n28396 , n28394 , n28395 );
not ( n28397 , n28380 );
or ( n28398 , n28397 , n12634 );
or ( n28399 , n12632 , n12653 );
nand ( n28400 , n28398 , n28399 );
nand ( n28401 , n27500 , n489 );
xor ( n28402 , n28400 , n28401 );
xor ( n28403 , n28402 , n28389 );
xor ( n28404 , n28400 , n28401 );
and ( n28405 , n28404 , n28389 );
and ( n28406 , n28400 , n28401 );
or ( n28407 , n28405 , n28406 );
not ( n28408 , n28346 );
not ( n28409 , n28370 );
nand ( n28410 , n28408 , n28409 );
nand ( n28411 , n27598 , n28410 );
nor ( n28412 , n28374 , n28392 );
nor ( n28413 , n28411 , n28412 );
and ( n28414 , n28413 , n27541 );
nand ( n28415 , n28414 , n25689 );
nand ( n28416 , n27489 , n27551 );
not ( n28417 , n28412 );
not ( n28418 , n28417 );
not ( n28419 , n28410 );
or ( n28420 , n28419 , n27601 );
not ( n28421 , n28409 );
nand ( n28422 , n28421 , n28346 );
nand ( n28423 , n28420 , n28422 );
not ( n28424 , n28423 );
or ( n28425 , n28418 , n28424 );
nand ( n28426 , n28374 , n28392 );
nand ( n28427 , n28425 , n28426 );
not ( n28428 , n28427 );
nand ( n28429 , n28410 , n28422 );
not ( n28430 , n15068 );
not ( n28431 , n15021 );
nand ( n28432 , n28431 , n15071 );
not ( n28433 , n28432 );
or ( n28434 , n28430 , n28433 );
or ( n28435 , n28432 , n15068 );
nand ( n28436 , n28434 , n28435 );
nand ( n28437 , n28396 , n28403 );
xor ( n28438 , n15027 , n15037 );
xor ( n28439 , n28438 , n15065 );
or ( n28440 , n15045 , n15048 );
nand ( n28441 , n28440 , n15049 );
not ( n28442 , n28441 );
or ( n28443 , n12635 , n12882 );
nand ( n28444 , n28443 , n489 );
not ( n28445 , n28401 );
and ( n28446 , n489 , n24043 );
xor ( n28447 , n28444 , n28446 );
xor ( n28448 , n28447 , n28445 );
xor ( n28449 , n25840 , n25841 );
and ( n28450 , n28449 , n25843 );
and ( n28451 , n25840 , n25841 );
or ( n28452 , n28450 , n28451 );
xor ( n28453 , n25671 , n25675 );
and ( n28454 , n28453 , n25844 );
and ( n28455 , n25671 , n25675 );
or ( n28456 , n28454 , n28455 );
nand ( n28457 , n25836 , n25765 );
and ( n28458 , n28457 , n471 );
and ( n28459 , n25395 , n469 );
xor ( n28460 , n28458 , n28459 );
and ( n28461 , n25261 , n470 );
xor ( n28462 , n28460 , n28461 );
xor ( n28463 , n28458 , n28459 );
and ( n28464 , n28463 , n28461 );
and ( n28465 , n28458 , n28459 );
or ( n28466 , n28464 , n28465 );
not ( n28467 , n10190 );
not ( n28468 , n25756 );
not ( n28469 , n25691 );
or ( n28470 , n28468 , n28469 );
nand ( n28471 , n28470 , n25758 );
xnor ( n28472 , n28471 , n28416 );
not ( n28473 , n28472 );
or ( n28474 , n28467 , n28473 );
not ( n28475 , n27390 );
nand ( n28476 , n28475 , n27358 );
nand ( n28477 , n28476 , n454 );
not ( n28478 , n28477 );
nor ( n28479 , n27327 , n25821 );
not ( n28480 , n28479 );
not ( n28481 , n25409 );
not ( n28482 , n24691 );
or ( n28483 , n28481 , n28482 );
nand ( n28484 , n28483 , n25413 );
not ( n28485 , n28484 );
or ( n28486 , n28480 , n28485 );
and ( n28487 , n25770 , n25822 );
nor ( n28488 , n28487 , n25819 );
nand ( n28489 , n28486 , n28488 );
not ( n28490 , n28489 );
or ( n28491 , n28478 , n28490 );
not ( n28492 , n454 );
nor ( n28493 , n28492 , n28476 );
or ( n28494 , n28489 , n28493 );
nand ( n28495 , n28491 , n28494 );
nand ( n28496 , n28474 , n28495 );
and ( n28497 , n28496 , n472 );
xor ( n28498 , n28497 , n28452 );
xor ( n28499 , n28498 , n28462 );
xor ( n28500 , n28497 , n28452 );
and ( n28501 , n28500 , n28462 );
and ( n28502 , n28497 , n28452 );
or ( n28503 , n28501 , n28502 );
nand ( n28504 , n25836 , n25765 );
and ( n28505 , n28504 , n470 );
not ( n28506 , n25261 );
nor ( n28507 , n28506 , n16080 );
xor ( n28508 , n28505 , n28507 );
not ( n28509 , n27490 );
not ( n28510 , n28509 );
not ( n28511 , n25678 );
not ( n28512 , n24579 );
or ( n28513 , n28511 , n28512 );
nand ( n28514 , n28513 , n25690 );
not ( n28515 , n28514 );
or ( n28516 , n28510 , n28515 );
not ( n28517 , n27552 );
buf ( n28518 , n28517 );
nand ( n28519 , n28516 , n28518 );
nand ( n28520 , n27546 , n27555 );
nand ( n28521 , n28520 , n10190 );
and ( n28522 , n28519 , n28521 );
not ( n28523 , n28519 );
not ( n28524 , n28520 );
nand ( n28525 , n28524 , n10190 );
and ( n28526 , n28523 , n28525 );
or ( n28527 , n28522 , n28526 );
not ( n28528 , n25253 );
nand ( n28529 , n28528 , n27360 );
nand ( n28530 , n27391 , n28529 );
and ( n28531 , n27360 , n25252 );
or ( n28532 , n28530 , n28531 );
not ( n28533 , n28532 );
nor ( n28534 , n28530 , n25205 );
nand ( n28535 , n25200 , n25179 , n28534 );
not ( n28536 , n28535 );
or ( n28537 , n28533 , n28536 );
nand ( n28538 , n27378 , n27382 );
nand ( n28539 , n27383 , n28538 );
not ( n28540 , n28539 );
nand ( n28541 , n28537 , n28540 );
not ( n28542 , n28541 );
nand ( n28543 , n28542 , n454 );
not ( n28544 , n28535 );
and ( n28545 , n28539 , n454 );
nand ( n28546 , n28532 , n28545 );
nor ( n28547 , n28544 , n28546 );
not ( n28548 , n28547 );
nand ( n28549 , n28527 , n28543 , n28548 );
and ( n28550 , n28549 , n472 );
xor ( n28551 , n28508 , n28550 );
xor ( n28552 , n28505 , n28507 );
and ( n28553 , n28552 , n28550 );
and ( n28554 , n28505 , n28507 );
or ( n28555 , n28553 , n28554 );
and ( n28556 , n28496 , n471 );
xor ( n28557 , n28556 , n28466 );
xor ( n28558 , n28557 , n28551 );
xor ( n28559 , n28556 , n28466 );
and ( n28560 , n28559 , n28551 );
and ( n28561 , n28556 , n28466 );
or ( n28562 , n28560 , n28561 );
and ( n28563 , n28504 , n469 );
and ( n28564 , n28532 , n28535 );
nand ( n28565 , n28540 , n454 );
nor ( n28566 , n28564 , n28565 );
nor ( n28567 , n28566 , n28547 );
nand ( n28568 , n28567 , n28527 );
and ( n28569 , n28568 , n471 );
xor ( n28570 , n28563 , n28569 );
and ( n28571 , n28496 , n470 );
xor ( n28572 , n28570 , n28571 );
xor ( n28573 , n28563 , n28569 );
and ( n28574 , n28573 , n28571 );
and ( n28575 , n28563 , n28569 );
or ( n28576 , n28574 , n28575 );
and ( n28577 , n27609 , n472 );
xor ( n28578 , n28577 , n28555 );
xor ( n28579 , n28578 , n28572 );
xor ( n28580 , n28577 , n28555 );
and ( n28581 , n28580 , n28572 );
and ( n28582 , n28577 , n28555 );
or ( n28583 , n28581 , n28582 );
not ( n28584 , n10190 );
not ( n28585 , n28514 );
not ( n28586 , n27601 );
nor ( n28587 , n28586 , n28429 );
nand ( n28588 , n28585 , n27557 , n28587 );
and ( n28589 , n28429 , n27599 );
and ( n28590 , n28589 , n27541 );
and ( n28591 , n28514 , n28590 );
or ( n28592 , n28429 , n27599 );
and ( n28593 , n27601 , n28592 );
not ( n28594 , n27601 );
not ( n28595 , n28429 );
and ( n28596 , n28594 , n28595 );
nor ( n28597 , n28593 , n28596 );
nor ( n28598 , n28591 , n28597 );
nand ( n28599 , n28595 , n27601 );
nor ( n28600 , n28599 , n27542 );
and ( n28601 , n27557 , n28600 );
not ( n28602 , n27557 );
and ( n28603 , n28602 , n28589 );
nor ( n28604 , n28601 , n28603 );
nand ( n28605 , n28588 , n28598 , n28604 );
not ( n28606 , n28605 );
or ( n28607 , n28584 , n28606 );
xnor ( n28608 , n27613 , n27638 );
not ( n28609 , n28608 );
nand ( n28610 , n28609 , n454 );
nor ( n28611 , n27615 , n28610 );
and ( n28612 , n27614 , n28611 );
not ( n28613 , n27614 );
nand ( n28614 , n28608 , n454 );
not ( n28615 , n28614 );
and ( n28616 , n28613 , n28615 );
nor ( n28617 , n28612 , n28616 );
not ( n28618 , n28617 );
not ( n28619 , n27615 );
nor ( n28620 , n28619 , n28614 );
nor ( n28621 , n28618 , n28620 );
not ( n28622 , n28621 );
not ( n28623 , n27405 );
or ( n28624 , n28622 , n28623 );
nand ( n28625 , n27385 , n28484 );
not ( n28626 , n28610 );
nand ( n28627 , n28626 , n27614 );
and ( n28628 , n28617 , n28627 );
nand ( n28629 , n28625 , n27404 , n28628 );
nand ( n28630 , n28624 , n28629 );
nand ( n28631 , n28607 , n28630 );
and ( n28632 , n28631 , n472 );
and ( n28633 , n28496 , n469 );
xor ( n28634 , n28632 , n28633 );
and ( n28635 , n28549 , n470 );
xor ( n28636 , n28634 , n28635 );
xor ( n28637 , n28632 , n28633 );
and ( n28638 , n28637 , n28635 );
and ( n28639 , n28632 , n28633 );
or ( n28640 , n28638 , n28639 );
and ( n28641 , n27609 , n471 );
xor ( n28642 , n28641 , n28576 );
xor ( n28643 , n28642 , n28636 );
xor ( n28644 , n28641 , n28576 );
and ( n28645 , n28644 , n28636 );
and ( n28646 , n28641 , n28576 );
or ( n28647 , n28645 , n28646 );
nor ( n28648 , n28411 , n27540 );
not ( n28649 , n28648 );
not ( n28650 , n28519 );
or ( n28651 , n28649 , n28650 );
and ( n28652 , n28417 , n28426 );
not ( n28653 , n28652 );
not ( n28654 , n28411 );
not ( n28655 , n28654 );
not ( n28656 , n27555 );
not ( n28657 , n28656 );
or ( n28658 , n28655 , n28657 );
not ( n28659 , n28423 );
nand ( n28660 , n28658 , n28659 );
nor ( n28661 , n28653 , n28660 );
nand ( n28662 , n28651 , n28661 );
not ( n28663 , n28509 );
not ( n28664 , n28514 );
or ( n28665 , n28663 , n28664 );
nand ( n28666 , n28665 , n28517 );
not ( n28667 , n28648 );
nor ( n28668 , n28667 , n28652 );
and ( n28669 , n28666 , n28668 );
not ( n28670 , n28660 );
nor ( n28671 , n28670 , n28652 );
nor ( n28672 , n28669 , n28671 );
nand ( n28673 , n28662 , n28672 );
and ( n28674 , n28673 , n472 , n10190 );
and ( n28675 , n469 , n28568 );
xor ( n28676 , n28674 , n28675 );
and ( n28677 , n27609 , n470 );
xor ( n28678 , n28676 , n28677 );
xor ( n28679 , n28674 , n28675 );
and ( n28680 , n28679 , n28677 );
and ( n28681 , n28674 , n28675 );
or ( n28682 , n28680 , n28681 );
buf ( n28683 , n28631 );
and ( n28684 , n28683 , n471 );
xor ( n28685 , n28684 , n28640 );
xor ( n28686 , n28685 , n28678 );
xor ( n28687 , n28684 , n28640 );
and ( n28688 , n28687 , n28678 );
and ( n28689 , n28684 , n28640 );
or ( n28690 , n28688 , n28689 );
and ( n28691 , n28673 , n471 , n10190 );
not ( n28692 , n28413 );
not ( n28693 , n27556 );
or ( n28694 , n28692 , n28693 );
nand ( n28695 , n28694 , n28428 );
not ( n28696 , n28695 );
and ( n28697 , n28414 , n25678 );
not ( n28698 , n28697 );
not ( n28699 , n24555 );
nand ( n28700 , n28699 , n24578 );
not ( n28701 , n28700 );
buf ( n28702 , n24572 );
not ( n28703 , n28702 );
nand ( n28704 , n28701 , n28703 );
not ( n28705 , n28704 );
or ( n28706 , n28698 , n28705 );
nand ( n28707 , n28706 , n28415 );
not ( n28708 , n28707 );
nand ( n28709 , n28696 , n28708 );
or ( n28710 , n28396 , n28403 );
not ( n28711 , n28710 );
not ( n28712 , n28711 );
nand ( n28713 , n28712 , n28437 );
and ( n28714 , n10190 , n472 );
and ( n28715 , n28713 , n28714 );
and ( n28716 , n28709 , n28715 );
not ( n28717 , n28709 );
not ( n28718 , n28714 );
nor ( n28719 , n28718 , n28713 );
and ( n28720 , n28717 , n28719 );
or ( n28721 , n28716 , n28720 );
xor ( n28722 , n28691 , n28721 );
and ( n28723 , n28631 , n470 );
xor ( n28724 , n28722 , n28723 );
xor ( n28725 , n28691 , n28721 );
and ( n28726 , n28725 , n28723 );
and ( n28727 , n28691 , n28721 );
or ( n28728 , n28726 , n28727 );
and ( n28729 , n27609 , n469 );
xor ( n28730 , n28729 , n28724 );
xor ( n28731 , n28730 , n28682 );
xor ( n28732 , n28729 , n28724 );
and ( n28733 , n28732 , n28682 );
and ( n28734 , n28729 , n28724 );
or ( n28735 , n28733 , n28734 );
not ( n28736 , n28448 );
not ( n28737 , n28407 );
or ( n28738 , n28736 , n28737 );
or ( n28739 , n28448 , n28407 );
nand ( n28740 , n28738 , n28739 );
nand ( n28741 , n28740 , n10190 );
nor ( n28742 , n28741 , n28711 );
not ( n28743 , n28742 );
not ( n28744 , n28743 );
not ( n28745 , n28697 );
not ( n28746 , n28704 );
or ( n28747 , n28745 , n28746 );
nand ( n28748 , n28747 , n28415 );
not ( n28749 , n28748 );
or ( n28750 , n28744 , n28749 );
not ( n28751 , n10190 );
nor ( n28752 , n28751 , n28740 );
nand ( n28753 , n28752 , n28437 );
nor ( n28754 , n28695 , n28753 );
nand ( n28755 , n28750 , n28754 );
and ( n28756 , n28695 , n28742 );
or ( n28757 , n28741 , n28437 );
nand ( n28758 , n28752 , n28437 , n28711 );
nand ( n28759 , n28757 , n28758 );
nor ( n28760 , n28756 , n28759 );
nand ( n28761 , n28748 , n28742 );
nand ( n28762 , n28755 , n28760 , n28761 );
and ( n28763 , n28762 , n472 );
and ( n28764 , n28673 , n10190 );
and ( n28765 , n28764 , n470 );
xor ( n28766 , n28763 , n28765 );
not ( n28767 , n28708 );
nor ( n28768 , n28695 , n28713 , n454 );
not ( n28769 , n28768 );
or ( n28770 , n28767 , n28769 );
or ( n28771 , n28707 , n28695 );
and ( n28772 , n28713 , n10190 );
nand ( n28773 , n28771 , n28772 );
nand ( n28774 , n28770 , n28773 );
and ( n28775 , n28774 , n471 );
xor ( n28776 , n28766 , n28775 );
xor ( n28777 , n28763 , n28765 );
and ( n28778 , n28777 , n28775 );
and ( n28779 , n28763 , n28765 );
or ( n28780 , n28778 , n28779 );
and ( n28781 , n28683 , n469 );
xor ( n28782 , n28781 , n28776 );
xor ( n28783 , n28782 , n28728 );
xor ( n28784 , n28781 , n28776 );
and ( n28785 , n28784 , n28728 );
and ( n28786 , n28781 , n28776 );
or ( n28787 , n28785 , n28786 );
buf ( n28788 , n28774 );
and ( n28789 , n28788 , n470 );
not ( n28790 , n28710 );
not ( n28791 , n28707 );
or ( n28792 , n28790 , n28791 );
and ( n28793 , n28695 , n28710 );
not ( n28794 , n28437 );
nor ( n28795 , n28793 , n28794 );
nand ( n28796 , n28792 , n28795 );
and ( n28797 , n28796 , n28741 );
not ( n28798 , n28796 );
not ( n28799 , n28740 );
nand ( n28800 , n28799 , n10190 );
and ( n28801 , n28798 , n28800 );
nor ( n28802 , n28797 , n28801 );
and ( n28803 , n28802 , n471 );
and ( n28804 , n28764 , n469 );
xor ( n28805 , n28803 , n28804 );
xor ( n28806 , n28789 , n28805 );
xor ( n28807 , n28806 , n28780 );
not ( n28808 , n16771 );
not ( n28809 , n28808 );
nor ( n28810 , n17648 , n23854 );
not ( n28811 , n28810 );
not ( n28812 , n23862 );
or ( n28813 , n28811 , n28812 );
not ( n28814 , n17648 );
not ( n28815 , n23865 );
and ( n28816 , n28814 , n28815 );
nor ( n28817 , n28816 , n17680 );
nand ( n28818 , n28813 , n28817 );
not ( n28819 , n28818 );
or ( n28820 , n28809 , n28819 );
nand ( n28821 , n28820 , n17684 );
not ( n28822 , n28643 );
not ( n28823 , n28583 );
nand ( n28824 , n28822 , n28823 );
nor ( n28825 , n28579 , n28562 );
nor ( n28826 , n28558 , n28503 );
nor ( n28827 , n28825 , n28826 );
nand ( n28828 , n28824 , n28827 );
nor ( n28829 , n28686 , n28647 );
nor ( n28830 , n28828 , n28829 );
not ( n28831 , n28830 );
not ( n28832 , n28731 );
not ( n28833 , n28690 );
nand ( n28834 , n28832 , n28833 );
not ( n28835 , n28783 );
not ( n28836 , n28735 );
nand ( n28837 , n28835 , n28836 );
nand ( n28838 , n28834 , n28837 );
nor ( n28839 , n28831 , n28838 );
nand ( n28840 , n28787 , n28807 );
not ( n28841 , n25587 );
nand ( n28842 , n17104 , n17343 );
not ( n28843 , n28499 );
not ( n28844 , n28456 );
nand ( n28845 , n28843 , n28844 );
nand ( n28846 , n28499 , n28456 );
nand ( n28847 , n28845 , n28846 );
or ( n28848 , n28503 , n28558 );
nand ( n28849 , n28558 , n28503 );
and ( n28850 , n28848 , n28849 );
and ( n28851 , n25641 , n25643 );
not ( n28852 , n28851 );
xor ( n28853 , n17289 , n17291 );
xor ( n28854 , n28853 , n17308 );
nor ( n28855 , n28833 , n28832 );
not ( n28856 , n27162 );
and ( n28857 , n17282 , n17327 );
not ( n28858 , n17320 );
nand ( n28859 , n28858 , n17318 );
xnor ( n28860 , n17340 , n28842 );
and ( n28861 , n17063 , n17347 );
not ( n28862 , n28836 );
nand ( n28863 , n28862 , n28783 );
xor ( n28864 , n28291 , n28256 );
nor ( n28865 , n28499 , n28456 );
nor ( n28866 , n25845 , n25849 );
nor ( n28867 , n28865 , n28866 );
not ( n28868 , n28867 );
not ( n28869 , n25667 );
or ( n28870 , n28868 , n28869 );
not ( n28871 , n25851 );
and ( n28872 , n28845 , n28871 );
not ( n28873 , n28846 );
nor ( n28874 , n28872 , n28873 );
nand ( n28875 , n28870 , n28874 );
not ( n28876 , n28875 );
not ( n28877 , n25645 );
not ( n28878 , n27136 );
or ( n28879 , n28877 , n28878 );
nand ( n28880 , n28867 , n25516 );
nand ( n28881 , n25650 , n25653 , n25547 );
nor ( n28882 , n28880 , n28881 );
nand ( n28883 , n28879 , n28882 );
not ( n28884 , n28880 );
nand ( n28885 , n25592 , n28884 );
nand ( n28886 , n28876 , n28883 , n28885 );
buf ( n28887 , n28886 );
not ( n28888 , n28887 );
nand ( n28889 , n28837 , n28863 );
not ( n28890 , n28823 );
not ( n28891 , n28643 );
not ( n28892 , n28891 );
or ( n28893 , n28890 , n28892 );
nor ( n28894 , n28562 , n28579 );
or ( n28895 , n28894 , n28849 );
nand ( n28896 , n28579 , n28562 );
nand ( n28897 , n28895 , n28896 );
nand ( n28898 , n28893 , n28897 );
buf ( n28899 , n28643 );
nand ( n28900 , n28583 , n28899 );
nand ( n28901 , n28647 , n28686 );
nand ( n28902 , n28898 , n28900 , n28901 );
not ( n28903 , n28902 );
not ( n28904 , n28686 );
not ( n28905 , n28647 );
nand ( n28906 , n28904 , n28905 );
not ( n28907 , n28906 );
nor ( n28908 , n28903 , n28907 );
nand ( n28909 , n28832 , n28833 );
and ( n28910 , n28908 , n28909 );
nor ( n28911 , n28910 , n28855 );
nand ( n28912 , n28899 , n28583 );
nand ( n28913 , n28824 , n28912 );
not ( n28914 , n28240 );
nand ( n28915 , n28914 , n28031 );
buf ( n28916 , n28827 );
not ( n28917 , n28293 );
not ( n28918 , n27019 );
or ( n28919 , n28917 , n28918 );
not ( n28920 , n28292 );
and ( n28921 , n28920 , n28213 );
nor ( n28922 , n28921 , n28298 );
nand ( n28923 , n28919 , n28922 );
or ( n28924 , n28913 , n18007 );
not ( n28925 , n28916 );
not ( n28926 , n28887 );
or ( n28927 , n28925 , n28926 );
not ( n28928 , n28897 );
nand ( n28929 , n28927 , n28928 );
not ( n28930 , n28913 );
nor ( n28931 , n28930 , n18007 );
nand ( n28932 , n28929 , n28931 );
and ( n28933 , n28218 , n28147 );
xnor ( n28934 , n28215 , n28933 );
or ( n28935 , n28934 , n23837 );
not ( n28936 , n28825 );
nand ( n28937 , n28936 , n28896 );
not ( n28938 , n28937 );
nor ( n28939 , n28938 , n18007 );
or ( n28940 , n28686 , n28647 );
nand ( n28941 , n28940 , n28901 );
and ( n28942 , n28941 , n23837 );
not ( n28943 , n25850 );
nand ( n28944 , n25845 , n25849 );
nand ( n28945 , n28943 , n28944 );
not ( n28946 , n28831 );
or ( n28947 , n28852 , n18007 );
not ( n28948 , n27159 );
not ( n28949 , n28856 );
or ( n28950 , n28948 , n28949 );
not ( n28951 , n25640 );
nand ( n28952 , n28950 , n28951 );
or ( n28953 , n28947 , n28952 );
not ( n28954 , n28952 );
or ( n28955 , n28851 , n18007 );
or ( n28956 , n28954 , n28955 );
xor ( n28957 , n28287 , n26995 );
or ( n28958 , n28957 , n23837 );
nand ( n28959 , n28953 , n28956 , n28958 );
buf ( n28960 , n25650 );
nand ( n28961 , n28960 , n25586 );
or ( n28962 , n28961 , n18007 );
not ( n28963 , n25653 );
not ( n28964 , n27137 );
or ( n28965 , n28963 , n28964 );
nand ( n28966 , n28965 , n25584 );
or ( n28967 , n28962 , n28966 );
not ( n28968 , n28961 );
nor ( n28969 , n28968 , n18007 );
nand ( n28970 , n28966 , n28969 );
and ( n28971 , n28284 , n27002 );
not ( n28972 , n28284 );
and ( n28973 , n28972 , n28257 );
or ( n28974 , n28971 , n28973 );
or ( n28975 , n28974 , n23837 );
nand ( n28976 , n28967 , n28970 , n28975 );
nand ( n28977 , n25660 , n25666 );
or ( n28978 , n28977 , n18007 );
or ( n28979 , n27071 , n27067 );
nand ( n28980 , n28979 , n27069 );
or ( n28981 , n28978 , n28980 );
not ( n28982 , n28977 );
nor ( n28983 , n28982 , n18007 );
nand ( n28984 , n28980 , n28983 );
or ( n28985 , n28864 , n23837 );
nand ( n28986 , n28981 , n28984 , n28985 );
nand ( n28987 , n25591 , n25547 );
not ( n28988 , n28987 );
nand ( n28989 , n28988 , n23837 );
nand ( n28990 , n25653 , n28960 );
not ( n28991 , n28990 );
not ( n28992 , n28991 );
not ( n28993 , n27137 );
or ( n28994 , n28992 , n28993 );
nand ( n28995 , n28994 , n28841 );
or ( n28996 , n28989 , n28995 );
not ( n28997 , n28987 );
not ( n28998 , n23837 );
nor ( n28999 , n28997 , n28998 );
nand ( n29000 , n28995 , n28999 );
xnor ( n29001 , n28286 , n28259 );
nand ( n29002 , n29001 , n28998 );
nand ( n29003 , n28996 , n29000 , n29002 );
and ( n29004 , n28912 , n28901 );
or ( n29005 , n28643 , n28583 );
nand ( n29006 , n29005 , n28897 );
and ( n29007 , n29006 , n28912 );
not ( n29008 , n17297 );
or ( n29009 , n17307 , n29008 );
or ( n29010 , n29008 , n17303 );
and ( n29011 , n29008 , n17302 , n17300 );
nor ( n29012 , n17300 , n17297 , n17302 );
nor ( n29013 , n29011 , n29012 );
nand ( n29014 , n29009 , n29010 , n29013 );
and ( n29015 , n17247 , n472 );
not ( n29016 , n28850 );
nand ( n29017 , n29016 , n23837 );
or ( n29018 , n28888 , n29017 );
and ( n29019 , n28850 , n23837 );
nand ( n29020 , n28888 , n29019 );
buf ( n29021 , n28250 );
not ( n29022 , n29021 );
not ( n29023 , n28300 );
or ( n29024 , n29022 , n29023 );
or ( n29025 , n29021 , n28300 );
nand ( n29026 , n29024 , n29025 );
nand ( n29027 , n29026 , n18007 );
nand ( n29028 , n29018 , n29020 , n29027 );
nand ( n29029 , n28876 , n28883 , n28885 );
not ( n29030 , n28911 );
not ( n29031 , n28909 );
nor ( n29032 , n29031 , n28831 );
nand ( n29033 , n28887 , n29032 );
not ( n29034 , n29033 );
or ( n29035 , n29030 , n29034 );
and ( n29036 , n28889 , n23837 );
nand ( n29037 , n29035 , n29036 );
nor ( n29038 , n28889 , n18007 );
nand ( n29039 , n28911 , n29033 , n29038 );
not ( n29040 , n27960 );
not ( n29041 , n28156 );
not ( n29042 , n28215 );
or ( n29043 , n29041 , n29042 );
nand ( n29044 , n29043 , n28222 );
not ( n29045 , n29044 );
or ( n29046 , n29040 , n29045 );
nand ( n29047 , n29046 , n28226 );
xor ( n29048 , n29047 , n28301 );
nand ( n29049 , n29048 , n18007 );
nand ( n29050 , n29037 , n29039 , n29049 );
not ( n29051 , n28855 );
not ( n29052 , n28837 );
or ( n29053 , n29051 , n29052 );
nand ( n29054 , n29053 , n28863 );
not ( n29055 , n28236 );
and ( n29056 , n28329 , n28233 , n28231 );
nand ( n29057 , n28002 , n28021 );
nor ( n29058 , n29056 , n29057 );
nor ( n29059 , n29055 , n29058 );
xor ( n29060 , n28915 , n29059 );
nand ( n29061 , n29060 , n23844 );
nand ( n29062 , C1 , n29061 );
nor ( n29063 , n28838 , n28907 );
and ( n29064 , n28902 , n29063 );
nor ( n29065 , n29064 , n29054 );
and ( n29066 , n29006 , n29004 );
nor ( n29067 , n29066 , n28907 );
not ( n29068 , n29067 );
and ( n29069 , n28248 , n18007 );
nor ( n29070 , C0 , n29069 );
nand ( n29071 , n29070 , C1 , C1 , C1 );
and ( n29072 , n23698 , n23726 );
nor ( n29073 , n29072 , n23729 );
not ( n29074 , n29073 );
and ( n29075 , n29074 , n23738 );
nor ( n29076 , n29073 , n23740 );
nor ( n29077 , n29075 , n29076 );
not ( n29078 , n23737 );
nand ( n29079 , n29078 , n29073 , n23732 );
not ( n29080 , n23732 );
nand ( n29081 , n29080 , n29073 , n23737 );
nand ( n29082 , n29077 , n29079 , n29081 );
not ( n29083 , n28946 );
not ( n29084 , n28887 );
or ( n29085 , n29083 , n29084 );
nand ( n29086 , n29085 , n29068 );
or ( n29087 , n28924 , n28929 );
nand ( n29088 , n29087 , n28932 , n28935 );
not ( n29089 , n29007 );
not ( n29090 , n28828 );
nand ( n29091 , n28887 , n29090 );
not ( n29092 , n29091 );
or ( n29093 , n29089 , n29092 );
nand ( n29094 , n29093 , n28942 );
not ( n29095 , n23837 );
nor ( n29096 , n29095 , n28941 );
and ( n29097 , n29091 , n29007 , n29096 );
not ( n29098 , n28220 );
nor ( n29099 , n29098 , n28154 );
not ( n29100 , n29099 );
not ( n29101 , n28198 );
not ( n29102 , n27290 );
or ( n29103 , n29101 , n29102 );
nand ( n29104 , n29103 , n28214 );
and ( n29105 , n29104 , n28147 );
not ( n29106 , n28218 );
nor ( n29107 , n29105 , n29106 );
not ( n29108 , n29107 );
or ( n29109 , n29100 , n29108 );
or ( n29110 , n29107 , n29099 );
nand ( n29111 , n29109 , n29110 );
and ( n29112 , n29111 , n18007 );
nor ( n29113 , n29097 , n29112 );
nand ( n29114 , n29094 , n29113 );
not ( n29115 , n23837 );
nand ( n29116 , n29115 , n28334 );
nand ( n29117 , C1 , C1 , n29116 , C1 );
nand ( n29118 , n28848 , n29029 , n28939 );
not ( n29119 , n28253 );
nor ( n29120 , n28299 , n23837 );
nand ( n29121 , n29119 , n29120 );
and ( n29122 , n28299 , n18007 );
nand ( n29123 , n28253 , n29122 );
not ( n29124 , n28848 );
not ( n29125 , n28937 );
nand ( n29126 , n29124 , n29125 , n28849 , n23837 );
and ( n29127 , n29121 , n29123 , n29126 );
not ( n29128 , n28849 );
nand ( n29129 , n29128 , n28939 );
not ( n29130 , n29029 );
and ( n29131 , n29125 , n28849 , n23837 );
nand ( n29132 , n29130 , n29131 );
nand ( n29133 , n29118 , n29127 , n29129 , n29132 );
not ( n29134 , n28944 );
buf ( n29135 , n28847 );
not ( n29136 , n29135 );
or ( n29137 , n29134 , n29136 );
not ( n29138 , n28945 );
or ( n29139 , n29138 , n29135 );
nand ( n29140 , n29137 , n29139 );
not ( n29141 , n29140 );
not ( n29142 , n28847 );
nand ( n29143 , n29142 , n25669 , n28944 );
not ( n29144 , n29143 );
nand ( n29145 , n29144 , n25854 );
not ( n29146 , n29145 );
or ( n29147 , n29141 , n29146 );
nand ( n29148 , n29147 , n23837 );
and ( n29149 , n28847 , n25850 , n23837 );
nand ( n29150 , n25670 , n29149 );
nand ( n29151 , n29148 , n29150 , n27297 );
not ( n29152 , n28855 );
and ( n29153 , n28909 , n29152 );
nor ( n29154 , n29153 , n18007 );
nand ( n29155 , n29086 , n29154 );
nand ( n29156 , n28946 , n28887 );
not ( n29157 , n18007 );
nand ( n29158 , n29157 , n29152 , n28909 );
nor ( n29159 , n29067 , n29158 );
and ( n29160 , n29156 , n29159 );
xnor ( n29161 , n28304 , n29044 );
nor ( n29162 , n29161 , n23837 );
nor ( n29163 , n29160 , n29162 );
nand ( n29164 , n29155 , n29163 );
nand ( n29165 , n15063 , n15052 );
or ( n29166 , n15050 , n29165 );
not ( n29167 , n15052 );
and ( n29168 , n15050 , n15063 , n29167 );
not ( n29169 , n15063 );
and ( n29170 , n15053 , n29169 );
nor ( n29171 , n29168 , n29170 );
nand ( n29172 , n29166 , C1 , n29171 );
not ( n29173 , n17595 );
not ( n29174 , n23919 );
or ( n29175 , n29173 , n29174 );
nand ( n29176 , n29175 , n23921 );
not ( n29177 , n27304 );
xor ( n29178 , n17344 , n28861 );
nand ( n29179 , n23845 , n29178 );
nand ( n29180 , n29177 , n29179 );
xor ( n29181 , n28857 , n17324 );
not ( n29182 , n454 );
and ( n29183 , n27622 , n454 );
and ( n29184 , n28436 , n29182 );
nor ( n29185 , n29183 , n29184 );
not ( n29186 , n29185 );
not ( n29187 , n23845 );
not ( n29188 , n29015 );
or ( n29189 , n29187 , n29188 );
not ( n29190 , n23644 );
nand ( n29191 , n29190 , n23844 );
nand ( n29192 , n29189 , n29191 );
and ( n29193 , n27628 , n454 );
and ( n29194 , n28439 , n29182 );
nor ( n29195 , n29193 , n29194 );
not ( n29196 , n29195 );
and ( n29197 , n27632 , n454 );
and ( n29198 , n28442 , n29182 );
nor ( n29199 , n29197 , n29198 );
not ( n29200 , n29199 );
not ( n29201 , n23845 );
not ( n29202 , n28854 );
or ( n29203 , n29201 , n29202 );
nand ( n29204 , n28314 , n23844 );
nand ( n29205 , n29203 , n29204 );
and ( n29206 , n27630 , n454 );
and ( n29207 , n29172 , n29182 );
nor ( n29208 , n29206 , n29207 );
not ( n29209 , n17586 );
not ( n29210 , n23916 );
or ( n29211 , n29209 , n29210 );
not ( n29212 , n17621 );
nand ( n29213 , n29211 , n29212 );
not ( n29214 , n17623 );
and ( n29215 , n17620 , n29214 );
nand ( n29216 , n29215 , n23837 );
or ( n29217 , n29213 , n29216 );
not ( n29218 , n28280 );
or ( n29219 , n29218 , n23837 );
not ( n29220 , n29213 );
not ( n29221 , n29215 );
nand ( n29222 , n29221 , n23837 );
or ( n29223 , n29220 , n29222 );
nand ( n29224 , n29217 , n29219 , n29223 );
nand ( n29225 , n17594 , n17590 );
not ( n29226 , n29225 );
nand ( n29227 , n29226 , n23837 );
or ( n29228 , n29176 , n29227 );
xor ( n29229 , n28282 , n28278 );
or ( n29230 , n29229 , n23837 );
not ( n29231 , n29176 );
nand ( n29232 , n29225 , n23837 );
or ( n29233 , n29231 , n29232 );
nand ( n29234 , n29228 , n29230 , n29233 );
nand ( n29235 , n28324 , n23844 );
and ( n29236 , n28923 , n29235 );
not ( n29237 , n28923 );
not ( n29238 , n28324 );
nand ( n29239 , n29238 , n23844 );
and ( n29240 , n29237 , n29239 );
nor ( n29241 , n29236 , n29240 );
not ( n29242 , n23845 );
not ( n29243 , n28860 );
or ( n29244 , n29242 , n29243 );
nand ( n29245 , n28289 , n23844 );
nand ( n29246 , n29244 , n29245 );
not ( n29247 , n23845 );
not ( n29248 , n29181 );
or ( n29249 , n29247 , n29248 );
nand ( n29250 , n28310 , n23844 );
nand ( n29251 , n29249 , n29250 );
nand ( n29252 , n29082 , n23844 );
not ( n29253 , n16955 );
nand ( n29254 , n29253 , n16990 );
buf ( n29255 , n17353 );
or ( n29256 , n29254 , n29255 );
not ( n29257 , n16990 );
nand ( n29258 , n29257 , n16955 );
or ( n29259 , n29258 , n29255 );
not ( n29260 , n17356 );
not ( n29261 , n16991 );
or ( n29262 , n29260 , n29261 );
nand ( n29263 , n29262 , n29255 );
nand ( n29264 , n29256 , n29259 , n29263 );
nand ( n29265 , n23845 , n29264 );
nand ( n29266 , n29252 , n29265 );
not ( n29267 , n23948 );
not ( n29268 , n29014 );
or ( n29269 , n29267 , n29268 );
nand ( n29270 , n28326 , n23844 );
nand ( n29271 , n29269 , n29270 );
or ( n29272 , n28787 , n28807 );
nand ( n29273 , n29272 , n28840 );
not ( n29274 , n28839 );
not ( n29275 , n28887 );
or ( n29276 , n29274 , n29275 );
nand ( n29277 , n29276 , n29065 );
not ( n29278 , n29273 );
nor ( n29279 , n29278 , n18007 );
nand ( n29280 , n29277 , n29279 );
xor ( n29281 , n28330 , n28311 );
or ( n29282 , n29281 , n23837 );
nand ( n29283 , C1 , n29280 , n29282 );
not ( n29284 , n17690 );
nand ( n29285 , n29284 , n17688 );
not ( n29286 , n29285 );
nand ( n29287 , n29286 , n23837 );
or ( n29288 , n28821 , n29287 );
and ( n29289 , n29285 , n23837 );
nand ( n29290 , n28821 , n29289 );
nand ( n29291 , n28271 , n18007 );
nand ( n29292 , n29288 , n29290 , n29291 );
nand ( n29293 , n28808 , n17684 );
not ( n29294 , n29293 );
nand ( n29295 , n29294 , n23837 );
nand ( n29296 , n28276 , n18007 );
not ( n29297 , n23850 );
not ( n29298 , n29208 );
xor ( n29299 , n23609 , n23618 );
xor ( n29300 , n29299 , n23657 );
not ( n29301 , n17311 );
not ( n29302 , n28859 );
or ( n29303 , n29301 , n29302 );
or ( n29304 , n17311 , n28859 );
nand ( n29305 , n29303 , n29304 );
and ( n29306 , n23845 , n29305 );
and ( n29307 , n29300 , n23844 );
nor ( n29308 , n29306 , n29307 );
not ( n29309 , n29308 );
or ( n29310 , n29295 , n28818 );
and ( n29311 , n29293 , n23837 );
nand ( n29312 , n28818 , n29311 );
nand ( n29313 , n29310 , n29312 , n29296 );
nand ( n29314 , n17851 , n17984 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
