module mul_11s_11s_1s(a, b, c);
  input signed [10:0] a;
  input signed [10:0] b;
  output signed c;
  assign c = a * b;
endmodule
