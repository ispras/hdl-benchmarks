// IWLS benchmark module "i10" printed on Wed May 29 16:38:44 2002
module i10(\V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) , \V10(0) , \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) , \V248(0) , \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) , \V66(0) , \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) , \V45(0) , \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) , \V34(0) , \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) , \V293(0) , \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) , \V275(0) , \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) , \V257(4) , \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) , \V149(3) , \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) , \V165(6) , \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) , \V169(0) , \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) , \V165(3) , \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) , \V288(4) , \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) , \V229(3) , \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) , \V223(3) , \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) , \V189(3) , \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) , \V183(3) , \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) , \V239(2) , \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) , \V234(1) , \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) , \V199(0) , \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) , \V257(0) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) , \V32(10) , \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) , \V84(2) , \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) , \V14(0) , \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) , \V213(1) , \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) , \V8(0) , \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) , \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) , \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) , \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) , \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) , \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) , \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) , \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) , \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) , \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) , \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) , \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) , \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) , \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) , \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) , \V78(0) , \V94(0) , \V94(1) , \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) , \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) , V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546, V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) , \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587, \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630, \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) , \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) , \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) , \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) , \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) , \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) , \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378, V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428, V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) , \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) , \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539, \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) , \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) , \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) , V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) , \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) , \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) , \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832, \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) , \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) , \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) , \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) , \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653, V654, V655, V656, V1370, V1371, V1372, V1373, V1374);
input
  \V246(0) ,
  \V229(3) ,
  \V229(2) ,
  \V229(5) ,
  \V229(4) ,
  \V38(0) ,
  \V171(0) ,
  \V229(1) ,
  \V229(0) ,
  \V57(0) ,
  \V248(0) ,
  \V118(3) ,
  \V118(2) ,
  \V118(5) ,
  \V59(0) ,
  \V118(4) ,
  \V288(3) ,
  \V288(2) ,
  \V78(0) ,
  \V288(5) ,
  \V118(1) ,
  \V78(1) ,
  \V302(0) ,
  \V288(4) ,
  \V118(0) ,
  \V78(2) ,
  \V269(0) ,
  \V78(3) ,
  \V78(4) ,
  \V288(1) ,
  \V78(5) ,
  \V288(0) ,
  \V118(7) ,
  \V194(3) ,
  \V118(6) ,
  \V194(2) ,
  \V194(4) ,
  \V288(7) ,
  \V175(0) ,
  \V288(6) ,
  \V194(1) ,
  \V194(0) ,
  \V177(0) ,
  \V40(0) ,
  \V1(0) ,
  \V214(0) ,
  \V42(0) ,
  \V3(0) ,
  \V101(0) ,
  \V271(0) ,
  \V290(0) ,
  \V216(0) ,
  \V44(0) ,
  \V5(0) ,
  \V63(0) ,
  \V292(0) ,
  \V46(0) ,
  \V124(3) ,
  \V7(0) ,
  \V124(2) ,
  \V124(5) ,
  \V65(0) ,
  \V124(4) ,
  \V84(0) ,
  \V124(1) ,
  \V84(1) ,
  \V124(0) ,
  \V84(2) ,
  \V275(0) ,
  \V84(3) ,
  \V84(4) ,
  \V84(5) ,
  \V294(0) ,
  \V239(3) ,
  \V239(2) ,
  \V239(4) ,
  \V48(0) ,
  \V9(0) ,
  \V239(1) ,
  \V239(0) ,
  \V67(0) ,
  \V258(0) ,
  \V277(0) ,
  \V183(3) ,
  \V183(2) ,
  \V183(5) ,
  \V183(4) ,
  \V183(1) ,
  \V183(0) ,
  \V69(0) ,
  \V109(0) ,
  \V88(0) ,
  \V88(1) ,
  \V88(2) ,
  \V279(0) ,
  \V88(3) ,
  \V149(3) ,
  \V149(2) ,
  \V149(5) ,
  \V149(4) ,
  \V149(1) ,
  \V10(0) ,
  \V149(0) ,
  \V149(7) ,
  \V149(6) ,
  \V189(3) ,
  \V12(0) ,
  \V189(2) ,
  \V189(5) ,
  \V203(0) ,
  \V189(4) ,
  \V189(1) ,
  \V50(0) ,
  \V189(0) ,
  \V241(0) ,
  \V260(0) ,
  \V14(0) ,
  \V205(0) ,
  \V33(0) ,
  \V52(0) ,
  \V243(0) ,
  \V71(0) ,
  \V262(0) ,
  \V16(0) ,
  \V207(0) ,
  \V35(0) ,
  \V132(3) ,
  \V132(2) ,
  \V245(0) ,
  \V132(5) ,
  \V132(4) ,
  \V132(1) ,
  \V132(0) ,
  \V132(7) ,
  \V37(0) ,
  \V132(6) ,
  \V56(0) ,
  \V247(0) ,
  \V94(0) ,
  \V134(1) ,
  \V94(1) ,
  \V134(0) ,
  \V39(0) ,
  \V172(0) ,
  \V268(3) ,
  \V268(2) ,
  \V268(5) ,
  \V268(4) ,
  \V249(0) ,
  \V301(0) ,
  \V268(1) ,
  \V268(0) ,
  \V174(0) ,
  \V289(0) ,
  \V213(3) ,
  \V213(2) ,
  \V213(5) ,
  \V213(4) ,
  \V199(3) ,
  \V199(2) ,
  \V100(3) ,
  \V213(1) ,
  \V100(2) ,
  \V213(0) ,
  \V199(4) ,
  \V100(5) ,
  \V41(0) ,
  \V100(4) ,
  \V2(0) ,
  \V199(1) ,
  \V60(0) ,
  \V199(0) ,
  \V100(1) ,
  \V100(0) ,
  \V270(0) ,
  \V234(3) ,
  \V234(2) ,
  \V234(4) ,
  \V215(0) ,
  \V43(0) ,
  \V4(0) ,
  \V234(1) ,
  \V234(0) ,
  \V62(0) ,
  \V102(0) ,
  \V32(11) ,
  \V272(0) ,
  \V32(10) ,
  \V291(0) ,
  \V45(0) ,
  \V6(0) ,
  \V274(0) ,
  \V293(0) ,
  \V257(3) ,
  \V257(2) ,
  \V257(5) ,
  \V8(0) ,
  \V257(4) ,
  \V66(0) ,
  \V257(1) ,
  \V257(0) ,
  \V257(7) ,
  \V257(6) ,
  \V295(0) ,
  \V108(3) ,
  \V108(2) ,
  \V108(5) ,
  \V108(4) ,
  \V68(0) ,
  \V108(1) ,
  \V108(0) ,
  \V259(0) ,
  \V165(3) ,
  \V165(2) ,
  \V278(0) ,
  \V165(5) ,
  \V165(4) ,
  \V165(1) ,
  \V165(0) ,
  \V165(7) ,
  \V165(6) ,
  \V11(0) ,
  \V202(0) ,
  \V169(1) ,
  \V169(0) ,
  \V240(0) ,
  \V223(3) ,
  \V223(2) ,
  \V13(0) ,
  \V223(5) ,
  \V223(4) ,
  \V204(0) ,
  \V32(0) ,
  \V32(1) ,
  \V223(1) ,
  \V32(2) ,
  \V223(0) ,
  \V32(3) ,
  \V51(0) ,
  \V32(4) ,
  \V32(5) ,
  \V242(0) ,
  \V32(6) ,
  \V70(0) ,
  \V32(7) ,
  \V110(0) ,
  \V32(8) ,
  \V261(0) ,
  \V32(9) ,
  \V280(0) ,
  \V15(0) ,
  \V34(0) ,
  \V53(0) ,
  \V244(0) ,
  \V91(0) ,
  \V91(1) ,
  \V55(0) ;
output
  \V1213(10) ,
  \V1213(11) ,
  \V1440(0) ,
  \V1833(0) ,
  \V1536(0) ,
  \V321(2) ,
  \V585(0) ,
  \V1480(0) ,
  \V1741(0) ,
  \V1760(0) ,
  \V603(0) ,
  \V1781(1) ,
  \V1781(0) ,
  \V1726(0) ,
  V356,
  V357,
  \V1745(0) ,
  \V1896(0) ,
  \V1613(1) ,
  V373,
  V377,
  \V1613(0) ,
  \V511(0) ,
  \V1467(0) ,
  \V1709(1) ,
  \V1709(0) ,
  \V1709(3) ,
  \V1709(2) ,
  V432,
  \V1709(4) ,
  \V1898(0) ,
  \V1392(0) ,
  \V1243(7) ,
  \V1243(6) ,
  \V1243(9) ,
  V512,
  \V1243(8) ,
  \V609(0) ,
  V527,
  V537,
  V538,
  V539,
  V540,
  V541,
  V542,
  V543,
  V544,
  V545,
  V546,
  V547,
  V548,
  \V798(0) ,
  \V1243(1) ,
  V587,
  \V1243(0) ,
  \V1243(3) ,
  \V1243(2) ,
  \V572(3) ,
  \V1243(5) ,
  \V572(2) ,
  \V1243(4) ,
  \V572(5) ,
  \V572(4) ,
  \V1281(0) ,
  \V572(1) ,
  V620,
  V621,
  \V572(0) ,
  V630,
  \V1693(0) ,
  V650,
  V651,
  V652,
  V653,
  V654,
  V655,
  V656,
  V657,
  \V591(0) ,
  \V572(7) ,
  \V572(6) ,
  \V572(9) ,
  \V572(8) ,
  \V1992(1) ,
  \V1992(0) ,
  V707,
  \V423(0) ,
  V763,
  V775,
  V778,
  V779,
  V780,
  V781,
  V782,
  V783,
  V784,
  V787,
  V789,
  V801,
  \V1864(0) ,
  V966,
  \V597(0) ,
  V986,
  \V1492(0) ,
  \V500(0) ,
  \V1901(0) ,
  \V1717(0) ,
  \V634(0) ,
  \V1213(7) ,
  \V1439(0) ,
  \V1213(6) ,
  \V1213(9) ,
  \V1213(8) ,
  \V375(0) ,
  \V1213(1) ,
  \V1213(0) ,
  \V1213(3) ,
  \V1213(2) ,
  \V1757(0) ,
  \V1213(5) ,
  \V1960(1) ,
  \V1213(4) ,
  \V1960(0) ,
  \V1512(1) ,
  \V1512(3) ,
  \V410(0) ,
  \V1512(2) ,
  V1256,
  V1257,
  V1258,
  V1259,
  \V1759(0) ,
  V1260,
  V1261,
  V1262,
  V1263,
  V1264,
  V1265,
  V1266,
  V1267,
  \V1552(1) ,
  \V398(0) ,
  \V1552(0) ,
  V1365,
  V1370,
  V1371,
  \V508(0) ,
  V1372,
  V1373,
  V1374,
  V1375,
  V1378,
  V1380,
  V1382,
  V1384,
  V1386,
  \V1629(0) ,
  V1387,
  \V1274(0) ,
  V1423,
  V1426,
  V1428,
  V1429,
  V1431,
  V1432,
  \V826(0) ,
  V1470,
  \V435(0) ,
  V1537,
  V1539,
  \V1968(0) ,
  \V1297(1) ,
  \V1481(0) ,
  \V1297(0) ,
  \V1297(3) ,
  \V1297(2) ,
  \V1297(4) ,
  \V640(0) ,
  V1669,
  V1719,
  V1736,
  V1832,
  \V1897(0) ,
  \V1652(0) ,
  \V1671(0) ,
  \V1899(0) ,
  \V1953(7) ,
  \V1953(6) ,
  \V1953(1) ,
  \V1953(0) ,
  \V1953(3) ,
  \V1953(2) ,
  \V1953(5) ,
  \V1953(4) ,
  \V1451(0) ,
  \V1863(0) ,
  \V1679(0) ,
  \V1829(7) ,
  \V1829(6) ,
  \V1829(9) ,
  \V1829(8) ,
  \V1771(1) ,
  \V1620(0) ,
  \V1771(0) ,
  \V1829(1) ,
  \V1829(0) ,
  \V1829(3) ,
  \V1829(2) ,
  \V1829(5) ,
  \V1829(4) ,
  \V1900(0) ,
  \V1921(1) ,
  \V1495(0) ,
  \V1921(0) ,
  \V1921(3) ,
  \V393(0) ,
  \V1921(2) ,
  \V1921(5) ,
  \V1921(4) ,
  \V1459(0) ,
  \V802(0) ,
  \V821(0) ,
  \V1758(0) ,
  \V1645(0) ;
wire
  \[189] ,
  \[190] ,
  \[380] ,
  \V1647(0) ,
  \[191] ,
  \[381] ,
  \[192] ,
  \[382] ,
  \[193] ,
  \[383] ,
  \[194] ,
  \[384] ,
  \[195] ,
  \[385] ,
  \[196] ,
  \[386] ,
  \[197] ,
  \[387] ,
  \[198] ,
  \[388] ,
  \[199] ,
  \[389] ,
  \V1421(0) ,
  \V470(0) ,
  \[0] ,
  \[1] ,
  \[390] ,
  \[2] ,
  \[3] ,
  \V731(0) ,
  \[4] ,
  \[393] ,
  \[5] ,
  \V2019(0) ,
  \[394] ,
  \[6] ,
  \[7] ,
  \[396] ,
  \[8] ,
  \[9] ,
  \[399] ,
  \V2078(0) ,
  \V493(0) ,
  \V1463(0) ,
  \V1331(0) ,
  V379,
  \V2002(0) ,
  V411,
  \V758(0) ,
  V433,
  V437,
  V439,
  \V1354(0) ,
  V440,
  V441,
  V446,
  V451,
  V452,
  V454,
  V456,
  \V1653(0) ,
  V505,
  \V1337(0) ,
  \V812(0) ,
  \V2061(0) ,
  \[200] ,
  \[201] ,
  \[202] ,
  \[203] ,
  \[204] ,
  \[205] ,
  \V1674(0) ,
  \[206] ,
  \[207] ,
  \[208] ,
  V646,
  \[209] ,
  V687,
  V695,
  V697,
  \[210] ,
  \[400] ,
  \[211] ,
  \[401] ,
  \[212] ,
  \[402] ,
  \[213] ,
  \V404(0) ,
  V700,
  V701,
  V702,
  \[214] ,
  \[404] ,
  V710,
  \[215] ,
  V721,
  \[216] ,
  V725,
  V726,
  V727,
  \[217] ,
  V735,
  V736,
  V737,
  \[407] ,
  V738,
  V739,
  V740,
  V741,
  V742,
  V743,
  V744,
  \[218] ,
  V745,
  V746,
  V747,
  \[408] ,
  V749,
  V750,
  V751,
  \[219] ,
  \[409] ,
  V768,
  V769,
  V799,
  \V2084(0) ,
  \[220] ,
  \[221] ,
  \[222] ,
  \[412] ,
  \[223] ,
  \[413] ,
  \[224] ,
  \[414] ,
  \[225] ,
  \[415] ,
  \[226] ,
  \[416] ,
  \[227] ,
  \[417] ,
  \[228] ,
  \[418] ,
  \[229] ,
  V856,
  V866,
  V896,
  \[230] ,
  \[231] ,
  \[232] ,
  \[233] ,
  \[234] ,
  V906,
  \[235] ,
  \[236] ,
  \[237] ,
  V936,
  \[238] ,
  V946,
  V954,
  V955,
  V976,
  \[240] ,
  \[430] ,
  \[431] ,
  \[432] ,
  \[244] ,
  \[434] ,
  \[245] ,
  \[435] ,
  \[437] ,
  \[248] ,
  \[438] ,
  \V467(0) ,
  \[441] ,
  \[252] ,
  \[442] ,
  \[253] ,
  \[443] ,
  \[444] ,
  \[445] ,
  \[446] ,
  \[257] ,
  \[258] ,
  \[448] ,
  \[449] ,
  \[260] ,
  \[450] ,
  \[262] ,
  \[263] ,
  \[266] ,
  \[267] ,
  V1125,
  \[270] ,
  \[271] ,
  \[272] ,
  \[464] ,
  \[465] ,
  \V2033(0) ,
  \[277] ,
  \[279] ,
  V1298,
  \[280] ,
  \[281] ,
  \[471] ,
  \[282] ,
  \[472] ,
  \[285] ,
  \[475] ,
  V1300,
  V1301,
  V1302,
  V1307,
  \[286] ,
  V1312,
  V1318,
  \[287] ,
  V1320,
  \[288] ,
  \[478] ,
  \[289] ,
  \[479] ,
  V1366,
  \V1255(1) ,
  \V1255(0) ,
  \V1255(3) ,
  \[290] ,
  \[480] ,
  \V1255(2) ,
  \[291] ,
  \[481] ,
  \V730(0) ,
  \[292] ,
  \[482] ,
  \[293] ,
  \[483] ,
  \[294] ,
  \[484] ,
  \[295] ,
  V1402,
  \[486] ,
  \V807(0) ,
  V1445,
  \V1422(0) ,
  V1476,
  \V490(0) ,
  \[497] ,
  \[498] ,
  V1535,
  \[499] ,
  \V2058(0) ,
  V1587,
  V1588,
  V1589,
  \V473(0) ,
  V1590,
  V1606,
  V1607,
  V1608,
  V1609,
  V1643,
  V1644,
  V1646,
  \V1351(0) ,
  V1735,
  \V1334(0) ,
  \[10] ,
  \[11] ,
  \[12] ,
  V1842,
  V1844,
  V1846,
  V1848,
  \[13] ,
  V1850,
  V1852,
  \[14] ,
  V1867,
  \[15] ,
  V1871,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \V759(0) ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  V1978,
  V1979,
  \[26] ,
  \[27] ,
  \[28] ,
  \[100] ,
  \[29] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[30] ,
  \V1357(0) ,
  \[108] ,
  \[31] ,
  \[109] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \V1395(0) ,
  \[37] ,
  \V2081(0) ,
  \[38] ,
  \[110] ,
  \[39] ,
  \[300] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \[116] ,
  \[306] ,
  \[117] ,
  \[40] ,
  \[307] ,
  \[118] ,
  \[41] ,
  \[119] ,
  \[42] ,
  \[309] ,
  \[43] ,
  \[44] ,
  \V2064(0) ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[120] ,
  \[49] ,
  \[500] ,
  \[121] ,
  \[311] ,
  \[501] ,
  \[122] ,
  \[502] ,
  \[123] ,
  \[503] ,
  \[124] ,
  \[504] ,
  \[125] ,
  \[505] ,
  \[126] ,
  \[127] ,
  \[50] ,
  \[317] ,
  \[507] ,
  \[128] ,
  \[51] ,
  \[318] ,
  \[508] ,
  \[129] ,
  \[52] ,
  \[319] ,
  \[509] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[130] ,
  \[59] ,
  \[320] ,
  \[510] ,
  \[131] ,
  \[321] ,
  \[511] ,
  \[132] ,
  \[512] ,
  \[133] ,
  \[323] ,
  \[134] ,
  \[324] ,
  \[135] ,
  \[325] ,
  \[136] ,
  \[326] ,
  \[137] ,
  \[60] ,
  \[327] ,
  \[138] ,
  \[61] ,
  \[328] ,
  \[139] ,
  \[62] ,
  \[329] ,
  \V445(0) ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[140] ,
  \[69] ,
  \[330] ,
  \[141] ,
  \[142] ,
  \[143] ,
  \[333] ,
  \[523] ,
  \[144] ,
  \[334] ,
  \[145] ,
  \[335] ,
  \[146] ,
  \[147] ,
  \[70] ,
  \[337] ,
  \[527] ,
  \[148] ,
  \[71] ,
  \[338] ,
  \[149] ,
  \[72] ,
  \[339] ,
  \[73] ,
  \V1417(0) ,
  \[74] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[150] ,
  \[340] ,
  \V1455(0) ,
  \[151] ,
  \[341] ,
  \[152] ,
  \[342] ,
  \[153] ,
  \V1999(0) ,
  \[343] ,
  \[154] ,
  \[155] ,
  \[345] ,
  \[156] ,
  \[536] ,
  \[157] ,
  \[347] ,
  \[537] ,
  \[158] ,
  \[348] ,
  \[538] ,
  \[159] ,
  \[82] ,
  \[349] ,
  \[539] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \V336(0) ,
  \[160] ,
  \V487(0) ,
  \V1306(0) ,
  \[89] ,
  \[350] ,
  \[540] ,
  \[161] ,
  \[351] ,
  \[541] ,
  \[162] ,
  \[542] ,
  \[163] ,
  \[353] ,
  \[543] ,
  \[164] ,
  \[354] ,
  \[544] ,
  \[355] ,
  \[545] ,
  \[166] ,
  \[356] ,
  \[546] ,
  V2014,
  \[167] ,
  \[90] ,
  \[547] ,
  V2025,
  V2027,
  V2028,
  \[168] ,
  V2029,
  \[91] ,
  V2034,
  \[169] ,
  V2039,
  \[92] ,
  \[359] ,
  V2045,
  V2047,
  \[93] ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[170] ,
  \[99] ,
  \[171] ,
  \[361] ,
  \[172] ,
  \[362] ,
  \[173] ,
  \[174] ,
  \[364] ,
  \[175] ,
  \[365] ,
  V2106,
  \[176] ,
  V2109,
  \[366] ,
  \V1681(0) ,
  \[177] ,
  \[367] ,
  V2122,
  \[178] ,
  \[368] ,
  \[179] ,
  \[369] ,
  \[180] ,
  \[370] ,
  \[181] ,
  \[371] ,
  \[182] ,
  \[372] ,
  \[183] ,
  \[373] ,
  \[184] ,
  \[374] ,
  \[185] ,
  \[375] ,
  \[186] ,
  \[187] ,
  \[188] ;
assign
  \[189]  = (\[536]  & V725) | (\[330]  & \V108(2) ),
  \V1213(10)  = \[71] ,
  \V1213(11)  = \[70] ,
  \[190]  = (\[536]  & V700) | (\[330]  & \V108(3) ),
  \[380]  = (~\[286]  & ~\V78(1) ) | (\[286]  & \V78(1) ),
  \V1647(0)  = \[415]  | V726,
  \[191]  = (\[330]  & \V108(4) ) | ~\[388] ,
  \[381]  = (~\[287]  & ~\V78(5) ) | (\[287]  & \V78(5) ),
  \[192]  = (\[412]  & \V108(5) ) | \[538] ,
  \[382]  = (~\[288]  & ~\V84(3) ) | (\[288]  & \V84(3) ),
  \[193]  = (\[404]  & \V124(5) ) | ((\[399]  & \V213(5) ) | (\[393]  & \V100(5) )),
  \[383]  = (~\[289]  & ~\V88(1) ) | (\[289]  & \V88(1) ),
  \[194]  = (\[442]  & \V108(4) ) | ((\[404]  & \V124(4) ) | ((\[399]  & \V213(4) ) | (\[393]  & \V100(4) ))),
  \[384]  = (~\[290]  & ~\[197] ) | (\[290]  & \[197] ),
  \[195]  = (\[442]  & \V108(3) ) | ((\[404]  & \V124(3) ) | ((\[399]  & \V213(3) ) | (\[393]  & \V100(3) ))),
  \[385]  = (~\[291]  & ~\[199] ) | (\[291]  & \[199] ),
  \[196]  = (\[442]  & \V108(2) ) | ((\[404]  & \V124(2) ) | ((\[399]  & \V213(2) ) | (\[393]  & \V100(2) ))),
  \[386]  = (~\[292]  & ~\[204] ) | (\[292]  & \[204] ),
  \[197]  = (\[442]  & \V108(1) ) | ((\[404]  & \V124(1) ) | ((\[399]  & \V213(1) ) | (\[393]  & \V100(1) ))),
  \[387]  = (~\[293]  & ~\[207] ) | (\[293]  & \[207] ),
  \[198]  = (\[442]  & \V108(0) ) | ((\[404]  & \V124(0) ) | ((\[399]  & \V213(0) ) | (\[393]  & \V100(0) ))),
  \[388]  = ~\V15(0)  | \V16(0) ,
  \[199]  = \[359]  & \V132(1) ,
  \[389]  = \[328]  | ~\V199(2) ,
  \V1421(0)  = (\[415]  & V2122) | ((\[415]  & \V60(0) ) | ((V726 & ~\V174(0) ) | (\V1395(0)  & ~\V174(0) ))),
  \V470(0)  = (\[350]  & (V454 & ~V1852)) | ((~\[434]  & ~V1852) | (V1852 & V446)),
  \V1440(0)  = \[127] ,
  \[0]  = ~\[91] ,
  \[1]  = (~\[354]  & (~\[325]  & (~\[324]  & (~V954 & (\V1255(2)  & ~V433))))) | ((~\[418]  & (~\[354]  & (~\[325]  & (~\[324]  & ~V433)))) | ((~\[354]  & (~\[325]  & (~\[324]  & (\V1255(3)  & ~V433)))) | ((~\[354]  & (~\[325]  & (~\[324]  & (\V1255(0)  & ~V433)))) | (~\[354]  & (~\[325]  & (~\[324]  & \[238] )))))),
  \[390]  = \[329]  | ~\V194(3) ,
  \V1833(0)  = \[184] ,
  \[2]  = (~\[370]  & (~\[369]  & (~\[326]  & (~V955 & (\V1255(2)  & ~\V1681(0) ))))) | (~\[370]  & (~\[369]  & (\[341]  & (~\[326]  & ~\V1681(0) )))),
  \[3]  = \V10(0)  & \V13(0) ,
  \V731(0)  = \[374]  & (V701 & ~V721),
  \[4]  = \[120]  | (\[118]  | (\[99]  | (\[95]  | (\[94]  | (\[61]  | (\[56]  | \[54] )))))),
  \[393]  = V736,
  \[5]  = (\V203(0)  & \V35(0) ) | V697,
  \V2019(0)  = (\V1647(0)  & (~V1445 & ~\[65] )) | V2014,
  \[394]  = (~V1979 & (~V735 & \V14(0) )) | (~V1979 & (\V14(0)  & ~\V56(0) )),
  \[6]  = (\V1681(0)  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & (~\V248(0)  & (\V288(7)  & \V288(6) ))))))) | ((\[438]  & (~\[281]  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & ~\V248(0) )))))) | ((\[437]  & (~\[282]  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & ~\V248(0) )))))) | ((\[354]  & (~\[280]  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & ~\V248(0) )))))) | ((\[326]  & (~\[280]  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & ~\V248(0) )))))) | ((~\[318]  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & (~\V248(0)  & \V288(7) )))))) | ((~\[282]  & (\V1681(0)  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & ~\V248(0) )))))) | ((~\[281]  & (\V1681(0)  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & ~\V248(0) )))))) | ((\[160]  & (\V247(0)  & (\V246(0)  & (\V245(0)  & (\V244(0)  & (\V243(0)  & ~\V248(0) )))))) | (V1867 & (\[160]  & ~\V248(0) )))))))))),
  \[7]  = \[486]  | (~\[317]  | (~\[230]  | (~\[9]  | \[6] ))),
  \[396]  = V1646 & ~V695,
  \V1536(0)  = \[139] ,
  \[8]  = ~\[435]  | (V695 | \V15(0) ),
  \V321(2)  = \[0] ,
  \[9]  = (~V695 & (\[52]  & (\V66(0)  & ~\V215(0) ))) | ((\[539]  & \[65] ) | ((~\[365]  & \V56(0) ) | ((\[327]  & V411) | ((V710 & \[65] ) | ((\V1681(0)  & \[65] ) | ((\V1681(0)  & \V70(0) ) | ((\V1681(0)  & \V59(0) ) | ((\V731(0)  & \[65] ) | ((\V174(0)  & \V56(0) ) | (\[512]  | (\[355]  | \[160] ))))))))))),
  \V585(0)  = \[39] ,
  \[399]  = V735,
  \V1480(0)  = \[132] ,
  \V1741(0)  = \[163] ,
  \V1760(0)  = \[168] ,
  \V2078(0)  = 0,
  \V493(0)  = (\V473(0)  & (~V1850 & V437)) | ((V1850 & V441) | ~\[337] ),
  \V1463(0)  = (\V1455(0)  & (~\V259(0)  & ~\V258(0) )) | (\V1455(0)  & (\V259(0)  & \V258(0) )),
  \V1331(0)  = (\[471]  & V1320) | (V1312 & V1848),
  \V603(0)  = \[43] ,
  \V1781(1)  = \[171] ,
  \V1781(0)  = \[172] ,
  \V1726(0)  = \[161] ,
  V356 = \[1] ,
  V357 = \[2] ,
  \V1745(0)  = \[164] ,
  \V1896(0)  = \[187] ,
  \V1613(1)  = \[145] ,
  V373 = \[3] ,
  V377 = \[5] ,
  V379 = (\[484]  & \[65] ) | (V701 & \[65] ),
  \V1613(0)  = \[144] ,
  \V511(0)  = \[14] ,
  \V2002(0)  = (V1445 & (~\[65]  & (\V272(0)  & (\V134(0)  & (\V134(1)  & (\V242(0)  & ~\V275(0) )))))) | ((\[416]  & (\V1647(0)  & (~V1445 & (~\[65]  & \V242(0) )))) | ((~\[364]  & (~\[65]  & (\V272(0)  & ~\V275(0) ))) | ((~\[364]  & (~V1445 & ~\[65] )) | \V1999(0) ))),
  \V1467(0)  = \[130] ,
  \V1709(1)  = \[157] ,
  \V1709(0)  = \[158] ,
  \V1709(3)  = \[155] ,
  V411 = \[539]  & V687,
  \V1709(2)  = \[156] ,
  \V758(0)  = (\[475]  & (~V751 & (~V750 & ~V749))) | (\[545]  & (~V742 & ~V738)),
  V432 = \[10] ,
  V433 = V749 & ~\[65] ,
  V437 = (~V1298 & V1850) | (V1298 & ~V1850),
  V439 = (~V1302 & V1852) | (V1302 & ~V1852),
  \V1709(4)  = \[154] ,
  \V1354(0)  = (\[338]  & (\V1334(0)  & ~V1846)) | (V1846 & V1307),
  V440 = (~\[280]  & ~V1307) | (\[280]  & V1307),
  V441 = (~\[501]  & ~V439) | (\[501]  & V439),
  V446 = (~V440 & \V445(0) ) | (V440 & ~\V445(0) ),
  V451 = (~\[280]  & (~V440 & ~V1312)) | ((\[280]  & (~V440 & V1312)) | ((V440 & (~V1312 & \V445(0) )) | (V1312 & V446))),
  V452 = (V437 & V441) | ~\[414] ,
  V454 = (~\[414]  & ~V446) | (\[414]  & V446),
  V456 = \[509]  & V451,
  \V1898(0)  = \[189] ,
  \V1392(0)  = \[119] ,
  \V1653(0)  = \[353]  | (V746 | (V743 | (V744 | \[152] ))),
  \V1243(7)  = \[84] ,
  \V1243(6)  = \[85] ,
  V505 = (\[372]  & \V56(0) ) | ((~\[277]  & \V56(0) ) | ~\[416] ),
  \V1243(9)  = \[82] ,
  \V1337(0)  = (~V1848 & ~V1302) | (V1848 & V1302),
  V512 = \[15] ,
  \V1243(8)  = \[83] ,
  \V609(0)  = \[44] ,
  V527 = \[16] ,
  V537 = \[17] ,
  V538 = \[18] ,
  V539 = \[19] ,
  V540 = \[20] ,
  \V812(0)  = (\[502]  & \V62(0) ) | ((~V976 & \V56(0) ) | (V741 & \V65(0) )),
  V541 = \[21] ,
  V542 = \[22] ,
  V543 = \[23] ,
  V544 = \[24] ,
  V545 = \[25] ,
  V546 = \[26] ,
  V547 = \[27] ,
  V548 = \[28] ,
  \V2061(0)  = (~\[508]  & ~V2034) | (\[508]  & V2034),
  \V798(0)  = \[63] ,
  \V1243(1)  = \[90] ,
  V587 = \[40] ,
  \V1243(0)  = \[91] ,
  \V1243(3)  = \[88] ,
  \V1243(2)  = \[89] ,
  \V572(3)  = \[35] ,
  \[200]  = (\[400]  & \V118(5) ) | (\[359]  & \V132(7) ),
  \V1243(5)  = \[86] ,
  \V572(2)  = \[36] ,
  \[201]  = (\[400]  & \V118(4) ) | (\[359]  & \V132(6) ),
  \V1243(4)  = \[87] ,
  \V572(5)  = \[33] ,
  \[202]  = (\[400]  & \V118(3) ) | (\[359]  & \V132(5) ),
  \V572(4)  = \[34] ,
  \[203]  = (\[400]  & \V118(2) ) | (\[359]  & \V132(4) ),
  \V1281(0)  = \[105] ,
  \[204]  = (\[400]  & \V118(1) ) | (\[359]  & \V132(3) ),
  \[205]  = (\[400]  & \V118(0) ) | (\[359]  & \V132(2) ),
  \V1674(0)  = (\[537]  & (\V261(0)  & (\V165(3)  & (\V165(1)  & (\V165(7)  & (\V165(6)  & (\V165(5)  & (\V165(4)  & (\V165(2)  & \V165(0) ))))))))) | (\V261(0)  & (~\V204(0)  & (\V165(3)  & (\V165(1)  & (\V165(7)  & (\V165(6)  & (\V165(5)  & (\V165(4)  & (\V165(2)  & \V165(0) ))))))))),
  \V572(1)  = \[37] ,
  V620 = \[45] ,
  V621 = \[46] ,
  \[206]  = (\[359]  & \V132(0) ) | (V751 & \V108(5) ),
  \V572(0)  = \[38] ,
  V630 = \[47] ,
  \[207]  = (\[258]  & \V46(0) ) | (V743 & \V118(7) ),
  \[208]  = (\[258]  & \V48(0) ) | (V743 & \V118(6) ),
  \V1693(0)  = \[153] ,
  V646 = ~\[449]  & (\V257(4)  & (\V257(3)  & \V257(5) )),
  V650 = \[212] ,
  V651 = \[213] ,
  V652 = \[214] ,
  V653 = \[215] ,
  V654 = \[216] ,
  \[209]  = (\[388]  & (~V743 & (\V110(0)  & \V14(0) ))) | ((\[388]  & (\V110(0)  & (\V14(0)  & ~\V56(0) ))) | ((~V743 & (\V110(0)  & (\V108(4)  & \V14(0) ))) | ((~V743 & (\V110(0)  & (~\V101(0)  & \V14(0) ))) | ((\V110(0)  & (\V108(4)  & (\V14(0)  & ~\V56(0) ))) | ((\V110(0)  & (~\V101(0)  & (\V14(0)  & ~\V56(0) ))) | ((V700 & (\[166]  & ~\V110(0) )) | (V700 & (~\V110(0)  & \V102(0) )))))))),
  V655 = \[217] ,
  V656 = \[218] ,
  V657 = \[50] ,
  \V591(0)  = \[41] ,
  \V572(7)  = \[31] ,
  V687 = \V169(1)  & \V1395(0) ,
  \V572(6)  = \[32] ,
  V695 = \V165(1)  & (~\V165(2)  & \V165(0) ),
  V697 = \V165(1)  & (\V165(2)  & (~\V165(0)  & \V203(0) )),
  \V572(9)  = \[29] ,
  \V572(8)  = \[30] ,
  \[210]  = (~\[343]  & (~\[248]  & ~\V134(1) )) | (\[343]  & (~\[248]  & \V134(1) )),
  \[400]  = V743,
  \[211]  = (~\[343]  & (~\[248]  & (~\[210]  & ~\V134(0) ))) | ((\[343]  & (~\[248]  & \V134(0) )) | (\[210]  & \V134(0) )),
  \[401]  = (~V1978 & (~V736 & \V14(0) )) | (~V1978 & (\V14(0)  & ~\V56(0) )),
  \V1992(1)  = \[210] ,
  \[212]  = (~\[497]  & ~\V257(0) ) | (\[497]  & \V257(0) ),
  \[402]  = \[333] ,
  \V1992(0)  = \[211] ,
  \[213]  = (~\[498]  & ~\V257(1) ) | (\[498]  & \V257(1) ),
  \V404(0)  = (~\[374]  & (V701 & ~\V149(3) )) | (~V687 & \V730(0) ),
  V700 = ~\[371]  & ~\V149(0) ,
  V701 = \[479]  & ~\V149(1) ,
  V702 = ~\V149(2)  & (\V149(1)  & ~\V149(0) ),
  \[214]  = (~V646 & \V257(2) ) | (V646 & ~\V257(2) ),
  V707 = \[51] ,
  \[404]  = V742,
  V710 = \[484]  & \V149(3) ,
  \[215]  = (~V646 & (~\[216]  & \V257(4) )) | (~V646 & \V257(3) ),
  V721 = V701 & \V149(3) ,
  \[216]  = (~\[499]  & ~\V257(4) ) | (\[499]  & \V257(4) ),
  V725 = \[547]  & (~\V149(3)  & \V149(4) ),
  V726 = \[547]  & (~\V149(3)  & ~\V149(4) ),
  V727 = \[547]  & \V149(3) ,
  \V423(0)  = \[9] ,
  \[217]  = (~\[449]  & ~\V257(5) ) | (\[449]  & \V257(5) ),
  V735 = \[481]  & \[367] ,
  V736 = \[540]  & \[368] ,
  V737 = \[541]  & \[367] ,
  \[407]  = (~\V41(0)  & ~\V45(0) ) | (\V41(0)  & \V45(0) ),
  V738 = \[545]  & \[441] ,
  V739 = \[481]  & \[441] ,
  V740 = \[441]  & (\[368]  & ~\V149(7) ),
  V741 = \[541]  & \[441] ,
  V742 = \[545]  & \[482] ,
  V743 = \[482]  & \[481] ,
  V744 = \[482]  & (\[368]  & ~\V149(7) ),
  \[218]  = (~\V257(6)  & \V257(7) ) | (\V257(6)  & ~\V257(7) ),
  V745 = \[541]  & \[482] ,
  V746 = \[481]  & ~\[374] ,
  V747 = \V759(0)  & ~\V149(7) ,
  \[408]  = ~\V14(0)  | \V289(0) ,
  V749 = \[540]  & (\[475]  & ~\V149(6) ),
  V750 = \[475]  & (\[367]  & (~\V149(6)  & \V149(7) )),
  V751 = \[540]  & (\[475]  & \V149(6) ),
  \[219]  = (~V1366 & \V268(0) ) | (V1366 & ~\V268(0) ),
  \[409]  = ~\[371]  | ~\V149(0) ,
  V763 = \[52] ,
  V768 = \V759(0)  & (\V149(7)  & ~\V174(0) ),
  V769 = V725 & ~\V174(0) ,
  V775 = \[53] ,
  V778 = \[54] ,
  V779 = \[55] ,
  V780 = \[56] ,
  V781 = \[57] ,
  V782 = \[58] ,
  V783 = \[59] ,
  V784 = \[60] ,
  V787 = \[61] ,
  V789 = \[62] ,
  V799 = \[543]  & (\V165(3)  & (~\V165(6)  & \V70(0) )),
  \V2084(0)  = (\V2064(0)  & (~V1842 & V2025)) | ~\[339] ,
  \[220]  = (~V1366 & (~\[221]  & \V268(2) )) | (~V1366 & \V268(1) ),
  \[221]  = (~\[500]  & ~\V268(2) ) | (\[500]  & \V268(2) ),
  \[222]  = (~\[450]  & ~\V268(3) ) | (\[450]  & \V268(3) ),
  \[412]  = ~V751 | ~\V56(0) ,
  \[223]  = (~\V268(4)  & \V268(5) ) | (\V268(4)  & ~\V268(5) ),
  \[413]  = ~V2106 | V379,
  V801 = \[64] ,
  \[224]  = (~\V1255(3)  & V437) | (\V1255(3)  & ~V437),
  \[414]  = V437 | V441,
  \[225]  = (~V2025 & \V1255(3) ) | (V2025 & ~\V1255(3) ),
  \[415]  = V727 | V769,
  \[226]  = (~\V1255(3)  & V1298) | (\V1255(3)  & ~V1298),
  \[416]  = ~\[415]  | ~\V56(0) ,
  \[227]  = (~V2029 & ~\V1255(2) ) | (V2029 & \V1255(2) ),
  \[417]  = ~\V288(7)  | \V288(6) ,
  \[228]  = (~\V1255(2)  & V1302) | (\V1255(2)  & ~V1302),
  \[418]  = \V288(7)  | \V288(6) ,
  \[229]  = ~\V1417(0) ,
  V856 = (~\[295]  & (~\[282]  & (\[227]  & (~V2045 & (V2025 & ~\V1255(3) ))))) | ((\[544]  & (~\[282]  & (\[227]  & (V2045 & ~\V1255(3) )))) | (~\[295]  & (~\[282]  & (~\[227]  & (~V2025 & \V1255(3) ))))),
  V866 = (\[544]  & (~\[282]  & (\[227]  & (~\[225]  & V2034)))) | (~\[295]  & (~\[282]  & (\[227]  & (~\[225]  & ~V2034)))),
  V896 = (~\[281]  & (\[238]  & (~\[228]  & (V1320 & (V1318 & (~\V1255(3)  & (\V1255(0)  & V1298))))))) | ((~\[281]  & (\[238]  & (\[228]  & (V1320 & (V1318 & (\V1255(3)  & (\V1255(0)  & ~V1298))))))) | ((~\[281]  & (~\[232]  & (~\[228]  & (V1320 & (~V1318 & (~\V1255(3)  & (\V1255(0)  & V1298))))))) | ((~\[281]  & (~\[232]  & (\[228]  & (V1320 & (~V1318 & (\V1255(3)  & (\V1255(0)  & ~V1298))))))) | ((\[544]  & (~\[281]  & (~\[228]  & (~V1320 & (V1318 & (~\V1255(3)  & V1298)))))) | ((\[544]  & (~\[281]  & (\[228]  & (~V1320 & (V1318 & (\V1255(3)  & ~V1298)))))) | ((~\[295]  & (~\[281]  & (~\[228]  & (~V1320 & (~V1318 & (~\V1255(3)  & V1298)))))) | (~\[295]  & (~\[281]  & (\[228]  & (~V1320 & (~V1318 & (\V1255(3)  & ~V1298)))))))))))),
  \[230]  = (~V687 & ~\[52] ) | ~\[65] ,
  \[231]  = \[229]  & ~V1125,
  \[232]  = \V1255(1)  | V433,
  \[233]  = (~V1587 & \V94(0) ) | (V1587 & ~\V94(0) ),
  \[234]  = (~V1589 & \V94(1) ) | (V1589 & ~\V94(1) ),
  V906 = (~\[295]  & (~\[281]  & (~\[228]  & (~\[226]  & (~V1312 & ~V1307))))) | ((\[295]  & (~\[281]  & (~\[232]  & (~\[228]  & (~\[226]  & V1312))))) | (\[544]  & (~\[281]  & (~\[228]  & (~\[226]  & V1307))))),
  \[235]  = \[231]  & V2122,
  \V1864(0)  = \[186] ,
  \[236]  = (~V1646 & ~\V149(7) ) | ~V701,
  \[237]  = ~V695 | \V165(7) ,
  V936 = (~\[280]  & (\[238]  & (\[224]  & (V456 & (~\V1255(2)  & (\V1255(0)  & (V454 & ~V452))))))) | ((~\[280]  & (\[238]  & (\[224]  & (V456 & (\V1255(2)  & (\V1255(0)  & (V454 & V452))))))) | ((~\[280]  & (~\[232]  & (\[224]  & (V456 & (~\V1255(2)  & (\V1255(0)  & (~V454 & ~V452))))))) | ((~\[280]  & (~\[232]  & (\[224]  & (V456 & (\V1255(2)  & (\V1255(0)  & (~V454 & V452))))))) | ((\[544]  & (~\[280]  & (\[224]  & (~V456 & (~\V1255(2)  & (V454 & ~V452)))))) | ((\[544]  & (~\[280]  & (\[224]  & (~V456 & (\V1255(2)  & (V454 & V452)))))) | ((~\[295]  & (~\[280]  & (\[224]  & (~V456 & (~\V1255(2)  & (~V454 & ~V452)))))) | (~\[295]  & (~\[280]  & (\[224]  & (~V456 & (\V1255(2)  & (~V454 & V452)))))))))))),
  \[238]  = \V1255(1)  & ~V433,
  V946 = (~\[280]  & (\[238]  & (~\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~V441 & (V446 & ~V451))))))) | ((~\[280]  & (\[238]  & (~\[224]  & (~\V1255(2)  & (\V1255(0)  & (~V441 & (V446 & V451))))))) | ((~\[280]  & (\[238]  & (~\[224]  & (\V1255(2)  & (~\V1255(0)  & (V441 & (V446 & ~V451))))))) | ((~\[280]  & (\[238]  & (~\[224]  & (\V1255(2)  & (\V1255(0)  & (V441 & (V446 & V451))))))) | ((~\[280]  & (~\[232]  & (~\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~V441 & (~V446 & ~V451))))))) | ((~\[280]  & (~\[232]  & (~\[224]  & (~\V1255(2)  & (\V1255(0)  & (~V441 & (~V446 & V451))))))) | ((~\[280]  & (~\[232]  & (~\[224]  & (\V1255(2)  & (~\V1255(0)  & (V441 & (~V446 & ~V451))))))) | (~\[280]  & (~\[232]  & (~\[224]  & (\V1255(2)  & (\V1255(0)  & (V441 & (~V446 & V451))))))))))))),
  V954 = ~\[318]  & (\V1255(2)  & \V288(7) ),
  V955 = ~\[341]  & (\V1255(2)  & \V288(7) ),
  V966 = \[68] ,
  \V597(0)  = \[42] ,
  V976 = (~\[353]  & (\[319]  & (~V746 & (~V743 & ~V744)))) | (~\[353]  & (~V746 & (~V743 & (~\V1681(0)  & ~V744)))),
  V986 = \[69] ,
  \[240]  = \[235]  & (\V1421(0)  & ~\V1681(0) ),
  \[430]  = \[337]  | \V470(0) ,
  \[431]  = 0,
  \[432]  = 0,
  \[244]  = ~\V404(0)  | ~\V56(0) ,
  \[434]  = \[350]  | V454,
  \[245]  = ~V741 | ~\V62(0) ,
  \[435]  = (V411 & \V62(0) ) | \[355] ,
  \V1492(0)  = \[134] ,
  \[437]  = \[369]  | \[324] ,
  \[248]  = ~V2109 | ~V2106,
  \[438]  = \[370]  | \[325] ,
  \V500(0)  = \[12] ,
  \V467(0)  = (\[434]  & V456) | (V1852 & V451),
  \[441]  = ~\V149(4)  & \V149(5) ,
  \[252]  = ~\V807(0)  & \V14(0) ,
  \[442]  = V750,
  \[253]  = ~\V1647(0)  | ~\[65] ,
  \[443]  = ~\V13(0)  & \V10(0) ,
  \[444]  = ~\[237]  | \V302(0) ,
  \V1901(0)  = \[192] ,
  \V1717(0)  = \[159] ,
  \[445]  = \V731(0)  | V721,
  \[446]  = \V807(0)  | V697,
  \[257]  = \[229]  & V1125,
  \[258]  = V740 | V741,
  \[448]  = ~\V759(0)  | ~\V56(0) ,
  \[449]  = ~\V257(6)  | ~\V257(7) ,
  \V634(0)  = \[48] ,
  \V1213(7)  = \[74] ,
  \V1439(0)  = \[126] ,
  \V1213(6)  = \[75] ,
  \V1213(9)  = \[72] ,
  \[260]  = ~\V66(0)  | ~\V215(0) ,
  \[450]  = ~\V268(4)  | ~\V268(5) ,
  \V1213(8)  = \[73] ,
  \[262]  = ~\[248]  & \V2019(0) ,
  \[263]  = ~V710 | V687,
  \V375(0)  = \[4] ,
  \[266]  = ~V695 | \V290(0) ,
  \[267]  = \[266]  | ~\V165(7) ,
  \V1213(1)  = \V1255(1) ,
  V1125 = ~\V1681(0)  & \[52] ,
  \V1213(0)  = \V1255(0) ,
  \V1213(3)  = \V1255(3) ,
  \V1213(2)  = \V1255(2) ,
  \V1757(0)  = \V15(0) ,
  \V1213(5)  = \[76] ,
  \V1960(1)  = \[207] ,
  \V1213(4)  = \[77] ,
  \V1960(0)  = \[208] ,
  \[270]  = ~\V1422(0) ,
  \[271]  = \[240]  & \V1395(0) ,
  \V1512(1)  = \[138] ,
  \[272]  = \[240]  & ~\V1395(0) ,
  \V1512(3)  = \[136] ,
  \[464]  = \[372]  | \V1647(0) ,
  \V410(0)  = \[8] ,
  \V1512(2)  = \[137] ,
  \[465]  = (\V759(0)  & (\[52]  & ~\V174(0) )) | \V758(0) ,
  \V2033(0)  = (~V2027 & V1844) | (V2027 & V1842),
  \[277]  = ~V739 | V1476,
  \[279]  = ~V737 | ~\V66(0) ,
  V1256 = \[92] ,
  V1257 = \[93] ,
  V1258 = \[94] ,
  V1259 = \[95] ,
  \V1759(0)  = \[167] ,
  V1260 = \[96] ,
  V1261 = \[97] ,
  V1262 = \[98] ,
  V1263 = \[99] ,
  V1264 = \[100] ,
  V1265 = \[101] ,
  V1266 = \[102] ,
  V1267 = \[103] ,
  V1298 = (~V2025 & V1846) | (V2025 & ~V1846),
  \[280]  = ~\V288(1)  | ~\V288(0) ,
  \[281]  = ~\V288(3)  | ~\V288(2) ,
  \[471]  = V1318 | (V1302 | ~V1298),
  \[282]  = ~\V288(5)  | ~\V288(4) ,
  \[472]  = V2045,
  \[285]  = ~V1867 | ~\V194(0) ,
  \[475]  = V702 & \V149(3) ,
  V1300 = (~V2029 & V1848) | (V2029 & ~V1848),
  V1301 = (~\[281]  & ~V2034) | (\[281]  & V2034),
  V1302 = (~\[503]  & ~V1300) | (\[503]  & V1300),
  V1307 = (~V1301 & \V1306(0) ) | (V1301 & ~\V1306(0) ),
  \[286]  = (~\V78(3)  & \V78(2) ) | (\V78(3)  & ~\V78(2) ),
  V1312 = (~\[281]  & (~V1301 & ~V2039)) | ((V1301 & (~V2039 & \V1306(0) )) | (V2039 & V1307)),
  V1318 = (~\[504]  & ~V1307) | (\[504]  & V1307),
  \[287]  = (~\V84(0)  & \V84(1) ) | (\V84(0)  & ~\V84(1) ),
  V1320 = \[511]  & V1312,
  \V1552(1)  = \[142] ,
  \[288]  = (~\V84(4)  & \V84(5) ) | (\V84(4)  & ~\V84(5) ),
  \[478]  = ~V2122 & (~\V1421(0)  & ~\V1681(0) ),
  \V398(0)  = \[7] ,
  \V1552(0)  = \[143] ,
  \[289]  = (~\V88(3)  & \V88(2) ) | (\V88(3)  & ~\V88(2) ),
  \[479]  = \V149(2)  & ~\V149(0) ,
  V1365 = \[111] ,
  V1366 = ~\[450]  & (\V268(2)  & (\V268(1)  & \V268(3) )),
  V1370 = \[219] ,
  V1371 = \[220] ,
  \V508(0)  = \[13] ,
  V1372 = \[221] ,
  V1373 = \[222] ,
  V1374 = \[223] ,
  V1375 = \[112] ,
  V1378 = \[113] ,
  V1380 = \[114] ,
  V1382 = \[115] ,
  V1384 = \[116] ,
  V1386 = \[117] ,
  \V1629(0)  = \[147] ,
  V1387 = \[118] ,
  \V1255(1)  = (\[272]  & \V183(1) ) | ((\[271]  & \V223(1) ) | (\[270]  & \V32(1) )),
  \V1255(0)  = (\[272]  & \V183(0) ) | ((\[271]  & \V223(0) ) | (\[270]  & \V32(0) )),
  \V1255(3)  = (\[272]  & \V183(3) ) | ((\[271]  & \V223(3) ) | (\[270]  & \V32(3) )),
  \[290]  = (~\[196]  & \[195] ) | (\[196]  & ~\[195] ),
  \[480]  = ~V2109 & ~\V2019(0) ,
  \V1255(2)  = (\[272]  & \V183(2) ) | ((\[271]  & \V223(2) ) | (\[270]  & \V32(2) )),
  \[291]  = (~\[194]  & \[193] ) | (\[194]  & ~\[193] ),
  \[481]  = \[366]  & \V149(7) ,
  \V1274(0)  = \[104] ,
  \V730(0)  = (\[441]  & (\[51]  & (\V88(3)  & \V88(2) ))) | (\[367]  & (\[51]  & (~\V88(3)  & ~\V88(2) ))),
  \[292]  = (~\[203]  & \[202] ) | (\[203]  & ~\[202] ),
  \[482]  = \V149(4)  & ~\V149(5) ,
  \[293]  = (~\[201]  & \[200] ) | (\[201]  & ~\[200] ),
  \[483]  = \[333] ,
  \[294]  = V736 | V735,
  \[484]  = V700 & ~\V174(0) ,
  \[295]  = \[232]  | \V1255(0) ,
  V1402 = (\[505]  & \[52] ) | (\[52]  & \V59(0) ),
  \[486]  = \V214(0)  | \V43(0) ,
  \V807(0)  = \[444]  | (~\[266]  | \V2002(0) ),
  V1423 = \[120] ,
  V1426 = \[121] ,
  V1428 = \[122] ,
  V1429 = \[123] ,
  V1431 = \[124] ,
  V1432 = \[125] ,
  V1445 = (~V769 & \V278(0) ) | (\V278(0)  & ~\V277(0) ),
  \V826(0)  = \[67] ,
  \V1422(0)  = (V769 & \V60(0) ) | ((V721 & \V60(0) ) | ~\V1417(0) ),
  V1470 = \[131] ,
  V1476 = (~\[234]  & (~V1590 & (V745 & \V56(0) ))) | ((~\[234]  & (~V1590 & (V739 & \V56(0) ))) | ((~\[234]  & (~V1590 & (V744 & \V56(0) ))) | ((\[234]  & (V1590 & (V745 & \V56(0) ))) | ((\[234]  & (V1590 & (V739 & \V56(0) ))) | ((\[234]  & (V1590 & (V744 & \V56(0) ))) | ((~\[233]  & (~V1588 & (V745 & \V56(0) ))) | ((~\[233]  & (~V1588 & (V739 & \V56(0) ))) | ((~\[233]  & (~V1588 & (V744 & \V56(0) ))) | ((\[233]  & (V1588 & (V745 & \V56(0) ))) | ((\[233]  & (V1588 & (V739 & \V56(0) ))) | ((\[233]  & (V1588 & (V744 & \V56(0) ))) | ((\[413]  & (~\[234]  & ~V1590)) | ((\[413]  & (\[234]  & V1590)) | ((\[413]  & (~\[233]  & ~V1588)) | (\[413]  & (\[233]  & V1588)))))))))))))))),
  \V490(0)  = (\[337]  & (\V470(0)  & ~V1850)) | ((~\[430]  & ~V1850) | (V1850 & V446)),
  \[497]  = \[213]  | ~\V257(1) ,
  \V435(0)  = \[11] ,
  \[498]  = ~V646 | ~\V257(2) ,
  V1535 = (\[236]  & (~\V2002(0)  & (~\V1395(0)  & (~\V1647(0)  & (~\V172(0)  & (\V177(0)  & ~\V248(0) )))))) | ((\[236]  & (~\V2002(0)  & (~\V1395(0)  & (~\V172(0)  & (\V177(0)  & (~\V278(0)  & ~\V248(0) )))))) | ((\[236]  & (~\V2002(0)  & (~\V1647(0)  & (~\V171(0)  & (~\V172(0)  & (\V177(0)  & ~\V248(0) )))))) | ((\[236]  & (~\V2002(0)  & (~\V171(0)  & (~\V172(0)  & (\V177(0)  & (~\V278(0)  & ~\V248(0) )))))) | ((\[362]  & (~\V2002(0)  & (~\V1647(0)  & (\V177(0)  & (~\V248(0)  & ~\V56(0) ))))) | ((\[362]  & (~\V2002(0)  & (\V177(0)  & (~\V278(0)  & (~\V248(0)  & ~\V56(0) ))))) | ((\[307]  & (~\V2002(0)  & (V687 & (\V730(0)  & \V59(0) )))) | ((\[307]  & (~\V2002(0)  & (~\V274(0)  & ~\V271(0) ))) | (~\[244]  & (\[236]  & (~\V2002(0)  & ~\V172(0) )))))))))),
  V1537 = \[140] ,
  V1539 = \[141] ,
  \[499]  = \[217]  | ~\V257(5) ,
  \V2058(0)  = ~\[472]  | V2047,
  V1587 = (~\[380]  & ~\V78(0) ) | (\[380]  & \V78(0) ),
  V1588 = (~\[381]  & ~\V78(4) ) | (\[381]  & \V78(4) ),
  V1589 = (~\[382]  & ~\V84(2) ) | (\[382]  & \V84(2) ),
  \V473(0)  = (~V1852 & ~V441) | (V1852 & V441),
  \V1968(0)  = \[209] ,
  V1590 = (~\[383]  & ~\V88(0) ) | (\[383]  & \V88(0) ),
  \V1297(1)  = \[109] ,
  \V1481(0)  = \[133] ,
  \V1297(0)  = \[110] ,
  V1606 = (~\[384]  & ~\[198] ) | (\[384]  & \[198] ),
  V1607 = (~\[385]  & ~\[206] ) | (\[385]  & \[206] ),
  V1608 = (~\[386]  & ~\[205] ) | (\[386]  & \[205] ),
  V1609 = (~\[387]  & ~\[208] ) | (\[387]  & \[208] ),
  \V1297(3)  = \[107] ,
  \V1297(2)  = \[108] ,
  \V1297(4)  = \[106] ,
  V1643 = (\[413]  & (\V336(0)  & ~\[52] )) | ((\[351]  & (\V336(0)  & \V56(0) )) | ((V768 & (\V336(0)  & \V56(0) )) | ((\V336(0)  & (\[52]  & \V66(0) )) | (~\[279]  & \V336(0) )))),
  V1644 = (\[484]  & (~\[408]  & (\[396]  & V687))) | ((~\[408]  & (~\[362]  & (~V695 & ~\V302(0) ))) | ((~\[408]  & (\[396]  & V768)) | (~\[408]  & (\[396]  & V738)))),
  V1646 = (\V207(0)  & ~\V172(0) ) | (\V207(0)  & ~\V56(0) ),
  \V640(0)  = \[49] ,
  V1669 = \[150] ,
  V1719 = \[160] ,
  \V1351(0)  = (\V1331(0)  & ~V1846) | (V1312 & V1846),
  V1735 = (~V726 & ~\V241(0) ) | ~\V1647(0) ,
  V1736 = \[162] ,
  \V1334(0)  = (\V1337(0)  & (~V1848 & ~V1307)) | ((~\V1337(0)  & V1307) | (V1307 & V1302)),
  \[10]  = ~\[486]  & (\[317]  & (\[260]  & (\[230]  & (~V1646 & (~V1643 & (~\V1681(0)  & (~V1476 & (\[9]  & (~\[6]  & ~\V15(0) ))))))))),
  \[11]  = \[10]  | \[47] ,
  V1832 = \[183] ,
  \[12]  = ~\V14(0)  | \V271(0) ,
  V1842 = \V288(5)  & ~\V288(4) ,
  V1844 = ~\V288(5)  & \V288(4) ,
  V1846 = \V288(3)  & ~\V288(2) ,
  V1848 = ~\V288(3)  & \V288(2) ,
  \V1897(0)  = \[188] ,
  \[13]  = (~\[365]  & \V59(0) ) | ((\[258]  & \V56(0) ) | (~\[245]  | V505)),
  V1850 = \V288(1)  & ~\V288(0) ,
  V1852 = ~\V288(1)  & \V288(0) ,
  \[14]  = (\V45(0)  & ~\V43(0) ) | \V40(0) ,
  V1867 = ~\[390]  & (\V194(1)  & \V194(2) ),
  \[15]  = (~\V44(0)  & (~\V42(0)  & (~\V38(0)  & ~\V39(0) ))) | ((~\V44(0)  & (~\V42(0)  & (\V38(0)  & \V39(0) ))) | ((\V44(0)  & (\V42(0)  & (~\V38(0)  & ~\V39(0) ))) | (\V44(0)  & (\V42(0)  & (\V38(0)  & \V39(0) ))))),
  V1871 = ~\[389]  & (\V199(0)  & \V199(1) ),
  \[16]  = ~\[486]  & (\[435]  & (~V1646 & ~V695)),
  \[17]  = \V1255(0)  & V769,
  \[18]  = \V1255(1)  & V769,
  \[19]  = \V1255(2)  & V769,
  \V1652(0)  = \[149] ,
  \V1671(0)  = \[151] ,
  \V759(0)  = ~\[374]  & \[368] ,
  \[20]  = \V1255(3)  & V769,
  \[21]  = V769 & \[77] ,
  \[22]  = V769 & \[76] ,
  \[23]  = V769 & \[75] ,
  \V1899(0)  = \[190] ,
  \[24]  = V769 & \[74] ,
  \[25]  = V769 & \[73] ,
  V1978 = \[546]  & \[349] ,
  V1979 = \[546]  & V725,
  \[26]  = V769 & \[72] ,
  \[27]  = V769 & \[71] ,
  \[28]  = V769 & \[70] ,
  \[100]  = \V12(0)  & \V4(0) ,
  \[29]  = (\[402]  & \[82] ) | (\[262]  & ~\V199(4) ),
  \[101]  = \[100]  & \V52(0) ,
  \V1953(7)  = \[200] ,
  \[102]  = \V11(0)  & \V4(0) ,
  \V1953(6)  = \[201] ,
  \[103]  = \V11(0)  & \V2(0) ,
  \[104]  = (~\[464]  & (\[252]  & (~V768 & (~V747 & (~V749 & (~\V404(0)  & (~\[160]  & \V59(0) ))))))) | ((~\[464]  & (\[252]  & (~V768 & (~V749 & (~\V404(0)  & (~\[160]  & (\V174(0)  & \V59(0) ))))))) | (\[542]  & ~\[365] )),
  \[105]  = (\[396]  & V725) | ((\[394]  & \V213(0) ) | (\[348]  & V1979)),
  \[106]  = (\[394]  & \V213(5) ) | (V1979 & \V165(7) ),
  \[107]  = (\[394]  & \V213(4) ) | (V1979 & \V165(6) ),
  \[30]  = (\[262]  & (~\V199(3)  & \V199(4) )) | ((\[262]  & (\V199(3)  & ~\V199(4) )) | (\[402]  & \[83] )),
  \V1357(0)  = (\V1337(0)  & (~V1846 & V1298)) | ((V1846 & V1302) | ~\[338] ),
  \[108]  = (\[394]  & \V213(3) ) | (V1979 & \V165(5) ),
  \[31]  = (~\[328]  & (\[262]  & ~\V199(2) )) | ((\[328]  & (\[262]  & \V199(2) )) | (\[402]  & \[84] )),
  \[109]  = (\[394]  & \V213(2) ) | (V1979 & \V165(4) ),
  \[32]  = (~\[389]  & (\[262]  & ~\V199(1) )) | ((\[389]  & (\[262]  & \V199(1) )) | (\[402]  & \[85] )),
  \[33]  = (~\[389]  & (\[262]  & (~V1871 & \V199(1) ))) | ((\[262]  & (~V1871 & \V199(0) )) | (\[402]  & \[86] )),
  \[34]  = (\[262]  & (~V1871 & \V194(4) )) | ((\[262]  & (V1871 & ~\V194(4) )) | (\[402]  & \[87] )),
  \V1953(1)  = \[199] ,
  \[35]  = (~\[329]  & (\[262]  & ~\V194(3) )) | ((\[329]  & (\[262]  & \V194(3) )) | ((\[483]  & \[88] ) | (\[480]  & \V149(7) ))),
  \V1953(0)  = \[206] ,
  \[36]  = (~\[390]  & (\[262]  & ~\V194(2) )) | ((\[390]  & (\[262]  & \V194(2) )) | ((\[483]  & \[89] ) | (\[480]  & \V149(6) ))),
  \V1953(3)  = \[204] ,
  \V1395(0)  = V700 | V701,
  \[37]  = (~\[390]  & (\[262]  & (~V1867 & \V194(2) ))) | ((\[262]  & (~V1867 & \V194(1) )) | ((\[483]  & \[90] ) | (\[480]  & \V149(5) ))),
  \V2081(0)  = (\V2061(0)  & ~V1842) | (V1842 & V2034),
  \V1953(2)  = \[205] ,
  \[38]  = (\[262]  & (~V1867 & \V194(0) )) | ((\[262]  & (V1867 & ~\V194(0) )) | ((\[483]  & \[91] ) | (\[480]  & \V149(4) ))),
  \V1953(5)  = \[202] ,
  \[110]  = (\[394]  & \V213(1) ) | (V1979 & \V165(3) ),
  \[39]  = ~\V34(0) ,
  \[300]  = \[257]  & V1402,
  \V1953(4)  = \[203] ,
  \[111]  = \[542]  & (~\[502]  & (~\[323]  & (~V738 & ~\V1681(0) ))),
  \[112]  = ~\V268(5) ,
  \[113]  = \[248]  & \[58] ,
  \[114]  = (\[364]  & (\[285]  & (\V2019(0)  & (\[58]  & ~\V248(0) )))) | ((V2014 & \[58] ) | \[113] ),
  \[115]  = (V379 & \[58] ) | (V721 & \[58] ),
  \[116]  = V744 & (~V695 & (~V1476 & (\[58]  & \V56(0) ))),
  \[306]  = V702 & ~\V149(3) ,
  \[117]  = ~\[373]  & \[58] ,
  \[40]  = \[253]  & ~\V243(0) ,
  \[307]  = (~V1646 & ~\V56(0) ) | \[236] ,
  \[118]  = \V8(0)  & \V9(0) ,
  \[41]  = (\[253]  & (~\[40]  & ~\V244(0) )) | (\[40]  & \V244(0) ),
  \[119]  = (\[543]  & (\[537]  & (\[252]  & \V165(3) ))) | (\[252]  & (~V411 & (~V741 & \V65(0) ))),
  \[42]  = (\[253]  & (~\V245(0)  & (\V244(0)  & \V243(0) ))) | ((\[253]  & (\V245(0)  & ~\V244(0) )) | (\[40]  & \V245(0) )),
  \[309]  = (\[238]  & (~\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~\V493(0)  & (\V490(0)  & (~\V487(0)  & V1850))))))) | ((\[238]  & (~\[224]  & (~\V1255(2)  & (\V1255(0)  & (~\V493(0)  & (\V490(0)  & (\V487(0)  & V1850))))))) | ((\[238]  & (~\[224]  & (\V1255(2)  & (~\V1255(0)  & (\V493(0)  & (\V490(0)  & (~\V487(0)  & V1850))))))) | ((\[238]  & (~\[224]  & (\V1255(2)  & (\V1255(0)  & (\V493(0)  & (\V490(0)  & (\V487(0)  & V1850))))))) | ((\[238]  & (\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~\V493(0)  & (\V490(0)  & (~\V487(0)  & \V288(0) ))))))) | ((\[238]  & (\[224]  & (~\V1255(2)  & (\V1255(0)  & (~\V493(0)  & (\V490(0)  & (\V487(0)  & \V288(0) ))))))) | ((\[238]  & (\[224]  & (\V1255(2)  & (~\V1255(0)  & (\V493(0)  & (\V490(0)  & (~\V487(0)  & \V288(0) ))))))) | ((\[238]  & (\[224]  & (\V1255(2)  & (\V1255(0)  & (\V493(0)  & (\V490(0)  & (\V487(0)  & \V288(0) ))))))) | ((~\[232]  & (~\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~\V493(0)  & (~\V490(0)  & (~\V487(0)  & V1850))))))) | ((~\[232]  & (~\[224]  & (~\V1255(2)  & (\V1255(0)  & (~\V493(0)  & (~\V490(0)  & (\V487(0)  & V1850))))))) | ((~\[232]  & (~\[224]  & (\V1255(2)  & (~\V1255(0)  & (\V493(0)  & (~\V490(0)  & (~\V487(0)  & V1850))))))) | ((~\[232]  & (~\[224]  & (\V1255(2)  & (\V1255(0)  & (\V493(0)  & (~\V490(0)  & (\V487(0)  & V1850))))))) | ((~\[232]  & (\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~\V493(0)  & (~\V490(0)  & (~\V487(0)  & \V288(0) ))))))) | ((~\[232]  & (\[224]  & (~\V1255(2)  & (\V1255(0)  & (~\V493(0)  & (~\V490(0)  & (\V487(0)  & \V288(0) ))))))) | ((~\[232]  & (\[224]  & (\V1255(2)  & (~\V1255(0)  & (\V493(0)  & (~\V490(0)  & (~\V487(0)  & \V288(0) ))))))) | ((~\[232]  & (\[224]  & (\V1255(2)  & (\V1255(0)  & (\V493(0)  & (~\V490(0)  & (\V487(0)  & \V288(0) ))))))) | V936))))))))))))))),
  \[43]  = (\[253]  & (~\[42]  & (~\V246(0)  & \V245(0) ))) | ((\[253]  & (\V246(0)  & ~\V245(0) )) | (\[42]  & \V246(0) )),
  \[44]  = (\[253]  & (~\[43]  & (~\V247(0)  & \V246(0) ))) | ((\[253]  & (\V247(0)  & ~\V246(0) )) | (\[43]  & \V247(0) )),
  \V2064(0)  = (V1844 & V2029) | ~\[508] ,
  \[45]  = (\[365]  & (\[277]  & (\[245]  & ~V505))) | ((\[365]  & (\[277]  & (\[245]  & V1646))) | ((\[245]  & (~V505 & ~\V59(0) )) | ((\[245]  & (V1646 & ~\V59(0) )) | (V695 | \V214(0) )))),
  \[46]  = \[407]  & \V293(0) ,
  \[47]  = (~V1735 & (V1445 & (~\V302(0)  & \V59(0) ))) | ((V745 & (~\V302(0)  & (~\V62(0)  & \V56(0) ))) | ((~\[253]  & (V1445 & ~\V302(0) )) | ((~V745 & (\V270(0)  & ~\V302(0) )) | (\V270(0)  & (~\V302(0)  & ~\V62(0) ))))),
  \[48]  = (~\V202(0)  & ~\V271(0) ) | ((~\V274(0)  & ~\V271(0) ) | (~\V269(0)  & \V271(0) )),
  \[120]  = \V9(0)  & \V1(0) ,
  \[49]  = (~\V202(0)  & \V274(0) ) | \V271(0) ,
  \[500]  = \[222]  | ~\V268(3) ,
  \[121]  = \[443]  & \V1(0) ,
  \[311]  = ~V721 | ~\[65] ,
  \[501]  = ~V1298 | ~V1850,
  \[122]  = \V1(0)  & \V11(0) ,
  \[502]  = V739 | V740,
  \[123]  = \V1(0)  & \V12(0) ,
  \[503]  = ~V2025 | ~V1846,
  \[124]  = (\[120]  & ~\V109(0) ) | (\[120]  & \V13(0) ),
  \[504]  = V1302 | V1298,
  \[125]  = \[252]  & \V66(0) ,
  \[505]  = \V60(0)  | \V56(0) ,
  \[126]  = (~V769 & (\V277(0)  & \V14(0) )) | V746,
  \[127]  = V1445 | ~\V14(0) ,
  \[50]  = ~\V257(7) ,
  \[317]  = (~\[444]  & ~V697) | ~\[160] ,
  \[507]  = V2025,
  \[128]  = (\[373]  & (~\V1455(0)  & (\V14(0)  & \V258(0) ))) | ((V1366 & (~\[219]  & (\V14(0)  & ~\V258(0) ))) | (\V1455(0)  & (\V14(0)  & ~\V258(0) ))),
  \[51]  = \[484]  & ~\V149(3) ,
  \[318]  = \[295]  | ~\V288(6) ,
  \[508]  = V1844 | V2029,
  \[129]  = (~\V1455(0)  & (\V259(0)  & \V14(0) )) | (\V1455(0)  & (~\V259(0)  & \V14(0) )),
  \[52]  = (~V799 & (\V759(0)  & (~\[65]  & (~\V291(0)  & (~\V292(0)  & (\V169(0)  & ~\V55(0) )))))) | (\[347]  & (~V799 & (~\V291(0)  & (~\V292(0)  & \V169(0) )))),
  \[319]  = \V260(0)  | (\V259(0)  | (~\V258(0)  | \V59(0) )),
  \[509]  = ~V454 | V446,
  \[53]  = \[537]  & (\[252]  & \V1674(0) ),
  \[54]  = \V9(0)  & \V5(0) ,
  \[55]  = \[443]  & \V6(0) ,
  \[56]  = \V6(0)  & \V9(0) ,
  \[57]  = (~\[448]  & (\V12(0)  & (\V6(0)  & ~\V174(0) ))) | (\V12(0)  & (\V6(0)  & \V52(0) )),
  \[58]  = \[443]  & \V7(0) ,
  \[130]  = (~\V1463(0)  & (\V260(0)  & \V14(0) )) | (\V1463(0)  & (~\V260(0)  & \V14(0) )),
  \[59]  = \V11(0)  & \V5(0) ,
  \V1451(0)  = \[128] ,
  \[320]  = 0,
  \[510]  = V2034,
  \[131]  = \[252]  & (~V737 & \V67(0) ),
  \[321]  = V768 | V687,
  \[511]  = ~V1318,
  \[132]  = (~V701 & \V15(0) ) | ((\[65]  & \V15(0) ) | V1476),
  \[512]  = (~\[253]  & ~V1445) | ~\[311] ,
  \[133]  = ~\V214(0) ,
  \[323]  = (\[539]  & ~V687) | ((V687 & \V730(0) ) | \V731(0) ),
  \[134]  = (~\V1999(0)  & (\V69(0)  & (\V14(0)  & \V215(0) ))) | ((~\V1999(0)  & (\V68(0)  & (\V14(0)  & \V215(0) ))) | ((~\V1999(0)  & (\V14(0)  & (\V70(0)  & \V215(0) ))) | ((~\[260]  & (~\V1999(0)  & \V14(0) )) | (\V216(0)  & ~\V214(0) )))),
  \[324]  = (~\[295]  & (~\[225]  & (~\V2084(0)  & (~\V2081(0)  & (V1842 & ~\V1255(2) ))))) | ((~\[295]  & (\[225]  & (~\V2084(0)  & (~\V2081(0)  & (~\V1255(2)  & \V288(4) ))))) | ((\[544]  & (~\[225]  & (\V2081(0)  & (V1842 & ~\V1255(2) )))) | ((\[544]  & (\[225]  & (\V2081(0)  & (~\V1255(2)  & \V288(4) )))) | ((~\[295]  & (~\[225]  & (\V2084(0)  & (V1842 & \V1255(2) )))) | ((~\[295]  & (\[225]  & (\V2084(0)  & (\V1255(2)  & \V288(4) )))) | V856))))),
  \[135]  = ~\V175(0) ,
  \V1863(0)  = \[185] ,
  \[325]  = (\[238]  & (~\[226]  & (~\V1357(0)  & (\V1354(0)  & (~\V1351(0)  & (V1846 & (~\V1255(2)  & ~\V1255(0) ))))))) | ((\[238]  & (~\[226]  & (~\V1357(0)  & (\V1354(0)  & (\V1351(0)  & (V1846 & (~\V1255(2)  & \V1255(0) ))))))) | ((\[238]  & (~\[226]  & (\V1357(0)  & (\V1354(0)  & (~\V1351(0)  & (V1846 & (\V1255(2)  & ~\V1255(0) ))))))) | ((\[238]  & (~\[226]  & (\V1357(0)  & (\V1354(0)  & (\V1351(0)  & (V1846 & (\V1255(2)  & \V1255(0) ))))))) | ((\[238]  & (\[226]  & (~\V1357(0)  & (\V1354(0)  & (~\V1351(0)  & (~\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((\[238]  & (\[226]  & (~\V1357(0)  & (\V1354(0)  & (\V1351(0)  & (~\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | ((\[238]  & (\[226]  & (\V1357(0)  & (\V1354(0)  & (~\V1351(0)  & (\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((\[238]  & (\[226]  & (\V1357(0)  & (\V1354(0)  & (\V1351(0)  & (\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (~\[226]  & (~\V1357(0)  & (~\V1354(0)  & (~\V1351(0)  & (V1846 & (~\V1255(2)  & ~\V1255(0) ))))))) | ((~\[232]  & (~\[226]  & (~\V1357(0)  & (~\V1354(0)  & (\V1351(0)  & (V1846 & (~\V1255(2)  & \V1255(0) ))))))) | ((~\[232]  & (~\[226]  & (\V1357(0)  & (~\V1354(0)  & (~\V1351(0)  & (V1846 & (\V1255(2)  & ~\V1255(0) ))))))) | ((~\[232]  & (~\[226]  & (\V1357(0)  & (~\V1354(0)  & (\V1351(0)  & (V1846 & (\V1255(2)  & \V1255(0) ))))))) | ((~\[232]  & (\[226]  & (~\V1357(0)  & (~\V1354(0)  & (~\V1351(0)  & (~\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (\[226]  & (~\V1357(0)  & (~\V1354(0)  & (\V1351(0)  & (~\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (\[226]  & (\V1357(0)  & (~\V1354(0)  & (~\V1351(0)  & (\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (\[226]  & (\V1357(0)  & (~\V1354(0)  & (\V1351(0)  & (\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | V896))))))))))))))),
  \V1679(0)  = \[152] ,
  \[136]  = (~V1535 & ~\V2002(0) ) | ((V1535 & V955) | ((V1535 & V954) | ((V1535 & V946) | ((V1535 & V936) | ((V1535 & V906) | ((V1535 & V896) | ((V1535 & V866) | (V1535 & V856)))))))),
  \[326]  = (\[238]  & (~\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~\V473(0)  & (\V470(0)  & (~\V467(0)  & \V288(0) ))))))) | ((\[238]  & (~\[224]  & (~\V1255(2)  & (\V1255(0)  & (~\V473(0)  & (\V470(0)  & (\V467(0)  & \V288(0) ))))))) | ((\[238]  & (~\[224]  & (\V1255(2)  & (~\V1255(0)  & (\V473(0)  & (\V470(0)  & (~\V467(0)  & \V288(0) ))))))) | ((\[238]  & (~\[224]  & (\V1255(2)  & (\V1255(0)  & (\V473(0)  & (\V470(0)  & (\V467(0)  & \V288(0) ))))))) | ((~\[232]  & (~\[224]  & (~\V1255(2)  & (~\V1255(0)  & (~\V473(0)  & (~\V470(0)  & (~\V467(0)  & \V288(0) ))))))) | ((~\[232]  & (~\[224]  & (~\V1255(2)  & (\V1255(0)  & (~\V473(0)  & (~\V470(0)  & (\V467(0)  & \V288(0) ))))))) | ((~\[232]  & (~\[224]  & (\V1255(2)  & (~\V1255(0)  & (\V473(0)  & (~\V470(0)  & (~\V467(0)  & \V288(0) ))))))) | ((~\[232]  & (~\[224]  & (\V1255(2)  & (\V1255(0)  & (\V473(0)  & (~\V470(0)  & (\V467(0)  & \V288(0) ))))))) | V946))))))),
  \[137]  = (\[437]  & V1535) | ((\[307]  & ~V1535) | \[527] ),
  \[60]  = \V11(0)  & \V7(0) ,
  \[327]  = \V62(0)  | \V56(0) ,
  \[138]  = (\[448]  & ~V1535) | ((\[438]  & V1535) | \[527] ),
  \[61]  = \V9(0)  & \V7(0) ,
  \[328]  = ~\V199(3)  | ~\V199(4) ,
  \[139]  = ~V1535,
  \[62]  = (\[99]  & ~\V71(0) ) | ((\[99]  & ~\V202(0) ) | (\[99]  & \V13(0) )),
  \[329]  = ~V1871 | ~\V194(4) ,
  \V445(0)  = V1302 & ~V441,
  \[63]  = (\[237]  & (\V812(0)  & ~\[163] )) | ((\[446]  & ~V1735) | ((~\[409]  & ~\V1681(0) ) | ((~V695 & \V290(0) ) | (\[408]  | (~\[267]  | (\V302(0)  | \V214(0) )))))),
  \[64]  = V799 & ~\V759(0) ,
  \[65]  = \V51(0)  | \V52(0) ,
  \[66]  = (~\[311]  & \V149(5) ) | (\[311]  & ~\V279(0) ),
  \[67]  = (\[311]  & (~\V280(0)  & ~\V279(0) )) | ((\[311]  & (\V280(0)  & \V279(0) )) | (~\[311]  & \V149(4) )),
  \[68]  = (\[465]  & (\[252]  & \V56(0) )) | ((\[409]  & (\[252]  & \[65] )) | ((\[252]  & (V799 & \V759(0) )) | (\[252]  & (\V1681(0)  & \[65] )))),
  \[140]  = \[252]  & \V68(0) ,
  \[69]  = (~\[465]  & (\[252]  & (V976 & \V56(0) ))) | ((\[464]  & (\[252]  & \V59(0) )) | (\[542]  & \V1681(0) )),
  \[330]  = ~V750 | ~\V56(0) ,
  \[141]  = (\[252]  & \V50(0) ) | (\[252]  & \V69(0) ),
  \[142]  = (~\[335]  & ~\V239(4) ) | (V379 & \[82] ),
  \[143]  = (~\[335]  & (~\V239(3)  & \V239(4) )) | ((~\[335]  & (\V239(3)  & ~\V239(4) )) | (V379 & \[83] )),
  \[333]  = ~V2106 & ~\V2019(0) ,
  \[523]  = (~V1445 & V769) | \[445] ,
  \[144]  = (~V1607 & ~V1606) | (V1607 & V1606),
  \[334]  = \[257]  & ~V1402,
  \V1829(7)  = \[175] ,
  \[145]  = (~V1609 & ~V1608) | (V1609 & V1608),
  \[335]  = ~V721 | \[65] ,
  \V1829(6)  = \[176] ,
  \[146]  = (\V2002(0)  & \V174(0) ) | ((V695 & \V174(0) ) | ((\V292(0)  & ~\V302(0) ) | V799)),
  \V1829(9)  = \[173] ,
  \[147]  = (\[277]  & (~V741 & ~\V294(0) )) | ((V739 & (\V91(1)  & \V62(0) )) | ((V739 & (\V91(0)  & \V59(0) )) | ~\[407] )),
  \[70]  = (\[345]  & \V257(6) ) | ((\[334]  & \V32(4) ) | ((\[300]  & \V32(1) ) | ((\[272]  & \V189(5) ) | ((\[271]  & \V229(5) ) | (\[270]  & \V32(11) ))))),
  \[337]  = \V473(0)  | V437,
  \[527]  = (\[326]  & V1535) | ((\[309]  & V1535) | \V2002(0) ),
  \V1829(8)  = \[174] ,
  \[148]  = (V701 & (\[65]  & \V149(7) )) | (V1644 | V1643),
  \[71]  = (\[345]  & \V257(5) ) | ((\[334]  & \V32(3) ) | ((\[300]  & \V32(0) ) | ((\[272]  & \V189(4) ) | ((\[271]  & \V229(4) ) | (\[270]  & \V32(10) ))))),
  \[338]  = \V1337(0)  | V1298,
  \[149]  = (\V1647(0)  & V1445) | (\V1681(0)  | (~\V295(0)  | (\V290(0)  | (\V249(0)  | \V289(0) )))),
  \[72]  = (\[345]  & \V257(4) ) | ((\[272]  & \V189(3) ) | ((\[271]  & \V229(3) ) | ((\[270]  & \V32(9) ) | ((\[257]  & \V32(2) ) | \[300] )))),
  \[339]  = \V2064(0)  | V2025,
  \[73]  = (\[345]  & \V257(3) ) | ((\[272]  & \V189(2) ) | ((\[271]  & \V229(2) ) | ((\[270]  & \V32(8) ) | ((\[257]  & \V32(1) ) | \[300] )))),
  \V1417(0)  = (~V726 & (~V727 & (~\V1681(0)  & (\V53(0)  & ~\V56(0) )))) | ((\[539]  & (~V411 & \V57(0) )) | ((\[539]  & (~V411 & \V53(0) )) | ((\[539]  & (~V411 & \V56(0) )) | ((~\[505]  & (\[361]  & \V57(0) )) | ((~\[505]  & (\[361]  & \V53(0) )) | ((\[523]  & \V57(0) ) | ((\[523]  & \V53(0) ) | ((\[523]  & \V56(0) ) | ((~\[263]  & \V57(0) ) | ((~\[263]  & \V53(0) ) | ((~\[263]  & \V56(0) ) | V745))))))))))),
  \[74]  = (\[345]  & \V257(2) ) | ((\[272]  & \V189(1) ) | ((\[271]  & \V229(1) ) | ((\[270]  & \V32(7) ) | ((\[257]  & \V32(0) ) | \[300] )))),
  \[75]  = (\[345]  & \V257(1) ) | ((\[272]  & \V189(0) ) | ((\[271]  & \V229(0) ) | ((\[270]  & \V32(6) ) | \[300] ))),
  \V1771(1)  = \[169] ,
  \V1620(0)  = \[146] ,
  \[76]  = (\[345]  & \V257(0) ) | ((\[272]  & \V183(5) ) | ((\[271]  & \V223(5) ) | ((\[270]  & \V32(5) ) | \[334] ))),
  \V1771(0)  = \[170] ,
  \[77]  = (\[345]  & \V257(6) ) | ((\[272]  & \V183(4) ) | ((\[271]  & \V223(4) ) | (\[270]  & \V32(4) ))),
  \V1829(1)  = \[181] ,
  \V1829(0)  = \[182] ,
  \[150]  = (~\[351]  & (\[340]  & (\[279]  & (~\V1653(0)  & ~\[163] )))) | ((\[340]  & (\[279]  & (\V1653(0)  & \V812(0) ))) | ((\[340]  & (\[279]  & (\V1653(0)  & \V2002(0) ))) | ((\[340]  & (\[279]  & (\V812(0)  & ~\[163] ))) | ((\[340]  & (\[279]  & (\V2002(0)  & ~\[163] ))) | ((\[279]  & (~\[267]  & ~\[163] )) | (\[279]  & \V289(0) )))))),
  \[340]  = \[237]  | \[65] ,
  \V1829(3)  = \[179] ,
  \V1455(0)  = (V1366 & (\V268(0)  & \V258(0) )) | (~\[373]  & ~\V258(0) ),
  \[151]  = ~\V205(0) ,
  \[341]  = \[318]  | ~\V1255(3) ,
  \V1829(2)  = \[180] ,
  \[152]  = (\[319]  & (\V262(0)  & \V14(0) )) | \V1674(0) ,
  \[342]  = (~\[321]  & ~V738) | (\[321]  & \V59(0) ),
  \V1829(5)  = \[177] ,
  \[153]  = (\[396]  & (\[349]  & (~V1644 & ~V747))) | ((\[401]  & \V100(0) ) | (\[348]  & V1978)),
  \V1999(0)  = (\[342]  & (V1646 & ~V701)) | ((V738 & (V1646 & \V62(0) )) | (\[536]  | \V214(0) )),
  \[343]  = V745 | (\V274(0)  | ~\V271(0) ),
  \V1829(4)  = \[178] ,
  \[154]  = (\[401]  & \V100(5) ) | (V1978 & \V165(7) ),
  \V1900(0)  = \[191] ,
  \[155]  = (\[401]  & \V100(4) ) | (V1978 & \V165(6) ),
  \[345]  = \[235]  & (~\V1421(0)  & \V1681(0) ),
  \[156]  = (\[401]  & \V100(3) ) | (V1978 & \V165(5) ),
  \[536]  = \V172(0)  & (\V67(0)  & \V215(0) ),
  \[157]  = (\[401]  & \V100(2) ) | (V1978 & \V165(4) ),
  \[347]  = V725 | V700,
  \[537]  = \[52]  & \V70(0) ,
  \[158]  = (\[401]  & \V100(1) ) | (V1978 & \V165(3) ),
  \[348]  = (\[543]  & (~\V165(3)  & (~\V165(7)  & ~\V165(6) ))) | V1646,
  \[538]  = ~\V15(0)  & \V16(0) ,
  \[159]  = (~\[446]  & (~V721 & \[160] )) | ((~\[446]  & (\[160]  & \V280(0) )) | \[512] ),
  \[82]  = (\[300]  & \V32(11) ) | ((\[272]  & \V199(4) ) | ((\[271]  & \V239(4) ) | (\[270]  & \V88(1) ))),
  \[349]  = V702 | V700,
  \[539]  = ~\V730(0)  & \[51] ,
  \[83]  = (\[300]  & \V32(10) ) | ((\[272]  & \V199(3) ) | ((\[271]  & \V239(3) ) | (\[270]  & \V88(0) ))),
  \[84]  = (\[300]  & \V32(9) ) | ((\[272]  & \V199(2) ) | ((\[271]  & \V239(2) ) | (\[270]  & \V84(5) ))),
  \[85]  = (\[334]  & \V32(11) ) | ((\[300]  & \V32(8) ) | ((\[272]  & \V199(1) ) | ((\[271]  & \V239(1) ) | (\[270]  & \V84(4) )))),
  \[86]  = (\[334]  & \V32(10) ) | ((\[300]  & \V32(7) ) | ((\[272]  & \V199(0) ) | ((\[271]  & \V239(0) ) | (\[270]  & \V84(3) )))),
  \[87]  = (\[334]  & \V32(9) ) | ((\[300]  & \V32(6) ) | ((\[272]  & \V194(4) ) | ((\[271]  & \V234(4) ) | (\[270]  & \V84(2) )))),
  \[88]  = (\[478]  & \V149(7) ) | ((\[334]  & \V32(8) ) | ((\[300]  & \V32(5) ) | ((\[272]  & \V194(3) ) | ((\[271]  & \V234(3) ) | (\[270]  & \V84(1) ))))),
  \V336(0)  = (~V452 & (~V446 & (~V451 & (\V32(3)  & (\V32(2)  & ~\V32(0) ))))) | ((~V452 & (~V446 & (V451 & (\V32(3)  & (\V32(2)  & \V32(0) ))))) | ((~V452 & (~V451 & (\V32(3)  & (\V32(2)  & (\V32(1)  & ~\V32(0) ))))) | ((~V452 & (V451 & (\V32(3)  & (\V32(2)  & (\V32(1)  & \V32(0) ))))) | ((~\[414]  & (~V446 & (~V451 & (\V32(3)  & ~\V32(0) )))) | ((~\[414]  & (~V446 & (V451 & (\V32(3)  & \V32(0) )))) | ((~\[414]  & (~V451 & (\V32(3)  & (\V32(1)  & ~\V32(0) )))) | ((~\[414]  & (V451 & (\V32(3)  & (\V32(1)  & \V32(0) )))) | ((~V441 & (~V446 & (~V451 & (\V32(2)  & ~\V32(0) )))) | ((~V441 & (~V446 & (V451 & (\V32(2)  & \V32(0) )))) | ((~V441 & (~V451 & (\V32(2)  & (\V32(1)  & ~\V32(0) )))) | ((~V441 & (V451 & (\V32(2)  & (\V32(1)  & \V32(0) )))) | ((~V446 & (~V451 & (\V32(1)  & ~\V32(0) ))) | ((~V446 & (V451 & (\V32(1)  & \V32(0) ))) | (~V451 & \V32(0) )))))))))))))),
  \[160]  = ~V695 & (\V240(0)  & ~\V172(0) ),
  \V487(0)  = (\[430]  & (\V467(0)  & ~V1850)) | (V1850 & V451),
  \V1306(0)  = V2029 & ~V1302,
  \[89]  = (\[478]  & \V149(6) ) | ((\[334]  & \V32(7) ) | ((\[300]  & \V32(4) ) | ((\[272]  & \V194(2) ) | ((\[271]  & \V234(2) ) | (\[270]  & \V84(0) ))))),
  \[350]  = V452 | ~V437,
  \[540]  = \[367]  & ~\V149(7) ,
  \[161]  = (~\[415]  & (\V242(0)  & \V14(0) )) | (~\[285]  & (V1535 & \V1647(0) )),
  \[351]  = \[258]  | V739,
  \[541]  = \[368]  & \V149(7) ,
  \[162]  = ~\[340]  & (V1735 & (~\V290(0)  & ~\V289(0) )),
  \[542]  = \[252]  & \V62(0) ,
  \[163]  = (\[396]  & (\[342]  & ~V701)) | ((V738 & (V1646 & \V62(0) )) | \[546] ),
  \[353]  = \[294]  | V742,
  \[543]  = ~\V165(5)  & ~\V165(4) ,
  \[164]  = V747 | (V725 | (~\V33(0)  | ~\V289(0) )),
  \[354]  = \[309]  | \V1681(0) ,
  \[544]  = \[238]  & ~\V1255(0) ,
  \[355]  = (\[323]  & \V59(0) ) | ~\[244] ,
  \[545]  = \[366]  & ~\V149(7) ,
  \[166]  = \[538]  | ~\[388] ,
  \[356]  = \[327]  | \V50(0) ,
  \[546]  = V695 & \V290(0) ,
  \V1921(1)  = \[197] ,
  \V1495(0)  = \[135] ,
  V2014 = ~\[343]  & (\[285]  & (V1445 & (\V134(0)  & \V134(1) ))),
  \[167]  = (\[412]  & (\V101(0)  & \V14(0) )) | (\[538]  & \[347] ),
  \[90]  = (\[478]  & \V149(5) ) | ((\[334]  & \V32(6) ) | ((\[300]  & \V32(3) ) | ((\[272]  & \V194(1) ) | ((\[271]  & \V234(1) ) | (\[270]  & \V78(5) ))))),
  \[547]  = \[479]  & \V149(1) ,
  \V1921(0)  = \[198] ,
  V2025 = (~\[417]  & V1842) | (\[417]  & ~V1842),
  V2027 = (~\[375]  & ~V1844) | (\[375]  & V1844),
  V2028 = (~\[418]  & \[282] ) | (\[418]  & ~\[282] ),
  \[168]  = ~\V101(0) ,
  V2029 = (~V2027 & (V1842 & ~V2025)) | (V2027 & ~V1842),
  \[91]  = (\[478]  & \V149(4) ) | ((\[345]  & \V257(7) ) | ((\[334]  & \V32(5) ) | ((\[300]  & \V32(2) ) | ((\[272]  & \V194(0) ) | ((\[271]  & \V234(0) ) | (\[270]  & \V78(4) )))))),
  \V1921(3)  = \[195] ,
  \V393(0)  = \[6] ,
  V2034 = (~V2028 & \V2033(0) ) | (V2028 & ~\V2033(0) ),
  \[169]  = (~V745 & ~\V134(1) ) | (V745 & ~\V88(3) ),
  V2039 = ~\[418]  & V2034,
  \[92]  = \[443]  & \V2(0) ,
  \[359]  = V742,
  \V1921(2)  = \[196] ,
  V2045 = (~\[507]  & ~V2034) | (\[507]  & V2034),
  V2047 = ~\[510]  | V2039,
  \[93]  = (~\[445]  & (~V745 & (~V769 & (~V710 & (~\[51]  & (\V57(0)  & (\V2(0)  & (\V12(0)  & (~\V174(0)  & ~\V35(0) ))))))))) | ((~V745 & (~V739 & (~\V57(0)  & (\V2(0)  & (\V12(0)  & (~\V174(0)  & ~\V35(0) )))))) | (V745 & (~\V63(0)  & (~\V60(0)  & (\V2(0)  & (\V12(0)  & (~\V174(0)  & ~\V35(0) ))))))),
  \V1921(5)  = \[193] ,
  \[94]  = \V9(0)  & \V2(0) ,
  \V1921(4)  = \[194] ,
  \[95]  = \V9(0)  & \V3(0) ,
  \[96]  = \V11(0)  & \V3(0) ,
  \[97]  = \[96]  & ~\V62(0) ,
  \[98]  = \[443]  & \V4(0) ,
  \[170]  = (~V745 & ~\V134(0) ) | (V745 & ~\V88(2) ),
  \[99]  = \V9(0)  & \V4(0) ,
  \V1459(0)  = \[129] ,
  \[171]  = (~V745 & ~\[70] ) | (V745 & ~\V78(3) ),
  \[361]  = V710 | V411,
  \[172]  = (~V745 & ~\[71] ) | (V745 & ~\V78(2) ),
  \[362]  = ~V1646 | ~V701,
  \[173]  = (~\[91]  & ~\V37(0) ) | (~\[82]  & \V37(0) ),
  \[174]  = (~\[83]  & \V37(0) ) | (~\[70]  & ~\V37(0) ),
  \[364]  = V1735 | ~\V261(0) ,
  \[175]  = (~\[84]  & \V37(0) ) | (~\[71]  & ~\V37(0) ),
  \[365]  = ~V710 | ~V687,
  V2106 = ~\[65]  | ~V769,
  \[176]  = (~\[85]  & \V37(0) ) | (~\[72]  & ~\V37(0) ),
  V2109 = ~\[65]  | ~V727,
  \[366]  = \[306]  & ~\V149(6) ,
  \V802(0)  = \[65] ,
  \V1681(0)  = \V262(0)  | \V1674(0) ,
  \[177]  = (~\[86]  & \V37(0) ) | (~\[73]  & ~\V37(0) ),
  \[367]  = ~\V149(4)  & ~\V149(5) ,
  V2122 = V1445 | (~V727 | \V59(0) ),
  \[178]  = (~\[87]  & \V37(0) ) | (~\[74]  & ~\V37(0) ),
  \[368]  = \[306]  & \V149(6) ,
  \[179]  = (~\[88]  & \V37(0) ) | (~\[75]  & ~\V37(0) ),
  \[369]  = (~\[295]  & (~\[225]  & (~\V2064(0)  & (~\V2061(0)  & (~\V1255(2)  & \V288(4) ))))) | ((\[544]  & (~\[225]  & (\V2061(0)  & (~\V2058(0)  & ~\V1255(2) )))) | ((~\[295]  & (~\[225]  & (\V2064(0)  & (\V1255(2)  & \V288(4) )))) | V866)),
  \V821(0)  = \[66] ,
  \V1758(0)  = \[166] ,
  \[180]  = (~\[89]  & \V37(0) ) | (~\[76]  & ~\V37(0) ),
  \[370]  = (\[238]  & (~\[226]  & (~\V1337(0)  & (\V1334(0)  & (~\V1331(0)  & (~\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((\[238]  & (~\[226]  & (~\V1337(0)  & (\V1334(0)  & (\V1331(0)  & (~\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | ((\[238]  & (~\[226]  & (\V1337(0)  & (\V1334(0)  & (~\V1331(0)  & (\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((\[238]  & (~\[226]  & (\V1337(0)  & (\V1334(0)  & (\V1331(0)  & (\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (~\[226]  & (~\V1337(0)  & (~\V1334(0)  & (~\V1331(0)  & (~\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (~\[226]  & (~\V1337(0)  & (~\V1334(0)  & (\V1331(0)  & (~\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (~\[226]  & (\V1337(0)  & (~\V1334(0)  & (~\V1331(0)  & (\V1255(2)  & (~\V1255(0)  & \V288(2) ))))))) | ((~\[232]  & (~\[226]  & (\V1337(0)  & (~\V1334(0)  & (\V1331(0)  & (\V1255(2)  & (\V1255(0)  & \V288(2) ))))))) | V906))))))),
  \V1645(0)  = \[148] ,
  \[181]  = (~\[90]  & \V37(0) ) | (~\[77]  & ~\V37(0) ),
  \[371]  = \V149(2)  | \V149(1) ,
  \[182]  = (~\V1255(2)  & \V37(0) ) | (~\[91]  & ~\V37(0) ),
  \[372]  = ~\[263]  | V721,
  \[183]  = (~\[356]  & (\V261(0)  & \V14(0) )) | ((\[319]  & (\V261(0)  & \V14(0) )) | ((V1366 & (\V268(0)  & \V14(0) )) | (~\V262(0)  & (\V261(0)  & \V14(0) )))),
  \[373]  = ~\[356]  | ~\V1681(0) ,
  \[184]  = ~\V261(0) ,
  \[374]  = ~\V149(4)  | ~\V149(5) ,
  \[185]  = ~\V301(0) ,
  \[375]  = (~\V288(7)  & \V288(6) ) | ~\[417] ,
  \[186]  = ~\V302(0) ,
  \[187]  = (\[330]  & \V108(0) ) | ((\V15(0)  & \V16(0) ) | V1476),
  \[188]  = (\[330]  & \V108(1) ) | (V769 & V1476);
endmodule

