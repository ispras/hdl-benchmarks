module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 ;
output g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 ;
wire t_0 , t_1 , t_2 , t_3 ;
buf ( n1  , g0 );
buf ( n2  , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9  , g8 );
buf ( n10  , g9 );
buf ( n11  , g10 );
buf ( n12  , g11 );
buf ( n13  , g12 );
buf ( n14  , g13 );
buf ( n15  , g14 );
buf ( n16  , g15 );
buf ( n17  , g16 );
buf ( n18  , g17 );
buf ( n19  , g18 );
buf ( n20  , g19 );
buf ( n21  , g20 );
buf ( n22  , g21 );
buf ( n23  , g22 );
buf ( n24  , g23 );
buf ( n25  , g24 );
buf ( n26  , g25 );
buf ( n27  , g26 );
buf ( n28  , g27 );
buf ( n29  , g28 );
buf ( n30  , g29 );
buf ( n31  , g30 );
buf ( n32  , g31 );
buf ( n33  , g32 );
buf ( n34  , g33 );
buf ( n35  , g34 );
buf ( n36  , g35 );
buf ( n37  , g36 );
buf ( n38  , g37 );
buf ( n39  , g38 );
buf ( n40  , g39 );
buf ( n41  , g40 );
buf ( n42  , g41 );
buf ( n43  , g42 );
buf ( n44  , g43 );
buf ( n45  , g44 );
buf ( n46  , g45 );
buf ( n47  , g46 );
buf ( n48  , g47 );
buf ( n49  , g48 );
buf ( n50  , g49 );
buf ( n51  , g50 );
buf ( n52  , g51 );
buf ( n53  , g52 );
buf ( n54  , g53 );
buf ( n55  , g54 );
buf ( n56  , g55 );
buf ( n57  , g56 );
buf ( n58  , g57 );
buf ( n59  , g58 );
buf ( n60  , g59 );
buf ( n61  , g60 );
buf ( n62  , g61 );
buf ( n63  , g62 );
buf ( n64  , g63 );
buf ( n65  , g64 );
buf ( n66  , g65 );
buf ( n67  , g66 );
buf ( n68  , g67 );
buf ( n69  , g68 );
buf ( n70  , g69 );
buf ( n71  , g70 );
buf ( n72  , g71 );
buf ( n73  , g72 );
buf ( n74  , g73 );
buf ( n75  , g74 );
buf ( n76  , g75 );
buf ( n77  , g76 );
buf ( n78  , g77 );
buf ( n79  , g78 );
buf ( n80  , g79 );
buf ( n81  , g80 );
buf ( n82  , g81 );
buf ( n83  , g82 );
buf ( n84  , g83 );
buf ( n85  , g84 );
buf ( n86  , g85 );
buf ( n87  , g86 );
buf ( n88  , g87 );
buf ( n89  , g88 );
buf ( n90  , g89 );
buf ( n91  , g90 );
buf ( n92  , g91 );
buf ( n93  , g92 );
buf ( n94  , g93 );
buf ( n95  , g94 );
buf ( n96  , g95 );
buf ( n97  , g96 );
buf ( n98  , g97 );
buf ( n99  , g98 );
buf ( n100  , g99 );
buf ( n101  , g100 );
buf ( n102  , g101 );
buf ( n103  , g102 );
buf ( n104  , g103 );
buf ( n105  , g104 );
buf ( n106  , g105 );
buf ( n107  , g106 );
buf ( n108  , g107 );
buf ( n109  , g108 );
buf ( n110  , g109 );
buf ( n111  , g110 );
buf ( n112  , g111 );
buf ( n113  , g112 );
buf ( n114  , g113 );
buf ( n115  , g114 );
buf ( n116  , g115 );
buf ( n117  , g116 );
buf ( n118  , g117 );
buf ( n119  , g118 );
buf ( n120  , g119 );
buf ( n121  , g120 );
buf ( n122  , g121 );
buf ( n123  , g122 );
buf ( n124  , g123 );
buf ( n125  , g124 );
buf ( n126  , g125 );
buf ( n127  , g126 );
buf ( n128  , g127 );
buf ( n129  , g128 );
buf ( n130  , g129 );
buf ( n131  , g130 );
buf ( n132  , g131 );
buf ( n133  , g132 );
buf ( n134  , g133 );
buf ( n135  , g134 );
buf ( n136  , g135 );
buf ( n137  , g136 );
buf ( n138  , g137 );
buf ( n139  , g138 );
buf ( n140  , g139 );
buf ( n141  , g140 );
buf ( n142  , g141 );
buf ( n143  , g142 );
buf ( n144  , g143 );
buf ( n145  , g144 );
buf ( n146  , g145 );
buf ( n147  , g146 );
buf ( n148  , g147 );
buf ( n149  , g148 );
buf ( n150  , g149 );
buf ( n151  , g150 );
buf ( n152  , g151 );
buf ( n153  , g152 );
buf ( n154  , g153 );
buf ( n155  , g154 );
buf ( n156  , g155 );
buf ( n157  , g156 );
buf ( n158  , g157 );
buf ( n159  , g158 );
buf ( n160  , g159 );
buf ( n161  , g160 );
buf ( n162  , g161 );
buf ( n163  , g162 );
buf ( n164  , g163 );
buf ( n165  , g164 );
buf ( n166  , g165 );
buf ( n167  , g166 );
buf ( n168  , g167 );
buf ( n169  , g168 );
buf ( n170  , g169 );
buf ( n171  , g170 );
buf ( n172  , g171 );
buf ( n173  , g172 );
buf ( n174  , g173 );
buf ( n175  , g174 );
buf ( n176  , g175 );
buf ( n177  , g176 );
buf ( n178  , g177 );
buf ( n179  , g178 );
buf ( n180  , g179 );
buf ( n181  , g180 );
buf ( n182  , g181 );
buf ( n183  , g182 );
buf ( n184  , g183 );
buf ( n185  , g184 );
buf ( n186  , g185 );
buf ( n187  , g186 );
buf ( n188  , g187 );
buf ( n189  , g188 );
buf ( n190  , g189 );
buf ( n191  , g190 );
buf ( n192  , g191 );
buf ( n193  , g192 );
buf ( n194  , g193 );
buf ( n195  , g194 );
buf ( n196  , g195 );
buf ( n197  , g196 );
buf ( n198  , g197 );
buf ( n199  , g198 );
buf ( n200  , g199 );
buf ( n201  , g200 );
buf ( n202  , g201 );
buf ( n203  , g202 );
buf ( n204  , g203 );
buf ( n205  , g204 );
buf ( n206  , g205 );
buf ( n207  , g206 );
buf ( n208  , g207 );
buf ( n209  , g208 );
buf ( n210  , g209 );
buf ( n211  , g210 );
buf ( n212  , g211 );
buf ( n213  , g212 );
buf ( n214  , g213 );
buf ( n215  , g214 );
buf ( n216  , g215 );
buf ( n217  , g216 );
buf ( n218  , g217 );
buf ( n219  , g218 );
buf ( n220  , g219 );
buf ( n221  , g220 );
buf ( n222  , g221 );
buf ( n223  , g222 );
buf ( n224  , g223 );
buf ( n225  , g224 );
buf ( n226  , g225 );
buf ( n227  , g226 );
buf ( n228  , g227 );
buf ( n229  , g228 );
buf ( n230  , g229 );
buf ( n231  , g230 );
buf ( n232  , g231 );
buf ( n233  , g232 );
buf ( n234  , g233 );
buf ( n235  , g234 );
buf ( n236  , g235 );
buf ( n237  , g236 );
buf ( n238  , g237 );
buf ( n239  , g238 );
buf ( n240  , g239 );
buf ( n241  , g240 );
buf ( n242  , g241 );
buf ( n243  , g242 );
buf ( n244  , g243 );
buf ( n245  , g244 );
buf ( n246  , g245 );
buf ( n247  , g246 );
buf ( n248  , g247 );
buf ( n249  , g248 );
buf ( n250  , g249 );
buf ( n251  , g250 );
buf ( n252  , g251 );
buf ( n253  , g252 );
buf ( n254  , g253 );
buf ( n255  , g254 );
buf ( n256  , g255 );
buf ( g256 , n257  );
buf ( g257 , n258  );
buf ( g258 , n259  );
buf ( g259 , n260  );
buf ( g260 , n261  );
buf ( g261 , n262  );
buf ( g262 , n263  );
buf ( g263 , n264  );
buf ( g264 , n265  );
buf ( g265 , n266  );
buf ( g266 , n267  );
buf ( g267 , n268  );
buf ( g268 , n269  );
buf ( g269 , n270  );
buf ( g270 , n271  );
buf ( g271 , n272  );
buf ( g272 , n273  );
buf ( g273 , n274  );
buf ( g274 , n275  );
buf ( g275 , n276  );
buf ( g276 , n277  );
buf ( g277 , n278  );
buf ( g278 , n279  );
buf ( g279 , n280  );
buf ( g280 , n281  );
buf ( g281 , n282  );
buf ( g282 , n283  );
buf ( g283 , n284  );
buf ( g284 , n285  );
buf ( g285 , n286  );
buf ( g286 , n287  );
buf ( g287 , n288  );
buf ( g288 , n289  );
buf ( g289 , n290  );
buf ( g290 , n291  );
buf ( g291 , n292  );
buf ( g292 , n293  );
buf ( g293 , n294  );
buf ( g294 , n295  );
buf ( g295 , n296  );
buf ( g296 , n297  );
buf ( g297 , n298  );
buf ( g298 , n299  );
buf ( g299 , n300  );
buf ( g300 , n301  );
buf ( g301 , n302  );
buf ( g302 , n303  );
buf ( g303 , n304  );
buf ( g304 , n305  );
buf ( g305 , n306  );
buf ( g306 , n307  );
buf ( g307 , n308  );
buf ( g308 , n309  );
buf ( g309 , n310  );
buf ( g310 , n311  );
buf ( g311 , n312  );
buf ( g312 , n313  );
buf ( g313 , n314  );
buf ( g314 , n315  );
buf ( g315 , n316  );
buf ( g316 , n317  );
buf ( g317 , n318  );
buf ( g318 , n319  );
buf ( g319 , n320  );
buf ( g320 , n321  );
buf ( g321 , n322  );
buf ( g322 , n323  );
buf ( g323 , n324  );
buf ( g324 , n325  );
buf ( g325 , n326  );
buf ( g326 , n327  );
buf ( g327 , n328  );
buf ( g328 , n329  );
buf ( g329 , n330  );
buf ( g330 , n331  );
buf ( g331 , n332  );
buf ( g332 , n333  );
buf ( g333 , n334  );
buf ( g334 , n335  );
buf ( g335 , n336  );
buf ( g336 , n337  );
buf ( g337 , n338  );
buf ( g338 , n339  );
buf ( g339 , n340  );
buf ( g340 , n341  );
buf ( g341 , n342  );
buf ( g342 , n343  );
buf ( g343 , n344  );
buf ( g344 , n345  );
buf ( g345 , n346  );
buf ( g346 , n347  );
buf ( g347 , n348  );
buf ( g348 , n349  );
buf ( g349 , n350  );
buf ( g350 , n351  );
buf ( g351 , n352  );
buf ( g352 , n353  );
buf ( g353 , n354  );
buf ( g354 , n355  );
buf ( g355 , n356  );
buf ( g356 , n357  );
buf ( g357 , n358  );
buf ( g358 , n359  );
buf ( g359 , n360  );
buf ( g360 , n361  );
buf ( g361 , n362  );
buf ( g362 , n363  );
buf ( g363 , n364  );
buf ( g364 , n365  );
buf ( g365 , n366  );
buf ( g366 , n367  );
buf ( g367 , n368  );
buf ( g368 , n369  );
buf ( g369 , n370  );
buf ( g370 , n371  );
buf ( g371 , n372  );
buf ( g372 , n373  );
buf ( g373 , n374  );
buf ( g374 , n375  );
buf ( g375 , n376  );
buf ( g376 , n377  );
buf ( g377 , n378  );
buf ( g378 , n379  );
buf ( g379 , n380  );
buf ( g380 , n381  );
buf ( g381 , n382  );
buf ( g382 , n383  );
buf ( g383 , n384  );
buf ( g384 , n385  );
buf ( g385 , n386  );
buf ( g386 , n387  );
buf ( g387 , n388  );
buf ( g388 , n389  );
buf ( g389 , n390  );
buf ( g390 , n391  );
buf ( g391 , n392  );
buf ( g392 , n393  );
buf ( g393 , n394  );
buf ( g394 , n395  );
buf ( g395 , n396  );
buf ( g396 , n397  );
buf ( g397 , n398  );
buf ( g398 , n399  );
buf ( g399 , n400  );
buf ( g400 , n401  );
buf ( g401 , n402  );
buf ( g402 , n403  );
buf ( g403 , n404  );
buf ( g404 , n405  );
buf ( g405 , n406  );
buf ( g406 , n407  );
buf ( g407 , n408  );
buf ( g408 , n409  );
buf ( g409 , n410  );
buf ( g410 , n411  );
buf ( g411 , n412  );
buf ( g412 , n413  );
buf ( g413 , n414  );
buf ( g414 , n415  );
buf ( g415 , n416  );
buf ( g416 , n417  );
buf ( g417 , n418  );
buf ( g418 , n419  );
buf ( g419 , n420  );
buf ( g420 , n421  );
buf ( g421 , n422  );
buf ( g422 , n423  );
buf ( g423 , n424  );
buf ( g424 , n425  );
buf ( g425 , n426  );
buf ( g426 , n427  );
buf ( g427 , n428  );
buf ( g428 , n429  );
buf ( g429 , n430  );
buf ( g430 , n431  );
buf ( g431 , n432  );
buf ( g432 , n433  );
buf ( g433 , n434  );
buf ( g434 , n435  );
buf ( g435 , n436  );
buf ( g436 , n437  );
buf ( g437 , n438  );
buf ( g438 , n439  );
buf ( g439 , n440  );
buf ( g440 , n441  );
buf ( g441 , n442  );
buf ( g442 , n443  );
buf ( g443 , n444  );
buf ( g444 , n445  );
buf ( g445 , n446  );
buf ( g446 , n447  );
buf ( g447 , n448  );
buf ( g448 , n449  );
buf ( g449 , n450  );
buf ( g450 , n451  );
buf ( g451 , n452  );
buf ( g452 , n453  );
buf ( g453 , n454  );
buf ( g454 , n455  );
buf ( g455 , n456  );
buf ( g456 , n457  );
buf ( g457 , n458  );
buf ( g458 , n459  );
buf ( g459 , n460  );
buf ( g460 , n461  );
buf ( g461 , n462  );
buf ( g462 , n463  );
buf ( g463 , n464  );
buf ( g464 , n465  );
buf ( g465 , n466  );
buf ( g466 , n467  );
buf ( g467 , n468  );
buf ( g468 , n469  );
buf ( g469 , n470  );
buf ( g470 , n471  );
buf ( g471 , n472  );
buf ( g472 , n473  );
buf ( g473 , n474  );
buf ( g474 , n475  );
buf ( g475 , n476  );
buf ( g476 , n477  );
buf ( g477 , n478  );
buf ( g478 , n479  );
buf ( g479 , n480  );
buf ( g480 , n481  );
buf ( g481 , n482  );
buf ( g482 , n483  );
buf ( g483 , n484  );
buf ( g484 , n485  );
buf ( g485 , n486  );
buf ( g486 , n487  );
buf ( g487 , n488  );
buf ( g488 , n489  );
buf ( g489 , n490  );
buf ( g490 , n491  );
buf ( g491 , n492  );
buf ( g492 , n493  );
buf ( g493 , n494  );
buf ( g494 , n495  );
buf ( g495 , n496  );
buf ( g496 , n497  );
buf ( g497 , n498  );
buf ( g498 , n499  );
buf ( g499 , n500  );
buf ( g500 , n501  );
buf ( n257 , n5542 );
buf ( n258 , n5352 );
buf ( n259 , n5527 );
buf ( n260 , n5532 );
buf ( n261 , n5507 );
buf ( n262 , n5512 );
buf ( n263 , n5517 );
buf ( n264 , n5522 );
buf ( n265 , n5497 );
buf ( n266 , n5502 );
buf ( n267 , n5347 );
buf ( n268 , n5567 );
buf ( n269 , n5342 );
buf ( n270 , n5492 );
buf ( n271 , n5482 );
buf ( n272 , n5472 );
buf ( n273 , n5487 );
buf ( n274 , n5477 );
buf ( n275 , n5602 );
buf ( n276 , n5572 );
buf ( n277 , n5332 );
buf ( n278 , n5462 );
buf ( n279 , n5467 );
buf ( n280 , n5437 );
buf ( n281 , n5326 );
buf ( n282 , n5457 );
buf ( n283 , n5562 );
buf ( n284 , n5337 );
buf ( n285 , n5447 );
buf ( n286 , n5452 );
buf ( n287 , n5432 );
buf ( n288 , n5442 );
buf ( n289 , n5547 );
buf ( n290 , n5382 );
buf ( n291 , n5552 );
buf ( n292 , n5387 );
buf ( n293 , n5417 );
buf ( n294 , n5422 );
buf ( n295 , n5557 );
buf ( n296 , n5427 );
buf ( n297 , n5537 );
buf ( n298 , n5372 );
buf ( n299 , n5367 );
buf ( n300 , n5597 );
buf ( n301 , n5357 );
buf ( n302 , n5582 );
buf ( n303 , n5412 );
buf ( n304 , n5407 );
buf ( n305 , n5587 );
buf ( n306 , n5577 );
buf ( n307 , n5392 );
buf ( n308 , n5402 );
buf ( n309 , n5362 );
buf ( n310 , n5592 );
buf ( n311 , n5397 );
buf ( n312 , n5377 );
buf ( n313 , n2315 );
buf ( n314 , n4969 );
buf ( n315 , n942 );
buf ( n316 , n4974 );
buf ( n317 , n1678 );
buf ( n318 , n4995 );
buf ( n319 , n2827 );
buf ( n320 , n4964 );
buf ( n321 , n3631 );
buf ( n322 , n5051 );
buf ( n323 , n1551 );
buf ( n324 , n5070 );
buf ( n325 , n2511 );
buf ( n326 , n5248 );
buf ( n327 , n1610 );
buf ( n328 , n5083 );
buf ( n329 , n2559 );
buf ( n330 , n5212 );
buf ( n331 , n3279 );
buf ( n332 , n4952 );
buf ( n333 , n3340 );
buf ( n334 , n5206 );
buf ( n335 , n3678 );
buf ( n336 , n5094 );
buf ( n337 , n1136 );
buf ( n338 , n5268 );
buf ( n339 , n3389 );
buf ( n340 , n4980 );
buf ( n341 , n1471 );
buf ( n342 , n5230 );
buf ( n343 , n3444 );
buf ( n344 , n5218 );
buf ( n345 , n3500 );
buf ( n346 , n4990 );
buf ( n347 , n721 );
buf ( n348 , n5140 );
buf ( n349 , n2605 );
buf ( n350 , n5044 );
buf ( n351 , n1279 );
buf ( n352 , n5037 );
buf ( n353 , n1878 );
buf ( n354 , n5013 );
buf ( n355 , n2658 );
buf ( n356 , n5284 );
buf ( n357 , n3059 );
buf ( n358 , n5224 );
buf ( n359 , n2983 );
buf ( n360 , n5237 );
buf ( n361 , n1998 );
buf ( n362 , n5100 );
buf ( n363 , n2699 );
buf ( n364 , n4958 );
buf ( n365 , n1204 );
buf ( n366 , n5060 );
buf ( n367 , n1939 );
buf ( n368 , n5302 );
buf ( n369 , n2751 );
buf ( n370 , n5314 );
buf ( n371 , n2111 );
buf ( n372 , n5106 );
buf ( n373 , n2914 );
buf ( n374 , n5007 );
buf ( n375 , n3552 );
buf ( n376 , n5255 );
buf ( n377 , n2837 );
buf ( n378 , n1986 );
buf ( n379 , n2014 );
buf ( n380 , n3557 );
buf ( n381 , n1210 );
buf ( n382 , n2843 );
buf ( n383 , n3683 );
buf ( n384 , n2848 );
buf ( n385 , n2853 );
buf ( n386 , n2832 );
buf ( n387 , n2919 );
buf ( n388 , n727 );
buf ( n389 , n3562 );
buf ( n390 , n3567 );
buf ( n391 , n2003 );
buf ( n392 , n1216 );
buf ( n393 , n2924 );
buf ( n394 , n1222 );
buf ( n395 , n3572 );
buf ( n396 , n2929 );
buf ( n397 , n2009 );
buf ( n398 , n3577 );
buf ( n399 , n2935 );
buf ( n400 , n1991 );
buf ( n401 , n3582 );
buf ( n402 , n2020 );
buf ( n403 , n3587 );
buf ( n404 , n2026 );
buf ( n405 , n3592 );
buf ( n406 , n3688 );
buf ( n407 , n2031 );
buf ( n408 , n2940 );
buf ( n409 , n5017 );
buf ( n410 , n5130 );
buf ( n411 , n5076 );
buf ( n412 , n4946 );
buf ( n413 , n5134 );
buf ( n414 , n5088 );
buf ( n415 , n5200 );
buf ( n416 , n5143 );
buf ( n417 , n5110 );
buf ( n418 , n5278 );
buf ( n419 , n5150 );
buf ( n420 , n5154 );
buf ( n421 , n5241 );
buf ( n422 , n5160 );
buf ( n423 , n5167 );
buf ( n424 , n5272 );
buf ( n425 , n5064 );
buf ( n426 , n5290 );
buf ( n427 , n5262 );
buf ( n428 , n5171 );
buf ( n429 , n4999 );
buf ( n430 , n5308 );
buf ( n431 , n5177 );
buf ( n432 , n5025 );
buf ( n433 , n5021 );
buf ( n434 , n5296 );
buf ( n435 , n5183 );
buf ( n436 , n5318 );
buf ( n437 , n4984 );
buf ( n438 , n5190 );
buf ( n439 , n5125 );
buf ( n440 , n5321 );
buf ( n441 , n5054 );
buf ( n442 , n5029 );
buf ( n443 , n5195 );
buf ( n444 , n5249 );
buf ( n445 , n4030 );
buf ( n446 , n4054 );
buf ( n447 , n3745 );
buf ( n448 , n4076 );
buf ( n449 , n4099 );
buf ( n450 , n4121 );
buf ( n451 , n4142 );
buf ( n452 , n4161 );
buf ( n453 , n4182 );
buf ( n454 , n4202 );
buf ( n455 , n4223 );
buf ( n456 , n3804 );
buf ( n457 , n4245 );
buf ( n458 , n4265 );
buf ( n459 , n4286 );
buf ( n460 , n3933 );
buf ( n461 , n4308 );
buf ( n462 , n4328 );
buf ( n463 , n4347 );
buf ( n464 , n3860 );
buf ( n465 , n4367 );
buf ( n466 , n4388 );
buf ( n467 , n3776 );
buf ( n468 , n4938 );
buf ( n469 , n4408 );
buf ( n470 , n4428 );
buf ( n471 , n4446 );
buf ( n472 , n3885 );
buf ( n473 , n4469 );
buf ( n474 , n4492 );
buf ( n475 , n4515 );
buf ( n476 , n3980 );
buf ( n477 , n4535 );
buf ( n478 , n4556 );
buf ( n479 , n4577 );
buf ( n480 , n4004 );
buf ( n481 , n4598 );
buf ( n482 , n4619 );
buf ( n483 , n4640 );
buf ( n484 , n4659 );
buf ( n485 , n4681 );
buf ( n486 , n4701 );
buf ( n487 , n4722 );
buf ( n488 , n3834 );
buf ( n489 , n4743 );
buf ( n490 , n4763 );
buf ( n491 , n4784 );
buf ( n492 , n3955 );
buf ( n493 , n4805 );
buf ( n494 , n4825 );
buf ( n495 , n4846 );
buf ( n496 , n3911 );
buf ( n497 , n4865 );
buf ( n498 , n4884 );
buf ( n499 , n4902 );
buf ( n500 , n4920 );
buf ( n501 , n5117 );
and ( n504 , n196 , n197 , n198 , n199 );
buf ( n505 , n504 );
not ( n506 , n505 );
buf ( n507 , n506 );
buf ( n508 , n507 );
not ( n509 , n199 );
and ( n510 , n102 , n509 );
and ( n511 , n94 , n199 );
nor ( n512 , n510 , n511 );
and ( n513 , n508 , n512 );
not ( n514 , n508 );
and ( n515 , n135 , n242 );
not ( n516 , n135 );
not ( n517 , n242 );
and ( n518 , n516 , n517 );
or ( n519 , n515 , n518 );
buf ( n520 , n519 );
not ( n521 , n520 );
not ( n522 , n521 );
not ( n523 , n522 );
xor ( n524 , n134 , n234 );
buf ( n525 , n524 );
buf ( n526 , n525 );
not ( n527 , n526 );
not ( n528 , n527 );
xor ( n529 , n136 , n238 );
not ( n530 , n529 );
not ( n531 , n530 );
xor ( n532 , n132 , n255 );
not ( n533 , n532 );
not ( n534 , n533 );
xor ( n535 , n163 , n252 );
buf ( n536 , n535 );
not ( n537 , n536 );
xor ( n538 , n133 , n248 );
nand ( n539 , n537 , n538 );
not ( n540 , n538 );
nand ( n541 , n536 , n540 );
nand ( n542 , n539 , n541 );
nand ( n543 , n534 , n542 );
and ( n544 , n531 , n543 );
not ( n545 , n531 );
not ( n546 , n532 );
nand ( n547 , n546 , n536 );
not ( n548 , n547 );
xor ( n549 , n133 , n248 );
not ( n550 , n549 );
nand ( n551 , n548 , n550 );
and ( n552 , n545 , n551 );
nor ( n553 , n544 , n552 );
not ( n554 , n553 );
or ( n555 , n528 , n554 );
not ( n556 , n529 );
not ( n557 , n556 );
not ( n558 , n557 );
and ( n559 , n134 , n234 );
not ( n560 , n134 );
not ( n561 , n234 );
and ( n562 , n560 , n561 );
nor ( n563 , n559 , n562 );
nand ( n564 , n563 , n532 );
nor ( n565 , n539 , n564 );
nand ( n566 , n558 , n565 );
nand ( n567 , n555 , n566 );
not ( n568 , n567 );
or ( n569 , n523 , n568 );
nor ( n570 , n535 , n532 );
and ( n571 , n538 , n570 );
not ( n572 , n571 );
not ( n573 , n524 );
not ( n574 , n573 );
nor ( n575 , n572 , n574 );
nand ( n576 , n558 , n521 , n575 );
nand ( n577 , n569 , n576 );
not ( n578 , n577 );
not ( n579 , n529 );
buf ( n580 , n579 );
buf ( n581 , n519 );
not ( n582 , n581 );
not ( n583 , n524 );
not ( n584 , n535 );
nand ( n585 , n584 , n532 );
nor ( n586 , n549 , n585 );
nand ( n587 , n583 , n586 );
not ( n588 , n587 );
nand ( n589 , n580 , n582 , n588 );
not ( n590 , n589 );
buf ( n591 , n520 );
not ( n592 , n591 );
buf ( n593 , n524 );
not ( n594 , n549 );
buf ( n595 , n570 );
and ( n596 , n593 , n594 , n595 );
not ( n597 , n596 );
not ( n598 , n579 );
nor ( n599 , n597 , n598 );
nand ( n600 , n592 , n599 );
not ( n601 , n600 );
nor ( n602 , n590 , n601 );
not ( n603 , n585 );
nand ( n604 , n549 , n603 );
not ( n605 , n604 );
nor ( n606 , n573 , n519 );
nand ( n607 , n605 , n579 , n606 );
not ( n608 , n520 );
not ( n609 , n608 );
not ( n610 , n530 );
not ( n611 , n593 );
nand ( n612 , n535 , n532 );
nor ( n613 , n538 , n612 );
nand ( n614 , n611 , n613 );
nor ( n615 , n610 , n614 );
nand ( n616 , n609 , n615 );
and ( n617 , n607 , n616 );
nand ( n618 , n579 , n520 , n525 , n586 );
not ( n619 , n582 );
not ( n620 , n579 );
nand ( n621 , n574 , n571 );
nor ( n622 , n620 , n621 );
nand ( n623 , n619 , n622 );
not ( n624 , n593 );
and ( n625 , n556 , n624 , n594 , n595 );
nand ( n626 , n619 , n625 );
and ( n627 , n618 , n623 , n626 );
nand ( n628 , n578 , n602 , n617 , n627 );
not ( n629 , n521 );
not ( n630 , n612 );
nand ( n631 , n549 , n630 );
not ( n632 , n631 );
nand ( n633 , n557 , n574 , n632 );
nor ( n634 , n629 , n633 );
not ( n635 , n634 );
not ( n636 , n579 );
not ( n637 , n613 );
nor ( n638 , n611 , n637 );
nand ( n639 , n636 , n638 );
not ( n640 , n639 );
not ( n641 , n629 );
nand ( n642 , n640 , n641 );
not ( n643 , n550 );
not ( n644 , n547 );
nand ( n645 , n557 , n583 , n643 , n644 );
not ( n646 , n645 );
nand ( n647 , n641 , n646 );
not ( n648 , n558 );
nor ( n649 , n551 , n583 );
nand ( n650 , n592 , n648 , n649 );
nand ( n651 , n635 , n642 , n647 , n650 );
nor ( n652 , n628 , n651 );
and ( n653 , n557 , n574 , n586 );
nand ( n654 , n641 , n653 );
not ( n655 , n520 );
buf ( n656 , n531 );
and ( n657 , n655 , n656 , n596 );
not ( n658 , n657 );
nand ( n659 , n654 , n658 );
nor ( n660 , n525 , n604 );
nand ( n661 , n656 , n655 , n660 );
not ( n662 , n661 );
nor ( n663 , n659 , n662 );
not ( n664 , n551 );
not ( n665 , n520 );
not ( n666 , n525 );
nand ( n667 , n664 , n610 , n665 , n666 );
nand ( n668 , n581 , n636 , n526 , n632 );
and ( n669 , n667 , n668 );
not ( n670 , n669 );
buf ( n671 , n521 );
nand ( n672 , n656 , n596 );
nor ( n673 , n671 , n672 );
not ( n674 , n631 );
nand ( n675 , n674 , n636 , n581 , n666 );
buf ( n676 , n608 );
buf ( n677 , n530 );
nor ( n678 , n621 , n677 );
nand ( n679 , n676 , n678 );
nand ( n680 , n675 , n679 );
nor ( n681 , n670 , n673 , n680 );
nand ( n682 , n663 , n681 );
and ( n683 , n676 , n615 );
not ( n684 , n676 );
not ( n685 , n594 );
nand ( n686 , n644 , n685 , n525 );
nor ( n687 , n686 , n620 );
and ( n688 , n684 , n687 );
nor ( n689 , n683 , n688 );
nand ( n690 , n644 , n643 , n583 );
nor ( n691 , n690 , n598 );
nand ( n692 , n522 , n691 );
not ( n693 , n692 );
nor ( n694 , n677 , n587 );
nand ( n695 , n609 , n694 );
not ( n696 , n695 );
nor ( n697 , n693 , n696 );
and ( n698 , n530 , n593 , n613 );
not ( n699 , n698 );
nor ( n700 , n582 , n699 );
not ( n701 , n700 );
not ( n702 , n591 );
nand ( n703 , n702 , n687 );
nand ( n704 , n701 , n703 );
and ( n705 , n666 , n632 );
nand ( n706 , n580 , n582 , n705 );
nand ( n707 , n550 , n595 );
nor ( n708 , n525 , n707 );
nand ( n709 , n620 , n581 , n708 );
nand ( n710 , n706 , n709 );
nor ( n711 , n704 , n710 );
nand ( n712 , n689 , n697 , n711 );
nor ( n713 , n682 , n712 );
nand ( n714 , n652 , n713 );
not ( n715 , n175 );
and ( n716 , n714 , n715 );
not ( n717 , n714 );
and ( n718 , n717 , n175 );
nor ( n719 , n716 , n718 );
and ( n720 , n514 , n719 );
nor ( n721 , n513 , n720 );
not ( n722 , n508 );
not ( n723 , n47 );
and ( n724 , n722 , n723 );
not ( n725 , n722 );
and ( n726 , n725 , n719 );
nor ( n727 , n724 , n726 );
not ( n728 , n163 );
and ( n729 , n211 , n728 );
not ( n730 , n211 );
and ( n731 , n730 , n163 );
or ( n732 , n729 , n731 );
not ( n733 , n732 );
not ( n734 , n733 );
not ( n735 , n734 );
xor ( n736 , n161 , n204 );
not ( n737 , n736 );
not ( n738 , n737 );
not ( n739 , n738 );
not ( n740 , n739 );
not ( n741 , n159 );
nand ( n742 , n741 , n223 );
not ( n743 , n223 );
nand ( n744 , n743 , n159 );
nand ( n745 , n742 , n744 );
not ( n746 , n160 );
nand ( n747 , n746 , n227 );
not ( n748 , n227 );
nand ( n749 , n748 , n160 );
nand ( n750 , n747 , n749 );
nand ( n751 , n745 , n750 );
not ( n752 , n751 );
nand ( n753 , n740 , n752 );
xnor ( n754 , n132 , n214 );
not ( n755 , n754 );
not ( n756 , n755 );
not ( n757 , n756 );
xor ( n758 , n162 , n217 );
buf ( n759 , n758 );
not ( n760 , n759 );
not ( n761 , n760 );
or ( n762 , n753 , n757 , n761 );
nor ( n763 , n745 , n758 );
not ( n764 , n763 );
nand ( n765 , n758 , n745 );
nand ( n766 , n764 , n765 );
buf ( n767 , n750 );
not ( n768 , n767 );
not ( n769 , n754 );
not ( n770 , n769 );
not ( n771 , n770 );
and ( n772 , n766 , n768 , n771 );
not ( n773 , n758 );
not ( n774 , n773 );
buf ( n775 , n754 );
xor ( n776 , n160 , n227 );
xor ( n777 , n159 , n223 );
not ( n778 , n777 );
nand ( n779 , n776 , n778 );
not ( n780 , n779 );
nand ( n781 , n775 , n780 );
nor ( n782 , n774 , n781 );
nor ( n783 , n772 , n782 );
or ( n784 , n783 , n740 );
nand ( n785 , n762 , n784 );
nand ( n786 , n735 , n785 );
not ( n787 , n755 );
buf ( n788 , n758 );
nor ( n789 , n779 , n736 );
and ( n790 , n787 , n788 , n789 );
nand ( n791 , n733 , n790 );
not ( n792 , n791 );
not ( n793 , n732 );
not ( n794 , n793 );
not ( n795 , n794 );
buf ( n796 , n755 );
not ( n797 , n796 );
not ( n798 , n758 );
not ( n799 , n736 );
nor ( n800 , n777 , n776 );
nand ( n801 , n799 , n800 );
nor ( n802 , n798 , n801 );
not ( n803 , n802 );
nor ( n804 , n797 , n803 );
nand ( n805 , n795 , n804 );
not ( n806 , n805 );
nor ( n807 , n792 , n806 );
not ( n808 , n776 );
nand ( n809 , n808 , n737 , n745 );
not ( n810 , n809 );
not ( n811 , n758 );
nand ( n812 , n810 , n811 );
buf ( n813 , n775 );
nor ( n814 , n812 , n813 );
not ( n815 , n732 );
not ( n816 , n815 );
nand ( n817 , n814 , n816 );
not ( n818 , n817 );
not ( n819 , n733 );
not ( n820 , n788 );
nand ( n821 , n777 , n776 );
nor ( n822 , n738 , n821 );
nand ( n823 , n820 , n822 );
nor ( n824 , n771 , n823 );
nand ( n825 , n819 , n824 );
not ( n826 , n769 );
not ( n827 , n788 );
not ( n828 , n776 );
and ( n829 , n738 , n745 , n828 );
and ( n830 , n826 , n827 , n829 );
nand ( n831 , n816 , n830 );
nand ( n832 , n825 , n831 );
not ( n833 , n775 );
not ( n834 , n799 );
nor ( n835 , n777 , n776 );
and ( n836 , n833 , n811 , n834 , n835 );
nand ( n837 , n795 , n836 );
not ( n838 , n837 );
nor ( n839 , n818 , n832 , n838 );
and ( n840 , n786 , n807 , n839 );
not ( n841 , n755 );
and ( n842 , n841 , n798 , n834 , n835 );
not ( n843 , n842 );
nor ( n844 , n735 , n843 );
not ( n845 , n815 );
not ( n846 , n759 );
nand ( n847 , n834 , n780 );
nor ( n848 , n846 , n847 );
nand ( n849 , n797 , n845 , n848 );
not ( n850 , n732 );
buf ( n851 , n850 );
not ( n852 , n801 );
nand ( n853 , n852 , n826 , n827 );
not ( n854 , n853 );
nand ( n855 , n851 , n854 );
nand ( n856 , n849 , n855 );
nor ( n857 , n844 , n856 );
not ( n858 , n826 );
not ( n859 , n850 );
nor ( n860 , n774 , n847 );
nand ( n861 , n858 , n859 , n860 );
not ( n862 , n801 );
not ( n863 , n756 );
nand ( n864 , n862 , n863 , n794 , n760 );
nand ( n865 , n861 , n864 );
not ( n866 , n865 );
not ( n867 , n851 );
not ( n868 , n830 );
or ( n869 , n867 , n868 );
nand ( n870 , n851 , n824 );
nand ( n871 , n869 , n870 );
not ( n872 , n871 );
nor ( n873 , n813 , n823 );
nand ( n874 , n851 , n873 );
buf ( n875 , n788 );
nand ( n876 , n875 , n789 );
nor ( n877 , n813 , n876 );
nand ( n878 , n795 , n877 );
and ( n879 , n874 , n878 );
not ( n880 , n821 );
nand ( n881 , n880 , n834 , n788 , n755 );
not ( n882 , n881 );
nand ( n883 , n882 , n859 );
not ( n884 , n883 );
not ( n885 , n881 );
nand ( n886 , n733 , n885 );
not ( n887 , n886 );
nor ( n888 , n884 , n887 );
nand ( n889 , n866 , n872 , n879 , n888 );
not ( n890 , n809 );
nand ( n891 , n890 , n846 , n796 , n793 );
not ( n892 , n891 );
and ( n893 , n770 , n774 , n829 );
nand ( n894 , n851 , n893 );
and ( n895 , n770 , n759 , n810 );
nand ( n896 , n851 , n895 );
nand ( n897 , n894 , n896 );
nor ( n898 , n892 , n897 );
not ( n899 , n863 );
not ( n900 , n899 );
buf ( n901 , n732 );
not ( n902 , n822 );
nor ( n903 , n827 , n902 );
and ( n904 , n901 , n903 );
not ( n905 , n904 );
or ( n906 , n900 , n905 );
not ( n907 , n901 );
nand ( n908 , n907 , n842 );
nand ( n909 , n906 , n908 );
not ( n910 , n909 );
not ( n911 , n738 );
nor ( n912 , n788 , n911 , n821 );
nand ( n913 , n858 , n845 , n912 );
and ( n914 , n759 , n829 );
nand ( n915 , n914 , n845 , n858 );
nand ( n916 , n913 , n915 );
nand ( n917 , n797 , n794 , n860 );
not ( n918 , n789 );
nor ( n919 , n875 , n918 );
nand ( n920 , n757 , n901 , n919 );
nand ( n921 , n917 , n920 );
not ( n922 , n835 );
nor ( n923 , n922 , n798 , n739 );
nand ( n924 , n863 , n901 , n923 );
nand ( n925 , n813 , n901 , n802 );
nand ( n926 , n924 , n925 );
nor ( n927 , n916 , n921 , n926 );
nand ( n928 , n898 , n910 , n927 );
nor ( n929 , n889 , n928 );
nand ( n930 , n840 , n857 , n929 );
not ( n931 , n179 );
and ( n932 , n930 , n931 );
not ( n933 , n930 );
and ( n934 , n933 , n179 );
nor ( n935 , n932 , n934 );
buf ( n936 , n507 );
buf ( n937 , n936 );
or ( n938 , n935 , n937 );
buf ( n939 , n507 );
nand ( n940 , n70 , n939 );
or ( n941 , n199 , n940 );
nand ( n942 , n938 , n941 );
and ( n943 , n92 , n509 );
and ( n944 , n84 , n199 );
nor ( n945 , n943 , n944 );
and ( n946 , n939 , n945 );
not ( n947 , n939 );
xor ( n948 , n155 , n218 );
buf ( n949 , n948 );
buf ( n950 , n949 );
xor ( n951 , n156 , n207 );
buf ( n952 , n951 );
not ( n953 , n952 );
not ( n954 , n953 );
not ( n955 , n954 );
xor ( n956 , n160 , n225 );
not ( n957 , n956 );
buf ( n958 , n957 );
not ( n959 , n958 );
xor ( n960 , n159 , n200 );
not ( n961 , n960 );
not ( n962 , n961 );
xor ( n963 , n157 , n222 );
not ( n964 , n963 );
xor ( n965 , n158 , n213 );
nor ( n966 , n964 , n965 );
nand ( n967 , n962 , n966 );
not ( n968 , n967 );
nand ( n969 , n959 , n968 );
nor ( n970 , n955 , n969 );
nand ( n971 , n950 , n970 );
not ( n972 , n949 );
not ( n973 , n972 );
not ( n974 , n952 );
not ( n975 , n974 );
not ( n976 , n956 );
not ( n977 , n976 );
not ( n978 , n963 );
nand ( n979 , n978 , n965 );
nor ( n980 , n962 , n979 );
nand ( n981 , n977 , n980 );
not ( n982 , n981 );
nand ( n983 , n973 , n975 , n982 );
not ( n984 , n952 );
not ( n985 , n984 );
nor ( n986 , n985 , n969 );
nand ( n987 , n950 , n986 );
not ( n988 , n972 );
buf ( n989 , n960 );
nor ( n990 , n965 , n963 );
nand ( n991 , n989 , n990 );
nor ( n992 , n958 , n991 );
and ( n993 , n988 , n985 , n992 );
not ( n994 , n993 );
nand ( n995 , n971 , n983 , n987 , n994 );
not ( n996 , n995 );
not ( n997 , n990 );
not ( n998 , n997 );
buf ( n999 , n952 );
not ( n1000 , n999 );
not ( n1001 , n958 );
buf ( n1002 , n961 );
not ( n1003 , n1002 );
nand ( n1004 , n998 , n1000 , n1001 , n1003 );
not ( n1005 , n949 );
not ( n1006 , n1005 );
or ( n1007 , n1004 , n1006 );
nor ( n1008 , n951 , n948 );
not ( n1009 , n1008 );
not ( n1010 , n1009 );
not ( n1011 , n978 );
and ( n1012 , n1011 , n965 , n961 );
nand ( n1013 , n1001 , n1010 , n1012 );
nand ( n1014 , n1007 , n1013 );
not ( n1015 , n1014 );
not ( n1016 , n966 );
not ( n1017 , n951 );
nand ( n1018 , n948 , n1017 , n957 );
or ( n1019 , n1016 , n1018 );
not ( n1020 , n1019 );
not ( n1021 , n953 );
nand ( n1022 , n1011 , n956 );
xnor ( n1023 , n155 , n218 );
nor ( n1024 , n1022 , n1023 );
not ( n1025 , n1024 );
or ( n1026 , n1021 , n1025 );
not ( n1027 , n1011 );
not ( n1028 , n957 );
or ( n1029 , n1027 , n1028 );
not ( n1030 , n963 );
nand ( n1031 , n956 , n1030 );
nand ( n1032 , n1029 , n1031 );
nand ( n1033 , n1023 , n952 , n1032 );
nand ( n1034 , n1026 , n1033 );
nand ( n1035 , n965 , n1034 );
not ( n1036 , n1035 );
or ( n1037 , n1020 , n1036 );
nand ( n1038 , n1037 , n1002 );
nand ( n1039 , n1015 , n1038 );
buf ( n1040 , n1023 );
buf ( n1041 , n1040 );
nor ( n1042 , n1016 , n989 );
nand ( n1043 , n959 , n1042 );
nor ( n1044 , n1043 , n985 );
nand ( n1045 , n1041 , n1044 );
not ( n1046 , n984 );
not ( n1047 , n960 );
nand ( n1048 , n1047 , n990 );
nor ( n1049 , n958 , n1048 );
nand ( n1050 , n1046 , n1040 , n1049 );
nand ( n1051 , n1045 , n1050 );
nor ( n1052 , n1039 , n1051 );
nand ( n1053 , n950 , n955 , n1049 );
not ( n1054 , n1053 );
and ( n1055 , n960 , n965 , n963 );
and ( n1056 , n999 , n959 , n1055 );
not ( n1057 , n1056 );
nor ( n1058 , n950 , n1057 );
nor ( n1059 , n1054 , n1058 );
nand ( n1060 , n1041 , n970 );
nand ( n1061 , n1041 , n986 );
and ( n1062 , n1060 , n1061 );
nand ( n1063 , n996 , n1052 , n1059 , n1062 );
and ( n1064 , n958 , n1012 );
nand ( n1065 , n1064 , n985 , n988 );
not ( n1066 , n976 );
nor ( n1067 , n1048 , n1066 );
nand ( n1068 , n973 , n975 , n1067 );
nand ( n1069 , n1065 , n1068 );
buf ( n1070 , n1023 );
nand ( n1071 , n958 , n1055 );
nor ( n1072 , n954 , n1071 );
and ( n1073 , n1070 , n1072 );
not ( n1074 , n1070 );
not ( n1075 , n999 );
nor ( n1076 , n977 , n991 );
nand ( n1077 , n1075 , n1076 );
not ( n1078 , n1077 );
and ( n1079 , n1074 , n1078 );
nor ( n1080 , n1073 , n1079 );
not ( n1081 , n952 );
nor ( n1082 , n1081 , n1071 );
nand ( n1083 , n988 , n1082 );
nor ( n1084 , n979 , n1047 );
nand ( n1085 , n958 , n1084 );
nor ( n1086 , n954 , n1085 );
nand ( n1087 , n973 , n1086 );
and ( n1088 , n1083 , n1087 );
nand ( n1089 , n999 , n958 , n1042 );
nor ( n1090 , n1070 , n1089 );
not ( n1091 , n1090 );
not ( n1092 , n979 );
buf ( n1093 , n976 );
nand ( n1094 , n1092 , n1081 , n1093 , n1002 );
not ( n1095 , n1094 );
nand ( n1096 , n950 , n1095 );
nand ( n1097 , n1080 , n1088 , n1091 , n1096 );
nor ( n1098 , n1069 , n1097 );
not ( n1099 , n1075 );
nand ( n1100 , n1070 , n1099 , n1076 );
not ( n1101 , n1100 );
not ( n1102 , n1070 );
not ( n1103 , n1086 );
or ( n1104 , n1102 , n1103 );
nand ( n1105 , n952 , n976 );
nor ( n1106 , n1105 , n967 );
nand ( n1107 , n1040 , n1106 );
nand ( n1108 , n1104 , n1107 );
nor ( n1109 , n1101 , n1108 );
not ( n1110 , n1005 );
not ( n1111 , n954 );
not ( n1112 , n1055 );
nor ( n1113 , n1093 , n1112 );
nand ( n1114 , n1110 , n1111 , n1113 );
not ( n1115 , n1114 );
not ( n1116 , n1084 );
nor ( n1117 , n1116 , n1093 );
nand ( n1118 , n975 , n1117 );
nor ( n1119 , n1041 , n1118 );
nor ( n1120 , n1115 , n1119 );
nor ( n1121 , n950 , n1094 );
not ( n1122 , n1121 );
nor ( n1123 , n950 , n1089 );
nand ( n1124 , n974 , n1067 );
nor ( n1125 , n1110 , n1124 );
nor ( n1126 , n1123 , n1125 );
and ( n1127 , n1109 , n1120 , n1122 , n1126 );
nand ( n1128 , n1098 , n1127 );
nor ( n1129 , n1063 , n1128 );
not ( n1130 , n1129 );
not ( n1131 , n168 );
and ( n1132 , n1130 , n1131 );
and ( n1133 , n168 , n1129 );
nor ( n1134 , n1132 , n1133 );
and ( n1135 , n947 , n1134 );
nor ( n1136 , n946 , n1135 );
and ( n1137 , n120 , n509 );
and ( n1138 , n112 , n199 );
nor ( n1139 , n1137 , n1138 );
and ( n1140 , n508 , n1139 );
not ( n1141 , n508 );
not ( n1142 , n524 );
nand ( n1143 , n1142 , n533 );
nor ( n1144 , n541 , n1143 );
nor ( n1145 , n565 , n1144 );
or ( n1146 , n1145 , n677 );
nor ( n1147 , n529 , n538 );
nor ( n1148 , n563 , n536 );
nand ( n1149 , n1147 , n534 , n1148 );
nand ( n1150 , n1146 , n1149 );
nand ( n1151 , n1150 , n609 );
not ( n1152 , n1151 );
nor ( n1153 , n1152 , n634 );
nand ( n1154 , n526 , n580 , n582 , n632 );
nand ( n1155 , n619 , n599 );
nand ( n1156 , n1153 , n1154 , n1155 );
nand ( n1157 , n618 , n623 );
nor ( n1158 , n1156 , n1157 );
nand ( n1159 , n522 , n687 );
nand ( n1160 , n592 , n625 );
nand ( n1161 , n607 , n1160 );
not ( n1162 , n581 );
nand ( n1163 , n1162 , n579 , n660 );
nand ( n1164 , n649 , n591 , n580 );
nand ( n1165 , n1163 , n1164 );
not ( n1166 , n700 );
nand ( n1167 , n1166 , n576 );
nor ( n1168 , n1161 , n1165 , n1167 );
and ( n1169 , n1158 , n1159 , n616 , n1168 );
nand ( n1170 , n521 , n698 );
and ( n1171 , n1170 , n709 );
not ( n1172 , n582 );
nand ( n1173 , n1172 , n678 );
and ( n1174 , n1173 , n695 );
not ( n1175 , n706 );
nand ( n1176 , n656 , n655 , n575 );
not ( n1177 , n1176 );
nor ( n1178 , n1175 , n1177 );
not ( n1179 , n629 );
nand ( n1180 , n1179 , n691 );
nand ( n1181 , n702 , n694 );
and ( n1182 , n1180 , n1181 );
nand ( n1183 , n1171 , n1174 , n1178 , n1182 );
not ( n1184 , n686 );
nand ( n1185 , n648 , n676 , n1184 );
nand ( n1186 , n1185 , n654 , n658 );
nand ( n1187 , n650 , n667 );
not ( n1188 , n1187 );
not ( n1189 , n639 );
nand ( n1190 , n1189 , n1172 );
not ( n1191 , n591 );
nor ( n1192 , n1191 , n645 );
not ( n1193 , n675 );
nor ( n1194 , n1192 , n1193 );
nand ( n1195 , n1188 , n1190 , n1194 );
nor ( n1196 , n1183 , n1186 , n1195 );
nand ( n1197 , n1169 , n1196 );
not ( n1198 , n181 );
and ( n1199 , n1197 , n1198 );
not ( n1200 , n1197 );
and ( n1201 , n1200 , n181 );
nor ( n1202 , n1199 , n1201 );
and ( n1203 , n1141 , n1202 );
nor ( n1204 , n1140 , n1203 );
not ( n1205 , n507 );
not ( n1206 , n37 );
and ( n1207 , n1205 , n1206 );
not ( n1208 , n1205 );
and ( n1209 , n1208 , n1134 );
nor ( n1210 , n1207 , n1209 );
not ( n1211 , n936 );
not ( n1212 , n15 );
and ( n1213 , n1211 , n1212 );
not ( n1214 , n1211 );
and ( n1215 , n1214 , n935 );
nor ( n1216 , n1213 , n1215 );
not ( n1217 , n939 );
not ( n1218 , n65 );
and ( n1219 , n1217 , n1218 );
not ( n1220 , n1217 );
and ( n1221 , n1220 , n1202 );
nor ( n1222 , n1219 , n1221 );
buf ( n1223 , n507 );
and ( n1224 , n106 , n509 );
and ( n1225 , n98 , n199 );
nor ( n1226 , n1224 , n1225 );
and ( n1227 , n1223 , n1226 );
not ( n1228 , n1223 );
not ( n1229 , n614 );
nand ( n1230 , n598 , n655 , n1229 );
nand ( n1231 , n635 , n647 , n1230 , n667 );
nand ( n1232 , n671 , n622 );
not ( n1233 , n1232 );
not ( n1234 , n1160 );
nor ( n1235 , n1233 , n1234 );
nor ( n1236 , n573 , n556 );
not ( n1237 , n1236 );
and ( n1238 , n519 , n547 );
not ( n1239 , n519 );
and ( n1240 , n1239 , n585 );
nor ( n1241 , n1238 , n1240 );
not ( n1242 , n1241 );
or ( n1243 , n1237 , n1242 );
nor ( n1244 , n524 , n529 );
not ( n1245 , n595 );
not ( n1246 , n630 );
nand ( n1247 , n1245 , n1246 );
nand ( n1248 , n1244 , n581 , n1247 );
nand ( n1249 , n1243 , n1248 );
nand ( n1250 , n643 , n1249 );
and ( n1251 , n616 , n589 , n1163 , n1250 );
nand ( n1252 , n627 , n1235 , n1251 );
nor ( n1253 , n1231 , n1252 );
not ( n1254 , n1192 );
nand ( n1255 , n1190 , n1254 );
nand ( n1256 , n1172 , n653 );
nand ( n1257 , n1256 , n1173 );
not ( n1258 , n668 );
not ( n1259 , n1258 );
and ( n1260 , n661 , n1176 );
nand ( n1261 , n1259 , n1260 , n658 );
nor ( n1262 , n1255 , n1257 , n1261 );
nor ( n1263 , n551 , n526 );
nand ( n1264 , n671 , n558 , n1263 );
nand ( n1265 , n706 , n1264 );
not ( n1266 , n1170 );
not ( n1267 , n703 );
nor ( n1268 , n1266 , n1267 );
nor ( n1269 , n696 , n673 );
nand ( n1270 , n1268 , n1269 , n692 , n1164 );
nor ( n1271 , n1265 , n1270 );
nand ( n1272 , n1253 , n1262 , n1271 );
not ( n1273 , n191 );
and ( n1274 , n1272 , n1273 );
not ( n1275 , n1272 );
and ( n1276 , n1275 , n191 );
nor ( n1277 , n1274 , n1276 );
and ( n1278 , n1228 , n1277 );
nor ( n1279 , n1227 , n1278 );
and ( n1280 , n96 , n509 );
and ( n1281 , n88 , n199 );
nor ( n1282 , n1280 , n1281 );
and ( n1283 , n1223 , n1282 );
not ( n1284 , n1223 );
not ( n1285 , n139 );
and ( n1286 , n235 , n1285 );
not ( n1287 , n235 );
and ( n1288 , n1287 , n139 );
or ( n1289 , n1286 , n1288 );
buf ( n1290 , n1289 );
buf ( n1291 , n1290 );
not ( n1292 , n1291 );
xor ( n1293 , n140 , n240 );
not ( n1294 , n1293 );
not ( n1295 , n1294 );
not ( n1296 , n1295 );
xor ( n1297 , n138 , n245 );
buf ( n1298 , n1297 );
not ( n1299 , n1298 );
xor ( n1300 , n137 , n228 );
xor ( n1301 , n136 , n250 );
not ( n1302 , n1301 );
not ( n1303 , n1302 );
xor ( n1304 , n135 , n231 );
not ( n1305 , n1304 );
nand ( n1306 , n1300 , n1303 , n1305 );
nor ( n1307 , n1299 , n1306 );
nand ( n1308 , n1292 , n1296 , n1307 );
not ( n1309 , n1293 );
buf ( n1310 , n1309 );
buf ( n1311 , n1290 );
not ( n1312 , n1298 );
xor ( n1313 , n137 , n228 );
not ( n1314 , n1304 );
nand ( n1315 , n1313 , n1314 , n1302 );
nor ( n1316 , n1312 , n1315 );
nand ( n1317 , n1310 , n1311 , n1316 );
and ( n1318 , n1308 , n1317 );
not ( n1319 , n1291 );
not ( n1320 , n1319 );
not ( n1321 , n1297 );
not ( n1322 , n1300 );
not ( n1323 , n1301 );
not ( n1324 , n1323 );
and ( n1325 , n1321 , n1322 , n1324 , n1305 );
not ( n1326 , n1325 );
buf ( n1327 , n1293 );
buf ( n1328 , n1327 );
nor ( n1329 , n1326 , n1328 );
nand ( n1330 , n1320 , n1329 );
not ( n1331 , n1291 );
not ( n1332 , n1331 );
not ( n1333 , n1294 );
not ( n1334 , n1313 );
nand ( n1335 , n1321 , n1334 , n1304 , n1323 );
nor ( n1336 , n1333 , n1335 );
nand ( n1337 , n1332 , n1336 );
and ( n1338 , n1330 , n1337 );
not ( n1339 , n1290 );
not ( n1340 , n1339 );
not ( n1341 , n1340 );
not ( n1342 , n1309 );
not ( n1343 , n1298 );
and ( n1344 , n1313 , n1304 , n1301 );
nand ( n1345 , n1343 , n1344 );
nor ( n1346 , n1342 , n1345 );
nand ( n1347 , n1341 , n1346 );
not ( n1348 , n1340 );
nand ( n1349 , n1348 , n1336 );
nand ( n1350 , n1318 , n1338 , n1347 , n1349 );
not ( n1351 , n1339 );
buf ( n1352 , n1327 );
not ( n1353 , n1345 );
nand ( n1354 , n1351 , n1352 , n1353 );
not ( n1355 , n1304 );
not ( n1356 , n1355 );
not ( n1357 , n1300 );
not ( n1358 , n1297 );
nand ( n1359 , n1356 , n1357 , n1358 , n1324 );
nor ( n1360 , n1310 , n1359 );
nand ( n1361 , n1291 , n1360 );
nand ( n1362 , n1354 , n1361 );
nand ( n1363 , n1311 , n1342 , n1325 );
not ( n1364 , n1339 );
not ( n1365 , n1315 );
nand ( n1366 , n1312 , n1365 );
nor ( n1367 , n1366 , n1310 );
nand ( n1368 , n1364 , n1367 );
nand ( n1369 , n1363 , n1368 );
nor ( n1370 , n1362 , n1369 );
buf ( n1371 , n1290 );
not ( n1372 , n1371 );
not ( n1373 , n1372 );
not ( n1374 , n1309 );
not ( n1375 , n1313 );
not ( n1376 , n1302 );
nand ( n1377 , n1375 , n1376 , n1355 );
nor ( n1378 , n1343 , n1377 );
nand ( n1379 , n1374 , n1378 );
not ( n1380 , n1379 );
nand ( n1381 , n1373 , n1380 );
nand ( n1382 , n1304 , n1323 );
not ( n1383 , n1313 );
nor ( n1384 , n1382 , n1383 );
nand ( n1385 , n1312 , n1384 );
not ( n1386 , n1385 );
nand ( n1387 , n1319 , n1352 , n1386 );
nand ( n1388 , n1381 , n1387 );
not ( n1389 , n1358 );
and ( n1390 , n1327 , n1389 , n1344 );
nand ( n1391 , n1292 , n1390 );
not ( n1392 , n1311 );
not ( n1393 , n1335 );
nand ( n1394 , n1295 , n1393 );
not ( n1395 , n1394 );
nand ( n1396 , n1392 , n1395 );
nand ( n1397 , n1391 , n1396 );
nor ( n1398 , n1388 , n1397 );
nand ( n1399 , n1370 , n1398 );
nor ( n1400 , n1350 , n1399 );
buf ( n1401 , n1311 );
not ( n1402 , n1401 );
not ( n1403 , n1402 );
nor ( n1404 , n1304 , n1301 );
nand ( n1405 , n1357 , n1404 );
nor ( n1406 , n1343 , n1405 );
nand ( n1407 , n1296 , n1406 );
not ( n1408 , n1407 );
and ( n1409 , n1403 , n1408 );
not ( n1410 , n1374 );
not ( n1411 , n1358 );
nor ( n1412 , n1411 , n1306 );
nand ( n1413 , n1410 , n1412 );
nor ( n1414 , n1348 , n1413 );
nor ( n1415 , n1409 , n1414 );
not ( n1416 , n1300 );
not ( n1417 , n1416 );
and ( n1418 , n1293 , n1303 );
not ( n1419 , n1293 );
and ( n1420 , n1419 , n1323 );
nor ( n1421 , n1418 , n1420 );
nor ( n1422 , n1417 , n1421 );
not ( n1423 , n1305 );
not ( n1424 , n1321 );
or ( n1425 , n1423 , n1424 );
not ( n1426 , n1355 );
nand ( n1427 , n1426 , n1297 );
nand ( n1428 , n1425 , n1427 );
and ( n1429 , n1422 , n1331 , n1428 );
not ( n1430 , n1293 );
nor ( n1431 , n1430 , n1321 );
nor ( n1432 , n1300 , n1382 );
nand ( n1433 , n1431 , n1290 , n1432 );
not ( n1434 , n1433 );
nor ( n1435 , n1429 , n1434 );
not ( n1436 , n1390 );
nor ( n1437 , n1341 , n1436 );
not ( n1438 , n1437 );
nor ( n1439 , n1401 , n1413 );
not ( n1440 , n1291 );
and ( n1441 , n1440 , n1410 , n1406 );
nor ( n1442 , n1439 , n1441 );
and ( n1443 , n1435 , n1438 , n1442 );
not ( n1444 , n1291 );
nand ( n1445 , n1352 , n1444 , n1412 );
nand ( n1446 , n1342 , n1372 , n1406 );
nand ( n1447 , n1445 , n1446 );
nand ( n1448 , n1311 , n1346 );
nor ( n1449 , n1333 , n1385 );
not ( n1450 , n1321 );
nand ( n1451 , n1450 , n1344 );
nor ( n1452 , n1333 , n1451 );
nand ( n1453 , n1304 , n1301 );
nor ( n1454 , n1300 , n1453 );
nand ( n1455 , n1450 , n1294 , n1454 );
nor ( n1456 , n1339 , n1455 );
not ( n1457 , n1456 );
not ( n1458 , n1311 );
nand ( n1459 , n1328 , n1458 , n1307 );
not ( n1460 , n1311 );
not ( n1461 , n1309 );
and ( n1462 , n1461 , n1450 , n1365 );
nor ( n1463 , n1447 , t_0 );
nand ( n1464 , n1400 , n1415 , n1443 , n1463 );
not ( n1465 , n184 );
and ( n1466 , n1464 , n1465 );
not ( n1467 , n1464 );
and ( n1468 , n1467 , n184 );
nor ( n1469 , n1466 , n1468 );
and ( n1470 , n1284 , n1469 );
nor ( n1471 , n1283 , n1470 );
not ( n1472 , n507 );
not ( n1473 , n1472 );
and ( n1474 , n78 , n509 );
and ( n1475 , n70 , n199 );
nor ( n1476 , n1474 , n1475 );
and ( n1477 , n1473 , n1476 );
not ( n1478 , n1473 );
not ( n1479 , n1118 );
nand ( n1480 , n1041 , n1479 );
nand ( n1481 , n1010 , n1117 );
nand ( n1482 , n1480 , n1481 );
nor ( n1483 , n985 , n981 );
nand ( n1484 , n950 , n1483 );
nand ( n1485 , n987 , n1484 );
nor ( n1486 , n1482 , n1485 );
not ( n1487 , n950 );
not ( n1488 , n1004 );
not ( n1489 , n1488 );
or ( n1490 , n1487 , n1489 );
nand ( n1491 , n1490 , n983 );
not ( n1492 , n1491 );
nand ( n1493 , n1486 , n1492 , n1059 );
not ( n1494 , n1075 );
not ( n1495 , n1043 );
nand ( n1496 , n1070 , n1494 , n1495 );
not ( n1497 , n965 );
nor ( n1498 , n963 , n956 );
and ( n1499 , n1023 , n1498 );
nor ( n1500 , n1499 , n1024 );
or ( n1501 , n1500 , n974 , n1003 );
not ( n1502 , n1011 );
or ( n1503 , n1018 , n1002 , n1502 );
nand ( n1504 , n1501 , n1503 );
nand ( n1505 , n1497 , n1504 );
and ( n1506 , n1496 , n1505 );
not ( n1507 , n1075 );
nand ( n1508 , n1507 , n1041 , n1001 , n1012 );
nand ( n1509 , n1506 , n1015 , n1508 , n1045 );
nor ( n1510 , n1493 , n1509 );
not ( n1511 , n1085 );
nand ( n1512 , n988 , n985 , n1511 );
nand ( n1513 , n1512 , n1096 );
not ( n1514 , n1513 );
and ( n1515 , n1091 , n1068 );
nand ( n1516 , n1070 , n1072 );
not ( n1517 , n1516 );
not ( n1518 , n1124 );
nand ( n1519 , n950 , n1518 );
not ( n1520 , n1519 );
nor ( n1521 , n1517 , n1520 );
not ( n1522 , n1083 );
nand ( n1523 , n1006 , n1072 );
not ( n1524 , n1523 );
nor ( n1525 , n1522 , n1524 );
nand ( n1526 , n1514 , n1515 , n1521 , n1525 );
not ( n1527 , n980 );
nor ( n1528 , n959 , n1527 );
nand ( n1529 , n1507 , n1070 , n1528 );
not ( n1530 , n1125 );
nand ( n1531 , n1529 , n1530 );
not ( n1532 , n1531 );
not ( n1533 , n1100 );
nor ( n1534 , n1533 , n1119 );
nand ( n1535 , n950 , n1056 );
not ( n1536 , n1535 );
not ( n1537 , n1107 );
nor ( n1538 , n1536 , n1537 );
and ( n1539 , n1010 , n1064 );
nor ( n1540 , n950 , n1077 );
nor ( n1541 , n1539 , n1540 );
nand ( n1542 , n1532 , n1534 , n1538 , n1541 );
nor ( n1543 , n1526 , n1542 );
nand ( n1544 , n1510 , n1543 );
not ( n1545 , n178 );
and ( n1546 , n1544 , n1545 );
not ( n1547 , n1544 );
and ( n1548 , n1547 , n178 );
nor ( n1549 , n1546 , n1548 );
and ( n1550 , n1478 , n1549 );
nor ( n1551 , n1477 , n1550 );
not ( n1552 , n507 );
not ( n1553 , n1552 );
and ( n1554 , n82 , n509 );
and ( n1555 , n74 , n199 );
nor ( n1556 , n1554 , n1555 );
and ( n1557 , n1553 , n1556 );
not ( n1558 , n1553 );
nand ( n1559 , n1041 , n1483 );
and ( n1560 , n1060 , n1559 );
or ( n1561 , n1002 , n1022 , n1009 );
nand ( n1562 , n952 , n949 );
not ( n1563 , n1498 );
nand ( n1564 , n1563 , n1022 );
nand ( n1565 , n1002 , n1564 );
or ( n1566 , n1562 , n1565 );
nand ( n1567 , n1561 , n1566 );
nand ( n1568 , n965 , n1567 );
and ( n1569 , n1496 , n1568 );
nand ( n1570 , n976 , n1008 );
not ( n1571 , n1570 );
nand ( n1572 , n1571 , n968 );
nand ( n1573 , n1560 , n1569 , n1572 , n1045 );
not ( n1574 , n1480 );
nor ( n1575 , n1491 , n1574 );
nand ( n1576 , n950 , n1044 );
not ( n1577 , n1576 );
not ( n1578 , n1484 );
nor ( n1579 , n1577 , n1578 );
not ( n1580 , n1058 );
not ( n1581 , n987 );
nor ( n1582 , n1581 , n993 );
nand ( n1583 , n1575 , n1579 , n1580 , n1582 );
nor ( n1584 , n1573 , n1583 );
and ( n1585 , n1065 , n1096 );
nand ( n1586 , n950 , n1106 );
and ( n1587 , n1586 , n1523 );
not ( n1588 , n1090 );
nand ( n1589 , n1588 , n1050 );
nand ( n1590 , n1087 , n1519 );
nor ( n1591 , n1589 , n1590 );
nand ( n1592 , n1585 , n1587 , n1591 );
not ( n1593 , n1530 );
nor ( n1594 , n1593 , n1115 );
not ( n1595 , n1082 );
nor ( n1596 , n1006 , n1595 );
nor ( n1597 , n1596 , n1539 );
not ( n1598 , n1529 );
nor ( n1599 , n1598 , n1101 );
nor ( n1600 , n1123 , n1121 );
nand ( n1601 , n1594 , n1597 , n1599 , n1600 );
nor ( n1602 , n1592 , n1601 );
nand ( n1603 , n1584 , n1602 );
not ( n1604 , n194 );
and ( n1605 , n1603 , n1604 );
not ( n1606 , n1603 );
and ( n1607 , n1606 , n194 );
nor ( n1608 , n1605 , n1607 );
and ( n1609 , n1558 , n1608 );
nor ( n1610 , n1557 , n1609 );
not ( n1611 , n831 );
nand ( n1612 , n734 , n790 );
not ( n1613 , n1612 );
nor ( n1614 , n1611 , n1613 );
not ( n1615 , n897 );
nand ( n1616 , n1614 , n870 , n1615 );
not ( n1617 , n1616 );
not ( n1618 , n765 );
nand ( n1619 , n1618 , n732 , n770 , n767 );
not ( n1620 , n1619 );
not ( n1621 , n788 );
or ( n1622 , n1621 , n781 );
nor ( n1623 , n745 , n750 );
not ( n1624 , n1623 );
nand ( n1625 , n1624 , n751 );
not ( n1626 , n1625 );
nand ( n1627 , n1626 , n811 , n769 );
nand ( n1628 , n1622 , n1627 );
nand ( n1629 , n1628 , n733 );
not ( n1630 , n1629 );
or ( n1631 , n1620 , n1630 );
nand ( n1632 , n1631 , n740 );
not ( n1633 , n863 );
nand ( n1634 , n1633 , n851 , n923 );
nand ( n1635 , n899 , n816 , n919 );
nand ( n1636 , n1632 , n1634 , n1635 );
nand ( n1637 , n917 , n855 );
nor ( n1638 , n1636 , n1637 );
and ( n1639 , n913 , n791 );
not ( n1640 , n812 );
nand ( n1641 , n1640 , n901 , n813 );
not ( n1642 , n1641 );
not ( n1643 , n859 );
not ( n1644 , n895 );
or ( n1645 , n1643 , n1644 );
nand ( n1646 , n813 , n901 , n912 );
nand ( n1647 , n1645 , n1646 );
nor ( n1648 , n1642 , n1647 );
nand ( n1649 , n1617 , n1638 , n1639 , n1648 );
nand ( n1650 , n734 , n873 );
nand ( n1651 , n883 , n1650 );
nand ( n1652 , n771 , n815 , n903 );
nor ( n1653 , n1621 , n809 );
nand ( n1654 , n757 , n901 , n1653 );
nand ( n1655 , n1652 , n1654 );
not ( n1656 , n1655 );
nand ( n1657 , n1656 , n874 , n891 );
nor ( n1658 , n1651 , n1657 );
and ( n1659 , n920 , n864 );
nand ( n1660 , n819 , n877 );
not ( n1661 , n1660 );
not ( n1662 , n836 );
nor ( n1663 , n735 , n1662 );
nor ( n1664 , n1661 , n1663 );
nand ( n1665 , n757 , n733 , n848 );
and ( n1666 , n1665 , n805 , n837 , n908 );
nand ( n1667 , n1658 , n1659 , n1664 , n1666 );
nor ( n1668 , n1649 , n1667 );
not ( n1669 , n1668 );
not ( n1670 , n187 );
and ( n1671 , n1669 , n1670 );
nor ( n1672 , n1667 , n1649 );
and ( n1673 , n187 , n1672 );
nor ( n1674 , n1671 , n1673 );
or ( n1675 , n1674 , n937 );
nand ( n1676 , n72 , n936 );
or ( n1677 , n199 , n1676 );
nand ( n1678 , n1675 , n1677 );
and ( n1679 , n108 , n509 );
and ( n1680 , n100 , n199 );
nor ( n1681 , n1679 , n1680 );
and ( n1682 , n508 , n1681 );
not ( n1683 , n508 );
xor ( n1684 , n154 , n216 );
buf ( n1685 , n1684 );
buf ( n1686 , n1685 );
xor ( n1687 , n153 , n224 );
not ( n1688 , n1687 );
not ( n1689 , n1688 );
xor ( n1690 , n152 , n202 );
not ( n1691 , n1690 );
xor ( n1692 , n151 , n220 );
nand ( n1693 , n1691 , n1692 );
nor ( n1694 , n1689 , n1693 );
nand ( n1695 , n1686 , n1694 );
xor ( n1696 , n156 , n205 );
not ( n1697 , n1696 );
buf ( n1698 , n1697 );
nor ( n1699 , n1695 , n1698 );
xor ( n1700 , n155 , n209 );
buf ( n1701 , n1700 );
not ( n1702 , n1701 );
not ( n1703 , n1702 );
nand ( n1704 , n1699 , n1703 );
not ( n1705 , n1704 );
not ( n1706 , n1705 );
not ( n1707 , n1690 );
nor ( n1708 , n1707 , n1692 );
nand ( n1709 , n1689 , n1708 );
not ( n1710 , n1684 );
buf ( n1711 , n1710 );
not ( n1712 , n1711 );
nor ( n1713 , n1709 , n1712 );
nand ( n1714 , n1713 , n1698 );
nor ( n1715 , n1714 , n1703 );
not ( n1716 , n1715 );
not ( n1717 , n1686 );
buf ( n1718 , n1692 );
not ( n1719 , n1690 );
not ( n1720 , n1719 );
not ( n1721 , n1687 );
not ( n1722 , n1721 );
and ( n1723 , n1718 , n1720 , n1722 );
and ( n1724 , n1717 , n1723 );
buf ( n1725 , n1696 );
not ( n1726 , n1725 );
not ( n1727 , n1726 );
nand ( n1728 , n1724 , n1703 , n1727 );
nand ( n1729 , n1706 , n1716 , n1728 );
not ( n1730 , n1685 );
nor ( n1731 , n1692 , n1690 );
and ( n1732 , n1688 , n1731 );
nand ( n1733 , n1730 , n1732 );
not ( n1734 , n1733 );
not ( n1735 , n1697 );
not ( n1736 , n1735 );
buf ( n1737 , n1700 );
not ( n1738 , n1737 );
nand ( n1739 , n1734 , n1736 , n1738 );
not ( n1740 , n1719 );
not ( n1741 , n1740 );
not ( n1742 , n1741 );
nor ( n1743 , n1702 , n1742 );
not ( n1744 , n1721 );
not ( n1745 , n1744 );
not ( n1746 , n1745 );
not ( n1747 , n1746 );
buf ( n1748 , n1692 );
not ( n1749 , n1748 );
not ( n1750 , n1710 );
and ( n1751 , n156 , n205 );
not ( n1752 , n156 );
not ( n1753 , n205 );
and ( n1754 , n1752 , n1753 );
nor ( n1755 , n1751 , n1754 );
not ( n1756 , n1755 );
nand ( n1757 , n1749 , n1750 , n1756 );
not ( n1758 , n1710 );
not ( n1759 , n1692 );
not ( n1760 , n1759 );
or ( n1761 , n1758 , n1760 );
nand ( n1762 , n1684 , n1718 );
nand ( n1763 , n1761 , n1762 );
nand ( n1764 , n1725 , n1763 );
nand ( n1765 , n1757 , n1764 );
not ( n1766 , n1765 );
or ( n1767 , n1747 , n1766 );
nor ( n1768 , n1722 , n1759 );
not ( n1769 , n1685 );
nand ( n1770 , n1768 , n1697 , n1769 );
nand ( n1771 , n1767 , n1770 );
nand ( n1772 , n1743 , n1771 );
nand ( n1773 , n1739 , n1772 );
nor ( n1774 , n1729 , n1773 );
buf ( n1775 , n1701 );
not ( n1776 , n1775 );
nor ( n1777 , n1714 , n1776 );
not ( n1778 , n1777 );
buf ( n1779 , n1725 );
nor ( n1780 , n1779 , n1695 );
not ( n1781 , n1780 );
not ( n1782 , n1738 );
nor ( n1783 , n1781 , n1782 );
not ( n1784 , n1783 );
not ( n1785 , n1737 );
not ( n1786 , n1693 );
nand ( n1787 , n1744 , n1786 );
not ( n1788 , n1755 );
nand ( n1789 , n1685 , n1788 );
nor ( n1790 , n1787 , n1789 );
nand ( n1791 , n1785 , n1790 );
nor ( n1792 , n1755 , n1700 );
not ( n1793 , n1750 );
nand ( n1794 , n1718 , n1690 );
nor ( n1795 , n1794 , n1689 );
nand ( n1796 , n1793 , n1795 );
not ( n1797 , n1796 );
nand ( n1798 , n1792 , n1797 );
nand ( n1799 , n1791 , n1798 );
not ( n1800 , n1737 );
not ( n1801 , n1800 );
not ( n1802 , n1731 );
not ( n1803 , n1802 );
nand ( n1804 , n1803 , n1712 , n1697 , n1745 );
not ( n1805 , n1804 );
nand ( n1806 , n1801 , n1805 );
buf ( n1807 , n1785 );
nand ( n1808 , n1807 , n1805 );
nand ( n1809 , n1806 , n1808 );
not ( n1810 , n1775 );
nand ( n1811 , n1688 , n1708 );
nor ( n1812 , n1711 , n1811 );
nand ( n1813 , n1810 , n1736 , n1812 );
not ( n1814 , n1735 );
not ( n1815 , n1802 );
nand ( n1816 , n1815 , n1689 );
nor ( n1817 , n1816 , n1730 );
nand ( n1818 , n1814 , n1800 , n1817 );
nand ( n1819 , n1813 , n1818 );
nor ( n1820 , n1799 , n1809 , n1819 );
and ( n1821 , n1774 , n1778 , n1784 , n1820 );
nor ( n1822 , n1796 , n1736 );
nand ( n1823 , n1782 , n1822 );
not ( n1824 , n1701 );
not ( n1825 , n1824 );
not ( n1826 , n1685 );
and ( n1827 , n1826 , n1744 , n1786 );
nand ( n1828 , n1735 , n1827 );
not ( n1829 , n1828 );
nand ( n1830 , n1825 , n1829 );
and ( n1831 , n1823 , n1830 );
nand ( n1832 , n1779 , n1812 );
nor ( n1833 , n1832 , n1810 );
not ( n1834 , n1737 );
not ( n1835 , n1697 );
nand ( n1836 , n1835 , n1817 );
nor ( n1837 , n1834 , n1836 );
nor ( n1838 , n1833 , n1837 );
nand ( n1839 , n1712 , n1723 );
nor ( n1840 , n1698 , n1839 );
nand ( n1841 , n1807 , n1840 );
nand ( n1842 , n1776 , n1822 );
nor ( n1843 , n1730 , n1709 );
nand ( n1844 , n1835 , n1737 , n1843 );
nand ( n1845 , n1776 , n1699 );
and ( n1846 , n1841 , n1842 , n1844 , n1845 );
nand ( n1847 , n1831 , n1838 , n1846 );
nor ( n1848 , n1733 , n1726 );
nand ( n1849 , n1848 , n1782 );
not ( n1850 , n1849 );
not ( n1851 , n1839 );
and ( n1852 , n1738 , n1736 , n1851 );
nor ( n1853 , n1850 , n1852 );
not ( n1854 , n1725 );
and ( n1855 , n1854 , n1793 , n1723 );
nand ( n1856 , n1825 , n1855 );
not ( n1857 , n1856 );
nor ( n1858 , n1836 , n1825 );
nor ( n1859 , n1857 , n1858 );
not ( n1860 , n1769 );
nand ( n1861 , n1726 , n1737 , n1860 , n1795 );
not ( n1862 , n1824 );
nand ( n1863 , n1862 , n1790 );
and ( n1864 , n1861 , n1863 );
and ( n1865 , n1702 , n1835 , n1812 );
nor ( n1866 , n1686 , n1811 );
and ( n1867 , n1727 , n1702 , n1866 );
nor ( n1868 , n1865 , n1867 );
nand ( n1869 , n1853 , n1859 , n1864 , n1868 );
nor ( n1870 , n1847 , n1869 );
nand ( n1871 , n1821 , n1870 );
not ( n1872 , n166 );
and ( n1873 , n1871 , n1872 );
not ( n1874 , n1871 );
and ( n1875 , n1874 , n166 );
nor ( n1876 , n1873 , n1875 );
and ( n1877 , n1683 , n1876 );
nor ( n1878 , n1682 , n1877 );
and ( n1879 , n122 , n509 );
and ( n1880 , n114 , n199 );
nor ( n1881 , n1879 , n1880 );
and ( n1882 , n939 , n1881 );
not ( n1883 , n939 );
not ( n1884 , n1455 );
nand ( n1885 , n1392 , n1884 );
and ( n1886 , n1347 , n1885 );
not ( n1887 , n1366 );
nand ( n1888 , n1296 , n1311 , n1887 );
not ( n1889 , n1374 );
nor ( n1890 , n1411 , n1405 );
nand ( n1891 , n1889 , n1291 , n1890 );
and ( n1892 , n1888 , n1891 );
nand ( n1893 , n1348 , n1449 );
nand ( n1894 , n1886 , n1892 , n1893 , n1349 );
nor ( n1895 , n1460 , n1394 );
nor ( n1896 , n1895 , n1362 );
not ( n1897 , n1381 );
not ( n1898 , n1462 );
not ( n1899 , n1371 );
nor ( n1900 , n1898 , n1899 );
nor ( n1901 , n1897 , n1900 );
not ( n1902 , n1291 );
nand ( n1903 , n1902 , n1360 );
and ( n1904 , n1391 , n1903 , n1387 );
nand ( n1905 , n1896 , n1901 , n1904 );
nor ( n1906 , n1894 , n1905 );
not ( n1907 , n1441 );
not ( n1908 , n1324 );
nor ( n1909 , n1908 , n1352 );
not ( n1910 , n1299 );
and ( n1911 , n1313 , n1355 );
nand ( n1912 , n1909 , n1910 , n1401 , n1911 );
nand ( n1913 , n1907 , n1308 , n1912 );
nand ( n1914 , n1293 , n1297 );
not ( n1915 , n1384 );
nor ( n1916 , n1914 , n1915 );
not ( n1917 , n1916 );
nor ( n1918 , n1917 , n1341 );
not ( n1919 , n1918 );
nand ( n1920 , n1348 , n1329 );
or ( n1921 , n1295 , n1416 , n1427 );
nand ( n1922 , n1428 , n1327 , n1416 );
nand ( n1923 , n1921 , n1922 );
nand ( n1924 , n1923 , n1341 , n1908 );
nand ( n1925 , n1919 , n1920 , n1924 );
nor ( n1926 , n1913 , n1925 );
nand ( n1927 , n1341 , n1367 );
not ( n1928 , n1359 );
nand ( n1929 , n1340 , n1410 , n1928 );
nand ( n1930 , n1929 , n1445 );
nor ( n1931 , t_2 , n1930 );
nand ( n1932 , n1906 , n1415 , n1926 , n1931 );
not ( n1933 , n189 );
and ( n1934 , n1932 , n1933 );
not ( n1935 , n1932 );
and ( n1936 , n1935 , n189 );
nor ( n1937 , n1934 , n1936 );
and ( n1938 , n1883 , n1937 );
nor ( n1939 , n1882 , n1938 );
not ( n1940 , n61 );
and ( n1941 , n1211 , n1940 );
not ( n1942 , n1211 );
nor ( n1943 , n733 , n853 );
not ( n1944 , n1943 );
not ( n1945 , n771 );
or ( n1946 , n765 , n750 , n739 );
nand ( n1947 , n763 , n750 , n911 );
nand ( n1948 , n1946 , n1947 );
not ( n1949 , n1948 );
or ( n1950 , n1945 , n1949 );
not ( n1951 , n739 );
nand ( n1952 , n766 , n826 , n767 , n1951 );
nand ( n1953 , n1950 , n1952 );
nand ( n1954 , n907 , n1953 );
nand ( n1955 , n1944 , n1954 , n1634 );
nand ( n1956 , n1612 , n925 );
nor ( n1957 , n1955 , n1956 );
and ( n1958 , n760 , n829 );
nand ( n1959 , n858 , n734 , n1958 );
and ( n1960 , n1650 , n1959 );
nor ( n1961 , n1647 , n909 );
nand ( n1962 , n849 , n894 );
nor ( n1963 , n1962 , n871 );
nand ( n1964 , n1957 , n1960 , n1961 , n1963 );
and ( n1965 , n883 , n817 );
and ( n1966 , n886 , n791 );
and ( n1967 , n891 , n1652 );
and ( n1968 , n1965 , n1966 , n1967 );
and ( n1969 , n861 , n924 );
nand ( n1970 , n819 , n804 );
not ( n1971 , n1970 );
nor ( n1972 , n1663 , n1971 );
not ( n1973 , n805 );
nand ( n1974 , n1665 , n864 );
not ( n1975 , n893 );
nor ( n1976 , n1975 , n1643 );
nor ( n1977 , n1973 , n1974 , n1976 );
nand ( n1978 , n1968 , n1969 , n1972 , n1977 );
nor ( n1979 , n1964 , n1978 );
not ( n1980 , n1979 );
not ( n1981 , n165 );
and ( n1982 , n1980 , n1981 );
and ( n1983 , n165 , n1979 );
nor ( n1984 , n1982 , n1983 );
and ( n1985 , n1942 , n1984 );
nor ( n1986 , n1941 , n1985 );
not ( n1987 , n17 );
and ( n1988 , n722 , n1987 );
not ( n1989 , n722 );
and ( n1990 , n1989 , n1674 );
nor ( n1991 , n1988 , n1990 );
and ( n1992 , n116 , n509 );
and ( n1993 , n108 , n199 );
nor ( n1994 , n1992 , n1993 );
and ( n1995 , n937 , n1994 );
not ( n1996 , n937 );
and ( n1997 , n1996 , n1984 );
nor ( n1998 , n1995 , n1997 );
not ( n1999 , n23 );
and ( n2000 , n1472 , n1999 );
not ( n2001 , n1472 );
and ( n2002 , n2001 , n1549 );
nor ( n2003 , n2000 , n2002 );
not ( n2004 , n936 );
not ( n2005 , n41 );
and ( n2006 , n2004 , n2005 );
not ( n2007 , n2004 );
and ( n2008 , n2007 , n1469 );
nor ( n2009 , n2006 , n2008 );
not ( n2010 , n53 );
and ( n2011 , n1217 , n2010 );
not ( n2012 , n1217 );
and ( n2013 , n2012 , n1876 );
nor ( n2014 , n2011 , n2013 );
not ( n2015 , n936 );
not ( n2016 , n67 );
and ( n2017 , n2015 , n2016 );
not ( n2018 , n2015 );
and ( n2019 , n2018 , n1937 );
nor ( n2020 , n2017 , n2019 );
not ( n2021 , n936 );
not ( n2022 , n51 );
and ( n2023 , n2021 , n2022 );
not ( n2024 , n2021 );
and ( n2025 , n2024 , n1277 );
nor ( n2026 , n2023 , n2025 );
not ( n2027 , n27 );
and ( n2028 , n1205 , n2027 );
not ( n2029 , n1205 );
and ( n2030 , n2029 , n1608 );
nor ( n2031 , n2028 , n2030 );
and ( n2032 , n126 , n509 );
and ( n2033 , n118 , n199 );
nor ( n2034 , n2032 , n2033 );
and ( n2035 , n1223 , n2034 );
not ( n2036 , n1223 );
not ( n2037 , n1708 );
not ( n2038 , n2037 );
nand ( n2039 , n2038 , n1717 , n1725 , n1746 );
nor ( n2040 , n2039 , n1834 );
nor ( n2041 , n2040 , n1833 );
not ( n2042 , n1865 );
nand ( n2043 , n2041 , n2042 , n1849 );
not ( n2044 , n2039 );
nand ( n2045 , n1807 , n2044 );
nand ( n2046 , n1810 , n1848 );
nand ( n2047 , n1864 , n2045 , n2046 );
nor ( n2048 , n2043 , n2047 );
nand ( n2049 , n1801 , n1840 );
nand ( n2050 , n2049 , n1704 );
not ( n2051 , n1837 );
not ( n2052 , n1737 );
not ( n2053 , n2052 );
nor ( n2054 , n1828 , n2053 );
nand ( n2055 , n1725 , n1860 , n1795 );
nor ( n2056 , n1775 , n2055 );
nor ( n2057 , n2054 , n2056 );
nand ( n2058 , n2051 , n2057 , n1842 );
nor ( n2059 , n2050 , n2058 );
nand ( n2060 , n2048 , n1831 , n2059 );
nand ( n2061 , n1818 , n1716 );
not ( n2062 , n1860 );
not ( n2063 , n2062 );
not ( n2064 , n1740 );
nor ( n2065 , n2064 , n1688 );
not ( n2066 , n1700 );
nor ( n2067 , n2066 , n1748 );
nand ( n2068 , n2065 , n1697 , n2067 );
nor ( n2069 , n1756 , n1700 );
not ( n2070 , n1718 );
not ( n2071 , n1722 );
or ( n2072 , n2070 , n2071 );
or ( n2073 , n1748 , n1689 );
nand ( n2074 , n2072 , n2073 );
nand ( n2075 , n2069 , n1741 , n2074 );
nand ( n2076 , n2068 , n2075 );
nand ( n2077 , n2063 , n2076 );
not ( n2078 , n1816 );
nand ( n2079 , n2078 , n1717 , n1854 );
or ( n2080 , n1775 , n2079 );
not ( n2081 , n1770 );
not ( n2082 , n1742 );
not ( n2083 , n2082 );
nand ( n2084 , n2081 , n2083 , n2053 );
nand ( n2085 , n2077 , n2080 , n1739 , n2084 );
nor ( n2086 , n2061 , n2085 );
not ( n2087 , n2052 );
and ( n2088 , n1698 , n2087 , n1866 );
not ( n2089 , n1801 );
not ( n2090 , n1780 );
or ( n2091 , n2089 , n2090 );
nand ( n2092 , n2091 , n1856 );
nor ( n2093 , n2088 , n2092 );
nor ( n2094 , n1834 , n2079 );
nor ( n2095 , n1852 , n2094 );
nor ( n2096 , n1755 , n1685 );
not ( n2097 , n1701 );
nand ( n2098 , n2096 , n2097 , n1694 );
nand ( n2099 , n1806 , n2098 );
not ( n2100 , n1855 );
nor ( n2101 , n2100 , n1782 );
nor ( n2102 , n2099 , n2101 );
nand ( n2103 , n2086 , n2093 , n2095 , n2102 );
nor ( n2104 , n2060 , n2103 );
not ( n2105 , n2104 );
not ( n2106 , n172 );
and ( n2107 , n2105 , n2106 );
and ( n2108 , n172 , n2104 );
nor ( n2109 , n2107 , n2108 );
and ( n2110 , n2036 , n2109 );
nor ( n2111 , n2035 , n2110 );
not ( n2112 , n171 );
xor ( n2113 , n147 , n232 );
buf ( n2114 , n2113 );
xor ( n2115 , n148 , n243 );
not ( n2116 , n2115 );
buf ( n2117 , n2116 );
not ( n2118 , n2117 );
xor ( n2119 , n146 , n253 );
not ( n2120 , n2119 );
xor ( n2121 , n145 , n247 );
buf ( n2122 , n2121 );
not ( n2123 , n2122 );
not ( n2124 , n2123 );
xor ( n2125 , n143 , n229 );
xor ( n2126 , n144 , n237 );
nand ( n2127 , n2125 , n2126 );
not ( n2128 , n2127 );
nand ( n2129 , n2120 , n2124 , n2128 );
nor ( n2130 , n2118 , n2129 );
nand ( n2131 , n2114 , n2130 );
buf ( n2132 , n2115 );
not ( n2133 , n2132 );
buf ( n2134 , n2133 );
buf ( n2135 , n2121 );
not ( n2136 , n2126 );
and ( n2137 , n2135 , n2125 , n2136 );
not ( n2138 , n2137 );
not ( n2139 , n2120 );
nor ( n2140 , n2138 , n2139 );
nand ( n2141 , n2114 , n2134 , n2140 );
and ( n2142 , n2131 , n2141 );
buf ( n2143 , n2113 );
not ( n2144 , n2125 );
and ( n2145 , n2122 , n2126 , n2144 );
not ( n2146 , n2145 );
not ( n2147 , n2146 );
not ( n2148 , n2133 );
buf ( n2149 , n2119 );
not ( n2150 , n2149 );
nand ( n2151 , n2147 , n2148 , n2150 );
nor ( n2152 , n2143 , n2151 );
not ( n2153 , n2143 );
xor ( n2154 , n143 , n229 );
nor ( n2155 , n2154 , n2126 );
not ( n2156 , n2155 );
not ( n2157 , n2156 );
not ( n2158 , n2116 );
not ( n2159 , n2119 );
not ( n2160 , n2159 );
not ( n2161 , n2121 );
not ( n2162 , n2161 );
not ( n2163 , n2162 );
nand ( n2164 , n2157 , n2158 , n2160 , n2163 );
not ( n2165 , n2164 );
nand ( n2166 , n2153 , n2165 );
not ( n2167 , n2166 );
nor ( n2168 , n2152 , n2167 );
not ( n2169 , n2127 );
not ( n2170 , n2123 );
nand ( n2171 , n2169 , n2149 , n2170 );
not ( n2172 , n2171 );
not ( n2173 , n2132 );
nand ( n2174 , n2172 , n2173 , n2143 );
not ( n2175 , n2143 );
buf ( n2176 , n2132 );
not ( n2177 , n2149 );
nor ( n2178 , n2154 , n2126 );
nand ( n2179 , n2162 , n2178 );
nor ( n2180 , n2177 , n2179 );
nand ( n2181 , n2175 , n2176 , n2180 );
nand ( n2182 , n2174 , n2181 );
not ( n2183 , n2126 );
and ( n2184 , n2161 , n2125 , n2183 );
not ( n2185 , n2184 );
nor ( n2186 , n2177 , n2185 );
nand ( n2187 , n2143 , n2173 , n2186 );
not ( n2188 , n2122 );
and ( n2189 , n2188 , n2178 );
not ( n2190 , n2113 );
nor ( n2191 , n2190 , n2119 );
nand ( n2192 , n2189 , n2118 , n2191 );
nand ( n2193 , n2187 , n2192 );
nor ( n2194 , n2182 , n2193 );
and ( n2195 , n2142 , n2168 , n2194 );
not ( n2196 , n2143 );
not ( n2197 , n2117 );
not ( n2198 , n2160 );
nand ( n2199 , n2163 , n2128 );
nor ( n2200 , n2198 , n2199 );
nand ( n2201 , n2196 , n2197 , n2200 );
not ( n2202 , n2201 );
not ( n2203 , n2143 );
not ( n2204 , n2203 );
not ( n2205 , n2127 );
not ( n2206 , n2163 );
nand ( n2207 , n2205 , n2206 , n2150 , n2176 );
nor ( n2208 , n2204 , n2207 );
nor ( n2209 , n2202 , n2208 );
buf ( n2210 , n2143 );
buf ( n2211 , n2126 );
not ( n2212 , n2154 );
nand ( n2213 , n2188 , n2149 , n2211 , n2212 );
nor ( n2214 , n2213 , n2173 );
nand ( n2215 , n2210 , n2214 );
buf ( n2216 , n2114 );
nand ( n2217 , n2159 , n2184 );
nor ( n2218 , n2117 , n2217 );
nand ( n2219 , n2216 , n2218 );
and ( n2220 , n2215 , n2219 );
nand ( n2221 , n2149 , n2145 );
not ( n2222 , n2221 );
not ( n2223 , n2117 );
nand ( n2224 , n2222 , n2223 , n2114 );
buf ( n2225 , n2158 );
and ( n2226 , n2120 , n2188 , n2128 );
nand ( n2227 , n2143 , n2225 , n2226 );
nand ( n2228 , n2224 , n2227 );
not ( n2229 , n2143 );
nor ( n2230 , n2229 , n2164 );
not ( n2231 , n2230 );
not ( n2232 , n2114 );
nand ( n2233 , n2232 , n2218 );
nand ( n2234 , n2231 , n2233 );
nor ( n2235 , n2228 , n2234 );
nand ( n2236 , n2195 , n2209 , n2220 , n2235 );
not ( n2237 , n2113 );
and ( n2238 , n2237 , n2116 );
not ( n2239 , n2238 );
or ( n2240 , n2239 , n2213 );
nor ( n2241 , n2134 , n2171 );
nand ( n2242 , n2210 , n2241 );
nand ( n2243 , n2114 , n2223 , n2186 );
nand ( n2244 , n2240 , n2242 , n2243 );
and ( n2245 , n2149 , n2188 , n2155 );
nand ( n2246 , n2245 , n2173 );
nor ( n2247 , n2246 , n2216 );
not ( n2248 , n2247 );
not ( n2249 , n2211 );
not ( n2250 , n2249 );
not ( n2251 , n2250 );
not ( n2252 , n2132 );
not ( n2253 , n2154 );
not ( n2254 , n2135 );
or ( n2255 , n2253 , n2254 );
or ( n2256 , n2154 , n2162 );
nand ( n2257 , n2255 , n2256 );
nand ( n2258 , n2251 , n2252 , n2198 , n2257 );
not ( n2259 , n2258 );
not ( n2260 , n2135 );
nand ( n2261 , n2125 , n2119 );
nor ( n2262 , n2260 , n2261 );
or ( n2263 , n2250 , n2262 );
not ( n2264 , n2249 );
not ( n2265 , n2122 );
nor ( n2266 , n2154 , n2119 );
nand ( n2267 , n2265 , n2266 );
nand ( n2268 , n2264 , n2267 );
nand ( n2269 , n2263 , n2268 , n2176 );
not ( n2270 , n2269 );
or ( n2271 , n2259 , n2270 );
not ( n2272 , n2114 );
nand ( n2273 , n2271 , n2272 );
nand ( n2274 , n2248 , n2273 );
nor ( n2275 , n2244 , n2274 );
nor ( n2276 , n2225 , n2221 );
nand ( n2277 , n2203 , n2276 );
and ( n2278 , n2133 , n2160 , n2124 , n2155 );
nand ( n2279 , n2272 , n2278 );
and ( n2280 , n2277 , n2279 );
not ( n2281 , n2146 );
nand ( n2282 , n2281 , n2143 , n2173 , n2198 );
not ( n2283 , n2179 );
nand ( n2284 , n2177 , n2283 );
not ( n2285 , n2284 );
nand ( n2286 , n2285 , n2143 , n2134 );
nand ( n2287 , n2282 , n2286 );
not ( n2288 , n2287 );
not ( n2289 , n2114 );
not ( n2290 , n2289 );
not ( n2291 , n2127 );
not ( n2292 , n2124 );
nand ( n2293 , n2291 , n2252 , n2139 , n2292 );
not ( n2294 , n2293 );
not ( n2295 , n2294 );
or ( n2296 , n2290 , n2295 );
nand ( n2297 , n2238 , n2226 );
nand ( n2298 , n2296 , n2297 );
and ( n2299 , n2117 , n2159 , n2184 );
and ( n2300 , n2153 , n2299 );
not ( n2301 , n2153 );
and ( n2302 , n2301 , n2278 );
nor ( n2303 , n2300 , n2302 );
not ( n2304 , n2303 );
nor ( n2305 , n2298 , n2304 );
nand ( n2306 , n2275 , n2280 , n2288 , n2305 );
nor ( n2307 , n2236 , n2306 );
not ( n2308 , n2307 );
and ( n2309 , n2112 , n2308 );
and ( n2310 , n171 , n2307 );
nor ( n2311 , n2309 , n2310 );
or ( n2312 , n508 , n2311 );
nand ( n2313 , n68 , n936 );
or ( n2314 , n199 , n2313 );
nand ( n2315 , n2312 , n2314 );
and ( n2316 , n80 , n509 );
and ( n2317 , n72 , n199 );
nor ( n2318 , n2316 , n2317 );
and ( n2319 , n939 , n2318 );
not ( n2320 , n939 );
xor ( n2321 , n149 , n208 );
not ( n2322 , n2321 );
xor ( n2323 , n148 , n215 );
xor ( n2324 , n147 , n226 );
nor ( n2325 , n2323 , n2324 );
nand ( n2326 , n2322 , n2325 );
xor ( n2327 , n150 , n201 );
not ( n2328 , n2327 );
not ( n2329 , n2328 );
nor ( n2330 , n2326 , n2329 );
not ( n2331 , n2330 );
xor ( n2332 , n152 , n212 );
not ( n2333 , n2332 );
xor ( n2334 , n151 , n221 );
not ( n2335 , n2334 );
nand ( n2336 , n2333 , n2335 );
nor ( n2337 , n2331 , n2336 );
not ( n2338 , n2324 );
not ( n2339 , n2338 );
not ( n2340 , n2323 );
and ( n2341 , n2321 , n2339 , n2340 );
not ( n2342 , n2341 );
xor ( n2343 , n149 , n208 );
not ( n2344 , n2324 );
nand ( n2345 , n2323 , n2344 );
nor ( n2346 , n2343 , n2345 );
not ( n2347 , n2346 );
and ( n2348 , n2342 , n2347 );
buf ( n2349 , n2334 );
not ( n2350 , n2328 );
not ( n2351 , n2332 );
not ( n2352 , n2351 );
or ( n2353 , n2350 , n2352 );
xor ( n2354 , n152 , n212 );
nand ( n2355 , n2327 , n2354 );
nand ( n2356 , n2353 , n2355 );
nand ( n2357 , n2349 , n2356 );
nor ( n2358 , n2348 , n2357 );
nor ( n2359 , n2337 , n2358 );
not ( n2360 , n2327 );
not ( n2361 , n2343 );
not ( n2362 , n2361 );
and ( n2363 , n2360 , n2362 , n2325 );
not ( n2364 , n2333 );
not ( n2365 , n2364 );
not ( n2366 , n2349 );
nand ( n2367 , n2363 , n2365 , n2366 );
not ( n2368 , n2351 );
buf ( n2369 , n2368 );
not ( n2370 , n2366 );
nand ( n2371 , n2323 , n2324 );
not ( n2372 , n2371 );
nand ( n2373 , n2372 , n2362 , n2329 );
not ( n2374 , n2373 );
nand ( n2375 , n2369 , n2370 , n2374 );
buf ( n2376 , n2327 );
not ( n2377 , n2376 );
not ( n2378 , n2377 );
nor ( n2379 , n2343 , n2371 );
nand ( n2380 , n2378 , n2379 );
not ( n2381 , n2380 );
not ( n2382 , n2334 );
not ( n2383 , n2382 );
buf ( n2384 , n2383 );
buf ( n2385 , n2364 );
nand ( n2386 , n2381 , n2384 , n2385 );
and ( n2387 , n2359 , n2367 , n2375 , n2386 );
not ( n2388 , n2324 );
nand ( n2389 , n2388 , n2321 , n2323 );
not ( n2390 , n2389 );
buf ( n2391 , n2376 );
not ( n2392 , n2391 );
not ( n2393 , n2392 );
not ( n2394 , n2332 );
not ( n2395 , n2394 );
not ( n2396 , n2395 );
not ( n2397 , n2366 );
nand ( n2398 , n2390 , n2393 , n2396 , n2397 );
not ( n2399 , n2334 );
buf ( n2400 , n2399 );
nand ( n2401 , n2378 , n2346 );
nor ( n2402 , n2369 , n2401 );
nand ( n2403 , n2400 , n2402 );
nand ( n2404 , n2398 , n2403 );
not ( n2405 , n2342 );
not ( n2406 , n2382 );
nor ( n2407 , n2368 , n2406 );
nand ( n2408 , n2405 , n2407 , n2392 );
not ( n2409 , n2332 );
not ( n2410 , n2409 );
nor ( n2411 , n2329 , n2389 );
not ( n2412 , n2411 );
nor ( n2413 , n2410 , n2412 );
nand ( n2414 , n2400 , n2413 );
nand ( n2415 , n2408 , n2414 );
nor ( n2416 , n2404 , n2415 );
buf ( n2417 , n2366 );
nor ( n2418 , n2410 , n2380 );
nand ( n2419 , n2417 , n2418 );
not ( n2420 , n2349 );
not ( n2421 , n2343 );
nor ( n2422 , n2344 , n2323 );
and ( n2423 , n2329 , n2421 , n2422 );
nand ( n2424 , n2396 , n2420 , n2423 );
nand ( n2425 , n2419 , n2424 );
not ( n2426 , n2425 );
not ( n2427 , n2417 );
not ( n2428 , n2395 );
not ( n2429 , n2391 );
nor ( n2430 , n2429 , n2389 );
nand ( n2431 , n2428 , n2430 );
or ( n2432 , n2427 , n2431 );
not ( n2433 , n2326 );
and ( n2434 , n2378 , n2433 );
nand ( n2435 , n2428 , n2384 , n2434 );
nand ( n2436 , n2432 , n2435 );
not ( n2437 , n2436 );
and ( n2438 , n2387 , n2416 , n2426 , n2437 );
not ( n2439 , n2409 );
not ( n2440 , n2349 );
not ( n2441 , n2338 );
nor ( n2442 , n2321 , n2340 , n2441 );
nand ( n2443 , n2360 , n2442 );
not ( n2444 , n2443 );
nand ( n2445 , n2439 , n2440 , n2444 );
not ( n2446 , n2445 );
buf ( n2447 , n2383 );
not ( n2448 , n2447 );
not ( n2449 , n2418 );
or ( n2450 , n2448 , n2449 );
nor ( n2451 , n2399 , n2368 );
nand ( n2452 , n2451 , n2391 , n2341 );
nand ( n2453 , n2450 , n2452 );
nor ( n2454 , n2446 , n2453 );
nor ( n2455 , n2439 , n2373 );
nand ( n2456 , n2400 , n2455 );
not ( n2457 , n2344 );
and ( n2458 , n2377 , n2421 , n2323 , n2457 );
nand ( n2459 , n2428 , n2447 , n2458 );
and ( n2460 , n2456 , n2459 );
nand ( n2461 , n2395 , n2330 );
not ( n2462 , n2461 );
nand ( n2463 , n2400 , n2462 );
not ( n2464 , n2463 );
buf ( n2465 , n2399 );
not ( n2466 , n2401 );
nand ( n2467 , n2385 , n2465 , n2466 );
not ( n2468 , n2376 );
nand ( n2469 , n2343 , n2325 );
nor ( n2470 , n2468 , n2469 );
nand ( n2471 , n2369 , n2440 , n2470 );
nand ( n2472 , n2467 , n2471 );
nor ( n2473 , n2464 , n2472 );
nand ( n2474 , n2454 , n2460 , n2473 );
and ( n2475 , n2360 , n2421 , n2457 , n2340 );
nand ( n2476 , n2439 , n2475 );
nor ( n2477 , n2427 , n2476 );
not ( n2478 , n2477 );
not ( n2479 , n2384 );
nand ( n2480 , n2439 , n2423 );
not ( n2481 , n2480 );
and ( n2482 , n2479 , n2481 );
not ( n2483 , n2479 );
not ( n2484 , n2364 );
nor ( n2485 , n2322 , n2371 );
nand ( n2486 , n2468 , n2485 );
nor ( n2487 , n2484 , n2486 );
and ( n2488 , n2483 , n2487 );
nor ( n2489 , n2482 , n2488 );
nand ( n2490 , n2478 , n2489 );
nand ( n2491 , n2465 , n2487 );
nand ( n2492 , n2439 , n2420 , n2458 );
nand ( n2493 , n2491 , n2492 );
not ( n2494 , n2493 );
not ( n2495 , n2363 );
nor ( n2496 , n2396 , n2495 );
nand ( n2497 , n2427 , n2496 );
nand ( n2498 , n2410 , n2383 , n2411 );
not ( n2499 , n2498 );
nor ( n2500 , n2465 , n2461 );
nor ( n2501 , n2499 , n2500 );
nand ( n2502 , n2494 , n2497 , n2501 );
nor ( n2503 , n2474 , n2490 , n2502 );
nand ( n2504 , n2438 , n2503 );
not ( n2505 , n186 );
and ( n2506 , n2504 , n2505 );
not ( n2507 , n2504 );
and ( n2508 , n2507 , n186 );
nor ( n2509 , n2506 , n2508 );
and ( n2510 , n2320 , n2509 );
nor ( n2511 , n2319 , n2510 );
and ( n2512 , n84 , n509 );
and ( n2513 , n76 , n199 );
nor ( n2514 , n2512 , n2513 );
and ( n2515 , n508 , n2514 );
not ( n2516 , n508 );
or ( n2517 , n522 , n639 );
not ( n2518 , n1148 );
nand ( n2519 , n563 , n536 );
not ( n2520 , n2519 );
not ( n2521 , n2520 );
nand ( n2522 , n2518 , n2521 );
nor ( n2523 , n550 , n529 );
nand ( n2524 , n2522 , n534 , n2523 );
not ( n2525 , n594 );
or ( n2526 , n2525 , n2520 );
nor ( n2527 , n556 , n534 );
not ( n2528 , n1148 );
nand ( n2529 , n685 , n2528 );
nand ( n2530 , n2526 , n2527 , n2529 );
nand ( n2531 , n2524 , n2530 );
nand ( n2532 , n2531 , n629 );
nand ( n2533 , n2517 , n2532 , n1230 );
not ( n2534 , n1185 );
not ( n2535 , n626 );
nor ( n2536 , n2533 , n2534 , n2535 );
nand ( n2537 , n1163 , n618 );
not ( n2538 , n2537 );
nand ( n2539 , n2538 , n607 , n1155 );
nand ( n2540 , n1232 , n600 );
nor ( n2541 , n2539 , n2540 );
nand ( n2542 , n2536 , n616 , n692 , n2541 );
nand ( n2543 , n1256 , n1264 , n1173 );
nand ( n2544 , n689 , n1180 , n1171 );
nor ( n2545 , n2543 , n2544 );
not ( n2546 , n679 );
nor ( n2547 , n2546 , n662 );
not ( n2548 , n1181 );
nor ( n2549 , n2548 , n657 );
and ( n2550 , n2549 , n669 , n1194 );
nand ( n2551 , n2545 , n2547 , n2550 );
nor ( n2552 , n2542 , n2551 );
not ( n2553 , n2552 );
not ( n2554 , n169 );
and ( n2555 , n2553 , n2554 );
and ( n2556 , n169 , n2552 );
nor ( n2557 , n2555 , n2556 );
and ( n2558 , n2516 , n2557 );
nor ( n2559 , n2515 , n2558 );
and ( n2560 , n104 , n509 );
and ( n2561 , n96 , n199 );
nor ( n2562 , n2560 , n2561 );
and ( n2563 , n1223 , n2562 );
not ( n2564 , n1223 );
not ( n2565 , n1497 );
not ( n2566 , n1002 );
or ( n2567 , n1502 , n2566 , n1570 );
not ( n2568 , n1031 );
nand ( n2569 , n989 , n948 );
nand ( n2570 , n1047 , n1023 );
nand ( n2571 , n952 , n2568 , n2569 , n2570 );
nand ( n2572 , n2567 , n2571 );
not ( n2573 , n2572 );
or ( n2574 , n2565 , n2573 );
nand ( n2575 , n2574 , n1496 );
not ( n2576 , n1018 );
nand ( n2577 , n2576 , n1012 );
and ( n2578 , n2577 , n1050 );
nand ( n2579 , n2578 , n1013 , n1559 );
nor ( n2580 , n2575 , n2579 );
nand ( n2581 , n1061 , n1576 );
nand ( n2582 , n971 , n1481 );
nor ( n2583 , n2581 , n2582 );
and ( n2584 , n2580 , n2583 , n1492 , n1059 );
not ( n2585 , n1586 );
nor ( n2586 , n2585 , n1524 );
nand ( n2587 , n950 , n1078 );
not ( n2588 , n2587 );
nand ( n2589 , n1068 , n1512 );
nor ( n2590 , n2588 , n2589 , n1596 );
and ( n2591 , n1585 , n2586 , n2590 );
or ( n2592 , n1598 , n1108 );
and ( n2593 , n1535 , n1114 );
not ( n2594 , n1540 );
not ( n2595 , n1123 );
nand ( n2596 , n2593 , n2594 , n2595 , n1530 );
nor ( n2597 , n2592 , n2596 );
nand ( n2598 , n2584 , n2591 , n2597 );
not ( n2599 , n183 );
and ( n2600 , n2598 , n2599 );
not ( n2601 , n2598 );
and ( n2602 , n2601 , n183 );
nor ( n2603 , n2600 , n2602 );
and ( n2604 , n2564 , n2603 );
nor ( n2605 , n2563 , n2604 );
and ( n2606 , n110 , n509 );
and ( n2607 , n102 , n199 );
nor ( n2608 , n2606 , n2607 );
and ( n2609 , n1473 , n2608 );
not ( n2610 , n1473 );
not ( n2611 , n1347 );
nor ( n2612 , n2611 , n1414 );
nand ( n2613 , n1296 , n1291 , n1378 );
nand ( n2614 , n2613 , n1891 );
not ( n2615 , n2614 );
and ( n2616 , n2615 , n1317 , n1893 );
nand ( n2617 , n2612 , n2616 );
not ( n2618 , n1354 );
nor ( n2619 , n2618 , n1369 );
nand ( n2620 , n1331 , n1916 );
not ( n2621 , n2620 );
nor ( n2622 , n2621 , n1434 );
and ( n2623 , n1391 , n1903 , n1396 );
nand ( n2624 , n2619 , n2622 , n2623 );
nor ( n2625 , n2617 , n2624 );
not ( n2626 , n1340 );
and ( n2627 , n2626 , n1452 );
not ( n2628 , n2626 );
and ( n2629 , n2628 , n1336 );
nor ( n2630 , n2627 , n2629 );
not ( n2631 , n1910 );
nand ( n2632 , n1402 , n2631 , n1911 , n1420 );
nand ( n2633 , n2632 , n1442 );
not ( n2634 , n1918 );
nor ( n2635 , n1305 , n1300 );
not ( n2636 , n2635 );
not ( n2637 , n1420 );
or ( n2638 , n2636 , n2637 );
or ( n2639 , n2635 , n1911 );
nand ( n2640 , n2639 , n1418 );
nand ( n2641 , n2638 , n2640 );
not ( n2642 , n1331 );
nand ( n2643 , n2641 , n2642 , n1910 );
nand ( n2644 , n2634 , n1920 , n2643 );
nor ( n2645 , n2633 , n2644 );
nand ( n2646 , n1459 , n1457 );
nand ( n2647 , n1328 , n1371 , n1890 );
and ( n2648 , n1929 , n2647 );
nand ( n2649 , n2648 , t_3 , t_1 );
nor ( n2650 , n2646 , n2649 );
nand ( n2651 , n2625 , n2630 , n2645 , n2650 );
not ( n2652 , n174 );
and ( n2653 , n2651 , n2652 );
not ( n2654 , n2651 );
and ( n2655 , n2654 , n174 );
nor ( n2656 , n2653 , n2655 );
and ( n2657 , n2610 , n2656 );
nor ( n2658 , n2609 , n2657 );
and ( n2659 , n118 , n509 );
and ( n2660 , n110 , n199 );
nor ( n2661 , n2659 , n2660 );
and ( n2662 , n937 , n2661 );
not ( n2663 , n937 );
and ( n2664 , n1641 , n1646 );
nand ( n2665 , n2664 , n825 , n896 );
not ( n2666 , n2665 );
nand ( n2667 , n2666 , n872 , n857 );
nand ( n2668 , n875 , n739 , n756 , n1625 );
not ( n2669 , n2668 );
and ( n2670 , n773 , n821 );
not ( n2671 , n773 );
not ( n2672 , n835 );
and ( n2673 , n2671 , n2672 );
nor ( n2674 , n2670 , n2673 );
nand ( n2675 , n2674 , n740 , n796 );
not ( n2676 , n2675 );
or ( n2677 , n2669 , n2676 );
nand ( n2678 , n2677 , n907 );
and ( n2679 , n1635 , n2678 );
not ( n2680 , n1943 );
nand ( n2681 , n2679 , n1634 , n2680 );
nor ( n2682 , n2667 , n2681 );
and ( n2683 , n886 , n1654 );
nand ( n2684 , n2683 , n891 , n913 , n791 );
nand ( n2685 , n915 , n1650 , n1959 );
nor ( n2686 , n2684 , n2685 );
not ( n2687 , n1976 );
nand ( n2688 , n2687 , n878 , n837 );
nand ( n2689 , n1660 , n861 , n864 );
nand ( n2690 , n1665 , n1970 );
nor ( n2691 , n2688 , n2689 , n2690 );
nand ( n2692 , n2682 , n2686 , n2691 );
not ( n2693 , n173 );
and ( n2694 , n2692 , n2693 );
not ( n2695 , n2692 );
and ( n2696 , n2695 , n173 );
nor ( n2697 , n2694 , n2696 );
and ( n2698 , n2663 , n2697 );
nor ( n2699 , n2662 , n2698 );
and ( n2700 , n124 , n509 );
and ( n2701 , n116 , n199 );
nor ( n2702 , n2700 , n2701 );
and ( n2703 , n1223 , n2702 );
not ( n2704 , n1223 );
nand ( n2705 , n1903 , n1927 );
buf ( n2706 , n1330 );
nand ( n2707 , n2706 , n1920 );
nand ( n2708 , n1893 , n1349 );
nor ( n2709 , n2705 , n2707 , n2708 );
not ( n2710 , n1448 );
nor ( n2711 , n2710 , n1439 );
not ( n2712 , n1457 );
nor ( n2713 , n1437 , n2712 );
nor ( n2714 , n1900 , n1895 );
and ( n2715 , n2630 , n2711 , n2713 , n2714 );
not ( n2716 , n1417 );
not ( n2717 , n2716 );
not ( n2718 , n1356 );
and ( n2719 , n2718 , n1291 );
not ( n2720 , n2718 );
and ( n2721 , n2720 , n1339 );
nor ( n2722 , n2719 , n2721 );
and ( n2723 , n2722 , n1910 , n1420 );
and ( n2724 , n1290 , n1356 );
not ( n2725 , n1290 );
and ( n2726 , n2725 , n2718 );
nor ( n2727 , n2724 , n2726 );
and ( n2728 , n2727 , n1299 , n1418 );
nor ( n2729 , n2723 , n2728 );
not ( n2730 , n2729 );
and ( n2731 , n2717 , n2730 );
nand ( n2732 , n1308 , n1907 );
nor ( n2733 , n2731 , n2732 );
and ( n2734 , n1445 , n1446 );
and ( n2735 , n1354 , n1387 );
and ( n2736 , n1459 , n1363 );
nand ( n2737 , n2734 , n2735 , n2736 );
and ( n2738 , n1885 , n2613 );
nand ( n2739 , n1433 , n2620 );
nand ( n2740 , n1888 , n2647 );
nor ( n2741 , n2739 , n2740 );
nand ( n2742 , n2738 , n2741 );
nor ( n2743 , n2737 , n2742 );
nand ( n2744 , n2709 , n2715 , n2733 , n2743 );
not ( n2745 , n164 );
and ( n2746 , n2744 , n2745 );
not ( n2747 , n2744 );
and ( n2748 , n2747 , n164 );
nor ( n2749 , n2746 , n2748 );
and ( n2750 , n2704 , n2749 );
nor ( n2751 , n2703 , n2750 );
nand ( n2752 , n2365 , n2420 , n2470 );
and ( n2753 , n2752 , n2435 );
not ( n2754 , n2398 );
nor ( n2755 , n2332 , n2334 );
nand ( n2756 , n2755 , n2475 );
nand ( n2757 , n2408 , n2756 );
nor ( n2758 , n2754 , n2757 );
nand ( n2759 , n2447 , n2413 );
nand ( n2760 , n2394 , n2335 );
nor ( n2761 , n2760 , n2443 );
nor ( n2762 , n2337 , n2761 );
and ( n2763 , n2759 , n2414 , n2762 );
nand ( n2764 , n2753 , n2758 , n2763 );
not ( n2765 , n2344 );
nand ( n2766 , n2376 , n2765 );
nor ( n2767 , n2327 , n2339 );
not ( n2768 , n2767 );
nand ( n2769 , n2766 , n2768 );
not ( n2770 , n2354 );
and ( n2771 , n2770 , n2340 );
nand ( n2772 , n2769 , n2383 , n2771 );
not ( n2773 , n2772 );
or ( n2774 , n2335 , n2767 );
and ( n2775 , n2354 , n2323 );
nand ( n2776 , n2399 , n2766 );
nand ( n2777 , n2774 , n2775 , n2776 );
not ( n2778 , n2777 );
or ( n2779 , n2773 , n2778 );
not ( n2780 , n2421 );
not ( n2781 , n2780 );
nand ( n2782 , n2779 , n2781 );
nand ( n2783 , n2468 , n2341 );
not ( n2784 , n2783 );
nand ( n2785 , n2784 , n2385 , n2397 );
nand ( n2786 , n2427 , n2487 );
nand ( n2787 , n2782 , n2785 , n2386 , n2786 );
nor ( n2788 , n2764 , n2787 );
nand ( n2789 , n2400 , n2496 );
nand ( n2790 , n2789 , n2460 );
not ( n2791 , n2400 );
nor ( n2792 , n2439 , n2486 );
not ( n2793 , n2792 );
nor ( n2794 , n2791 , n2793 );
not ( n2795 , n2794 );
nand ( n2796 , n2791 , n2455 );
not ( n2797 , n2472 );
nand ( n2798 , n2795 , n2419 , n2796 , n2797 );
nor ( n2799 , n2790 , n2798 );
not ( n2800 , n2476 );
and ( n2801 , n2791 , n2800 );
nand ( n2802 , n2368 , n2335 );
nand ( n2803 , n2391 , n2341 );
nor ( n2804 , n2802 , n2803 );
nor ( n2805 , n2801 , n2804 );
nand ( n2806 , n2492 , n2805 );
not ( n2807 , n2420 );
and ( n2808 , n2364 , n2391 , n2433 );
nand ( n2809 , n2807 , n2808 );
not ( n2810 , n2809 );
nor ( n2811 , n2810 , n2477 );
nor ( n2812 , n2394 , n2406 );
nand ( n2813 , n2812 , n2430 );
not ( n2814 , n2813 );
nor ( n2815 , n2814 , n2500 );
nand ( n2816 , n2811 , n2497 , n2815 );
nor ( n2817 , n2806 , n2816 );
nand ( n2818 , n2788 , n2799 , n2817 );
not ( n2819 , n195 );
and ( n2820 , n2818 , n2819 );
not ( n2821 , n2818 );
and ( n2822 , n2821 , n195 );
nor ( n2823 , n2820 , n2822 );
or ( n2824 , n2823 , n508 );
nand ( n2825 , n74 , n936 );
or ( n2826 , n199 , n2825 );
nand ( n2827 , n2824 , n2826 );
not ( n2828 , n63 );
and ( n2829 , n1211 , n2828 );
not ( n2830 , n1211 );
and ( n2831 , n2830 , n2697 );
nor ( n2832 , n2829 , n2831 );
not ( n2833 , n2 );
and ( n2834 , n2004 , n2833 );
not ( n2835 , n2004 );
and ( n2836 , n2835 , n2749 );
nor ( n2837 , n2834 , n2836 );
not ( n2838 , n508 );
not ( n2839 , n29 );
and ( n2840 , n2838 , n2839 );
not ( n2841 , n2838 );
and ( n2842 , n2841 , n2557 );
nor ( n2843 , n2840 , n2842 );
not ( n2844 , n13 );
and ( n2845 , n1472 , n2844 );
not ( n2846 , n1472 );
and ( n2847 , n2846 , n2311 );
nor ( n2848 , n2845 , n2847 );
not ( n2849 , n4 );
and ( n2850 , n2021 , n2849 );
not ( n2851 , n2021 );
and ( n2852 , n2851 , n2109 );
nor ( n2853 , n2850 , n2852 );
and ( n2854 , n128 , n509 );
and ( n2855 , n120 , n199 );
nor ( n2856 , n2854 , n2855 );
and ( n2857 , n1473 , n2856 );
not ( n2858 , n1473 );
not ( n2859 , n1746 );
not ( n2860 , n1697 );
nor ( n2861 , n1793 , n2860 );
or ( n2862 , n1749 , n1700 );
not ( n2863 , n2067 );
nand ( n2864 , n2862 , n2863 );
nand ( n2865 , n2083 , n2859 , n2861 , n2864 );
and ( n2866 , n1818 , n2865 );
not ( n2867 , n2049 );
nor ( n2868 , n1825 , n1804 );
nor ( n2869 , n2867 , n2868 );
not ( n2870 , n1700 );
not ( n2871 , n1768 );
or ( n2872 , n2870 , n2871 );
nand ( n2873 , n1749 , n1689 , n2066 );
nand ( n2874 , n2872 , n2873 );
and ( n2875 , n1727 , n2062 , n2082 , n2874 );
nor ( n2876 , n1715 , n2875 );
nand ( n2877 , n2866 , n2869 , n2876 );
nand ( n2878 , n1698 , n1862 , n1827 );
nand ( n2879 , n1791 , n2878 );
nand ( n2880 , n1843 , n1698 , n1785 );
nand ( n2881 , n1798 , n2880 );
nor ( n2882 , n2879 , n2881 );
not ( n2883 , n2098 );
nor ( n2884 , n2094 , n2883 );
nor ( n2885 , n1777 , n2088 );
nand ( n2886 , n2882 , n2884 , n2885 );
nor ( n2887 , n2877 , n2886 );
not ( n2888 , n2092 );
nand ( n2889 , n1863 , n2888 );
not ( n2890 , n2046 );
nor ( n2891 , n2890 , n2040 );
not ( n2892 , n1732 );
nor ( n2893 , n1793 , n2892 );
nand ( n2894 , n1727 , n1775 , n2893 );
nand ( n2895 , n2891 , n2894 , n1868 );
nor ( n2896 , n2889 , n2895 );
not ( n2897 , n1845 );
not ( n2898 , n2897 );
not ( n2899 , n1837 );
nand ( n2900 , n2898 , n2899 );
not ( n2901 , n2055 );
nand ( n2902 , n1801 , n2901 );
not ( n2903 , n1844 );
nor ( n2904 , n2903 , n2054 );
nand ( n2905 , n1841 , n2902 , n2904 );
nor ( n2906 , n2900 , n2905 );
nand ( n2907 , n2887 , n2896 , n1831 , n2906 );
not ( n2908 , n180 );
and ( n2909 , n2907 , n2908 );
not ( n2910 , n2907 );
and ( n2911 , n2910 , n180 );
nor ( n2912 , n2909 , n2911 );
and ( n2913 , n2858 , n2912 );
nor ( n2914 , n2857 , n2913 );
not ( n2915 , n55 );
and ( n2916 , n2015 , n2915 );
not ( n2917 , n2015 );
and ( n2918 , n2917 , n2656 );
nor ( n2919 , n2916 , n2918 );
not ( n2920 , n6 );
and ( n2921 , n1472 , n2920 );
not ( n2922 , n1472 );
and ( n2923 , n2922 , n2912 );
nor ( n2924 , n2921 , n2923 );
not ( n2925 , n49 );
and ( n2926 , n2021 , n2925 );
not ( n2927 , n2021 );
and ( n2928 , n2927 , n2603 );
nor ( n2929 , n2926 , n2928 );
not ( n2930 , n936 );
not ( n2931 , n25 );
and ( n2932 , n2930 , n2931 );
not ( n2933 , n2930 );
and ( n2934 , n2933 , n2509 );
nor ( n2935 , n2932 , n2934 );
not ( n2936 , n19 );
and ( n2937 , n2015 , n2936 );
not ( n2938 , n2015 );
and ( n2939 , n2938 , n2823 );
nor ( n2940 , n2937 , n2939 );
and ( n2941 , n114 , n509 );
and ( n2942 , n106 , n199 );
nor ( n2943 , n2941 , n2942 );
and ( n2944 , n508 , n2943 );
not ( n2945 , n508 );
and ( n2946 , n2080 , n1813 );
not ( n2947 , n1737 );
or ( n2948 , n1725 , n2947 , n1802 );
or ( n2949 , n1786 , n1700 );
nand ( n2950 , n1700 , n2037 );
nand ( n2951 , n2949 , n2950 , n1725 );
nand ( n2952 , n2948 , n2951 );
and ( n2953 , n2952 , n2062 , n2859 );
not ( n2954 , n1762 );
nand ( n2955 , n1742 , n1701 , n2954 );
nor ( n2956 , n2859 , n2955 , n1779 );
nor ( n2957 , n2953 , n2956 );
nand ( n2958 , n2946 , n2957 , n2880 , n1818 );
nand ( n2959 , n2878 , n1798 );
nor ( n2960 , n2101 , n1783 );
not ( n2961 , n2099 );
nand ( n2962 , n2960 , n2961 , n2885 );
nor ( n2963 , n2958 , n2959 , n2962 );
and ( n2964 , n1728 , n1823 );
not ( n2965 , n2056 );
and ( n2966 , n1841 , n2965 );
and ( n2967 , n2902 , n1704 );
nand ( n2968 , n2964 , n2966 , n2967 , n2904 );
not ( n2969 , n1864 );
nand ( n2970 , n2045 , n2046 );
nor ( n2971 , n2969 , n2970 );
nor ( n2972 , n1865 , n1858 );
and ( n2973 , n2972 , n2894 , n1849 );
nand ( n2974 , n2971 , n2973 );
nor ( n2975 , n2968 , n2974 );
nand ( n2976 , n2963 , n2975 );
not ( n2977 , n190 );
and ( n2978 , n2976 , n2977 );
not ( n2979 , n2976 );
and ( n2980 , n2979 , n190 );
nor ( n2981 , n2978 , n2980 );
and ( n2982 , n2945 , n2981 );
nor ( n2983 , n2944 , n2982 );
and ( n2984 , n112 , n509 );
and ( n2985 , n104 , n199 );
nor ( n2986 , n2984 , n2985 );
and ( n2987 , n939 , n2986 );
not ( n2988 , n939 );
not ( n2989 , n2219 );
nand ( n2990 , n2241 , n2289 );
not ( n2991 , n2990 );
nor ( n2992 , n2989 , n2991 );
nand ( n2993 , n2224 , n2227 );
and ( n2994 , n2149 , n2137 );
nand ( n2995 , n2114 , n2197 , n2994 );
not ( n2996 , n2114 );
nand ( n2997 , n2140 , n2225 , n2996 );
nand ( n2998 , n2995 , n2997 );
nor ( n2999 , n2993 , n2998 );
and ( n3000 , n2209 , n2992 , n2999 );
nand ( n3001 , n2203 , n2214 );
not ( n3002 , n3001 );
not ( n3003 , n2181 );
nor ( n3004 , n3002 , n3003 );
not ( n3005 , n3004 );
nor ( n3006 , n2289 , n2151 );
nor ( n3007 , n3006 , n2230 );
and ( n3008 , n2174 , n2141 );
not ( n3009 , n2284 );
and ( n3010 , n2114 , n2197 , n3009 );
not ( n3011 , n2192 );
nor ( n3012 , n3010 , n3011 );
nand ( n3013 , n3007 , n3008 , n3012 );
nor ( n3014 , n3005 , n3013 );
not ( n3015 , n2154 );
nand ( n3016 , n2265 , n2211 , n3015 );
nor ( n3017 , n2149 , n3016 );
nand ( n3018 , n2252 , n3017 );
nor ( n3019 , n2114 , n3018 );
nor ( n3020 , n3019 , n2247 );
not ( n3021 , n2277 );
nor ( n3022 , n2272 , n3018 );
nor ( n3023 , n3021 , n3022 );
not ( n3024 , n2239 );
not ( n3025 , n2284 );
and ( n3026 , n3024 , n3025 );
not ( n3027 , n2206 );
not ( n3028 , n2261 );
nand ( n3029 , n2251 , n3028 , n2238 );
not ( n3030 , n2127 );
nand ( n3031 , n3030 , n2149 , n2113 );
nand ( n3032 , n2190 , n2249 , n2266 );
nand ( n3033 , n3031 , n3032 );
nand ( n3034 , n2223 , n3033 );
nand ( n3035 , n3029 , n3034 );
and ( n3036 , n3027 , n3035 );
nor ( n3037 , n3026 , n3036 );
and ( n3038 , n3020 , n3023 , n3037 );
not ( n3039 , n2130 );
nor ( n3040 , n2216 , n3039 );
nor ( n3041 , n2210 , n2293 );
nor ( n3042 , n3040 , n3041 );
and ( n3043 , n2204 , n2299 );
not ( n3044 , n2994 );
nor ( n3045 , n2239 , n3044 );
nor ( n3046 , n3043 , n3045 );
not ( n3047 , n2282 );
not ( n3048 , n2143 );
nor ( n3049 , n2246 , n3048 );
nor ( n3050 , n3047 , n3049 );
and ( n3051 , n3042 , n3046 , n3050 , n2303 );
nand ( n3052 , n3000 , n3014 , n3038 , n3051 );
not ( n3053 , n182 );
and ( n3054 , n3052 , n3053 );
not ( n3055 , n3052 );
and ( n3056 , n3055 , n182 );
nor ( n3057 , n3054 , n3056 );
and ( n3058 , n2988 , n3057 );
nor ( n3059 , n2987 , n3058 );
and ( n3060 , n86 , n509 );
and ( n3061 , n78 , n199 );
nor ( n3062 , n3060 , n3061 );
and ( n3063 , n939 , n3062 );
not ( n3064 , n939 );
xor ( n3065 , n139 , n236 );
xor ( n3066 , n140 , n251 );
nand ( n3067 , n3065 , n3066 );
xor ( n3068 , n141 , n239 );
buf ( n3069 , n3068 );
nor ( n3070 , n3067 , n3069 );
not ( n3071 , n3070 );
not ( n3072 , n3071 );
xor ( n3073 , n143 , n244 );
buf ( n3074 , n3073 );
not ( n3075 , n3074 );
not ( n3076 , n3075 );
and ( n3077 , n144 , n254 );
not ( n3078 , n144 );
not ( n3079 , n254 );
and ( n3080 , n3078 , n3079 );
nor ( n3081 , n3077 , n3080 );
buf ( n3082 , n3081 );
buf ( n3083 , n3082 );
not ( n3084 , n3083 );
xor ( n3085 , n142 , n233 );
not ( n3086 , n3085 );
buf ( n3087 , n3086 );
not ( n3088 , n3087 );
nand ( n3089 , n3072 , n3076 , n3084 , n3088 );
not ( n3090 , n3089 );
buf ( n3091 , n3074 );
not ( n3092 , n3091 );
not ( n3093 , n3092 );
buf ( n3094 , n3082 );
not ( n3095 , n3070 );
not ( n3096 , n3085 );
not ( n3097 , n3096 );
nor ( n3098 , n3095 , n3097 );
nand ( n3099 , n3094 , n3098 );
nor ( n3100 , n3093 , n3099 );
nor ( n3101 , n3090 , n3100 );
buf ( n3102 , n3074 );
not ( n3103 , n3102 );
not ( n3104 , n3103 );
not ( n3105 , n3082 );
not ( n3106 , n3069 );
nor ( n3107 , n3106 , n3067 );
nand ( n3108 , n3086 , n3107 );
nor ( n3109 , n3105 , n3108 );
nand ( n3110 , n3104 , n3109 );
not ( n3111 , n3110 );
not ( n3112 , n3085 );
nor ( n3113 , n3065 , n3066 );
nand ( n3114 , n3069 , n3113 );
nor ( n3115 , n3112 , n3114 );
nand ( n3116 , n3094 , n3115 );
nor ( n3117 , n3092 , n3116 );
nor ( n3118 , n3111 , n3117 );
not ( n3119 , n3067 );
not ( n3120 , n3069 );
not ( n3121 , n3120 );
nand ( n3122 , n3119 , n3083 , n3097 , n3121 );
buf ( n3123 , n3074 );
not ( n3124 , n3123 );
nor ( n3125 , n3122 , n3124 );
not ( n3126 , n3082 );
not ( n3127 , n3085 );
nand ( n3128 , n3126 , n3127 , n3070 );
xor ( n3129 , n140 , n251 );
not ( n3130 , n3129 );
nand ( n3131 , n3082 , n3130 );
not ( n3132 , n3131 );
not ( n3133 , n3112 );
xor ( n3134 , n139 , n236 );
not ( n3135 , n3134 );
not ( n3136 , n3135 );
and ( n3137 , n3136 , n3069 );
not ( n3138 , n3137 );
or ( n3139 , n3133 , n3138 );
not ( n3140 , n3136 );
nand ( n3141 , n3140 , n3085 , n3120 );
nand ( n3142 , n3139 , n3141 );
nand ( n3143 , n3132 , n3142 );
and ( n3144 , n3128 , n3143 );
not ( n3145 , n3102 );
not ( n3146 , n3145 );
not ( n3147 , n3146 );
nor ( n3148 , n3144 , n3147 );
nor ( n3149 , n3125 , n3148 );
and ( n3150 , n3101 , n3118 , n3149 );
not ( n3151 , n3082 );
not ( n3152 , n3151 );
not ( n3153 , n3152 );
nand ( n3154 , n3097 , n3070 );
nor ( n3155 , n3123 , n3154 );
not ( n3156 , n3155 );
or ( n3157 , n3153 , n3156 );
not ( n3158 , n3120 );
not ( n3159 , n3065 );
nor ( n3160 , n3159 , n3066 );
nand ( n3161 , n3158 , n3160 );
not ( n3162 , n3085 );
nor ( n3163 , n3161 , n3162 );
nand ( n3164 , n3152 , n3103 , n3163 );
nand ( n3165 , n3157 , n3164 );
not ( n3166 , n3071 );
nor ( n3167 , n3074 , n3082 );
nand ( n3168 , n3166 , n3167 , n3087 );
not ( n3169 , n3073 );
not ( n3170 , n3169 );
not ( n3171 , n3170 );
not ( n3172 , n3069 );
nand ( n3173 , n3172 , n3160 );
nor ( n3174 , n3127 , n3173 );
nand ( n3175 , n3171 , n3084 , n3174 );
nand ( n3176 , n3168 , n3175 );
nor ( n3177 , n3165 , n3176 );
not ( n3178 , n3082 );
not ( n3179 , n3178 );
not ( n3180 , n3068 );
nand ( n3181 , n3180 , n3129 , n3135 );
nor ( n3182 , n3162 , n3181 );
nand ( n3183 , n3179 , n3170 , n3182 );
not ( n3184 , n3183 );
and ( n3185 , n3068 , n3129 , n3135 );
not ( n3186 , n3185 );
nor ( n3187 , n3162 , n3186 );
nand ( n3188 , n3084 , n3102 , n3187 );
not ( n3189 , n3188 );
nor ( n3190 , n3184 , n3189 );
not ( n3191 , n3107 );
nor ( n3192 , n3086 , n3191 );
and ( n3193 , n3103 , n3084 , n3192 );
not ( n3194 , n3082 );
not ( n3195 , n3085 );
not ( n3196 , n3195 );
not ( n3197 , n3135 );
nor ( n3198 , n3197 , n3129 );
nand ( n3199 , n3194 , n3196 , n3172 , n3198 );
not ( n3200 , n3199 );
not ( n3201 , n3170 );
nand ( n3202 , n3200 , n3201 );
not ( n3203 , n3202 );
nor ( n3204 , n3193 , n3203 );
nor ( n3205 , n3169 , n3085 );
not ( n3206 , n3161 );
nand ( n3207 , n3205 , n3126 , n3206 );
not ( n3208 , n3178 );
not ( n3209 , n3195 );
nor ( n3210 , n3209 , n3114 );
nand ( n3211 , n3208 , n3075 , n3210 );
not ( n3212 , n3211 );
not ( n3213 , n3212 );
nand ( n3214 , n3190 , n3204 , n3207 , n3213 );
not ( n3215 , n3171 );
nand ( n3216 , n3152 , n3187 );
or ( n3217 , n3215 , n3216 );
and ( n3218 , n3082 , n3096 , n3172 , n3198 );
nand ( n3219 , n3104 , n3218 );
nand ( n3220 , n3217 , n3219 );
nor ( n3221 , n3214 , n3220 );
not ( n3222 , n3082 );
nand ( n3223 , n3222 , n3163 );
nor ( n3224 , n3215 , n3223 );
not ( n3225 , n3145 );
not ( n3226 , n3218 );
nor ( n3227 , n3225 , n3226 );
nor ( n3228 , n3224 , n3227 );
not ( n3229 , n3091 );
nor ( n3230 , n3229 , n3223 );
not ( n3231 , n3123 );
nand ( n3232 , n3105 , n3115 );
nor ( n3233 , n3231 , n3232 );
nor ( n3234 , n3230 , n3233 );
not ( n3235 , n3082 );
nand ( n3236 , n3112 , n3185 );
nor ( n3237 , n3235 , n3236 );
nand ( n3238 , n3201 , n3237 );
not ( n3239 , n3238 );
not ( n3240 , n3160 );
not ( n3241 , n3240 );
not ( n3242 , n3096 );
not ( n3243 , n3121 );
nand ( n3244 , n3241 , n3082 , n3242 , n3243 );
nor ( n3245 , n3104 , n3244 );
nor ( n3246 , n3239 , n3245 );
nand ( n3247 , n3228 , n3234 , n3246 );
nor ( n3248 , n3074 , n3082 );
not ( n3249 , n3236 );
nand ( n3250 , n3248 , n3249 );
not ( n3251 , n3250 );
not ( n3252 , n3114 );
and ( n3253 , n3151 , n3127 , n3252 );
not ( n3254 , n3253 );
nor ( n3255 , n3254 , n3229 );
nor ( n3256 , n3251 , n3255 );
nand ( n3257 , n3084 , n3091 , n3182 );
nor ( n3258 , n3173 , n3209 );
nand ( n3259 , n3094 , n3091 , n3258 );
nand ( n3260 , n3257 , n3259 );
nor ( n3261 , n3242 , n3181 );
nand ( n3262 , n3222 , n3091 , n3261 );
xor ( n3263 , n143 , n244 );
nor ( n3264 , n3065 , n3263 );
nand ( n3265 , n3129 , n3180 , n3264 );
not ( n3266 , n3265 );
nand ( n3267 , n3087 , n3105 , n3266 );
nand ( n3268 , n3262 , n3267 );
nor ( n3269 , n3260 , n3268 );
nand ( n3270 , n3256 , n3269 );
nor ( n3271 , n3247 , n3270 );
nand ( n3272 , n3150 , n3177 , n3221 , n3271 );
not ( n3273 , n177 );
and ( n3274 , n3272 , n3273 );
not ( n3275 , n3272 );
and ( n3276 , n3275 , n177 );
nor ( n3277 , n3274 , n3276 );
and ( n3278 , n3064 , n3277 );
nor ( n3279 , n3063 , n3278 );
and ( n3280 , n88 , n509 );
and ( n3281 , n80 , n199 );
nor ( n3282 , n3280 , n3281 );
and ( n3283 , n1553 , n3282 );
not ( n3284 , n1553 );
nand ( n3285 , n3231 , n3253 );
or ( n3286 , n3130 , n3082 );
nand ( n3287 , n3286 , n3131 );
nand ( n3288 , n3287 , n3092 , n3142 );
nand ( n3289 , n3285 , n3288 );
not ( n3290 , n3244 );
nand ( n3291 , n3225 , n3290 );
nand ( n3292 , n3250 , n3110 , n3291 );
nor ( n3293 , n3289 , n3292 );
nor ( n3294 , n3176 , n3255 );
not ( n3295 , n3199 );
nand ( n3296 , n3295 , n3076 );
nand ( n3297 , n3257 , n3296 );
nor ( n3298 , n3093 , n3232 );
not ( n3299 , n3171 );
nand ( n3300 , n3084 , n3258 );
or ( n3301 , n3299 , n3300 );
nand ( n3302 , n3301 , n3188 );
nor ( n3303 , n3297 , n3298 , n3302 );
and ( n3304 , n3293 , n3294 , n3303 );
not ( n3305 , n3146 );
nor ( n3306 , n3305 , n3216 );
not ( n3307 , n3164 );
or ( n3308 , n3306 , n3307 );
not ( n3309 , n3122 );
nand ( n3310 , n3231 , n3309 );
not ( n3311 , n3310 );
nor ( n3312 , n3311 , n3100 );
not ( n3313 , n3237 );
nor ( n3314 , n3124 , n3313 );
nor ( n3315 , n3314 , n3117 );
nor ( n3316 , n3124 , n3099 );
not ( n3317 , n3316 );
nand ( n3318 , n3312 , n3315 , n3317 , n3259 );
nor ( n3319 , n3308 , n3318 );
not ( n3320 , n3220 );
not ( n3321 , n3108 );
nand ( n3322 , n3321 , n3091 , n3222 );
not ( n3323 , n3322 );
not ( n3324 , n3089 );
nor ( n3325 , n3323 , n3324 );
nand ( n3326 , n3179 , n3171 , n3261 );
nand ( n3327 , n3326 , n3211 );
not ( n3328 , n3327 );
nand ( n3329 , n3320 , n3325 , n3328 );
nor ( n3330 , n3229 , n3300 );
or ( n3331 , n3230 , n3330 );
nor ( n3332 , n3329 , n3331 );
nand ( n3333 , n3304 , n3319 , n3332 );
not ( n3334 , n185 );
and ( n3335 , n3333 , n3334 );
not ( n3336 , n3333 );
and ( n3337 , n3336 , n185 );
nor ( n3338 , n3335 , n3337 );
and ( n3339 , n3284 , n3338 );
nor ( n3340 , n3283 , n3339 );
and ( n3341 , n94 , n509 );
and ( n3342 , n86 , n199 );
nor ( n3343 , n3341 , n3342 );
and ( n3344 , n1553 , n3343 );
not ( n3345 , n1553 );
nand ( n3346 , n2386 , n2785 );
not ( n3347 , n3346 );
and ( n3348 , n2459 , n2367 );
and ( n3349 , n2375 , n2452 );
nand ( n3350 , n3347 , n3348 , n3349 );
nor ( n3351 , n2493 , n3350 );
not ( n3352 , n2403 );
nor ( n3353 , n2794 , n3352 );
nand ( n3354 , n2807 , n2792 );
not ( n3355 , n3354 );
nor ( n3356 , n2479 , n2480 );
nor ( n3357 , n3355 , n3356 );
nand ( n3358 , n2417 , n2808 );
not ( n3359 , n3358 );
not ( n3360 , n2759 );
nor ( n3361 , n3359 , n3360 );
and ( n3362 , n3353 , n3357 , n3361 );
not ( n3363 , n2807 );
not ( n3364 , n2402 );
or ( n3365 , n3363 , n3364 );
nand ( n3366 , n3365 , n2398 );
nor ( n3367 , n2425 , n3366 );
nand ( n3368 , n2815 , n2762 );
nand ( n3369 , n2498 , n2445 );
not ( n3370 , n3369 );
and ( n3371 , n2471 , n2756 );
not ( n3372 , n2457 );
nand ( n3373 , n2362 , n2329 , n3372 );
nand ( n3374 , n2361 , n2765 , n2328 );
and ( n3375 , n3373 , n3374 );
or ( n3376 , n2771 , n2775 );
nand ( n3377 , n3376 , n2406 );
nor ( n3378 , n3375 , n3377 );
nor ( n3379 , n2804 , n3378 );
nand ( n3380 , n3370 , n2809 , n3371 , n3379 );
nor ( n3381 , n3368 , n3380 );
nand ( n3382 , n3351 , n3362 , n3367 , n3381 );
not ( n3383 , n176 );
and ( n3384 , n3382 , n3383 );
not ( n3385 , n3382 );
and ( n3386 , n3385 , n176 );
nor ( n3387 , n3384 , n3386 );
and ( n3388 , n3345 , n3387 );
nor ( n3389 , n3344 , n3388 );
and ( n3390 , n98 , n509 );
and ( n3391 , n90 , n199 );
nor ( n3392 , n3390 , n3391 );
and ( n3393 , n939 , n3392 );
not ( n3394 , n939 );
not ( n3395 , n3285 );
not ( n3396 , n3395 );
and ( n3397 , n3120 , n3113 );
nand ( n3398 , n3397 , n3235 , n3127 , n3075 );
not ( n3399 , n3398 );
nor ( n3400 , n3125 , n3399 );
not ( n3401 , n3264 );
not ( n3402 , n3135 );
nand ( n3403 , n3402 , n3073 );
nand ( n3404 , n3401 , n3403 );
nor ( n3405 , n3120 , n3130 );
nand ( n3406 , n3404 , n3126 , n3405 );
or ( n3407 , n3129 , n3180 , n3403 );
nand ( n3408 , n3407 , n3265 );
nand ( n3409 , n3179 , n3408 );
nand ( n3410 , n3406 , n3409 );
nand ( n3411 , n3088 , n3410 );
nand ( n3412 , n3396 , n3400 , n3317 , n3411 );
not ( n3413 , n3296 );
nor ( n3414 , n3413 , n3302 );
and ( n3415 , n3168 , n3262 );
nand ( n3416 , n3126 , n3097 , n3070 );
nor ( n3417 , n3093 , n3416 );
nand ( n3418 , n3250 , n3202 );
nor ( n3419 , n3417 , n3418 );
nand ( n3420 , n3414 , n3415 , n3419 );
nor ( n3421 , n3412 , n3420 );
not ( n3422 , n3310 );
nor ( n3423 , n3422 , n3314 );
nor ( n3424 , n3307 , n3245 );
nand ( n3425 , n3124 , n3109 );
not ( n3426 , n3117 );
nand ( n3427 , n3423 , n3424 , n3425 , n3426 );
nand ( n3428 , n3183 , n3259 );
nor ( n3429 , n3427 , n3428 );
nand ( n3430 , n3207 , n3326 );
nor ( n3431 , n3224 , n3227 );
nor ( n3432 , n3299 , n3116 );
nor ( n3433 , n3432 , n3212 );
not ( n3434 , n3324 );
nand ( n3435 , n3431 , n3433 , n3322 , n3434 );
nor ( n3436 , n3430 , n3435 );
nand ( n3437 , n3421 , n3429 , n3436 );
not ( n3438 , n192 );
and ( n3439 , n3437 , n3438 );
not ( n3440 , n3437 );
and ( n3441 , n3440 , n192 );
nor ( n3442 , n3439 , n3441 );
and ( n3443 , n3394 , n3442 );
nor ( n3444 , n3393 , n3443 );
and ( n3445 , n100 , n509 );
and ( n3446 , n92 , n199 );
nor ( n3447 , n3445 , n3446 );
and ( n3448 , n939 , n3447 );
not ( n3449 , n939 );
and ( n3450 , n3170 , n3405 );
not ( n3451 , n3152 );
and ( n3452 , n3450 , n3140 , n3451 );
not ( n3453 , n3169 );
not ( n3454 , n3137 );
or ( n3455 , n3453 , n3454 );
nand ( n3456 , n3455 , n3235 );
nand ( n3457 , n3130 , n3456 );
nand ( n3458 , n3068 , n3263 );
or ( n3459 , n3136 , n3458 );
not ( n3460 , n3073 );
nand ( n3461 , n3136 , n3180 , n3460 );
nand ( n3462 , n3459 , n3461 );
nor ( n3463 , n3126 , n3462 );
nor ( n3464 , n3457 , n3463 );
nor ( n3465 , n3452 , n3464 );
or ( n3466 , n3465 , n3088 );
not ( n3467 , n3165 );
nand ( n3468 , n3466 , n3467 );
not ( n3469 , n3468 );
not ( n3470 , n3291 );
not ( n3471 , n3219 );
nor ( n3472 , n3470 , n3471 );
not ( n3473 , n3425 );
nor ( n3474 , n3473 , n3330 );
nor ( n3475 , n3432 , n3298 );
nand ( n3476 , n3472 , n3474 , n3475 );
nor ( n3477 , n3306 , n3233 );
and ( n3478 , n3168 , n3250 );
not ( n3479 , n3417 );
nand ( n3480 , n3477 , n3478 , n3479 , n3262 );
nor ( n3481 , n3476 , n3480 );
nor ( n3482 , n3297 , n3327 );
not ( n3483 , n3238 );
nor ( n3484 , n3483 , n3316 );
nor ( n3485 , n3125 , n3111 );
nand ( n3486 , n3482 , n3484 , n3485 );
nand ( n3487 , n3322 , n3175 );
nand ( n3488 , n3183 , n3398 );
nor ( n3489 , n3487 , n3488 );
not ( n3490 , n3193 );
nand ( n3491 , n3489 , n3490 , n3207 );
nor ( n3492 , n3486 , n3491 );
nand ( n3493 , n3469 , n3481 , n3492 );
not ( n3494 , n167 );
and ( n3495 , n3493 , n3494 );
not ( n3496 , n3493 );
and ( n3497 , n3496 , n167 );
nor ( n3498 , n3495 , n3497 );
and ( n3499 , n3449 , n3498 );
nor ( n3500 , n3448 , n3499 );
and ( n3501 , n130 , n509 );
and ( n3502 , n122 , n199 );
nor ( n3503 , n3501 , n3502 );
and ( n3504 , n939 , n3503 );
not ( n3505 , n939 );
not ( n3506 , n188 );
nand ( n3507 , n2114 , n2197 , n3017 );
nand ( n3508 , n3507 , n2192 );
not ( n3509 , n3508 );
and ( n3510 , n2294 , n2204 );
nor ( n3511 , n3510 , n2152 );
nand ( n3512 , n3509 , n3511 );
and ( n3513 , n3001 , n2166 );
nand ( n3514 , n2142 , n3513 );
nor ( n3515 , n3512 , n3514 );
not ( n3516 , n3010 );
and ( n3517 , n2224 , n3516 );
nor ( n3518 , n2289 , n2207 );
not ( n3519 , n2227 );
nor ( n3520 , n3518 , n3519 );
and ( n3521 , n2997 , n2233 );
and ( n3522 , n3520 , n3521 , n2990 , n2201 );
nand ( n3523 , n3515 , n3517 , n3522 );
not ( n3524 , n2262 );
nand ( n3525 , n3524 , n2267 );
nand ( n3526 , n3525 , n2173 , n2251 , n2143 );
nand ( n3527 , n2243 , n3526 );
not ( n3528 , n3527 );
nand ( n3529 , n2250 , n2148 );
nand ( n3530 , n2135 , n3015 );
not ( n3531 , n3530 );
not ( n3532 , n2120 );
and ( n3533 , n3531 , n3532 );
not ( n3534 , n2135 );
nand ( n3535 , n3534 , n2154 );
not ( n3536 , n3535 );
and ( n3537 , n3536 , n2159 );
nor ( n3538 , n3533 , n3537 );
nor ( n3539 , n3529 , n2114 , n3538 );
nor ( n3540 , n3019 , n3539 );
and ( n3541 , n3528 , n3540 , n2240 , n2279 );
nor ( n3542 , n3045 , n3040 );
nand ( n3543 , n2210 , n2276 );
and ( n3544 , n3543 , n2297 , n2303 );
nand ( n3545 , n3541 , n3050 , n3542 , n3544 );
nor ( n3546 , n3523 , n3545 );
not ( n3547 , n3546 );
and ( n3548 , n3506 , n3547 );
and ( n3549 , n188 , n3546 );
nor ( n3550 , n3548 , n3549 );
and ( n3551 , n3505 , n3550 );
nor ( n3552 , n3504 , n3551 );
not ( n3553 , n45 );
and ( n3554 , n1552 , n3553 );
not ( n3555 , n1552 );
and ( n3556 , n3555 , n3498 );
nor ( n3557 , n3554 , n3556 );
not ( n3558 , n39 );
and ( n3559 , n1205 , n3558 );
not ( n3560 , n1205 );
and ( n3561 , n3560 , n3387 );
nor ( n3562 , n3559 , n3561 );
not ( n3563 , n31 );
and ( n3564 , n1205 , n3563 );
not ( n3565 , n1205 );
and ( n3566 , n3565 , n3277 );
nor ( n3567 , n3564 , n3566 );
not ( n3568 , n57 );
and ( n3569 , n1552 , n3568 );
not ( n3570 , n1552 );
and ( n3571 , n3570 , n3057 );
nor ( n3572 , n3569 , n3571 );
not ( n3573 , n33 );
and ( n3574 , n1205 , n3573 );
not ( n3575 , n1205 );
and ( n3576 , n3575 , n3338 );
nor ( n3577 , n3574 , n3576 );
not ( n3578 , n8 );
and ( n3579 , n1205 , n3578 );
not ( n3580 , n1205 );
and ( n3581 , n3580 , n3550 );
nor ( n3582 , n3579 , n3581 );
not ( n3583 , n59 );
and ( n3584 , n1217 , n3583 );
not ( n3585 , n1217 );
and ( n3586 , n3585 , n2981 );
nor ( n3587 , n3584 , n3586 );
not ( n3588 , n43 );
and ( n3589 , n1552 , n3588 );
not ( n3590 , n1552 );
and ( n3591 , n3590 , n3442 );
nor ( n3592 , n3589 , n3591 );
and ( n3593 , n76 , n509 );
and ( n3594 , n68 , n199 );
nor ( n3595 , n3593 , n3594 );
and ( n3596 , n939 , n3595 );
not ( n3597 , n939 );
not ( n3598 , n3374 );
nand ( n3599 , n2365 , n2440 , n2323 , n3598 );
nand ( n3600 , n3599 , n2752 , n2367 );
not ( n3601 , n2761 );
not ( n3602 , n2355 );
not ( n3603 , n2371 );
nand ( n3604 , n2399 , n3602 , n3603 );
and ( n3605 , n2334 , n2325 );
nand ( n3606 , n3605 , n2356 );
nand ( n3607 , n3604 , n3606 );
nand ( n3608 , n2780 , n3607 );
nand ( n3609 , n2375 , n3601 , n3608 );
nor ( n3610 , n3600 , n3609 );
nand ( n3611 , n3354 , n2419 );
nor ( n3612 , n3611 , n2436 );
nor ( n3613 , n3366 , n2757 );
and ( n3614 , n3610 , n3612 , n3613 );
nand ( n3615 , n2492 , n2489 );
not ( n3616 , n3356 );
nand ( n3617 , n2805 , n3616 , n2501 );
nor ( n3618 , n3615 , n3617 );
not ( n3619 , n2453 );
nand ( n3620 , n2813 , n3619 );
nand ( n3621 , n2467 , n2789 );
nand ( n3622 , n3358 , n2796 , n2463 );
nor ( n3623 , n3620 , n3621 , n3622 );
nand ( n3624 , n3614 , n3618 , n3623 );
not ( n3625 , n170 );
and ( n3626 , n3624 , n3625 );
not ( n3627 , n3624 );
and ( n3628 , n3627 , n170 );
nor ( n3629 , n3626 , n3628 );
and ( n3630 , n3597 , n3629 );
nor ( n3631 , n3596 , n3630 );
and ( n3632 , n90 , n509 );
and ( n3633 , n82 , n199 );
nor ( n3634 , n3632 , n3633 );
and ( n3635 , n1223 , n3634 );
not ( n3636 , n1223 );
not ( n3637 , n2247 );
and ( n3638 , n2242 , n3637 );
not ( n3639 , n3518 );
nand ( n3640 , n3639 , n2995 );
not ( n3641 , n2266 );
nand ( n3642 , n3641 , n2261 );
nand ( n3643 , n2250 , n2206 , n2117 , n3642 );
nor ( n3644 , n2133 , n2264 );
and ( n3645 , n2159 , n3530 );
not ( n3646 , n2159 );
and ( n3647 , n3646 , n3535 );
nor ( n3648 , n3645 , n3647 );
nand ( n3649 , n3644 , n3648 );
and ( n3650 , n3643 , n3649 );
nor ( n3651 , n3650 , n2143 );
nor ( n3652 , n3640 , n3651 );
nand ( n3653 , n3638 , n3652 );
not ( n3654 , n2298 );
nor ( n3655 , n3022 , n3049 );
not ( n3656 , n3543 );
nor ( n3657 , n3656 , n2287 );
nand ( n3658 , n3654 , n3655 , n2279 , n3657 );
nor ( n3659 , n3653 , n3658 );
nor ( n3660 , n3006 , n3508 );
not ( n3661 , n2215 );
not ( n3662 , n2233 );
nor ( n3663 , n3661 , n3662 );
not ( n3664 , n2208 );
not ( n3665 , n2227 );
nor ( n3666 , n3665 , n2991 );
nand ( n3667 , n3660 , n3663 , n3664 , n3666 );
and ( n3668 , n2141 , n2187 );
nand ( n3669 , n3668 , n3046 , n3511 , n3004 );
nor ( n3670 , n3667 , n3669 );
nand ( n3671 , n3659 , n3670 );
not ( n3672 , n193 );
and ( n3673 , n3671 , n3672 );
not ( n3674 , n3671 );
and ( n3675 , n3674 , n193 );
nor ( n3676 , n3673 , n3675 );
and ( n3677 , n3636 , n3676 );
nor ( n3678 , n3635 , n3677 );
not ( n3679 , n21 );
and ( n3680 , n2930 , n3679 );
not ( n3681 , n2930 );
and ( n3682 , n3681 , n3629 );
nor ( n3683 , n3680 , n3682 );
not ( n3684 , n35 );
and ( n3685 , n2004 , n3684 );
not ( n3686 , n2004 );
and ( n3687 , n3686 , n3676 );
nor ( n3688 , n3685 , n3687 );
not ( n3689 , n9 );
buf ( n3690 , n3689 );
not ( n3691 , n10 );
and ( n3692 , n24 , n3691 );
and ( n3693 , n10 , n32 );
nor ( n3694 , n3692 , n3693 );
nand ( n3695 , n11 , n504 );
buf ( n3696 , n3695 );
not ( n3697 , n3696 );
not ( n3698 , n3697 );
or ( n3699 , n3694 , n3698 );
nand ( n3700 , n198 , n196 , n197 );
and ( n3701 , n10 , n256 );
not ( n3702 , n10 );
not ( n3703 , n256 );
and ( n3704 , n3702 , n3703 );
nor ( n3705 , n3701 , n3704 );
nand ( n3706 , n199 , n3705 );
or ( n3707 , n3700 , n3706 );
not ( n3708 , n3707 );
not ( n3709 , n3708 );
or ( n3710 , n202 , n3709 );
buf ( n3711 , n3695 );
nand ( n3712 , n3710 , n3711 );
not ( n3713 , n3712 );
buf ( n3714 , n3707 );
buf ( n3715 , n3714 );
not ( n3716 , n200 );
not ( n3717 , n197 );
nor ( n3718 , n196 , n199 );
nand ( n3719 , n3717 , n3718 );
or ( n3720 , n198 , n3719 );
nand ( n3721 , n197 , n198 );
or ( n3722 , n3721 , n3718 );
nand ( n3723 , n3720 , n3722 );
buf ( n3724 , n3723 );
buf ( n3725 , n3724 );
nor ( n3726 , n3716 , n3725 );
not ( n3727 , n3726 );
buf ( n3728 , n3723 );
buf ( n3729 , n3728 );
nand ( n3730 , n201 , n3729 );
nand ( n3731 , n3727 , n3730 );
nand ( n3732 , n256 , n3731 );
not ( n3733 , n256 );
not ( n3734 , n204 );
buf ( n3735 , n3724 );
nor ( n3736 , n3734 , n3735 );
not ( n3737 , n3736 );
buf ( n3738 , n3728 );
nand ( n3739 , n203 , n3738 );
nand ( n3740 , n3737 , n3739 );
nand ( n3741 , n3733 , n3740 );
nand ( n3742 , n3715 , n3732 , n3741 );
nand ( n3743 , n3713 , n3742 );
nand ( n3744 , n3699 , n3743 );
and ( n3745 , n3690 , n3744 );
and ( n3746 , n59 , n3691 );
and ( n3747 , n10 , n67 );
nor ( n3748 , n3746 , n3747 );
not ( n3749 , n3696 );
not ( n3750 , n3749 );
or ( n3751 , n3748 , n3750 );
not ( n3752 , n3707 );
not ( n3753 , n3752 );
or ( n3754 , n222 , n3753 );
nand ( n3755 , n3754 , n3696 );
not ( n3756 , n3755 );
buf ( n3757 , n3714 );
not ( n3758 , n220 );
nor ( n3759 , n3758 , n3725 );
not ( n3760 , n3759 );
buf ( n3761 , n3728 );
nand ( n3762 , n221 , n3761 );
nand ( n3763 , n3760 , n3762 );
nand ( n3764 , n256 , n3763 );
not ( n3765 , n256 );
not ( n3766 , n224 );
nor ( n3767 , n3766 , n3725 );
not ( n3768 , n3767 );
buf ( n3769 , n3728 );
nand ( n3770 , n223 , n3769 );
nand ( n3771 , n3768 , n3770 );
nand ( n3772 , n3765 , n3771 );
nand ( n3773 , n3757 , n3764 , n3772 );
nand ( n3774 , n3756 , n3773 );
nand ( n3775 , n3751 , n3774 );
and ( n3776 , n3690 , n3775 );
and ( n3777 , n17 , n3691 );
and ( n3778 , n10 , n25 );
nor ( n3779 , n3777 , n3778 );
not ( n3780 , n3696 );
not ( n3781 , n3780 );
or ( n3782 , n3779 , n3781 );
or ( n3783 , n211 , n3753 );
nand ( n3784 , n3783 , n3711 );
not ( n3785 , n3784 );
buf ( n3786 , n3714 );
not ( n3787 , n209 );
buf ( n3788 , n3728 );
nor ( n3789 , n3787 , n3788 );
not ( n3790 , n3789 );
nand ( n3791 , n210 , n3761 );
nand ( n3792 , n3790 , n3791 );
nand ( n3793 , n256 , n3792 );
not ( n3794 , n256 );
not ( n3795 , n213 );
nor ( n3796 , n3795 , n3735 );
not ( n3797 , n3796 );
nand ( n3798 , n212 , n3738 );
nand ( n3799 , n3797 , n3798 );
nand ( n3800 , n3794 , n3799 );
nand ( n3801 , n3786 , n3793 , n3800 );
nand ( n3802 , n3785 , n3801 );
nand ( n3803 , n3782 , n3802 );
and ( n3804 , n3690 , n3803 );
and ( n3805 , n46 , n3691 );
and ( n3806 , n10 , n54 );
nor ( n3807 , n3805 , n3806 );
not ( n3808 , n3697 );
or ( n3809 , n3807 , n3808 );
not ( n3810 , n3708 );
or ( n3811 , n243 , n3810 );
nand ( n3812 , n3811 , n3696 );
not ( n3813 , n3812 );
buf ( n3814 , n3714 );
not ( n3815 , n241 );
buf ( n3816 , n3728 );
nor ( n3817 , n3815 , n3816 );
not ( n3818 , n3817 );
buf ( n3819 , n242 );
buf ( n3820 , n3819 );
nand ( n3821 , n3820 , n3729 );
nand ( n3822 , n3818 , n3821 );
nand ( n3823 , n256 , n3822 );
not ( n3824 , n256 );
not ( n3825 , n245 );
nor ( n3826 , n3825 , n3788 );
not ( n3827 , n3826 );
nand ( n3828 , n244 , n3769 );
nand ( n3829 , n3827 , n3828 );
nand ( n3830 , n3824 , n3829 );
nand ( n3831 , n3814 , n3823 , n3830 );
nand ( n3832 , n3813 , n3831 );
nand ( n3833 , n3809 , n3832 );
and ( n3834 , n3690 , n3833 );
and ( n3835 , n18 , n3691 );
and ( n3836 , n10 , n26 );
nor ( n3837 , n3835 , n3836 );
not ( n3838 , n3697 );
or ( n3839 , n3837 , n3838 );
not ( n3840 , n3752 );
or ( n3841 , n219 , n3840 );
nand ( n3842 , n3841 , n3711 );
not ( n3843 , n3842 );
not ( n3844 , n217 );
nor ( n3845 , n3844 , n3788 );
not ( n3846 , n3845 );
nand ( n3847 , n218 , n3761 );
nand ( n3848 , n3846 , n3847 );
nand ( n3849 , n256 , n3848 );
not ( n3850 , n256 );
not ( n3851 , n221 );
nor ( n3852 , n3851 , n3788 );
not ( n3853 , n3852 );
nand ( n3854 , n220 , n3738 );
nand ( n3855 , n3853 , n3854 );
nand ( n3856 , n3850 , n3855 );
nand ( n3857 , n3715 , n3849 , n3856 );
nand ( n3858 , n3843 , n3857 );
nand ( n3859 , n3839 , n3858 );
and ( n3860 , n3690 , n3859 );
and ( n3861 , n19 , n3691 );
and ( n3862 , n10 , n27 );
nor ( n3863 , n3861 , n3862 );
not ( n3864 , n3697 );
or ( n3865 , n3863 , n3864 );
or ( n3866 , n227 , n3810 );
nand ( n3867 , n3866 , n3711 );
not ( n3868 , n3867 );
not ( n3869 , n225 );
nor ( n3870 , n3869 , n3735 );
not ( n3871 , n3870 );
nand ( n3872 , n226 , n3738 );
nand ( n3873 , n3871 , n3872 );
nand ( n3874 , n256 , n3873 );
not ( n3875 , n256 );
not ( n3876 , n201 );
nor ( n3877 , n3876 , n3788 );
not ( n3878 , n3877 );
nand ( n3879 , n200 , n3729 );
nand ( n3880 , n3878 , n3879 );
nand ( n3881 , n3875 , n3880 );
nand ( n3882 , n3786 , n3874 , n3881 );
nand ( n3883 , n3868 , n3882 );
nand ( n3884 , n3865 , n3883 );
and ( n3885 , n3690 , n3884 );
and ( n3886 , n45 , n3691 );
and ( n3887 , n10 , n53 );
nor ( n3888 , n3886 , n3887 );
or ( n3889 , n3888 , n3838 );
not ( n3890 , n3707 );
not ( n3891 , n3890 );
or ( n3892 , n251 , n3891 );
nand ( n3893 , n3892 , n3711 );
not ( n3894 , n3893 );
not ( n3895 , n249 );
nor ( n3896 , n3895 , n3816 );
not ( n3897 , n3896 );
nand ( n3898 , n250 , n3761 );
nand ( n3899 , n3897 , n3898 );
nand ( n3900 , n256 , n3899 );
not ( n3901 , n256 );
not ( n3902 , n253 );
nor ( n3903 , n3902 , n3788 );
not ( n3904 , n3903 );
nand ( n3905 , n252 , n3761 );
nand ( n3906 , n3904 , n3905 );
nand ( n3907 , n3901 , n3906 );
nand ( n3908 , n3715 , n3900 , n3907 );
nand ( n3909 , n3894 , n3908 );
nand ( n3910 , n3889 , n3909 );
and ( n3911 , n3690 , n3910 );
and ( n3912 , n50 , n3691 );
and ( n3913 , n10 , n58 );
nor ( n3914 , n3912 , n3913 );
or ( n3915 , n3914 , n3808 );
not ( n3916 , n3707 );
not ( n3917 , n3916 );
or ( n3918 , n215 , n3917 );
nand ( n3919 , n3918 , n3711 );
not ( n3920 , n3919 );
not ( n3921 , n3796 );
nand ( n3922 , n214 , n3761 );
nand ( n3923 , n3921 , n3922 );
nand ( n3924 , n256 , n3923 );
not ( n3925 , n256 );
not ( n3926 , n3845 );
nand ( n3927 , n216 , n3729 );
nand ( n3928 , n3926 , n3927 );
nand ( n3929 , n3925 , n3928 );
nand ( n3930 , n3715 , n3924 , n3929 );
nand ( n3931 , n3920 , n3930 );
nand ( n3932 , n3915 , n3931 );
and ( n3933 , n3690 , n3932 );
and ( n3934 , n14 , n3691 );
and ( n3935 , n10 , n22 );
nor ( n3936 , n3934 , n3935 );
not ( n3937 , n3780 );
or ( n3938 , n3936 , n3937 );
not ( n3939 , n3916 );
or ( n3940 , n247 , n3939 );
nand ( n3941 , n3940 , n3696 );
not ( n3942 , n3941 );
not ( n3943 , n3826 );
nand ( n3944 , n246 , n3729 );
nand ( n3945 , n3943 , n3944 );
nand ( n3946 , n256 , n3945 );
not ( n3947 , n256 );
not ( n3948 , n3896 );
nand ( n3949 , n248 , n3761 );
nand ( n3950 , n3948 , n3949 );
nand ( n3951 , n3947 , n3950 );
nand ( n3952 , n3814 , n3946 , n3951 );
nand ( n3953 , n3942 , n3952 );
nand ( n3954 , n3938 , n3953 );
and ( n3955 , n3690 , n3954 );
and ( n3956 , n48 , n3691 );
and ( n3957 , n10 , n56 );
nor ( n3958 , n3956 , n3957 );
not ( n3959 , n3780 );
or ( n3960 , n3958 , n3959 );
or ( n3961 , n231 , n3891 );
nand ( n3962 , n3961 , n3711 );
not ( n3963 , n3962 );
not ( n3964 , n229 );
nor ( n3965 , n3964 , n3788 );
not ( n3966 , n3965 );
nand ( n3967 , n230 , n3761 );
nand ( n3968 , n3966 , n3967 );
nand ( n3969 , n256 , n3968 );
not ( n3970 , n256 );
not ( n3971 , n233 );
nor ( n3972 , n3971 , n3788 );
not ( n3973 , n3972 );
nand ( n3974 , n232 , n3738 );
nand ( n3975 , n3973 , n3974 );
nand ( n3976 , n3970 , n3975 );
nand ( n3977 , n3786 , n3969 , n3976 );
nand ( n3978 , n3963 , n3977 );
nand ( n3979 , n3960 , n3978 );
and ( n3980 , n3690 , n3979 );
and ( n3981 , n47 , n3691 );
and ( n3982 , n10 , n55 );
nor ( n3983 , n3981 , n3982 );
not ( n3984 , n3780 );
or ( n3985 , n3983 , n3984 );
not ( n3986 , n3890 );
or ( n3987 , n235 , n3986 );
nand ( n3988 , n3987 , n3696 );
not ( n3989 , n3988 );
not ( n3990 , n3972 );
nand ( n3991 , n234 , n3738 );
nand ( n3992 , n3990 , n3991 );
nand ( n3993 , n256 , n3992 );
not ( n3994 , n256 );
not ( n3995 , n237 );
nor ( n3996 , n3995 , n3788 );
not ( n3997 , n3996 );
nand ( n3998 , n236 , n3738 );
nand ( n3999 , n3997 , n3998 );
nand ( n4000 , n3994 , n3999 );
nand ( n4001 , n3814 , n3993 , n4000 );
nand ( n4002 , n3989 , n4001 );
nand ( n4003 , n3985 , n4002 );
and ( n4004 , n3690 , n4003 );
and ( n4005 , n40 , n3691 );
and ( n4006 , n10 , n19 );
nor ( n4007 , n4005 , n4006 );
not ( n4008 , n3749 );
or ( n4009 , n4007 , n4008 );
not ( n4010 , n3708 );
or ( n4011 , n200 , n4010 );
nand ( n4012 , n4011 , n3711 );
not ( n4013 , n4012 );
buf ( n4014 , n3714 );
not ( n4015 , n226 );
nor ( n4016 , n4015 , n3788 );
not ( n4017 , n4016 );
nand ( n4018 , n227 , n3729 );
nand ( n4019 , n4017 , n4018 );
nand ( n4020 , n256 , n4019 );
not ( n4021 , n256 );
not ( n4022 , n202 );
nor ( n4023 , n4022 , n3788 );
not ( n4024 , n4023 );
nand ( n4025 , n4024 , n3730 );
nand ( n4026 , n4021 , n4025 );
nand ( n4027 , n4014 , n4020 , n4026 );
nand ( n4028 , n4013 , n4027 );
nand ( n4029 , n4009 , n4028 );
and ( n4030 , n3690 , n4029 );
and ( n4031 , n32 , n3691 );
and ( n4032 , n10 , n40 );
nor ( n4033 , n4031 , n4032 );
or ( n4034 , n4033 , n3864 );
not ( n4035 , n3752 );
or ( n4036 , n201 , n4035 );
nand ( n4037 , n4036 , n3696 );
not ( n4038 , n4037 );
not ( n4039 , n227 );
nor ( n4040 , n4039 , n3725 );
not ( n4041 , n4040 );
nand ( n4042 , n4041 , n3879 );
nand ( n4043 , n256 , n4042 );
not ( n4044 , n256 );
not ( n4045 , n203 );
nor ( n4046 , n4045 , n3816 );
not ( n4047 , n4046 );
nand ( n4048 , n202 , n3738 );
nand ( n4049 , n4047 , n4048 );
nand ( n4050 , n4044 , n4049 );
nand ( n4051 , n4014 , n4043 , n4050 );
nand ( n4052 , n4038 , n4051 );
nand ( n4053 , n4034 , n4052 );
and ( n4054 , n3690 , n4053 );
and ( n4055 , n16 , n3691 );
and ( n4056 , n10 , n24 );
nor ( n4057 , n4055 , n4056 );
or ( n4058 , n4057 , n3864 );
or ( n4059 , n203 , n4010 );
nand ( n4060 , n4059 , n3711 );
not ( n4061 , n4060 );
not ( n4062 , n3877 );
nand ( n4063 , n4062 , n4048 );
nand ( n4064 , n256 , n4063 );
not ( n4065 , n256 );
buf ( n4066 , n205 );
not ( n4067 , n4066 );
nor ( n4068 , n4067 , n3735 );
not ( n4069 , n4068 );
nand ( n4070 , n204 , n3761 );
nand ( n4071 , n4069 , n4070 );
nand ( n4072 , n4065 , n4071 );
nand ( n4073 , n3715 , n4064 , n4072 );
nand ( n4074 , n4061 , n4073 );
nand ( n4075 , n4058 , n4074 );
and ( n4076 , n3690 , n4075 );
and ( n4077 , n6 , n3691 );
and ( n4078 , n10 , n16 );
nor ( n4079 , n4077 , n4078 );
or ( n4080 , n4079 , n3698 );
not ( n4081 , n3752 );
or ( n4082 , n204 , n4081 );
nand ( n4083 , n4082 , n3711 );
not ( n4084 , n4083 );
not ( n4085 , n4023 );
nand ( n4086 , n4085 , n3739 );
nand ( n4087 , n256 , n4086 );
not ( n4088 , n256 );
not ( n4089 , n206 );
nor ( n4090 , n4089 , n3816 );
not ( n4091 , n4090 );
buf ( n4092 , n4066 );
nand ( n4093 , n4092 , n3738 );
nand ( n4094 , n4091 , n4093 );
nand ( n4095 , n4088 , n4094 );
nand ( n4096 , n4014 , n4087 , n4095 );
nand ( n4097 , n4084 , n4096 );
nand ( n4098 , n4080 , n4097 );
and ( n4099 , n3690 , n4098 );
and ( n4100 , n65 , n3691 );
and ( n4101 , n6 , n10 );
nor ( n4102 , n4100 , n4101 );
or ( n4103 , n4102 , n3781 );
not ( n4104 , n3916 );
or ( n4105 , n4092 , n4104 );
nand ( n4106 , n4105 , n3711 );
not ( n4107 , n4106 );
not ( n4108 , n4046 );
nand ( n4109 , n4108 , n4070 );
nand ( n4110 , n256 , n4109 );
not ( n4111 , n256 );
not ( n4112 , n207 );
nor ( n4113 , n4112 , n3735 );
not ( n4114 , n4113 );
nand ( n4115 , n206 , n3729 );
nand ( n4116 , n4114 , n4115 );
nand ( n4117 , n4111 , n4116 );
nand ( n4118 , n3715 , n4110 , n4117 );
nand ( n4119 , n4107 , n4118 );
nand ( n4120 , n4103 , n4119 );
and ( n4121 , n3690 , n4120 );
and ( n4122 , n57 , n3691 );
and ( n4123 , n10 , n65 );
nor ( n4124 , n4122 , n4123 );
or ( n4125 , n4124 , n3864 );
or ( n4126 , n206 , n3709 );
nand ( n4127 , n4126 , n3711 );
not ( n4128 , n4127 );
not ( n4129 , n3736 );
nand ( n4130 , n4129 , n4093 );
nand ( n4131 , n256 , n4130 );
not ( n4132 , n256 );
not ( n4133 , n208 );
nor ( n4134 , n4133 , n3725 );
not ( n4135 , n4134 );
nand ( n4136 , n207 , n3729 );
nand ( n4137 , n4135 , n4136 );
nand ( n4138 , n4132 , n4137 );
nand ( n4139 , n3715 , n4131 , n4138 );
nand ( n4140 , n4128 , n4139 );
nand ( n4141 , n4125 , n4140 );
and ( n4142 , n3690 , n4141 );
and ( n4143 , n49 , n3691 );
and ( n4144 , n10 , n57 );
nor ( n4145 , n4143 , n4144 );
or ( n4146 , n4145 , n3781 );
or ( n4147 , n207 , n3939 );
nand ( n4148 , n4147 , n3711 );
not ( n4149 , n4148 );
not ( n4150 , n4068 );
nand ( n4151 , n4150 , n4115 );
nand ( n4152 , n256 , n4151 );
not ( n4153 , n256 );
not ( n4154 , n3789 );
nand ( n4155 , n208 , n3769 );
nand ( n4156 , n4154 , n4155 );
nand ( n4157 , n4153 , n4156 );
nand ( n4158 , n4014 , n4152 , n4157 );
nand ( n4159 , n4149 , n4158 );
nand ( n4160 , n4146 , n4159 );
and ( n4161 , n3690 , n4160 );
and ( n4162 , n41 , n3691 );
and ( n4163 , n10 , n49 );
nor ( n4164 , n4162 , n4163 );
or ( n4165 , n4164 , n3750 );
or ( n4166 , n208 , n3986 );
nand ( n4167 , n4166 , n3696 );
not ( n4168 , n4167 );
not ( n4169 , n4090 );
nand ( n4170 , n4169 , n4136 );
nand ( n4171 , n256 , n4170 );
not ( n4172 , n256 );
not ( n4173 , n210 );
nor ( n4174 , n4173 , n3816 );
not ( n4175 , n4174 );
nand ( n4176 , n209 , n3738 );
nand ( n4177 , n4175 , n4176 );
nand ( n4178 , n4172 , n4177 );
nand ( n4179 , n4014 , n4171 , n4178 );
nand ( n4180 , n4168 , n4179 );
nand ( n4181 , n4165 , n4180 );
and ( n4182 , n3690 , n4181 );
and ( n4183 , n33 , n3691 );
and ( n4184 , n10 , n41 );
nor ( n4185 , n4183 , n4184 );
or ( n4186 , n4185 , n3750 );
or ( n4187 , n209 , n4081 );
nand ( n4188 , n4187 , n3696 );
not ( n4189 , n4188 );
not ( n4190 , n4113 );
nand ( n4191 , n4190 , n4155 );
nand ( n4192 , n256 , n4191 );
not ( n4193 , n256 );
not ( n4194 , n211 );
nor ( n4195 , n4194 , n3735 );
not ( n4196 , n4195 );
nand ( n4197 , n4196 , n3791 );
nand ( n4198 , n4193 , n4197 );
nand ( n4199 , n3715 , n4192 , n4198 );
nand ( n4200 , n4189 , n4199 );
nand ( n4201 , n4186 , n4200 );
and ( n4202 , n3690 , n4201 );
and ( n4203 , n25 , n3691 );
and ( n4204 , n10 , n33 );
nor ( n4205 , n4203 , n4204 );
or ( n4206 , n4205 , n3937 );
or ( n4207 , n210 , n3753 );
nand ( n4208 , n4207 , n3696 );
not ( n4209 , n4208 );
not ( n4210 , n4134 );
nand ( n4211 , n4210 , n4176 );
nand ( n4212 , n256 , n4211 );
not ( n4213 , n256 );
not ( n4214 , n212 );
nor ( n4215 , n4214 , n3725 );
not ( n4216 , n4215 );
nand ( n4217 , n211 , n3729 );
nand ( n4218 , n4216 , n4217 );
nand ( n4219 , n4213 , n4218 );
nand ( n4220 , n3715 , n4212 , n4219 );
nand ( n4221 , n4209 , n4220 );
nand ( n4222 , n4206 , n4221 );
and ( n4223 , n3690 , n4222 );
and ( n4224 , n7 , n3691 );
and ( n4225 , n10 , n17 );
nor ( n4226 , n4224 , n4225 );
not ( n4227 , n3749 );
or ( n4228 , n4226 , n4227 );
or ( n4229 , n212 , n3840 );
nand ( n4230 , n4229 , n3711 );
not ( n4231 , n4230 );
not ( n4232 , n4174 );
nand ( n4233 , n4232 , n4217 );
nand ( n4234 , n256 , n4233 );
not ( n4235 , n256 );
not ( n4236 , n214 );
nor ( n4237 , n4236 , n3725 );
not ( n4238 , n4237 );
nand ( n4239 , n213 , n3738 );
nand ( n4240 , n4238 , n4239 );
nand ( n4241 , n4235 , n4240 );
nand ( n4242 , n3786 , n4234 , n4241 );
nand ( n4243 , n4231 , n4242 );
nand ( n4244 , n4228 , n4243 );
and ( n4245 , n3690 , n4244 );
and ( n4246 , n66 , n3691 );
and ( n4247 , n7 , n10 );
nor ( n4248 , n4246 , n4247 );
or ( n4249 , n4248 , n4227 );
or ( n4250 , n213 , n4104 );
nand ( n4251 , n4250 , n3696 );
not ( n4252 , n4251 );
not ( n4253 , n4195 );
nand ( n4254 , n4253 , n3798 );
nand ( n4255 , n256 , n4254 );
not ( n4256 , n256 );
not ( n4257 , n215 );
nor ( n4258 , n4257 , n3725 );
not ( n4259 , n4258 );
nand ( n4260 , n4259 , n3922 );
nand ( n4261 , n4256 , n4260 );
nand ( n4262 , n4014 , n4255 , n4261 );
nand ( n4263 , n4252 , n4262 );
nand ( n4264 , n4249 , n4263 );
and ( n4265 , n3690 , n4264 );
and ( n4266 , n58 , n3691 );
and ( n4267 , n10 , n66 );
nor ( n4268 , n4266 , n4267 );
or ( n4269 , n4268 , n3808 );
or ( n4270 , n214 , n3753 );
nand ( n4271 , n4270 , n3711 );
not ( n4272 , n4271 );
not ( n4273 , n4215 );
nand ( n4274 , n4273 , n4239 );
nand ( n4275 , n256 , n4274 );
not ( n4276 , n256 );
not ( n4277 , n216 );
nor ( n4278 , n4277 , n3725 );
not ( n4279 , n4278 );
nand ( n4280 , n215 , n3738 );
nand ( n4281 , n4279 , n4280 );
nand ( n4282 , n4276 , n4281 );
nand ( n4283 , n4014 , n4275 , n4282 );
nand ( n4284 , n4272 , n4283 );
nand ( n4285 , n4269 , n4284 );
and ( n4286 , n3690 , n4285 );
and ( n4287 , n42 , n3691 );
and ( n4288 , n10 , n50 );
nor ( n4289 , n4287 , n4288 );
or ( n4290 , n4289 , n4227 );
not ( n4291 , n3916 );
or ( n4292 , n216 , n4291 );
nand ( n4293 , n4292 , n3711 );
not ( n4294 , n4293 );
not ( n4295 , n4237 );
nand ( n4296 , n4295 , n4280 );
nand ( n4297 , n256 , n4296 );
not ( n4298 , n256 );
not ( n4299 , n218 );
nor ( n4300 , n4299 , n3725 );
not ( n4301 , n4300 );
nand ( n4302 , n217 , n3729 );
nand ( n4303 , n4301 , n4302 );
nand ( n4304 , n4298 , n4303 );
nand ( n4305 , n3715 , n4297 , n4304 );
nand ( n4306 , n4294 , n4305 );
nand ( n4307 , n4290 , n4306 );
and ( n4308 , n3690 , n4307 );
and ( n4309 , n34 , n3691 );
and ( n4310 , n10 , n42 );
nor ( n4311 , n4309 , n4310 );
or ( n4312 , n4311 , n4227 );
or ( n4313 , n217 , n4035 );
nand ( n4314 , n4313 , n3711 );
not ( n4315 , n4314 );
not ( n4316 , n4258 );
nand ( n4317 , n4316 , n3927 );
nand ( n4318 , n256 , n4317 );
not ( n4319 , n256 );
not ( n4320 , n219 );
nor ( n4321 , n4320 , n3816 );
not ( n4322 , n4321 );
nand ( n4323 , n4322 , n3847 );
nand ( n4324 , n4319 , n4323 );
nand ( n4325 , n3757 , n4318 , n4324 );
nand ( n4326 , n4315 , n4325 );
nand ( n4327 , n4312 , n4326 );
and ( n4328 , n3690 , n4327 );
and ( n4329 , n26 , n3691 );
and ( n4330 , n10 , n34 );
nor ( n4331 , n4329 , n4330 );
or ( n4332 , n4331 , n3937 );
or ( n4333 , n218 , n3810 );
nand ( n4334 , n4333 , n3696 );
not ( n4335 , n4334 );
not ( n4336 , n4278 );
nand ( n4337 , n4336 , n4302 );
nand ( n4338 , n256 , n4337 );
not ( n4339 , n256 );
not ( n4340 , n3759 );
nand ( n4341 , n219 , n3761 );
nand ( n4342 , n4340 , n4341 );
nand ( n4343 , n4339 , n4342 );
nand ( n4344 , n3757 , n4338 , n4343 );
nand ( n4345 , n4335 , n4344 );
nand ( n4346 , n4332 , n4345 );
and ( n4347 , n3690 , n4346 );
and ( n4348 , n8 , n3691 );
and ( n4349 , n10 , n18 );
nor ( n4350 , n4348 , n4349 );
or ( n4351 , n4350 , n3937 );
or ( n4352 , n220 , n3810 );
nand ( n4353 , n4352 , n3711 );
not ( n4354 , n4353 );
not ( n4355 , n4300 );
nand ( n4356 , n4355 , n4341 );
nand ( n4357 , n256 , n4356 );
not ( n4358 , n256 );
not ( n4359 , n222 );
nor ( n4360 , n4359 , n3725 );
not ( n4361 , n4360 );
nand ( n4362 , n4361 , n3762 );
nand ( n4363 , n4358 , n4362 );
nand ( n4364 , n3715 , n4357 , n4363 );
nand ( n4365 , n4354 , n4364 );
nand ( n4366 , n4351 , n4365 );
and ( n4367 , n3690 , n4366 );
and ( n4368 , n67 , n3691 );
and ( n4369 , n8 , n10 );
nor ( n4370 , n4368 , n4369 );
or ( n4371 , n4370 , n3750 );
or ( n4372 , n221 , n4081 );
nand ( n4373 , n4372 , n3696 );
not ( n4374 , n4373 );
not ( n4375 , n4321 );
nand ( n4376 , n4375 , n3854 );
nand ( n4377 , n256 , n4376 );
not ( n4378 , n256 );
not ( n4379 , n223 );
nor ( n4380 , n4379 , n3735 );
not ( n4381 , n4380 );
nand ( n4382 , n222 , n3769 );
nand ( n4383 , n4381 , n4382 );
nand ( n4384 , n4378 , n4383 );
nand ( n4385 , n3757 , n4377 , n4384 );
nand ( n4386 , n4374 , n4385 );
nand ( n4387 , n4371 , n4386 );
and ( n4388 , n3690 , n4387 );
and ( n4389 , n43 , n3691 );
and ( n4390 , n10 , n51 );
nor ( n4391 , n4389 , n4390 );
or ( n4392 , n4391 , n3698 );
not ( n4393 , n3708 );
or ( n4394 , n224 , n4393 );
nand ( n4395 , n4394 , n3711 );
not ( n4396 , n4395 );
not ( n4397 , n4360 );
nand ( n4398 , n4397 , n3770 );
nand ( n4399 , n256 , n4398 );
not ( n4400 , n256 );
not ( n4401 , n4016 );
nand ( n4402 , n225 , n3729 );
nand ( n4403 , n4401 , n4402 );
nand ( n4404 , n4400 , n4403 );
nand ( n4405 , n3715 , n4399 , n4404 );
nand ( n4406 , n4396 , n4405 );
nand ( n4407 , n4392 , n4406 );
and ( n4408 , n3690 , n4407 );
and ( n4409 , n35 , n3691 );
and ( n4410 , n10 , n43 );
nor ( n4411 , n4409 , n4410 );
not ( n4412 , n3780 );
or ( n4413 , n4411 , n4412 );
or ( n4414 , n225 , n3986 );
nand ( n4415 , n4414 , n3696 );
not ( n4416 , n4415 );
not ( n4417 , n4380 );
nand ( n4418 , n224 , n3729 );
nand ( n4419 , n4417 , n4418 );
nand ( n4420 , n256 , n4419 );
not ( n4421 , n256 );
not ( n4422 , n4040 );
nand ( n4423 , n4422 , n3872 );
nand ( n4424 , n4421 , n4423 );
nand ( n4425 , n3715 , n4420 , n4424 );
nand ( n4426 , n4416 , n4425 );
nand ( n4427 , n4413 , n4426 );
and ( n4428 , n3690 , n4427 );
and ( n4429 , n27 , n3691 );
and ( n4430 , n10 , n35 );
nor ( n4431 , n4429 , n4430 );
or ( n4432 , n4431 , n4412 );
or ( n4433 , n226 , n4393 );
nand ( n4434 , n4433 , n3696 );
not ( n4435 , n4434 );
not ( n4436 , n3767 );
nand ( n4437 , n4436 , n4402 );
nand ( n4438 , n256 , n4437 );
not ( n4439 , n256 );
not ( n4440 , n3726 );
nand ( n4441 , n4440 , n4018 );
nand ( n4442 , n4439 , n4441 );
nand ( n4443 , n3786 , n4438 , n4442 );
nand ( n4444 , n4435 , n4443 );
nand ( n4445 , n4432 , n4444 );
and ( n4446 , n3690 , n4445 );
and ( n4447 , n5 , n3691 );
and ( n4448 , n10 , n13 );
nor ( n4449 , n4447 , n4448 );
or ( n4450 , n4449 , n3959 );
or ( n4451 , n228 , n4081 );
nand ( n4452 , n4451 , n3696 );
not ( n4453 , n4452 );
nor ( n4454 , n3079 , n3735 );
not ( n4455 , n4454 );
nand ( n4456 , n255 , n3769 );
nand ( n4457 , n4455 , n4456 );
nand ( n4458 , n256 , n4457 );
not ( n4459 , n256 );
not ( n4460 , n230 );
nor ( n4461 , n4460 , n3816 );
not ( n4462 , n4461 );
nand ( n4463 , n229 , n3761 );
nand ( n4464 , n4462 , n4463 );
nand ( n4465 , n4459 , n4464 );
nand ( n4466 , n3786 , n4458 , n4465 );
nand ( n4467 , n4453 , n4466 );
nand ( n4468 , n4450 , n4467 );
and ( n4469 , n3690 , n4468 );
and ( n4470 , n64 , n3691 );
and ( n4471 , n5 , n10 );
nor ( n4472 , n4470 , n4471 );
or ( n4473 , n4472 , n3959 );
or ( n4474 , n229 , n4010 );
nand ( n4475 , n4474 , n3711 );
not ( n4476 , n4475 );
not ( n4477 , n255 );
nor ( n4478 , n4477 , n3788 );
not ( n4479 , n4478 );
nand ( n4480 , n228 , n3761 );
nand ( n4481 , n4479 , n4480 );
nand ( n4482 , n256 , n4481 );
not ( n4483 , n256 );
not ( n4484 , n231 );
nor ( n4485 , n4484 , n3788 );
not ( n4486 , n4485 );
nand ( n4487 , n4486 , n3967 );
nand ( n4488 , n4483 , n4487 );
nand ( n4489 , n3814 , n4482 , n4488 );
nand ( n4490 , n4476 , n4489 );
nand ( n4491 , n4473 , n4490 );
and ( n4492 , n3690 , n4491 );
and ( n4493 , n56 , n3691 );
and ( n4494 , n10 , n64 );
nor ( n4495 , n4493 , n4494 );
or ( n4496 , n4495 , n3781 );
or ( n4497 , n230 , n3939 );
nand ( n4498 , n4497 , n3696 );
not ( n4499 , n4498 );
not ( n4500 , n228 );
nor ( n4501 , n4500 , n3735 );
not ( n4502 , n4501 );
nand ( n4503 , n4502 , n4463 );
nand ( n4504 , n256 , n4503 );
not ( n4505 , n256 );
not ( n4506 , n232 );
nor ( n4507 , n4506 , n3735 );
not ( n4508 , n4507 );
nand ( n4509 , n231 , n3761 );
nand ( n4510 , n4508 , n4509 );
nand ( n4511 , n4505 , n4510 );
nand ( n4512 , n3814 , n4504 , n4511 );
nand ( n4513 , n4499 , n4512 );
nand ( n4514 , n4496 , n4513 );
and ( n4515 , n3690 , n4514 );
and ( n4516 , n4 , n3691 );
and ( n4517 , n10 , n48 );
nor ( n4518 , n4516 , n4517 );
or ( n4519 , n4518 , n3959 );
or ( n4520 , n232 , n3917 );
nand ( n4521 , n4520 , n3711 );
not ( n4522 , n4521 );
not ( n4523 , n4461 );
nand ( n4524 , n4523 , n4509 );
nand ( n4525 , n256 , n4524 );
not ( n4526 , n256 );
nor ( n4527 , n561 , n3735 );
not ( n4528 , n4527 );
nand ( n4529 , n233 , n3738 );
nand ( n4530 , n4528 , n4529 );
nand ( n4531 , n4526 , n4530 );
nand ( n4532 , n3786 , n4525 , n4531 );
nand ( n4533 , n4522 , n4532 );
nand ( n4534 , n4519 , n4533 );
and ( n4535 , n3690 , n4534 );
and ( n4536 , n63 , n3691 );
and ( n4537 , n4 , n10 );
nor ( n4538 , n4536 , n4537 );
not ( n4539 , n3780 );
or ( n4540 , n4538 , n4539 );
or ( n4541 , n233 , n3840 );
nand ( n4542 , n4541 , n3711 );
not ( n4543 , n4542 );
not ( n4544 , n4485 );
nand ( n4545 , n4544 , n3974 );
nand ( n4546 , n256 , n4545 );
not ( n4547 , n256 );
not ( n4548 , n235 );
nor ( n4549 , n4548 , n3725 );
not ( n4550 , n4549 );
nand ( n4551 , n4550 , n3991 );
nand ( n4552 , n4547 , n4551 );
nand ( n4553 , n3814 , n4546 , n4552 );
nand ( n4554 , n4543 , n4553 );
nand ( n4555 , n4540 , n4554 );
and ( n4556 , n3690 , n4555 );
and ( n4557 , n55 , n3691 );
and ( n4558 , n10 , n63 );
nor ( n4559 , n4557 , n4558 );
or ( n4560 , n4559 , n4539 );
or ( n4561 , n234 , n3917 );
nand ( n4562 , n4561 , n3711 );
not ( n4563 , n4562 );
not ( n4564 , n4507 );
nand ( n4565 , n4564 , n4529 );
nand ( n4566 , n256 , n4565 );
not ( n4567 , n256 );
not ( n4568 , n236 );
nor ( n4569 , n4568 , n3725 );
not ( n4570 , n4569 );
nand ( n4571 , n235 , n3729 );
nand ( n4572 , n4570 , n4571 );
nand ( n4573 , n4567 , n4572 );
nand ( n4574 , n3814 , n4566 , n4573 );
nand ( n4575 , n4563 , n4574 );
nand ( n4576 , n4560 , n4575 );
and ( n4577 , n3690 , n4576 );
and ( n4578 , n39 , n3691 );
and ( n4579 , n10 , n47 );
nor ( n4580 , n4578 , n4579 );
or ( n4581 , n4580 , n4412 );
or ( n4582 , n236 , n3709 );
nand ( n4583 , n4582 , n3696 );
not ( n4584 , n4583 );
not ( n4585 , n4527 );
nand ( n4586 , n4585 , n4571 );
nand ( n4587 , n256 , n4586 );
not ( n4588 , n256 );
not ( n4589 , n238 );
nor ( n4590 , n4589 , n3725 );
not ( n4591 , n4590 );
nand ( n4592 , n237 , n3729 );
nand ( n4593 , n4591 , n4592 );
nand ( n4594 , n4588 , n4593 );
nand ( n4595 , n3814 , n4587 , n4594 );
nand ( n4596 , n4584 , n4595 );
nand ( n4597 , n4581 , n4596 );
and ( n4598 , n3690 , n4597 );
and ( n4599 , n31 , n3691 );
and ( n4600 , n10 , n39 );
nor ( n4601 , n4599 , n4600 );
or ( n4602 , n4601 , n4412 );
or ( n4603 , n237 , n4291 );
nand ( n4604 , n4603 , n3696 );
not ( n4605 , n4604 );
not ( n4606 , n4549 );
nand ( n4607 , n4606 , n3998 );
nand ( n4608 , n256 , n4607 );
not ( n4609 , n256 );
not ( n4610 , n239 );
nor ( n4611 , n4610 , n3735 );
not ( n4612 , n4611 );
nand ( n4613 , n238 , n3761 );
nand ( n4614 , n4612 , n4613 );
nand ( n4615 , n4609 , n4614 );
nand ( n4616 , n3715 , n4608 , n4615 );
nand ( n4617 , n4605 , n4616 );
nand ( n4618 , n4602 , n4617 );
and ( n4619 , n3690 , n4618 );
and ( n4620 , n23 , n3691 );
and ( n4621 , n10 , n31 );
nor ( n4622 , n4620 , n4621 );
or ( n4623 , n4622 , n3984 );
or ( n4624 , n238 , n4393 );
nand ( n4625 , n4624 , n3711 );
not ( n4626 , n4625 );
not ( n4627 , n4569 );
nand ( n4628 , n4627 , n4592 );
nand ( n4629 , n256 , n4628 );
not ( n4630 , n256 );
not ( n4631 , n240 );
nor ( n4632 , n4631 , n3735 );
not ( n4633 , n4632 );
nand ( n4634 , n239 , n3729 );
nand ( n4635 , n4633 , n4634 );
nand ( n4636 , n4630 , n4635 );
nand ( n4637 , n3715 , n4629 , n4636 );
nand ( n4638 , n4626 , n4637 );
nand ( n4639 , n4623 , n4638 );
and ( n4640 , n3690 , n4639 );
and ( n4641 , n15 , n3691 );
and ( n4642 , n10 , n23 );
nor ( n4643 , n4641 , n4642 );
or ( n4644 , n4643 , n3984 );
or ( n4645 , n239 , n3939 );
nand ( n4646 , n4645 , n3696 );
not ( n4647 , n4646 );
not ( n4648 , n3996 );
nand ( n4649 , n4648 , n4613 );
nand ( n4650 , n256 , n4649 );
not ( n4651 , n256 );
not ( n4652 , n3817 );
nand ( n4653 , n240 , n3738 );
nand ( n4654 , n4652 , n4653 );
nand ( n4655 , n4651 , n4654 );
nand ( n4656 , n3757 , n4650 , n4655 );
nand ( n4657 , n4647 , n4656 );
nand ( n4658 , n4644 , n4657 );
and ( n4659 , n3690 , n4658 );
and ( n4660 , n3 , n3691 );
and ( n4661 , n10 , n15 );
nor ( n4662 , n4660 , n4661 );
not ( n4663 , n3749 );
or ( n4664 , n4662 , n4663 );
or ( n4665 , n240 , n4035 );
nand ( n4666 , n4665 , n3711 );
not ( n4667 , n4666 );
not ( n4668 , n4590 );
nand ( n4669 , n4668 , n4634 );
nand ( n4670 , n256 , n4669 );
not ( n4671 , n256 );
not ( n4672 , n3819 );
nor ( n4673 , n4672 , n3735 );
not ( n4674 , n4673 );
nand ( n4675 , n241 , n3761 );
nand ( n4676 , n4674 , n4675 );
nand ( n4677 , n4671 , n4676 );
nand ( n4678 , n3757 , n4670 , n4677 );
nand ( n4679 , n4667 , n4678 );
nand ( n4680 , n4664 , n4679 );
and ( n4681 , n3690 , n4680 );
and ( n4682 , n62 , n3691 );
and ( n4683 , n3 , n10 );
nor ( n4684 , n4682 , n4683 );
or ( n4685 , n4684 , n4539 );
or ( n4686 , n241 , n3840 );
nand ( n4687 , n4686 , n3696 );
not ( n4688 , n4687 );
not ( n4689 , n4611 );
nand ( n4690 , n4689 , n4653 );
nand ( n4691 , n256 , n4690 );
not ( n4692 , n256 );
not ( n4693 , n243 );
nor ( n4694 , n4693 , n3725 );
not ( n4695 , n4694 );
nand ( n4696 , n4695 , n3821 );
nand ( n4697 , n4692 , n4696 );
nand ( n4698 , n3814 , n4691 , n4697 );
nand ( n4699 , n4688 , n4698 );
nand ( n4700 , n4685 , n4699 );
and ( n4701 , n3690 , n4700 );
and ( n4702 , n54 , n3691 );
and ( n4703 , n10 , n62 );
nor ( n4704 , n4702 , n4703 );
or ( n4705 , n4704 , n4663 );
or ( n4706 , n3820 , n3709 );
nand ( n4707 , n4706 , n3696 );
not ( n4708 , n4707 );
not ( n4709 , n4632 );
nand ( n4710 , n4709 , n4675 );
nand ( n4711 , n256 , n4710 );
not ( n4712 , n256 );
not ( n4713 , n244 );
nor ( n4714 , n4713 , n3788 );
not ( n4715 , n4714 );
nand ( n4716 , n243 , n3729 );
nand ( n4717 , n4715 , n4716 );
nand ( n4718 , n4712 , n4717 );
nand ( n4719 , n4014 , n4711 , n4718 );
nand ( n4720 , n4708 , n4719 );
nand ( n4721 , n4705 , n4720 );
and ( n4722 , n3690 , n4721 );
and ( n4723 , n38 , n3691 );
and ( n4724 , n10 , n46 );
nor ( n4725 , n4723 , n4724 );
or ( n4726 , n4725 , n4663 );
or ( n4727 , n244 , n4104 );
nand ( n4728 , n4727 , n3696 );
not ( n4729 , n4728 );
not ( n4730 , n4673 );
nand ( n4731 , n4730 , n4716 );
nand ( n4732 , n256 , n4731 );
not ( n4733 , n256 );
not ( n4734 , n246 );
nor ( n4735 , n4734 , n3816 );
not ( n4736 , n4735 );
nand ( n4737 , n245 , n3738 );
nand ( n4738 , n4736 , n4737 );
nand ( n4739 , n4733 , n4738 );
nand ( n4740 , n3814 , n4732 , n4739 );
nand ( n4741 , n4729 , n4740 );
nand ( n4742 , n4726 , n4741 );
and ( n4743 , n3690 , n4742 );
and ( n4744 , n30 , n3691 );
and ( n4745 , n10 , n38 );
nor ( n4746 , n4744 , n4745 );
or ( n4747 , n4746 , n3838 );
or ( n4748 , n245 , n4104 );
nand ( n4749 , n4748 , n3711 );
not ( n4750 , n4749 );
not ( n4751 , n4694 );
nand ( n4752 , n4751 , n3828 );
nand ( n4753 , n256 , n4752 );
not ( n4754 , n256 );
not ( n4755 , n247 );
nor ( n4756 , n4755 , n3735 );
not ( n4757 , n4756 );
nand ( n4758 , n4757 , n3944 );
nand ( n4759 , n4754 , n4758 );
nand ( n4760 , n3814 , n4753 , n4759 );
nand ( n4761 , n4750 , n4760 );
nand ( n4762 , n4747 , n4761 );
and ( n4763 , n3690 , n4762 );
and ( n4764 , n22 , n3691 );
and ( n4765 , n10 , n30 );
nor ( n4766 , n4764 , n4765 );
or ( n4767 , n4766 , n4663 );
or ( n4768 , n246 , n3986 );
nand ( n4769 , n4768 , n3696 );
not ( n4770 , n4769 );
not ( n4771 , n4714 );
nand ( n4772 , n4771 , n4737 );
nand ( n4773 , n256 , n4772 );
not ( n4774 , n256 );
not ( n4775 , n248 );
nor ( n4776 , n4775 , n3788 );
not ( n4777 , n4776 );
nand ( n4778 , n247 , n3738 );
nand ( n4779 , n4777 , n4778 );
nand ( n4780 , n4774 , n4779 );
nand ( n4781 , n3814 , n4773 , n4780 );
nand ( n4782 , n4770 , n4781 );
nand ( n4783 , n4767 , n4782 );
and ( n4784 , n3690 , n4783 );
and ( n4785 , n2 , n3691 );
and ( n4786 , n10 , n14 );
nor ( n4787 , n4785 , n4786 );
or ( n4788 , n4787 , n3808 );
or ( n4789 , n248 , n3891 );
nand ( n4790 , n4789 , n3711 );
not ( n4791 , n4790 );
not ( n4792 , n4735 );
nand ( n4793 , n4792 , n4778 );
nand ( n4794 , n256 , n4793 );
not ( n4795 , n256 );
not ( n4796 , n250 );
nor ( n4797 , n4796 , n3725 );
not ( n4798 , n4797 );
nand ( n4799 , n249 , n3769 );
nand ( n4800 , n4798 , n4799 );
nand ( n4801 , n4795 , n4800 );
nand ( n4802 , n3814 , n4794 , n4801 );
nand ( n4803 , n4791 , n4802 );
nand ( n4804 , n4788 , n4803 );
and ( n4805 , n3690 , n4804 );
and ( n4806 , n61 , n3691 );
and ( n4807 , n2 , n10 );
nor ( n4808 , n4806 , n4807 );
or ( n4809 , n4808 , n4539 );
or ( n4810 , n249 , n3917 );
nand ( n4811 , n4810 , n3696 );
not ( n4812 , n4811 );
not ( n4813 , n4756 );
nand ( n4814 , n4813 , n3949 );
nand ( n4815 , n256 , n4814 );
not ( n4816 , n256 );
not ( n4817 , n251 );
nor ( n4818 , n4817 , n3788 );
not ( n4819 , n4818 );
nand ( n4820 , n4819 , n3898 );
nand ( n4821 , n4816 , n4820 );
nand ( n4822 , n3786 , n4815 , n4821 );
nand ( n4823 , n4812 , n4822 );
nand ( n4824 , n4809 , n4823 );
and ( n4825 , n3690 , n4824 );
and ( n4826 , n53 , n3691 );
and ( n4827 , n10 , n61 );
nor ( n4828 , n4826 , n4827 );
or ( n4829 , n4828 , n3838 );
or ( n4830 , n250 , n3891 );
nand ( n4831 , n4830 , n3711 );
not ( n4832 , n4831 );
not ( n4833 , n4776 );
nand ( n4834 , n4833 , n4799 );
nand ( n4835 , n256 , n4834 );
not ( n4836 , n256 );
not ( n4837 , n252 );
nor ( n4838 , n4837 , n3735 );
not ( n4839 , n4838 );
nand ( n4840 , n251 , n3769 );
nand ( n4841 , n4839 , n4840 );
nand ( n4842 , n4836 , n4841 );
nand ( n4843 , n3814 , n4835 , n4842 );
nand ( n4844 , n4832 , n4843 );
nand ( n4845 , n4829 , n4844 );
and ( n4846 , n3690 , n4845 );
and ( n4847 , n37 , n3691 );
and ( n4848 , n10 , n45 );
nor ( n4849 , n4847 , n4848 );
or ( n4850 , n4849 , n4008 );
or ( n4851 , n252 , n4010 );
nand ( n4852 , n4851 , n3711 );
not ( n4853 , n4852 );
not ( n4854 , n4797 );
nand ( n4855 , n4854 , n4840 );
nand ( n4856 , n256 , n4855 );
not ( n4857 , n256 );
not ( n4858 , n4454 );
nand ( n4859 , n253 , n3769 );
nand ( n4860 , n4858 , n4859 );
nand ( n4861 , n4857 , n4860 );
nand ( n4862 , n3715 , n4856 , n4861 );
nand ( n4863 , n4853 , n4862 );
nand ( n4864 , n4850 , n4863 );
and ( n4865 , n3690 , n4864 );
and ( n4866 , n29 , n3691 );
and ( n4867 , n10 , n37 );
nor ( n4868 , n4866 , n4867 );
or ( n4869 , n4868 , n3984 );
or ( n4870 , n253 , n4291 );
nand ( n4871 , n4870 , n3711 );
not ( n4872 , n4871 );
not ( n4873 , n4818 );
nand ( n4874 , n4873 , n3905 );
nand ( n4875 , n256 , n4874 );
not ( n4876 , n256 );
not ( n4877 , n4478 );
nand ( n4878 , n254 , n3761 );
nand ( n4879 , n4877 , n4878 );
nand ( n4880 , n4876 , n4879 );
nand ( n4881 , n3757 , n4875 , n4880 );
nand ( n4882 , n4872 , n4881 );
nand ( n4883 , n4869 , n4882 );
and ( n4884 , n3690 , n4883 );
and ( n4885 , n21 , n3691 );
and ( n4886 , n10 , n29 );
nor ( n4887 , n4885 , n4886 );
or ( n4888 , n4887 , n4008 );
or ( n4889 , n254 , n4291 );
nand ( n4890 , n4889 , n3711 );
not ( n4891 , n4890 );
not ( n4892 , n4838 );
nand ( n4893 , n4892 , n4859 );
nand ( n4894 , n256 , n4893 );
not ( n4895 , n256 );
not ( n4896 , n4501 );
nand ( n4897 , n4896 , n4456 );
nand ( n4898 , n4895 , n4897 );
nand ( n4899 , n3814 , n4894 , n4898 );
nand ( n4900 , n4891 , n4899 );
nand ( n4901 , n4888 , n4900 );
and ( n4902 , n3690 , n4901 );
and ( n4903 , n13 , n3691 );
and ( n4904 , n10 , n21 );
nor ( n4905 , n4903 , n4904 );
or ( n4906 , n4905 , n4008 );
or ( n4907 , n255 , n4393 );
nand ( n4908 , n4907 , n3696 );
not ( n4909 , n4908 );
not ( n4910 , n3903 );
nand ( n4911 , n4910 , n4878 );
nand ( n4912 , n256 , n4911 );
not ( n4913 , n256 );
not ( n4914 , n3965 );
nand ( n4915 , n4914 , n4480 );
nand ( n4916 , n4913 , n4915 );
nand ( n4917 , n3814 , n4912 , n4916 );
nand ( n4918 , n4909 , n4917 );
nand ( n4919 , n4906 , n4918 );
and ( n4920 , n3690 , n4919 );
and ( n4921 , n51 , n3691 );
and ( n4922 , n10 , n59 );
nor ( n4923 , n4921 , n4922 );
or ( n4924 , n4923 , n3698 );
or ( n4925 , n223 , n4035 );
nand ( n4926 , n4925 , n3696 );
not ( n4927 , n4926 );
not ( n4928 , n3852 );
nand ( n4929 , n4928 , n4382 );
nand ( n4930 , n256 , n4929 );
not ( n4931 , n256 );
not ( n4932 , n3870 );
nand ( n4933 , n4932 , n4418 );
nand ( n4934 , n4931 , n4933 );
nand ( n4935 , n3757 , n4930 , n4934 );
nand ( n4936 , n4927 , n4935 );
nand ( n4937 , n4924 , n4936 );
and ( n4938 , n3690 , n4937 );
not ( n4939 , n135 );
buf ( n4940 , n504 );
buf ( n4941 , n4940 );
or ( n4942 , n4939 , n4941 );
not ( n4943 , n4940 );
not ( n4944 , n4943 );
nand ( n4945 , n44 , n4944 );
nand ( n4946 , n4942 , n4945 );
and ( n4947 , n87 , n509 );
and ( n4948 , n79 , n199 );
nor ( n4949 , n4947 , n4948 );
or ( n4950 , n4949 , n4941 );
nand ( n4951 , n145 , n4944 );
nand ( n4952 , n4950 , n4951 );
and ( n4953 , n119 , n509 );
and ( n4954 , n111 , n199 );
nor ( n4955 , n4953 , n4954 );
or ( n4956 , n4955 , n4941 );
nand ( n4957 , n141 , n4944 );
nand ( n4958 , n4956 , n4957 );
not ( n4959 , n163 );
buf ( n4960 , n4940 );
not ( n4961 , n4960 );
or ( n4962 , n4959 , n4961 );
nand ( n4963 , n509 , n75 , n4943 );
nand ( n4964 , n4962 , n4963 );
not ( n4965 , n139 );
not ( n4966 , n4960 );
or ( n4967 , n4965 , n4966 );
nand ( n4968 , n509 , n69 , n4943 );
nand ( n4969 , n4967 , n4968 );
not ( n4970 , n147 );
not ( n4971 , n4960 );
or ( n4972 , n4970 , n4971 );
nand ( n4973 , n509 , n71 , n4943 );
nand ( n4974 , n4972 , n4973 );
and ( n4975 , n95 , n509 );
and ( n4976 , n87 , n199 );
nor ( n4977 , n4975 , n4976 );
or ( n4978 , n4977 , n505 );
nand ( n4979 , n144 , n4944 );
nand ( n4980 , n4978 , n4979 );
not ( n4981 , n160 );
or ( n4982 , n4981 , n505 );
nand ( n4983 , n42 , n4944 );
nand ( n4984 , n4982 , n4983 );
and ( n4985 , n101 , n509 );
and ( n4986 , n93 , n199 );
nor ( n4987 , n4985 , n4986 );
or ( n4988 , n4987 , n4941 );
nand ( n4989 , n135 , n4944 );
nand ( n4990 , n4988 , n4989 );
not ( n4991 , n155 );
not ( n4992 , n4960 );
or ( n4993 , n4991 , n4992 );
nand ( n4994 , n509 , n73 , n4943 );
nand ( n4995 , n4993 , n4994 );
not ( n4996 , n152 );
or ( n4997 , n4996 , n4941 );
nand ( n4998 , n40 , n4944 );
nand ( n4999 , n4997 , n4998 );
and ( n5000 , n129 , n509 );
and ( n5001 , n121 , n199 );
nor ( n5002 , n5000 , n5001 );
not ( n5003 , n4943 );
or ( n5004 , n5002 , n5003 );
buf ( n5005 , n4940 );
nand ( n5006 , n148 , n5005 );
nand ( n5007 , n5004 , n5006 );
and ( n5008 , n109 , n509 );
and ( n5009 , n101 , n199 );
nor ( n5010 , n5008 , n5009 );
or ( n5011 , n5010 , n4941 );
nand ( n5012 , n134 , n4960 );
nand ( n5013 , n5011 , n5012 );
not ( n5014 , n132 );
or ( n5015 , n5014 , n4941 );
nand ( n5016 , n1 , n5005 );
nand ( n5017 , n5015 , n5016 );
not ( n5018 , n156 );
or ( n5019 , n5018 , n5003 );
nand ( n5020 , n7 , n5005 );
nand ( n5021 , n5019 , n5020 );
not ( n5022 , n155 );
or ( n5023 , n5022 , n505 );
nand ( n5024 , n16 , n4960 );
nand ( n5025 , n5023 , n5024 );
nand ( n5026 , n198 , n199 );
xor ( n5027 , n197 , n5026 );
nand ( n5028 , n3689 , n3695 );
nor ( n5029 , n5027 , n5028 );
not ( n5030 , n159 );
not ( n5031 , n505 );
or ( n5032 , n5030 , n5031 );
or ( n5033 , n509 , n99 );
or ( n5034 , n107 , n199 );
not ( n5035 , n4940 );
nand ( n5036 , n5033 , n5034 , n5035 );
nand ( n5037 , n5032 , n5036 );
not ( n5038 , n151 );
not ( n5039 , n505 );
or ( n5040 , n5038 , n5039 );
or ( n5041 , n509 , n97 );
or ( n5042 , n105 , n199 );
nand ( n5043 , n5041 , n5042 , n5035 );
nand ( n5044 , n5040 , n5043 );
not ( n5045 , n138 );
not ( n5046 , n505 );
or ( n5047 , n5045 , n5046 );
or ( n5048 , n509 , n69 );
or ( n5049 , n77 , n199 );
nand ( n5050 , n5048 , n5049 , n5035 );
nand ( n5051 , n5047 , n5050 );
nor ( n5052 , n3717 , n5026 );
xnor ( n5053 , n5052 , n196 );
nor ( n5054 , n5028 , n5053 );
and ( n5055 , n121 , n509 );
and ( n5056 , n113 , n199 );
nor ( n5057 , n5055 , n5056 );
or ( n5058 , n5057 , n4941 );
nand ( n5059 , n149 , n5005 );
nand ( n5060 , n5058 , n5059 );
not ( n5061 , n148 );
or ( n5062 , n5061 , n4941 );
nand ( n5063 , n5 , n4960 );
nand ( n5064 , n5062 , n5063 );
and ( n5065 , n79 , n509 );
and ( n5066 , n71 , n199 );
nor ( n5067 , n5065 , n5066 );
or ( n5068 , n5067 , n4941 );
nand ( n5069 , n146 , n4960 );
nand ( n5070 , n5068 , n5069 );
not ( n5071 , n134 );
not ( n5072 , n505 );
not ( n5073 , n5072 );
or ( n5074 , n5071 , n5073 );
nand ( n5075 , n52 , n4960 );
nand ( n5076 , n5074 , n5075 );
not ( n5077 , n162 );
not ( n5078 , n505 );
or ( n5079 , n5077 , n5078 );
or ( n5080 , n509 , n75 );
or ( n5081 , n83 , n199 );
nand ( n5082 , n5080 , n5081 , n5035 );
nand ( n5083 , n5079 , n5082 );
not ( n5084 , n137 );
not ( n5085 , n5072 );
or ( n5086 , n5084 , n5085 );
nand ( n5087 , n28 , n4960 );
nand ( n5088 , n5086 , n5087 );
and ( n5089 , n91 , n509 );
and ( n5090 , n83 , n199 );
nor ( n5091 , n5089 , n5090 );
or ( n5092 , n5091 , n4941 );
nand ( n5093 , n161 , n5005 );
nand ( n5094 , n5092 , n5093 );
and ( n5095 , n117 , n509 );
and ( n5096 , n109 , n199 );
nor ( n5097 , n5095 , n5096 );
or ( n5098 , n5097 , n5003 );
nand ( n5099 , n133 , n4960 );
nand ( n5100 , n5098 , n5099 );
and ( n5101 , n127 , n509 );
and ( n5102 , n119 , n199 );
nor ( n5103 , n5101 , n5102 );
or ( n5104 , n5103 , n505 );
nand ( n5105 , n140 , n5005 );
nand ( n5106 , n5104 , n5105 );
not ( n5107 , n140 );
or ( n5108 , n5107 , n4941 );
nand ( n5109 , n3 , n5005 );
nand ( n5110 , n5108 , n5109 );
not ( n5111 , n196 );
not ( n5112 , n5052 );
or ( n5113 , n5111 , n5112 );
nand ( n5114 , n5113 , n256 );
not ( n5115 , n3721 );
nand ( n5116 , n5115 , n196 , n199 , n10 );
nand ( n5117 , n5114 , n5116 );
not ( n5118 , n162 );
not ( n5119 , n4960 );
not ( n5120 , n5119 );
or ( n5121 , n5118 , n5120 );
not ( n5122 , n26 );
not ( n5123 , n505 );
or ( n5124 , n5122 , n5123 );
nand ( n5125 , n5121 , n5124 );
not ( n5126 , n133 );
not ( n5127 , n5072 );
or ( n5128 , n5126 , n5127 );
nand ( n5129 , n60 , n4960 );
nand ( n5130 , n5128 , n5129 );
not ( n5131 , n136 );
or ( n5132 , n5131 , n5003 );
nand ( n5133 , n36 , n5005 );
nand ( n5134 , n5132 , n5133 );
and ( n5135 , n103 , n509 );
and ( n5136 , n95 , n199 );
nor ( n5137 , n5135 , n5136 );
or ( n5138 , n5137 , n4941 );
nand ( n5139 , n143 , n5005 );
nand ( n5140 , n5138 , n5139 );
or ( n5141 , n1285 , n505 );
nand ( n5142 , n12 , n5005 );
nand ( n5143 , n5141 , n5142 );
not ( n5144 , n142 );
not ( n5145 , n5119 );
or ( n5146 , n5144 , n5145 );
not ( n5147 , n54 );
not ( n5148 , n505 );
or ( n5149 , n5147 , n5148 );
nand ( n5150 , n5146 , n5149 );
not ( n5151 , n143 );
or ( n5152 , n5151 , n5003 );
nand ( n5153 , n46 , n5005 );
nand ( n5154 , n5152 , n5153 );
not ( n5155 , n145 );
not ( n5156 , n5119 );
or ( n5157 , n5155 , n5156 );
not ( n5158 , n30 );
or ( n5159 , n5158 , n5148 );
nand ( n5160 , n5157 , n5159 );
not ( n5161 , n146 );
not ( n5162 , n4960 );
not ( n5163 , n5162 );
or ( n5164 , n5161 , n5163 );
not ( n5165 , n22 );
or ( n5166 , n5165 , n5123 );
nand ( n5167 , n5164 , n5166 );
not ( n5168 , n151 );
or ( n5169 , n5168 , n4941 );
nand ( n5170 , n48 , n5005 );
nand ( n5171 , n5169 , n5170 );
not ( n5172 , n154 );
not ( n5173 , n5162 );
or ( n5174 , n5172 , n5173 );
not ( n5175 , n24 );
or ( n5176 , n5175 , n5123 );
nand ( n5177 , n5174 , n5176 );
not ( n5178 , n158 );
not ( n5179 , n5162 );
or ( n5180 , n5178 , n5179 );
not ( n5181 , n58 );
or ( n5182 , n5181 , n5148 );
nand ( n5183 , n5180 , n5182 );
not ( n5184 , n161 );
not ( n5185 , n5119 );
or ( n5186 , n5184 , n5185 );
not ( n5187 , n34 );
not ( n5188 , n505 );
or ( n5189 , n5187 , n5188 );
nand ( n5190 , n5186 , n5189 );
and ( n5191 , n198 , n509 );
not ( n5192 , n198 );
and ( n5193 , n199 , n5192 );
nor ( n5194 , n5191 , n5193 );
nor ( n5195 , n5194 , n5028 );
not ( n5196 , n138 );
not ( n5197 , n5072 );
or ( n5198 , n5196 , n5197 );
nand ( n5199 , n20 , n4960 );
nand ( n5200 , n5198 , n5199 );
and ( n5201 , n89 , n509 );
and ( n5202 , n81 , n199 );
nor ( n5203 , n5201 , n5202 );
or ( n5204 , n5203 , n4941 );
nand ( n5205 , n153 , n5005 );
nand ( n5206 , n5204 , n5205 );
and ( n5207 , n85 , n509 );
and ( n5208 , n77 , n199 );
nor ( n5209 , n5207 , n5208 );
or ( n5210 , n5209 , n505 );
nand ( n5211 , n137 , n5005 );
nand ( n5212 , n5210 , n5211 );
and ( n5213 , n99 , n509 );
and ( n5214 , n91 , n199 );
nor ( n5215 , n5213 , n5214 );
or ( n5216 , n5215 , n4941 );
nand ( n5217 , n160 , n4960 );
nand ( n5218 , n5216 , n5217 );
and ( n5219 , n113 , n509 );
and ( n5220 , n105 , n199 );
nor ( n5221 , n5219 , n5220 );
or ( n5222 , n5221 , n4941 );
nand ( n5223 , n150 , n5005 );
nand ( n5224 , n5222 , n5223 );
and ( n5225 , n97 , n509 );
and ( n5226 , n89 , n199 );
nor ( n5227 , n5225 , n5226 );
or ( n5228 , n5227 , n4941 );
nand ( n5229 , n152 , n4960 );
nand ( n5230 , n5228 , n5229 );
not ( n5231 , n158 );
not ( n5232 , n505 );
or ( n5233 , n5231 , n5232 );
or ( n5234 , n509 , n107 );
or ( n5235 , n115 , n199 );
nand ( n5236 , n5234 , n5235 , n5035 );
nand ( n5237 , n5233 , n5236 );
not ( n5238 , n144 );
or ( n5239 , n5238 , n5003 );
nand ( n5240 , n38 , n505 );
nand ( n5241 , n5239 , n5240 );
not ( n5242 , n154 );
not ( n5243 , n505 );
or ( n5244 , n5242 , n5243 );
or ( n5245 , n509 , n73 );
or ( n5246 , n81 , n199 );
nand ( n5247 , n5245 , n5246 , n5035 );
nand ( n5248 , n5244 , n5247 );
nor ( n5249 , n199 , n5028 );
and ( n5250 , n131 , n509 );
and ( n5251 , n123 , n199 );
nor ( n5252 , n5250 , n5251 );
or ( n5253 , n5252 , n505 );
nand ( n5254 , n156 , n5005 );
nand ( n5255 , n5253 , n5254 );
not ( n5256 , n150 );
not ( n5257 , n505 );
not ( n5258 , n5257 );
or ( n5259 , n5256 , n5258 );
not ( n5260 , n56 );
or ( n5261 , n5260 , n5148 );
nand ( n5262 , n5259 , n5261 );
and ( n5263 , n93 , n509 );
and ( n5264 , n85 , n199 );
nor ( n5265 , n5263 , n5264 );
or ( n5266 , n5265 , n4941 );
nand ( n5267 , n136 , n505 );
nand ( n5268 , n5266 , n5267 );
not ( n5269 , n147 );
or ( n5270 , n5269 , n505 );
nand ( n5271 , n14 , n505 );
nand ( n5272 , n5270 , n5271 );
not ( n5273 , n141 );
not ( n5274 , n5257 );
or ( n5275 , n5273 , n5274 );
not ( n5276 , n62 );
or ( n5277 , n5276 , n5188 );
nand ( n5278 , n5275 , n5277 );
and ( n5279 , n111 , n509 );
and ( n5280 , n103 , n199 );
nor ( n5281 , n5279 , n5280 );
or ( n5282 , n5281 , n4941 );
nand ( n5283 , n142 , n505 );
nand ( n5284 , n5282 , n5283 );
not ( n5285 , n149 );
not ( n5286 , n5072 );
or ( n5287 , n5285 , n5286 );
not ( n5288 , n64 );
or ( n5289 , n5288 , n5188 );
nand ( n5290 , n5287 , n5289 );
not ( n5291 , n157 );
not ( n5292 , n5257 );
or ( n5293 , n5291 , n5292 );
not ( n5294 , n66 );
or ( n5295 , n5294 , n5188 );
nand ( n5296 , n5293 , n5295 );
and ( n5297 , n123 , n509 );
and ( n5298 , n115 , n199 );
nor ( n5299 , n5297 , n5298 );
or ( n5300 , n5299 , n4941 );
nand ( n5301 , n157 , n505 );
nand ( n5302 , n5300 , n5301 );
not ( n5303 , n153 );
not ( n5304 , n5257 );
or ( n5305 , n5303 , n5304 );
not ( n5306 , n32 );
or ( n5307 , n5306 , n506 );
nand ( n5308 , n5305 , n5307 );
and ( n5309 , n125 , n509 );
and ( n5310 , n117 , n199 );
nor ( n5311 , n5309 , n5310 );
or ( n5312 , n5311 , n4941 );
nand ( n5313 , n132 , n505 );
nand ( n5314 , n5312 , n5313 );
not ( n5315 , n159 );
or ( n5316 , n5315 , n4941 );
nand ( n5317 , n50 , n505 );
nand ( n5318 , n5316 , n5317 );
or ( n5319 , n728 , n4941 );
nand ( n5320 , n18 , n505 );
nand ( n5321 , n5319 , n5320 );
and ( n5322 , n199 , n44 );
not ( n5323 , n199 );
and ( n5324 , n5323 , n36 );
nor ( n5325 , n5322 , n5324 );
nor ( n5326 , n5325 , n4941 );
and ( n5327 , n199 , n40 );
not ( n5328 , n199 );
and ( n5329 , n5328 , n32 );
nor ( n5330 , n5327 , n5329 );
buf ( n5331 , n4940 );
nor ( n5332 , n5330 , n5331 );
and ( n5333 , n199 , n47 );
not ( n5334 , n199 );
and ( n5335 , n5334 , n39 );
nor ( n5336 , n5333 , n5335 );
nor ( n5337 , n5336 , n5331 );
and ( n5338 , n199 , n32 );
not ( n5339 , n199 );
and ( n5340 , n5339 , n24 );
nor ( n5341 , n5338 , n5340 );
nor ( n5342 , n5341 , n4941 );
and ( n5343 , n199 , n30 );
not ( n5344 , n199 );
and ( n5345 , n5344 , n22 );
nor ( n5346 , n5343 , n5345 );
nor ( n5347 , n5346 , n5331 );
and ( n5348 , n199 , n21 );
not ( n5349 , n199 );
and ( n5350 , n5349 , n13 );
nor ( n5351 , n5348 , n5350 );
nor ( n5352 , n5351 , n5331 );
and ( n5353 , n199 , n64 );
not ( n5354 , n199 );
and ( n5355 , n5354 , n56 );
nor ( n5356 , n5353 , n5355 );
nor ( n5357 , n5356 , n4941 );
and ( n5358 , n199 , n5 );
not ( n5359 , n199 );
and ( n5360 , n5359 , n64 );
nor ( n5361 , n5358 , n5360 );
nor ( n5362 , n5361 , n5331 );
and ( n5363 , n199 , n62 );
not ( n5364 , n199 );
and ( n5365 , n5364 , n54 );
nor ( n5366 , n5363 , n5365 );
nor ( n5367 , n5366 , n5331 );
and ( n5368 , n199 , n61 );
not ( n5369 , n199 );
and ( n5370 , n5369 , n53 );
nor ( n5371 , n5368 , n5370 );
nor ( n5372 , n5371 , n4941 );
and ( n5373 , n199 , n8 );
not ( n5374 , n199 );
and ( n5375 , n5374 , n67 );
nor ( n5376 , n5373 , n5375 );
nor ( n5377 , n5376 , n5331 );
and ( n5378 , n199 , n53 );
not ( n5379 , n199 );
and ( n5380 , n5379 , n45 );
nor ( n5381 , n5378 , n5380 );
nor ( n5382 , n5381 , n5331 );
and ( n5383 , n199 , n55 );
not ( n5384 , n199 );
and ( n5385 , n5384 , n47 );
nor ( n5386 , n5383 , n5385 );
nor ( n5387 , n5386 , n5331 );
and ( n5388 , n199 , n3 );
not ( n5389 , n199 );
and ( n5390 , n5389 , n62 );
nor ( n5391 , n5388 , n5390 );
nor ( n5392 , n5391 , n4941 );
and ( n5393 , n199 , n7 );
not ( n5394 , n199 );
and ( n5395 , n5394 , n66 );
nor ( n5396 , n5393 , n5395 );
nor ( n5397 , n5396 , n5331 );
and ( n5398 , n199 , n4 );
not ( n5399 , n199 );
and ( n5400 , n5399 , n63 );
nor ( n5401 , n5398 , n5400 );
nor ( n5402 , n5401 , n4941 );
and ( n5403 , n199 , n67 );
not ( n5404 , n199 );
and ( n5405 , n5404 , n59 );
nor ( n5406 , n5403 , n5405 );
nor ( n5407 , n5406 , n5331 );
and ( n5408 , n199 , n66 );
not ( n5409 , n199 );
and ( n5410 , n5409 , n58 );
nor ( n5411 , n5408 , n5410 );
nor ( n5412 , n5411 , n5331 );
and ( n5413 , n199 , n56 );
not ( n5414 , n199 );
and ( n5415 , n5414 , n48 );
nor ( n5416 , n5413 , n5415 );
nor ( n5417 , n5416 , n5331 );
and ( n5418 , n199 , n57 );
not ( n5419 , n199 );
and ( n5420 , n5419 , n49 );
nor ( n5421 , n5418 , n5420 );
nor ( n5422 , n5421 , n5331 );
and ( n5423 , n199 , n59 );
not ( n5424 , n199 );
and ( n5425 , n5424 , n51 );
nor ( n5426 , n5423 , n5425 );
nor ( n5427 , n5426 , n5331 );
and ( n5428 , n199 , n50 );
not ( n5429 , n199 );
and ( n5430 , n5429 , n42 );
nor ( n5431 , n5428 , n5430 );
nor ( n5432 , n5431 , n5331 );
and ( n5433 , n199 , n43 );
not ( n5434 , n199 );
and ( n5435 , n5434 , n35 );
nor ( n5436 , n5433 , n5435 );
nor ( n5437 , n5436 , n5331 );
and ( n5438 , n199 , n51 );
not ( n5439 , n199 );
and ( n5440 , n5439 , n43 );
nor ( n5441 , n5438 , n5440 );
nor ( n5442 , n5441 , n5331 );
and ( n5443 , n199 , n48 );
not ( n5444 , n199 );
and ( n5445 , n5444 , n40 );
nor ( n5446 , n5443 , n5445 );
nor ( n5447 , n5446 , n4941 );
and ( n5448 , n199 , n49 );
not ( n5449 , n199 );
and ( n5450 , n5449 , n41 );
nor ( n5451 , n5448 , n5450 );
nor ( n5452 , n5451 , n5331 );
and ( n5453 , n199 , n45 );
not ( n5454 , n199 );
and ( n5455 , n5454 , n37 );
nor ( n5456 , n5453 , n5455 );
nor ( n5457 , n5456 , n4941 );
and ( n5458 , n199 , n41 );
not ( n5459 , n199 );
and ( n5460 , n5459 , n33 );
nor ( n5461 , n5458 , n5460 );
nor ( n5462 , n5461 , n4941 );
and ( n5463 , n199 , n42 );
not ( n5464 , n199 );
and ( n5465 , n5464 , n34 );
nor ( n5466 , n5463 , n5465 );
nor ( n5467 , n5466 , n5331 );
and ( n5468 , n199 , n35 );
not ( n5469 , n199 );
and ( n5470 , n5469 , n27 );
nor ( n5471 , n5468 , n5470 );
nor ( n5472 , n5471 , n5331 );
and ( n5473 , n199 , n37 );
not ( n5474 , n199 );
and ( n5475 , n5474 , n29 );
nor ( n5476 , n5473 , n5475 );
nor ( n5477 , n5476 , n5331 );
and ( n5478 , n199 , n34 );
not ( n5479 , n199 );
and ( n5480 , n5479 , n26 );
nor ( n5481 , n5478 , n5480 );
nor ( n5482 , n5481 , n4941 );
and ( n5483 , n199 , n36 );
not ( n5484 , n199 );
and ( n5485 , n5484 , n28 );
nor ( n5486 , n5483 , n5485 );
nor ( n5487 , n5486 , n5331 );
and ( n5488 , n199 , n33 );
not ( n5489 , n199 );
and ( n5490 , n5489 , n25 );
nor ( n5491 , n5488 , n5490 );
nor ( n5492 , n5491 , n5331 );
and ( n5493 , n199 , n28 );
not ( n5494 , n199 );
and ( n5495 , n5494 , n20 );
nor ( n5496 , n5493 , n5495 );
nor ( n5497 , n5496 , n5331 );
and ( n5498 , n199 , n29 );
not ( n5499 , n199 );
and ( n5500 , n5499 , n21 );
nor ( n5501 , n5498 , n5500 );
nor ( n5502 , n5501 , n5331 );
and ( n5503 , n199 , n24 );
not ( n5504 , n199 );
and ( n5505 , n5504 , n16 );
nor ( n5506 , n5503 , n5505 );
nor ( n5507 , n5506 , n5331 );
and ( n5508 , n199 , n25 );
not ( n5509 , n199 );
and ( n5510 , n5509 , n17 );
nor ( n5511 , n5508 , n5510 );
nor ( n5512 , n5511 , n5331 );
and ( n5513 , n199 , n26 );
not ( n5514 , n199 );
and ( n5515 , n5514 , n18 );
nor ( n5516 , n5513 , n5515 );
nor ( n5517 , n5516 , n5331 );
and ( n5518 , n199 , n27 );
not ( n5519 , n199 );
and ( n5520 , n5519 , n19 );
nor ( n5521 , n5518 , n5520 );
nor ( n5522 , n5521 , n5331 );
and ( n5523 , n199 , n22 );
not ( n5524 , n199 );
and ( n5525 , n5524 , n14 );
nor ( n5526 , n5523 , n5525 );
nor ( n5527 , n5526 , n4941 );
and ( n5528 , n199 , n23 );
not ( n5529 , n199 );
and ( n5530 , n5529 , n15 );
nor ( n5531 , n5528 , n5530 );
nor ( n5532 , n5531 , n4941 );
and ( n5533 , n199 , n60 );
not ( n5534 , n199 );
and ( n5535 , n5534 , n52 );
nor ( n5536 , n5533 , n5535 );
nor ( n5537 , n5536 , n4941 );
and ( n5538 , n199 , n20 );
not ( n5539 , n199 );
and ( n5540 , n5539 , n12 );
nor ( n5541 , n5538 , n5540 );
nor ( n5542 , n5541 , n4941 );
and ( n5543 , n199 , n52 );
not ( n5544 , n199 );
and ( n5545 , n5544 , n44 );
nor ( n5546 , n5543 , n5545 );
nor ( n5547 , n5546 , n5331 );
and ( n5548 , n199 , n54 );
not ( n5549 , n199 );
and ( n5550 , n5549 , n46 );
nor ( n5551 , n5548 , n5550 );
nor ( n5552 , n5551 , n4941 );
and ( n5553 , n199 , n58 );
not ( n5554 , n199 );
and ( n5555 , n5554 , n50 );
nor ( n5556 , n5553 , n5555 );
nor ( n5557 , n5556 , n5331 );
and ( n5558 , n199 , n46 );
not ( n5559 , n199 );
and ( n5560 , n5559 , n38 );
nor ( n5561 , n5558 , n5560 );
nor ( n5562 , n5561 , n4941 );
and ( n5563 , n199 , n31 );
not ( n5564 , n199 );
and ( n5565 , n5564 , n23 );
nor ( n5566 , n5563 , n5565 );
nor ( n5567 , n5566 , n505 );
and ( n5568 , n199 , n39 );
not ( n5569 , n199 );
and ( n5570 , n5569 , n31 );
nor ( n5571 , n5568 , n5570 );
nor ( n5572 , n5571 , n505 );
and ( n5573 , n199 , n2 );
not ( n5574 , n199 );
and ( n5575 , n5574 , n61 );
nor ( n5576 , n5573 , n5575 );
nor ( n5577 , n5576 , n505 );
and ( n5578 , n199 , n65 );
not ( n5579 , n199 );
and ( n5580 , n5579 , n57 );
nor ( n5581 , n5578 , n5580 );
nor ( n5582 , n5581 , n505 );
and ( n5583 , n199 , n1 );
not ( n5584 , n199 );
and ( n5585 , n5584 , n60 );
nor ( n5586 , n5583 , n5585 );
nor ( n5587 , n5586 , n505 );
and ( n5588 , n199 , n6 );
not ( n5589 , n199 );
and ( n5590 , n5589 , n65 );
nor ( n5591 , n5588 , n5590 );
nor ( n5592 , n5591 , n505 );
and ( n5593 , n199 , n63 );
not ( n5594 , n199 );
and ( n5595 , n5594 , n55 );
nor ( n5596 , n5593 , n5595 );
nor ( n5597 , n5596 , n505 );
and ( n5598 , n199 , n38 );
not ( n5599 , n199 );
and ( n5600 , n5599 , n30 );
nor ( n5601 , n5598 , n5600 );
nor ( n5602 , n5601 , n505 );
endmodule
