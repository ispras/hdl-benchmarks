module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
output n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
 n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
 n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
 n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
 n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
 n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
 n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
 n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
 n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
 n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
 n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
 n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
 n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
wire n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
 n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
 n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
 n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
 n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
 n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
 n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
 n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
 n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
 n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
 n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
 n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
 n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
 n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
 n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
 n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
 n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
 n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
 n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
 n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
 n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , 
 n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
 n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , 
 n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , 
 n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , 
 n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , 
 n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , 
 n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , 
 n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , 
 n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , 
 n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , 
 n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , 
 n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , 
 n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , 
 n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , 
 n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , 
 n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , 
 n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , 
 n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
 n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , 
 n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
 n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , 
 n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , 
 n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , 
 n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
 n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
 n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
 n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , 
 n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , 
 n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , 
 n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
 n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , 
 n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , 
 n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , 
 n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
 n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
 n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
 n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , 
 n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , 
 n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
 n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , 
 n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , 
 n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , 
 n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
 n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
 n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , 
 n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
 n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
 n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , 
 n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , 
 n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , 
 n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , 
 n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , 
 n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , 
 n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , 
 n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
 n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , 
 n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , 
 n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , 
 n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , 
 n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , 
 n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , 
 n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , 
 n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , 
 n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , 
 n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , 
 n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
 n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , 
 n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , 
 n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , 
 n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
 n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
 n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , 
 n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , 
 n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , 
 n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , 
 n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , 
 n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , 
 n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , 
 n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , 
 n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , 
 n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , 
 n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , 
 n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
 n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
 n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
 n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
 n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
 n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
 n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , 
 n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , 
 n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , 
 n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
 n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
 n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
 n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
 n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
 n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
 n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
 n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
 n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
 n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
 n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
 n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
 n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
 n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , 
 n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , 
 n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , 
 n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , 
 n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , 
 n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
 n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , 
 n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , 
 n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , 
 n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , 
 n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
 n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
 n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
 n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , 
 n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , 
 n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , 
 n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , 
 n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
 n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , 
 n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , 
 n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , 
 n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , 
 n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , 
 n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , 
 n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , 
 n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , 
 n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , 
 n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , 
 n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , 
 n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
 n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , 
 n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , 
 n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , 
 n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , 
 n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , 
 n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , 
 n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , 
 n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , 
 n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , 
 n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , 
 n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , 
 n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , 
 n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , 
 n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , 
 n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
 n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , 
 n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
 n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , 
 n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , 
 n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , 
 n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , 
 n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
 n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , 
 n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , 
 n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , 
 n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , 
 n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , 
 n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , 
 n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
 n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
 n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , 
 n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , 
 n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , 
 n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , 
 n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , 
 n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
 n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , 
 n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , 
 n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , 
 n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , 
 n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , 
 n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , 
 n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , 
 n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , 
 n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , 
 n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
 n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
 n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , 
 n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , 
 n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , 
 n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , 
 n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , 
 n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , 
 n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , 
 n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , 
 n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
 n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
 n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , 
 n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , 
 n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
 n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
 n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
 n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
 n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , 
 n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , 
 n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , 
 n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , 
 n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , 
 n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , 
 n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , 
 n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , 
 n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , 
 n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , 
 n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , 
 n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , 
 n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , 
 n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , 
 n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , 
 n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , 
 n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , 
 n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , 
 n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , 
 n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , 
 n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , 
 n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , 
 n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , 
 n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , 
 n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , 
 n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , 
 n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , 
 n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , 
 n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , 
 n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , 
 n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , 
 n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , 
 n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , 
 n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , 
 n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , 
 n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , 
 n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , 
 n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , 
 n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , 
 n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , 
 n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , 
 n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , 
 n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , 
 n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , 
 n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
 n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
 n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , 
 n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , 
 n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , 
 n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , 
 n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , 
 n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , 
 n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , 
 n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , 
 n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , 
 n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , 
 n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , 
 n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , 
 n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , 
 n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , 
 n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , 
 n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , 
 n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , 
 n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , 
 n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , 
 n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , 
 n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , 
 n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , 
 n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , 
 n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , 
 n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , 
 n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , 
 n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , 
 n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
 n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , 
 n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
 n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
 n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
 n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
 n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , 
 n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
 n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , 
 n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
 n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , 
 n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , 
 n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , 
 n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , 
 n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , 
 n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , 
 n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , 
 n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , 
 n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , 
 n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , 
 n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , 
 n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , 
 n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , 
 n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , 
 n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , 
 n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
 n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
 n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
 n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , 
 n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , 
 n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , 
 n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , 
 n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , 
 n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , 
 n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , 
 n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
 n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , 
 n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
 n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
 n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
 n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
 n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
 n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
 n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
 n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , 
 n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , 
 n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
 n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , 
 n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
 n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
 n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
 n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
 n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
 n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , 
 n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , 
 n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , 
 n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , 
 n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , 
 n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
 n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , 
 n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , 
 n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , 
 n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , 
 n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , 
 n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , 
 n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , 
 n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , 
 n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , 
 n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
 n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , 
 n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , 
 n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , 
 n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , 
 n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , 
 n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , 
 n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , 
 n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , 
 n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , 
 n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , 
 n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , 
 n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , 
 n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , 
 n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , 
 n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , 
 n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , 
 n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , 
 n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , 
 n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , 
 n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , 
 n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , 
 n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , 
 n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , 
 n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , 
 n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , 
 n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , 
 n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , 
 n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , 
 n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , 
 n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , 
 n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , 
 n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , 
 n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , 
 n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , 
 n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , 
 n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , 
 n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , 
 n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , 
 n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , 
 n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , 
 n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , 
 n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , 
 n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , 
 n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , 
 n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , 
 n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , 
 n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , 
 n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , 
 n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , 
 n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , 
 n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , 
 n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , 
 n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , 
 n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , 
 n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , 
 n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , 
 n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , 
 n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , 
 n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , 
 n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , 
 n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , 
 n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , 
 n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , 
 n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , 
 n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , 
 n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , 
 n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
 n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , 
 n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , 
 n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , 
 n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , 
 n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , 
 n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , 
 n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
 n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , 
 n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , 
 n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
 n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
 n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , 
 n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , 
 n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , 
 n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , 
 n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , 
 n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , 
 n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , 
 n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , 
 n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , 
 n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , 
 n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , 
 n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
 n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , 
 n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , 
 n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , 
 n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , 
 n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , 
 n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , 
 n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , 
 n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , 
 n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , 
 n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , 
 n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , 
 n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , 
 n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , 
 n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , 
 n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , 
 n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , 
 n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , 
 n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , 
 n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , 
 n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , 
 n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , 
 n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , 
 n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , 
 n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , 
 n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , 
 n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , 
 n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , 
 n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , 
 n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , 
 n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , 
 n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , 
 n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , 
 n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , 
 n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , 
 n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , 
 n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , 
 n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , 
 n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , 
 n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , 
 n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , 
 n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , 
 n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , 
 n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , 
 n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , 
 n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , 
 n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , 
 n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , 
 n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , 
 n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , 
 n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , 
 n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , 
 n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , 
 n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , 
 n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , 
 n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , 
 n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , 
 n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , 
 n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , 
 n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , 
 n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , 
 n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , 
 n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , 
 n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , 
 n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , 
 n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , 
 n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , 
 n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , 
 n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , 
 n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , 
 n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , 
 n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
 n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
 n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , 
 n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , 
 n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , 
 n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , 
 n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , 
 n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , 
 n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , 
 n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , 
 n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , 
 n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , 
 n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , 
 n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , 
 n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , 
 n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , 
 n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , 
 n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , 
 n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , 
 n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , 
 n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , 
 n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , 
 n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , 
 n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , 
 n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , 
 n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , 
 n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , 
 n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , 
 n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , 
 n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , 
 n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , 
 n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , 
 n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , 
 n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , 
 n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , 
 n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , 
 n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , 
 n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , 
 n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , 
 n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , 
 n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , 
 n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , 
 n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , 
 n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , 
 n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , 
 n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , 
 n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , 
 n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , 
 n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , 
 n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , 
 n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , 
 n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , 
 n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , 
 n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , 
 n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , 
 n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , 
 n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , 
 n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , 
 n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , 
 n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , 
 n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , 
 n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , 
 n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , 
 n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , 
 n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , 
 n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , 
 n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , 
 n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , 
 n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , 
 n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
 n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , 
 n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , 
 n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , 
 n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , 
 n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , 
 n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , 
 n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , 
 n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , 
 n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
 n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
 n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
 n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
 n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
 n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , 
 n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , 
 n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , 
 n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , 
 n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , 
 n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , 
 n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , 
 n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , 
 n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , 
 n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , 
 n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , 
 n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , 
 n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , 
 n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , 
 n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , 
 n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , 
 n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
 n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
 n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , 
 n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , 
 n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , 
 n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , 
 n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , 
 n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , 
 n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , 
 n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , 
 n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , 
 n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , 
 n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , 
 n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , 
 n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , 
 n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , 
 n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , 
 n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , 
 n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , 
 n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , 
 n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , 
 n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , 
 n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , 
 n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , 
 n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , 
 n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , 
 n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , 
 n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , 
 n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , 
 n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , 
 n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , 
 n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , 
 n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , 
 n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , 
 n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , 
 n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , 
 n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , 
 n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , 
 n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
 n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
 n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
 n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , 
 n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , 
 n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , 
 n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , 
 n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , 
 n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , 
 n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , 
 n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , 
 n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , 
 n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , 
 n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , 
 n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , 
 n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , 
 n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
 n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , 
 n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , 
 n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , 
 n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , 
 n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , 
 n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , 
 n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , 
 n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
 n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
 n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
 n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
 n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , 
 n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , 
 n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
 n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
 n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
 n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
 n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
 n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
 n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
 n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
 n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
 n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
 n7645 , n7646 , C0n , C0 ;
buf ( n454 , n0 );
buf ( n455 , n1 );
buf ( n456 , n2 );
buf ( n457 , n3 );
buf ( n458 , n4 );
buf ( n459 , n5 );
buf ( n460 , n6 );
buf ( n461 , n7 );
buf ( n462 , n8 );
buf ( n463 , n9 );
buf ( n464 , n10 );
buf ( n465 , n11 );
buf ( n466 , n12 );
buf ( n467 , n13 );
buf ( n468 , n14 );
buf ( n469 , n15 );
buf ( n470 , n16 );
buf ( n471 , n17 );
buf ( n472 , n18 );
buf ( n473 , n19 );
buf ( n474 , n20 );
buf ( n475 , n21 );
buf ( n476 , n22 );
buf ( n477 , n23 );
buf ( n478 , n24 );
buf ( n479 , n25 );
buf ( n480 , n26 );
buf ( n481 , n27 );
buf ( n482 , n28 );
buf ( n483 , n29 );
buf ( n484 , n30 );
buf ( n485 , n31 );
buf ( n486 , n32 );
buf ( n487 , n33 );
buf ( n488 , n34 );
buf ( n489 , n35 );
buf ( n490 , n36 );
buf ( n491 , n37 );
buf ( n492 , n38 );
buf ( n493 , n39 );
buf ( n494 , n40 );
buf ( n495 , n41 );
buf ( n496 , n42 );
buf ( n497 , n43 );
buf ( n498 , n44 );
buf ( n499 , n45 );
buf ( n500 , n46 );
buf ( n501 , n47 );
buf ( n502 , n48 );
buf ( n503 , n49 );
buf ( n504 , n50 );
buf ( n505 , n51 );
buf ( n506 , n52 );
buf ( n507 , n53 );
buf ( n508 , n54 );
buf ( n509 , n55 );
buf ( n510 , n56 );
buf ( n511 , n57 );
buf ( n512 , n58 );
buf ( n513 , n59 );
buf ( n514 , n60 );
buf ( n515 , n61 );
buf ( n516 , n62 );
buf ( n517 , n63 );
buf ( n518 , n64 );
buf ( n519 , n65 );
buf ( n520 , n66 );
buf ( n521 , n67 );
buf ( n522 , n68 );
buf ( n523 , n69 );
buf ( n524 , n70 );
buf ( n525 , n71 );
buf ( n526 , n72 );
buf ( n527 , n73 );
buf ( n528 , n74 );
buf ( n529 , n75 );
buf ( n530 , n76 );
buf ( n531 , n77 );
buf ( n532 , n78 );
buf ( n533 , n79 );
buf ( n534 , n80 );
buf ( n535 , n81 );
buf ( n536 , n82 );
buf ( n537 , n83 );
buf ( n538 , n84 );
buf ( n539 , n85 );
buf ( n540 , n86 );
buf ( n541 , n87 );
buf ( n542 , n88 );
buf ( n543 , n89 );
buf ( n544 , n90 );
buf ( n545 , n91 );
buf ( n546 , n92 );
buf ( n547 , n93 );
buf ( n548 , n94 );
buf ( n549 , n95 );
buf ( n550 , n96 );
buf ( n551 , n97 );
buf ( n552 , n98 );
buf ( n99 , n553 );
buf ( n100 , n554 );
buf ( n101 , n555 );
buf ( n102 , n556 );
buf ( n103 , n557 );
buf ( n104 , n558 );
buf ( n105 , n559 );
buf ( n106 , n560 );
buf ( n107 , n561 );
buf ( n108 , n562 );
buf ( n109 , n563 );
buf ( n110 , n564 );
buf ( n111 , n565 );
buf ( n112 , n566 );
buf ( n113 , n567 );
buf ( n114 , n568 );
buf ( n115 , n569 );
buf ( n116 , n570 );
buf ( n117 , n571 );
buf ( n118 , n572 );
buf ( n119 , n573 );
buf ( n120 , n574 );
buf ( n121 , n575 );
buf ( n122 , n576 );
buf ( n123 , n577 );
buf ( n124 , n578 );
buf ( n125 , n579 );
buf ( n126 , n580 );
buf ( n127 , n581 );
buf ( n128 , n582 );
buf ( n129 , n583 );
buf ( n130 , n584 );
buf ( n131 , n585 );
buf ( n132 , n586 );
buf ( n133 , n587 );
buf ( n134 , n588 );
buf ( n135 , n589 );
buf ( n136 , n590 );
buf ( n137 , n591 );
buf ( n138 , n592 );
buf ( n139 , n593 );
buf ( n140 , n594 );
buf ( n141 , n595 );
buf ( n142 , n596 );
buf ( n143 , n597 );
buf ( n144 , n598 );
buf ( n145 , n599 );
buf ( n146 , n600 );
buf ( n147 , n601 );
buf ( n148 , n602 );
buf ( n149 , n603 );
buf ( n150 , n604 );
buf ( n151 , n605 );
buf ( n152 , n606 );
buf ( n153 , n607 );
buf ( n154 , n608 );
buf ( n155 , n609 );
buf ( n156 , n610 );
buf ( n157 , n611 );
buf ( n158 , n612 );
buf ( n159 , n613 );
buf ( n160 , n614 );
buf ( n161 , n615 );
buf ( n162 , n616 );
buf ( n163 , n617 );
buf ( n164 , n618 );
buf ( n165 , n619 );
buf ( n166 , n620 );
buf ( n167 , n621 );
buf ( n168 , n622 );
buf ( n169 , n623 );
buf ( n170 , n624 );
buf ( n171 , n625 );
buf ( n172 , n626 );
buf ( n173 , n627 );
buf ( n174 , n628 );
buf ( n175 , n629 );
buf ( n176 , n630 );
buf ( n177 , n631 );
buf ( n178 , n632 );
buf ( n179 , n633 );
buf ( n180 , n634 );
buf ( n181 , n635 );
buf ( n182 , n636 );
buf ( n183 , n637 );
buf ( n184 , n638 );
buf ( n185 , n639 );
buf ( n186 , n640 );
buf ( n187 , n641 );
buf ( n188 , n642 );
buf ( n189 , n643 );
buf ( n190 , n644 );
buf ( n191 , n645 );
buf ( n192 , n646 );
buf ( n193 , n647 );
buf ( n194 , n648 );
buf ( n195 , n649 );
buf ( n196 , n650 );
buf ( n197 , n651 );
buf ( n198 , n652 );
buf ( n199 , n653 );
buf ( n200 , n654 );
buf ( n201 , n655 );
buf ( n202 , n656 );
buf ( n203 , n657 );
buf ( n204 , n658 );
buf ( n205 , n659 );
buf ( n206 , n660 );
buf ( n207 , n661 );
buf ( n208 , n662 );
buf ( n209 , n663 );
buf ( n210 , n664 );
buf ( n211 , n665 );
buf ( n212 , n666 );
buf ( n213 , n667 );
buf ( n214 , n668 );
buf ( n215 , n669 );
buf ( n216 , n670 );
buf ( n217 , n671 );
buf ( n218 , n672 );
buf ( n219 , n673 );
buf ( n220 , n674 );
buf ( n221 , n675 );
buf ( n222 , n676 );
buf ( n223 , n677 );
buf ( n224 , n678 );
buf ( n225 , n679 );
buf ( n226 , n680 );
buf ( n553 , C0 );
buf ( n554 , C0 );
buf ( n555 , C0 );
buf ( n556 , C0 );
buf ( n557 , C0 );
buf ( n558 , C0 );
buf ( n559 , C0 );
buf ( n560 , C0 );
buf ( n561 , C0 );
buf ( n562 , C0 );
buf ( n563 , C0 );
buf ( n564 , C0 );
buf ( n565 , C0 );
buf ( n566 , C0 );
buf ( n567 , C0 );
buf ( n568 , C0 );
buf ( n569 , C0 );
buf ( n570 , C0 );
buf ( n571 , C0 );
buf ( n572 , C0 );
buf ( n573 , C0 );
buf ( n574 , C0 );
buf ( n575 , C0 );
buf ( n576 , C0 );
buf ( n577 , C0 );
buf ( n578 , C0 );
buf ( n579 , C0 );
buf ( n580 , C0 );
buf ( n581 , C0 );
buf ( n582 , C0 );
buf ( n583 , C0 );
buf ( n584 , n7547 );
buf ( n585 , n7496 );
buf ( n586 , n7433 );
buf ( n587 , n7360 );
buf ( n588 , n7275 );
buf ( n589 , n7178 );
buf ( n590 , n7071 );
buf ( n591 , n6954 );
buf ( n592 , n6827 );
buf ( n593 , n6690 );
buf ( n594 , n6546 );
buf ( n595 , n6400 );
buf ( n596 , n6247 );
buf ( n597 , n6085 );
buf ( n598 , n5925 );
buf ( n599 , n5753 );
buf ( n600 , n5594 );
buf ( n601 , n5426 );
buf ( n602 , n5257 );
buf ( n603 , n5098 );
buf ( n604 , n4949 );
buf ( n605 , n4810 );
buf ( n606 , n4681 );
buf ( n607 , n4559 );
buf ( n608 , n4445 );
buf ( n609 , n4341 );
buf ( n610 , n4249 );
buf ( n611 , n4170 );
buf ( n612 , n7646 );
buf ( n613 , n7637 );
buf ( n614 , n7628 );
buf ( n615 , n7619 );
buf ( n616 , n7610 );
buf ( n617 , C0 );
buf ( n618 , C0 );
buf ( n619 , C0 );
buf ( n620 , C0 );
buf ( n621 , C0 );
buf ( n622 , C0 );
buf ( n623 , C0 );
buf ( n624 , C0 );
buf ( n625 , C0 );
buf ( n626 , C0 );
buf ( n627 , C0 );
buf ( n628 , C0 );
buf ( n629 , C0 );
buf ( n630 , C0 );
buf ( n631 , C0 );
buf ( n632 , C0 );
buf ( n633 , C0 );
buf ( n634 , C0 );
buf ( n635 , C0 );
buf ( n636 , C0 );
buf ( n637 , C0 );
buf ( n638 , C0 );
buf ( n639 , C0 );
buf ( n640 , C0 );
buf ( n641 , C0 );
buf ( n642 , C0 );
buf ( n643 , C0 );
buf ( n644 , C0 );
buf ( n645 , C0 );
buf ( n646 , C0 );
buf ( n647 , C0 );
buf ( n648 , C0 );
buf ( n649 , C0 );
buf ( n650 , C0 );
buf ( n651 , n7602 );
buf ( n652 , n7583 );
buf ( n653 , n7555 );
buf ( n654 , n7504 );
buf ( n655 , n7441 );
buf ( n656 , n7368 );
buf ( n657 , n7283 );
buf ( n658 , n7186 );
buf ( n659 , n7079 );
buf ( n660 , n6962 );
buf ( n661 , n6835 );
buf ( n662 , n6698 );
buf ( n663 , n6554 );
buf ( n664 , n6408 );
buf ( n665 , n6255 );
buf ( n666 , n6093 );
buf ( n667 , n5933 );
buf ( n668 , n5761 );
buf ( n669 , n5602 );
buf ( n670 , n5434 );
buf ( n671 , n5265 );
buf ( n672 , n5106 );
buf ( n673 , n4957 );
buf ( n674 , n4818 );
buf ( n675 , n4689 );
buf ( n676 , n4570 );
buf ( n677 , n4458 );
buf ( n678 , n4354 );
buf ( n679 , n4259 );
buf ( n680 , n4180 );
buf ( n681 , n520 );
buf ( n682 , n681 );
buf ( n683 , n501 );
buf ( n684 , n683 );
buf ( n685 , n502 );
buf ( n686 , n685 );
xor ( n687 , n684 , n686 );
buf ( n688 , n503 );
buf ( n689 , n688 );
xor ( n690 , n686 , n689 );
not ( n691 , n690 );
and ( n692 , n687 , n691 );
and ( n693 , n682 , n692 );
buf ( n694 , n519 );
buf ( n695 , n694 );
and ( n696 , n695 , n690 );
nor ( n697 , n693 , n696 );
and ( n698 , n686 , n689 );
not ( n699 , n698 );
and ( n700 , n684 , n699 );
xnor ( n701 , n697 , n700 );
buf ( n702 , n518 );
buf ( n703 , n702 );
buf ( n704 , n504 );
buf ( n705 , n704 );
xor ( n706 , n689 , n705 );
not ( n707 , n705 );
and ( n708 , n706 , n707 );
and ( n709 , n703 , n708 );
buf ( n710 , n517 );
buf ( n711 , n710 );
and ( n712 , n711 , n705 );
nor ( n713 , n709 , n712 );
xnor ( n714 , n713 , n689 );
and ( n715 , n682 , n690 );
not ( n716 , n715 );
and ( n717 , n716 , n700 );
xor ( n718 , n714 , n717 );
xor ( n719 , n701 , n718 );
and ( n720 , n695 , n708 );
and ( n721 , n703 , n705 );
nor ( n722 , n720 , n721 );
xnor ( n723 , n722 , n689 );
and ( n724 , n723 , n715 );
xor ( n725 , n723 , n715 );
and ( n726 , n682 , n708 );
and ( n727 , n695 , n705 );
nor ( n728 , n726 , n727 );
xnor ( n729 , n728 , n689 );
and ( n730 , n682 , n705 );
not ( n731 , n730 );
and ( n732 , n731 , n689 );
and ( n733 , n729 , n732 );
and ( n734 , n725 , n733 );
or ( n735 , n724 , n734 );
xor ( n736 , n719 , n735 );
buf ( n737 , n736 );
not ( n738 , n456 );
and ( n739 , n738 , n488 );
and ( n740 , n472 , n456 );
or ( n741 , n739 , n740 );
buf ( n742 , n741 );
buf ( n743 , n742 );
buf ( n744 , n501 );
buf ( n745 , n744 );
buf ( n746 , n502 );
buf ( n747 , n746 );
xor ( n748 , n745 , n747 );
buf ( n749 , n503 );
buf ( n750 , n749 );
xor ( n751 , n747 , n750 );
not ( n752 , n751 );
and ( n753 , n748 , n752 );
and ( n754 , n743 , n753 );
not ( n755 , n456 );
and ( n756 , n755 , n487 );
and ( n757 , n471 , n456 );
or ( n758 , n756 , n757 );
buf ( n759 , n758 );
buf ( n760 , n759 );
and ( n761 , n760 , n751 );
nor ( n762 , n754 , n761 );
and ( n763 , n747 , n750 );
not ( n764 , n763 );
and ( n765 , n745 , n764 );
xnor ( n766 , n762 , n765 );
not ( n767 , n456 );
and ( n768 , n767 , n486 );
and ( n769 , n470 , n456 );
or ( n770 , n768 , n769 );
buf ( n771 , n770 );
buf ( n772 , n771 );
buf ( n773 , n504 );
buf ( n774 , n773 );
xor ( n775 , n750 , n774 );
not ( n776 , n774 );
and ( n777 , n775 , n776 );
and ( n778 , n772 , n777 );
not ( n779 , n456 );
and ( n780 , n779 , n485 );
and ( n781 , n469 , n456 );
or ( n782 , n780 , n781 );
buf ( n783 , n782 );
buf ( n784 , n783 );
and ( n785 , n784 , n774 );
nor ( n786 , n778 , n785 );
xnor ( n787 , n786 , n750 );
and ( n788 , n743 , n751 );
not ( n789 , n788 );
and ( n790 , n789 , n765 );
xor ( n791 , n787 , n790 );
xor ( n792 , n766 , n791 );
and ( n793 , n760 , n777 );
and ( n794 , n772 , n774 );
nor ( n795 , n793 , n794 );
xnor ( n796 , n795 , n750 );
and ( n797 , n796 , n788 );
xor ( n798 , n796 , n788 );
and ( n799 , n743 , n777 );
and ( n800 , n760 , n774 );
nor ( n801 , n799 , n800 );
xnor ( n802 , n801 , n750 );
and ( n803 , n743 , n774 );
not ( n804 , n803 );
and ( n805 , n804 , n750 );
and ( n806 , n802 , n805 );
and ( n807 , n798 , n806 );
or ( n808 , n797 , n807 );
xor ( n809 , n792 , n808 );
buf ( n810 , n809 );
not ( n811 , n455 );
and ( n812 , n811 , n737 );
and ( n813 , n810 , n455 );
or ( n814 , n812 , n813 );
and ( n815 , n711 , n708 );
buf ( n816 , n516 );
buf ( n817 , n816 );
and ( n818 , n817 , n705 );
nor ( n819 , n815 , n818 );
xnor ( n820 , n819 , n689 );
and ( n821 , n695 , n692 );
and ( n822 , n703 , n690 );
nor ( n823 , n821 , n822 );
xnor ( n824 , n823 , n700 );
xor ( n825 , n820 , n824 );
buf ( n826 , n500 );
buf ( n827 , n826 );
xor ( n828 , n827 , n684 );
and ( n829 , n682 , n828 );
xor ( n830 , n825 , n829 );
and ( n831 , n714 , n717 );
xor ( n832 , n830 , n831 );
and ( n833 , n701 , n718 );
and ( n834 , n719 , n735 );
or ( n835 , n833 , n834 );
xor ( n836 , n832 , n835 );
buf ( n837 , n836 );
and ( n838 , n784 , n777 );
not ( n839 , n456 );
and ( n840 , n839 , n484 );
and ( n841 , n468 , n456 );
or ( n842 , n840 , n841 );
buf ( n843 , n842 );
buf ( n844 , n843 );
and ( n845 , n844 , n774 );
nor ( n846 , n838 , n845 );
xnor ( n847 , n846 , n750 );
and ( n848 , n760 , n753 );
and ( n849 , n772 , n751 );
nor ( n850 , n848 , n849 );
xnor ( n851 , n850 , n765 );
xor ( n852 , n847 , n851 );
buf ( n853 , n500 );
buf ( n854 , n853 );
xor ( n855 , n854 , n745 );
and ( n856 , n743 , n855 );
xor ( n857 , n852 , n856 );
and ( n858 , n787 , n790 );
xor ( n859 , n857 , n858 );
and ( n860 , n766 , n791 );
and ( n861 , n792 , n808 );
or ( n862 , n860 , n861 );
xor ( n863 , n859 , n862 );
buf ( n864 , n863 );
not ( n865 , n455 );
and ( n866 , n865 , n837 );
and ( n867 , n864 , n455 );
or ( n868 , n866 , n867 );
and ( n869 , n820 , n824 );
and ( n870 , n824 , n829 );
and ( n871 , n820 , n829 );
or ( n872 , n869 , n870 , n871 );
and ( n873 , n817 , n708 );
buf ( n874 , n515 );
buf ( n875 , n874 );
and ( n876 , n875 , n705 );
nor ( n877 , n873 , n876 );
xnor ( n878 , n877 , n689 );
not ( n879 , n829 );
buf ( n880 , n499 );
buf ( n881 , n880 );
and ( n882 , n827 , n684 );
not ( n883 , n882 );
and ( n884 , n881 , n883 );
and ( n885 , n879 , n884 );
xor ( n886 , n878 , n885 );
and ( n887 , n703 , n692 );
and ( n888 , n711 , n690 );
nor ( n889 , n887 , n888 );
xnor ( n890 , n889 , n700 );
xor ( n891 , n886 , n890 );
xor ( n892 , n881 , n827 );
not ( n893 , n828 );
and ( n894 , n892 , n893 );
and ( n895 , n682 , n894 );
and ( n896 , n695 , n828 );
nor ( n897 , n895 , n896 );
xnor ( n898 , n897 , n884 );
xor ( n899 , n891 , n898 );
xor ( n900 , n872 , n899 );
and ( n901 , n830 , n831 );
and ( n902 , n832 , n835 );
or ( n903 , n901 , n902 );
xor ( n904 , n900 , n903 );
buf ( n905 , n904 );
and ( n906 , n847 , n851 );
and ( n907 , n851 , n856 );
and ( n908 , n847 , n856 );
or ( n909 , n906 , n907 , n908 );
and ( n910 , n844 , n777 );
not ( n911 , n456 );
and ( n912 , n911 , n483 );
and ( n913 , n467 , n456 );
or ( n914 , n912 , n913 );
buf ( n915 , n914 );
buf ( n916 , n915 );
and ( n917 , n916 , n774 );
nor ( n918 , n910 , n917 );
xnor ( n919 , n918 , n750 );
not ( n920 , n856 );
buf ( n921 , n499 );
buf ( n922 , n921 );
and ( n923 , n854 , n745 );
not ( n924 , n923 );
and ( n925 , n922 , n924 );
and ( n926 , n920 , n925 );
xor ( n927 , n919 , n926 );
and ( n928 , n772 , n753 );
and ( n929 , n784 , n751 );
nor ( n930 , n928 , n929 );
xnor ( n931 , n930 , n765 );
xor ( n932 , n927 , n931 );
xor ( n933 , n922 , n854 );
not ( n934 , n855 );
and ( n935 , n933 , n934 );
and ( n936 , n743 , n935 );
and ( n937 , n760 , n855 );
nor ( n938 , n936 , n937 );
xnor ( n939 , n938 , n925 );
xor ( n940 , n932 , n939 );
xor ( n941 , n909 , n940 );
and ( n942 , n857 , n858 );
and ( n943 , n859 , n862 );
or ( n944 , n942 , n943 );
xor ( n945 , n941 , n944 );
buf ( n946 , n945 );
not ( n947 , n455 );
and ( n948 , n947 , n905 );
and ( n949 , n946 , n455 );
or ( n950 , n948 , n949 );
and ( n951 , n878 , n885 );
and ( n952 , n695 , n894 );
and ( n953 , n703 , n828 );
nor ( n954 , n952 , n953 );
xnor ( n955 , n954 , n884 );
xor ( n956 , n951 , n955 );
and ( n957 , n875 , n708 );
buf ( n958 , n514 );
buf ( n959 , n958 );
and ( n960 , n959 , n705 );
nor ( n961 , n957 , n960 );
xnor ( n962 , n961 , n689 );
and ( n963 , n711 , n692 );
and ( n964 , n817 , n690 );
nor ( n965 , n963 , n964 );
xnor ( n966 , n965 , n700 );
xor ( n967 , n962 , n966 );
buf ( n968 , n498 );
buf ( n969 , n968 );
xor ( n970 , n969 , n881 );
and ( n971 , n682 , n970 );
xor ( n972 , n967 , n971 );
xor ( n973 , n956 , n972 );
and ( n974 , n886 , n890 );
and ( n975 , n890 , n898 );
and ( n976 , n886 , n898 );
or ( n977 , n974 , n975 , n976 );
xor ( n978 , n973 , n977 );
and ( n979 , n872 , n899 );
and ( n980 , n900 , n903 );
or ( n981 , n979 , n980 );
xor ( n982 , n978 , n981 );
buf ( n983 , n982 );
and ( n984 , n919 , n926 );
and ( n985 , n760 , n935 );
and ( n986 , n772 , n855 );
nor ( n987 , n985 , n986 );
xnor ( n988 , n987 , n925 );
xor ( n989 , n984 , n988 );
and ( n990 , n916 , n777 );
not ( n991 , n456 );
and ( n992 , n991 , n482 );
and ( n993 , n466 , n456 );
or ( n994 , n992 , n993 );
buf ( n995 , n994 );
buf ( n996 , n995 );
and ( n997 , n996 , n774 );
nor ( n998 , n990 , n997 );
xnor ( n999 , n998 , n750 );
and ( n1000 , n784 , n753 );
and ( n1001 , n844 , n751 );
nor ( n1002 , n1000 , n1001 );
xnor ( n1003 , n1002 , n765 );
xor ( n1004 , n999 , n1003 );
buf ( n1005 , n498 );
buf ( n1006 , n1005 );
xor ( n1007 , n1006 , n922 );
and ( n1008 , n743 , n1007 );
xor ( n1009 , n1004 , n1008 );
xor ( n1010 , n989 , n1009 );
and ( n1011 , n927 , n931 );
and ( n1012 , n931 , n939 );
and ( n1013 , n927 , n939 );
or ( n1014 , n1011 , n1012 , n1013 );
xor ( n1015 , n1010 , n1014 );
and ( n1016 , n909 , n940 );
and ( n1017 , n941 , n944 );
or ( n1018 , n1016 , n1017 );
xor ( n1019 , n1015 , n1018 );
buf ( n1020 , n1019 );
not ( n1021 , n455 );
and ( n1022 , n1021 , n983 );
and ( n1023 , n1020 , n455 );
or ( n1024 , n1022 , n1023 );
and ( n1025 , n959 , n708 );
buf ( n1026 , n513 );
buf ( n1027 , n1026 );
and ( n1028 , n1027 , n705 );
nor ( n1029 , n1025 , n1028 );
xnor ( n1030 , n1029 , n689 );
not ( n1031 , n971 );
buf ( n1032 , n497 );
buf ( n1033 , n1032 );
and ( n1034 , n969 , n881 );
not ( n1035 , n1034 );
and ( n1036 , n1033 , n1035 );
and ( n1037 , n1031 , n1036 );
xor ( n1038 , n1030 , n1037 );
and ( n1039 , n962 , n966 );
and ( n1040 , n966 , n971 );
and ( n1041 , n962 , n971 );
or ( n1042 , n1039 , n1040 , n1041 );
xor ( n1043 , n1038 , n1042 );
and ( n1044 , n817 , n692 );
and ( n1045 , n875 , n690 );
nor ( n1046 , n1044 , n1045 );
xnor ( n1047 , n1046 , n700 );
and ( n1048 , n703 , n894 );
and ( n1049 , n711 , n828 );
nor ( n1050 , n1048 , n1049 );
xnor ( n1051 , n1050 , n884 );
xor ( n1052 , n1047 , n1051 );
xor ( n1053 , n1033 , n969 );
not ( n1054 , n970 );
and ( n1055 , n1053 , n1054 );
and ( n1056 , n682 , n1055 );
and ( n1057 , n695 , n970 );
nor ( n1058 , n1056 , n1057 );
xnor ( n1059 , n1058 , n1036 );
xor ( n1060 , n1052 , n1059 );
xor ( n1061 , n1043 , n1060 );
and ( n1062 , n951 , n955 );
and ( n1063 , n955 , n972 );
and ( n1064 , n951 , n972 );
or ( n1065 , n1062 , n1063 , n1064 );
xor ( n1066 , n1061 , n1065 );
and ( n1067 , n973 , n977 );
and ( n1068 , n978 , n981 );
or ( n1069 , n1067 , n1068 );
xor ( n1070 , n1066 , n1069 );
buf ( n1071 , n1070 );
and ( n1072 , n999 , n1003 );
and ( n1073 , n1003 , n1008 );
and ( n1074 , n999 , n1008 );
or ( n1075 , n1072 , n1073 , n1074 );
and ( n1076 , n984 , n988 );
and ( n1077 , n988 , n1009 );
and ( n1078 , n984 , n1009 );
or ( n1079 , n1076 , n1077 , n1078 );
xor ( n1080 , n1075 , n1079 );
and ( n1081 , n996 , n777 );
not ( n1082 , n456 );
and ( n1083 , n1082 , n481 );
and ( n1084 , n465 , n456 );
or ( n1085 , n1083 , n1084 );
buf ( n1086 , n1085 );
buf ( n1087 , n1086 );
and ( n1088 , n1087 , n774 );
nor ( n1089 , n1081 , n1088 );
xnor ( n1090 , n1089 , n750 );
not ( n1091 , n1008 );
buf ( n1092 , n497 );
buf ( n1093 , n1092 );
and ( n1094 , n1006 , n922 );
not ( n1095 , n1094 );
and ( n1096 , n1093 , n1095 );
and ( n1097 , n1091 , n1096 );
xor ( n1098 , n1090 , n1097 );
and ( n1099 , n844 , n753 );
and ( n1100 , n916 , n751 );
nor ( n1101 , n1099 , n1100 );
xnor ( n1102 , n1101 , n765 );
and ( n1103 , n772 , n935 );
and ( n1104 , n784 , n855 );
nor ( n1105 , n1103 , n1104 );
xnor ( n1106 , n1105 , n925 );
xor ( n1107 , n1102 , n1106 );
xor ( n1108 , n1093 , n1006 );
not ( n1109 , n1007 );
and ( n1110 , n1108 , n1109 );
and ( n1111 , n743 , n1110 );
and ( n1112 , n760 , n1007 );
nor ( n1113 , n1111 , n1112 );
xnor ( n1114 , n1113 , n1096 );
xor ( n1115 , n1107 , n1114 );
xor ( n1116 , n1098 , n1115 );
xor ( n1117 , n1080 , n1116 );
and ( n1118 , n1010 , n1014 );
and ( n1119 , n1015 , n1018 );
or ( n1120 , n1118 , n1119 );
xor ( n1121 , n1117 , n1120 );
buf ( n1122 , n1121 );
not ( n1123 , n455 );
and ( n1124 , n1123 , n1071 );
and ( n1125 , n1122 , n455 );
or ( n1126 , n1124 , n1125 );
and ( n1127 , n1038 , n1042 );
and ( n1128 , n1042 , n1060 );
and ( n1129 , n1038 , n1060 );
or ( n1130 , n1127 , n1128 , n1129 );
and ( n1131 , n1047 , n1051 );
and ( n1132 , n1051 , n1059 );
and ( n1133 , n1047 , n1059 );
or ( n1134 , n1131 , n1132 , n1133 );
and ( n1135 , n1027 , n708 );
buf ( n1136 , n512 );
buf ( n1137 , n1136 );
and ( n1138 , n1137 , n705 );
nor ( n1139 , n1135 , n1138 );
xnor ( n1140 , n1139 , n689 );
and ( n1141 , n695 , n1055 );
and ( n1142 , n703 , n970 );
nor ( n1143 , n1141 , n1142 );
xnor ( n1144 , n1143 , n1036 );
xor ( n1145 , n1140 , n1144 );
buf ( n1146 , n496 );
buf ( n1147 , n1146 );
xor ( n1148 , n1147 , n1033 );
and ( n1149 , n682 , n1148 );
xor ( n1150 , n1145 , n1149 );
xor ( n1151 , n1134 , n1150 );
and ( n1152 , n1030 , n1037 );
and ( n1153 , n875 , n692 );
and ( n1154 , n959 , n690 );
nor ( n1155 , n1153 , n1154 );
xnor ( n1156 , n1155 , n700 );
xor ( n1157 , n1152 , n1156 );
and ( n1158 , n711 , n894 );
and ( n1159 , n817 , n828 );
nor ( n1160 , n1158 , n1159 );
xnor ( n1161 , n1160 , n884 );
xor ( n1162 , n1157 , n1161 );
xor ( n1163 , n1151 , n1162 );
xor ( n1164 , n1130 , n1163 );
and ( n1165 , n1061 , n1065 );
and ( n1166 , n1066 , n1069 );
or ( n1167 , n1165 , n1166 );
xor ( n1168 , n1164 , n1167 );
buf ( n1169 , n1168 );
and ( n1170 , n1075 , n1079 );
and ( n1171 , n1079 , n1116 );
and ( n1172 , n1075 , n1116 );
or ( n1173 , n1170 , n1171 , n1172 );
and ( n1174 , n1102 , n1106 );
and ( n1175 , n1106 , n1114 );
and ( n1176 , n1102 , n1114 );
or ( n1177 , n1174 , n1175 , n1176 );
and ( n1178 , n1090 , n1097 );
and ( n1179 , n1097 , n1115 );
and ( n1180 , n1090 , n1115 );
or ( n1181 , n1178 , n1179 , n1180 );
xor ( n1182 , n1177 , n1181 );
and ( n1183 , n1087 , n777 );
not ( n1184 , n456 );
and ( n1185 , n1184 , n480 );
and ( n1186 , n464 , n456 );
or ( n1187 , n1185 , n1186 );
buf ( n1188 , n1187 );
buf ( n1189 , n1188 );
and ( n1190 , n1189 , n774 );
nor ( n1191 , n1183 , n1190 );
xnor ( n1192 , n1191 , n750 );
and ( n1193 , n760 , n1110 );
and ( n1194 , n772 , n1007 );
nor ( n1195 , n1193 , n1194 );
xnor ( n1196 , n1195 , n1096 );
buf ( n1197 , n496 );
buf ( n1198 , n1197 );
xor ( n1199 , n1198 , n1093 );
and ( n1200 , n743 , n1199 );
xor ( n1201 , n1196 , n1200 );
xor ( n1202 , n1192 , n1201 );
and ( n1203 , n916 , n753 );
and ( n1204 , n996 , n751 );
nor ( n1205 , n1203 , n1204 );
xnor ( n1206 , n1205 , n765 );
and ( n1207 , n784 , n935 );
and ( n1208 , n844 , n855 );
nor ( n1209 , n1207 , n1208 );
xnor ( n1210 , n1209 , n925 );
xor ( n1211 , n1206 , n1210 );
xor ( n1212 , n1202 , n1211 );
xor ( n1213 , n1182 , n1212 );
xor ( n1214 , n1173 , n1213 );
and ( n1215 , n1117 , n1120 );
xor ( n1216 , n1214 , n1215 );
buf ( n1217 , n1216 );
not ( n1218 , n455 );
and ( n1219 , n1218 , n1169 );
and ( n1220 , n1217 , n455 );
or ( n1221 , n1219 , n1220 );
and ( n1222 , n1152 , n1156 );
and ( n1223 , n1156 , n1161 );
and ( n1224 , n1152 , n1161 );
or ( n1225 , n1222 , n1223 , n1224 );
and ( n1226 , n1137 , n708 );
buf ( n1227 , n511 );
buf ( n1228 , n1227 );
and ( n1229 , n1228 , n705 );
nor ( n1230 , n1226 , n1229 );
xnor ( n1231 , n1230 , n689 );
and ( n1232 , n703 , n1055 );
and ( n1233 , n711 , n970 );
nor ( n1234 , n1232 , n1233 );
xnor ( n1235 , n1234 , n1036 );
xor ( n1236 , n1231 , n1235 );
buf ( n1237 , n495 );
buf ( n1238 , n1237 );
xor ( n1239 , n1238 , n1147 );
not ( n1240 , n1148 );
and ( n1241 , n1239 , n1240 );
and ( n1242 , n682 , n1241 );
and ( n1243 , n695 , n1148 );
nor ( n1244 , n1242 , n1243 );
and ( n1245 , n1147 , n1033 );
not ( n1246 , n1245 );
and ( n1247 , n1238 , n1246 );
xnor ( n1248 , n1244 , n1247 );
xor ( n1249 , n1236 , n1248 );
xor ( n1250 , n1225 , n1249 );
and ( n1251 , n959 , n692 );
and ( n1252 , n1027 , n690 );
nor ( n1253 , n1251 , n1252 );
xnor ( n1254 , n1253 , n700 );
not ( n1255 , n1149 );
and ( n1256 , n1255 , n1247 );
xor ( n1257 , n1254 , n1256 );
and ( n1258 , n1140 , n1144 );
and ( n1259 , n1144 , n1149 );
and ( n1260 , n1140 , n1149 );
or ( n1261 , n1258 , n1259 , n1260 );
xor ( n1262 , n1257 , n1261 );
and ( n1263 , n817 , n894 );
and ( n1264 , n875 , n828 );
nor ( n1265 , n1263 , n1264 );
xnor ( n1266 , n1265 , n884 );
xor ( n1267 , n1262 , n1266 );
xor ( n1268 , n1250 , n1267 );
and ( n1269 , n1134 , n1150 );
and ( n1270 , n1150 , n1162 );
and ( n1271 , n1134 , n1162 );
or ( n1272 , n1269 , n1270 , n1271 );
xor ( n1273 , n1268 , n1272 );
and ( n1274 , n1130 , n1163 );
and ( n1275 , n1164 , n1167 );
or ( n1276 , n1274 , n1275 );
xor ( n1277 , n1273 , n1276 );
buf ( n1278 , n1277 );
and ( n1279 , n1177 , n1181 );
and ( n1280 , n1181 , n1212 );
and ( n1281 , n1177 , n1212 );
or ( n1282 , n1279 , n1280 , n1281 );
and ( n1283 , n844 , n935 );
and ( n1284 , n916 , n855 );
nor ( n1285 , n1283 , n1284 );
xnor ( n1286 , n1285 , n925 );
and ( n1287 , n996 , n753 );
and ( n1288 , n1087 , n751 );
nor ( n1289 , n1287 , n1288 );
xnor ( n1290 , n1289 , n765 );
not ( n1291 , n1200 );
buf ( n1292 , n495 );
buf ( n1293 , n1292 );
and ( n1294 , n1198 , n1093 );
not ( n1295 , n1294 );
and ( n1296 , n1293 , n1295 );
and ( n1297 , n1291 , n1296 );
xor ( n1298 , n1290 , n1297 );
xor ( n1299 , n1286 , n1298 );
and ( n1300 , n1192 , n1201 );
and ( n1301 , n1201 , n1211 );
and ( n1302 , n1192 , n1211 );
or ( n1303 , n1300 , n1301 , n1302 );
xor ( n1304 , n1299 , n1303 );
and ( n1305 , n1189 , n777 );
not ( n1306 , n456 );
and ( n1307 , n1306 , n479 );
and ( n1308 , n463 , n456 );
or ( n1309 , n1307 , n1308 );
buf ( n1310 , n1309 );
buf ( n1311 , n1310 );
and ( n1312 , n1311 , n774 );
nor ( n1313 , n1305 , n1312 );
xnor ( n1314 , n1313 , n750 );
and ( n1315 , n772 , n1110 );
and ( n1316 , n784 , n1007 );
nor ( n1317 , n1315 , n1316 );
xnor ( n1318 , n1317 , n1096 );
xor ( n1319 , n1314 , n1318 );
xor ( n1320 , n1293 , n1198 );
not ( n1321 , n1199 );
and ( n1322 , n1320 , n1321 );
and ( n1323 , n743 , n1322 );
and ( n1324 , n760 , n1199 );
nor ( n1325 , n1323 , n1324 );
xnor ( n1326 , n1325 , n1296 );
xor ( n1327 , n1319 , n1326 );
and ( n1328 , n1196 , n1200 );
xor ( n1329 , n1327 , n1328 );
and ( n1330 , n1206 , n1210 );
xor ( n1331 , n1329 , n1330 );
xor ( n1332 , n1304 , n1331 );
xor ( n1333 , n1282 , n1332 );
and ( n1334 , n1173 , n1213 );
and ( n1335 , n1214 , n1215 );
or ( n1336 , n1334 , n1335 );
xor ( n1337 , n1333 , n1336 );
buf ( n1338 , n1337 );
not ( n1339 , n455 );
and ( n1340 , n1339 , n1278 );
and ( n1341 , n1338 , n455 );
or ( n1342 , n1340 , n1341 );
and ( n1343 , n1257 , n1261 );
and ( n1344 , n1261 , n1266 );
and ( n1345 , n1257 , n1266 );
or ( n1346 , n1343 , n1344 , n1345 );
and ( n1347 , n1228 , n708 );
buf ( n1348 , n510 );
buf ( n1349 , n1348 );
and ( n1350 , n1349 , n705 );
nor ( n1351 , n1347 , n1350 );
xnor ( n1352 , n1351 , n689 );
and ( n1353 , n875 , n894 );
and ( n1354 , n959 , n828 );
nor ( n1355 , n1353 , n1354 );
xnor ( n1356 , n1355 , n884 );
xor ( n1357 , n1352 , n1356 );
and ( n1358 , n695 , n1241 );
and ( n1359 , n703 , n1148 );
nor ( n1360 , n1358 , n1359 );
xnor ( n1361 , n1360 , n1247 );
xor ( n1362 , n1357 , n1361 );
xor ( n1363 , n1346 , n1362 );
and ( n1364 , n1231 , n1235 );
and ( n1365 , n1235 , n1248 );
and ( n1366 , n1231 , n1248 );
or ( n1367 , n1364 , n1365 , n1366 );
and ( n1368 , n1254 , n1256 );
xor ( n1369 , n1367 , n1368 );
and ( n1370 , n1027 , n692 );
and ( n1371 , n1137 , n690 );
nor ( n1372 , n1370 , n1371 );
xnor ( n1373 , n1372 , n700 );
and ( n1374 , n711 , n1055 );
and ( n1375 , n817 , n970 );
nor ( n1376 , n1374 , n1375 );
xnor ( n1377 , n1376 , n1036 );
xor ( n1378 , n1373 , n1377 );
buf ( n1379 , n494 );
buf ( n1380 , n1379 );
xor ( n1381 , n1380 , n1238 );
and ( n1382 , n682 , n1381 );
xor ( n1383 , n1378 , n1382 );
xor ( n1384 , n1369 , n1383 );
xor ( n1385 , n1363 , n1384 );
and ( n1386 , n1225 , n1249 );
and ( n1387 , n1249 , n1267 );
and ( n1388 , n1225 , n1267 );
or ( n1389 , n1386 , n1387 , n1388 );
xor ( n1390 , n1385 , n1389 );
and ( n1391 , n1268 , n1272 );
and ( n1392 , n1273 , n1276 );
or ( n1393 , n1391 , n1392 );
xor ( n1394 , n1390 , n1393 );
buf ( n1395 , n1394 );
and ( n1396 , n1327 , n1328 );
and ( n1397 , n1328 , n1330 );
and ( n1398 , n1327 , n1330 );
or ( n1399 , n1396 , n1397 , n1398 );
and ( n1400 , n1299 , n1303 );
and ( n1401 , n1303 , n1331 );
and ( n1402 , n1299 , n1331 );
or ( n1403 , n1400 , n1401 , n1402 );
xor ( n1404 , n1399 , n1403 );
and ( n1405 , n1311 , n777 );
not ( n1406 , n456 );
and ( n1407 , n1406 , n478 );
and ( n1408 , n462 , n456 );
or ( n1409 , n1407 , n1408 );
buf ( n1410 , n1409 );
buf ( n1411 , n1410 );
and ( n1412 , n1411 , n774 );
nor ( n1413 , n1405 , n1412 );
xnor ( n1414 , n1413 , n750 );
and ( n1415 , n916 , n935 );
and ( n1416 , n996 , n855 );
nor ( n1417 , n1415 , n1416 );
xnor ( n1418 , n1417 , n925 );
xor ( n1419 , n1414 , n1418 );
and ( n1420 , n760 , n1322 );
and ( n1421 , n772 , n1199 );
nor ( n1422 , n1420 , n1421 );
xnor ( n1423 , n1422 , n1296 );
xor ( n1424 , n1419 , n1423 );
and ( n1425 , n1314 , n1318 );
and ( n1426 , n1318 , n1326 );
and ( n1427 , n1314 , n1326 );
or ( n1428 , n1425 , n1426 , n1427 );
and ( n1429 , n1290 , n1297 );
xor ( n1430 , n1428 , n1429 );
and ( n1431 , n1087 , n753 );
and ( n1432 , n1189 , n751 );
nor ( n1433 , n1431 , n1432 );
xnor ( n1434 , n1433 , n765 );
and ( n1435 , n784 , n1110 );
and ( n1436 , n844 , n1007 );
nor ( n1437 , n1435 , n1436 );
xnor ( n1438 , n1437 , n1096 );
xor ( n1439 , n1434 , n1438 );
buf ( n1440 , n494 );
buf ( n1441 , n1440 );
xor ( n1442 , n1441 , n1293 );
and ( n1443 , n743 , n1442 );
xor ( n1444 , n1439 , n1443 );
xor ( n1445 , n1430 , n1444 );
xor ( n1446 , n1424 , n1445 );
and ( n1447 , n1286 , n1298 );
xor ( n1448 , n1446 , n1447 );
xor ( n1449 , n1404 , n1448 );
and ( n1450 , n1282 , n1332 );
and ( n1451 , n1333 , n1336 );
or ( n1452 , n1450 , n1451 );
xor ( n1453 , n1449 , n1452 );
buf ( n1454 , n1453 );
not ( n1455 , n455 );
and ( n1456 , n1455 , n1395 );
and ( n1457 , n1454 , n455 );
or ( n1458 , n1456 , n1457 );
and ( n1459 , n1367 , n1368 );
and ( n1460 , n1368 , n1383 );
and ( n1461 , n1367 , n1383 );
or ( n1462 , n1459 , n1460 , n1461 );
and ( n1463 , n1137 , n692 );
and ( n1464 , n1228 , n690 );
nor ( n1465 , n1463 , n1464 );
xnor ( n1466 , n1465 , n700 );
not ( n1467 , n1382 );
buf ( n1468 , n493 );
buf ( n1469 , n1468 );
and ( n1470 , n1380 , n1238 );
not ( n1471 , n1470 );
and ( n1472 , n1469 , n1471 );
and ( n1473 , n1467 , n1472 );
xor ( n1474 , n1466 , n1473 );
and ( n1475 , n959 , n894 );
and ( n1476 , n1027 , n828 );
nor ( n1477 , n1475 , n1476 );
xnor ( n1478 , n1477 , n884 );
xor ( n1479 , n1474 , n1478 );
xor ( n1480 , n1469 , n1380 );
not ( n1481 , n1381 );
and ( n1482 , n1480 , n1481 );
and ( n1483 , n682 , n1482 );
and ( n1484 , n695 , n1381 );
nor ( n1485 , n1483 , n1484 );
xnor ( n1486 , n1485 , n1472 );
xor ( n1487 , n1479 , n1486 );
xor ( n1488 , n1462 , n1487 );
and ( n1489 , n1352 , n1356 );
and ( n1490 , n1356 , n1361 );
and ( n1491 , n1352 , n1361 );
or ( n1492 , n1489 , n1490 , n1491 );
and ( n1493 , n1373 , n1377 );
and ( n1494 , n1377 , n1382 );
and ( n1495 , n1373 , n1382 );
or ( n1496 , n1493 , n1494 , n1495 );
xor ( n1497 , n1492 , n1496 );
and ( n1498 , n1349 , n708 );
buf ( n1499 , n509 );
buf ( n1500 , n1499 );
and ( n1501 , n1500 , n705 );
nor ( n1502 , n1498 , n1501 );
xnor ( n1503 , n1502 , n689 );
and ( n1504 , n817 , n1055 );
and ( n1505 , n875 , n970 );
nor ( n1506 , n1504 , n1505 );
xnor ( n1507 , n1506 , n1036 );
xor ( n1508 , n1503 , n1507 );
and ( n1509 , n703 , n1241 );
and ( n1510 , n711 , n1148 );
nor ( n1511 , n1509 , n1510 );
xnor ( n1512 , n1511 , n1247 );
xor ( n1513 , n1508 , n1512 );
xor ( n1514 , n1497 , n1513 );
xor ( n1515 , n1488 , n1514 );
and ( n1516 , n1346 , n1362 );
and ( n1517 , n1362 , n1384 );
and ( n1518 , n1346 , n1384 );
or ( n1519 , n1516 , n1517 , n1518 );
xor ( n1520 , n1515 , n1519 );
and ( n1521 , n1385 , n1389 );
and ( n1522 , n1390 , n1393 );
or ( n1523 , n1521 , n1522 );
xor ( n1524 , n1520 , n1523 );
buf ( n1525 , n1524 );
and ( n1526 , n1424 , n1445 );
and ( n1527 , n1445 , n1447 );
and ( n1528 , n1424 , n1447 );
or ( n1529 , n1526 , n1527 , n1528 );
and ( n1530 , n1428 , n1429 );
and ( n1531 , n1429 , n1444 );
and ( n1532 , n1428 , n1444 );
or ( n1533 , n1530 , n1531 , n1532 );
and ( n1534 , n772 , n1322 );
and ( n1535 , n784 , n1199 );
nor ( n1536 , n1534 , n1535 );
xnor ( n1537 , n1536 , n1296 );
buf ( n1538 , n493 );
buf ( n1539 , n1538 );
xor ( n1540 , n1539 , n1441 );
not ( n1541 , n1442 );
and ( n1542 , n1540 , n1541 );
and ( n1543 , n743 , n1542 );
and ( n1544 , n760 , n1442 );
nor ( n1545 , n1543 , n1544 );
and ( n1546 , n1441 , n1293 );
not ( n1547 , n1546 );
and ( n1548 , n1539 , n1547 );
xnor ( n1549 , n1545 , n1548 );
xor ( n1550 , n1537 , n1549 );
and ( n1551 , n1189 , n753 );
and ( n1552 , n1311 , n751 );
nor ( n1553 , n1551 , n1552 );
xnor ( n1554 , n1553 , n765 );
not ( n1555 , n1443 );
and ( n1556 , n1555 , n1548 );
xor ( n1557 , n1554 , n1556 );
xor ( n1558 , n1550 , n1557 );
xor ( n1559 , n1533 , n1558 );
and ( n1560 , n1434 , n1438 );
and ( n1561 , n1438 , n1443 );
and ( n1562 , n1434 , n1443 );
or ( n1563 , n1560 , n1561 , n1562 );
and ( n1564 , n1414 , n1418 );
and ( n1565 , n1418 , n1423 );
and ( n1566 , n1414 , n1423 );
or ( n1567 , n1564 , n1565 , n1566 );
xor ( n1568 , n1563 , n1567 );
and ( n1569 , n1411 , n777 );
not ( n1570 , n456 );
and ( n1571 , n1570 , n477 );
and ( n1572 , n461 , n456 );
or ( n1573 , n1571 , n1572 );
buf ( n1574 , n1573 );
buf ( n1575 , n1574 );
and ( n1576 , n1575 , n774 );
nor ( n1577 , n1569 , n1576 );
xnor ( n1578 , n1577 , n750 );
and ( n1579 , n996 , n935 );
and ( n1580 , n1087 , n855 );
nor ( n1581 , n1579 , n1580 );
xnor ( n1582 , n1581 , n925 );
xor ( n1583 , n1578 , n1582 );
and ( n1584 , n844 , n1110 );
and ( n1585 , n916 , n1007 );
nor ( n1586 , n1584 , n1585 );
xnor ( n1587 , n1586 , n1096 );
xor ( n1588 , n1583 , n1587 );
xor ( n1589 , n1568 , n1588 );
xor ( n1590 , n1559 , n1589 );
xor ( n1591 , n1529 , n1590 );
and ( n1592 , n1399 , n1403 );
and ( n1593 , n1403 , n1448 );
and ( n1594 , n1399 , n1448 );
or ( n1595 , n1592 , n1593 , n1594 );
xor ( n1596 , n1591 , n1595 );
and ( n1597 , n1449 , n1452 );
xor ( n1598 , n1596 , n1597 );
buf ( n1599 , n1598 );
not ( n1600 , n455 );
and ( n1601 , n1600 , n1525 );
and ( n1602 , n1599 , n455 );
or ( n1603 , n1601 , n1602 );
and ( n1604 , n1462 , n1487 );
and ( n1605 , n1487 , n1514 );
and ( n1606 , n1462 , n1514 );
or ( n1607 , n1604 , n1605 , n1606 );
and ( n1608 , n1492 , n1496 );
and ( n1609 , n1496 , n1513 );
and ( n1610 , n1492 , n1513 );
or ( n1611 , n1608 , n1609 , n1610 );
and ( n1612 , n1503 , n1507 );
and ( n1613 , n1507 , n1512 );
and ( n1614 , n1503 , n1512 );
or ( n1615 , n1612 , n1613 , n1614 );
and ( n1616 , n1466 , n1473 );
xor ( n1617 , n1615 , n1616 );
and ( n1618 , n1027 , n894 );
and ( n1619 , n1137 , n828 );
nor ( n1620 , n1618 , n1619 );
xnor ( n1621 , n1620 , n884 );
xor ( n1622 , n1617 , n1621 );
xor ( n1623 , n1611 , n1622 );
and ( n1624 , n1474 , n1478 );
and ( n1625 , n1478 , n1486 );
and ( n1626 , n1474 , n1486 );
or ( n1627 , n1624 , n1625 , n1626 );
and ( n1628 , n1500 , n708 );
buf ( n1629 , n508 );
buf ( n1630 , n1629 );
and ( n1631 , n1630 , n705 );
nor ( n1632 , n1628 , n1631 );
xnor ( n1633 , n1632 , n689 );
and ( n1634 , n711 , n1241 );
and ( n1635 , n817 , n1148 );
nor ( n1636 , n1634 , n1635 );
xnor ( n1637 , n1636 , n1247 );
xor ( n1638 , n1633 , n1637 );
and ( n1639 , n695 , n1482 );
and ( n1640 , n703 , n1381 );
nor ( n1641 , n1639 , n1640 );
xnor ( n1642 , n1641 , n1472 );
xor ( n1643 , n1638 , n1642 );
xor ( n1644 , n1627 , n1643 );
and ( n1645 , n1228 , n692 );
and ( n1646 , n1349 , n690 );
nor ( n1647 , n1645 , n1646 );
xnor ( n1648 , n1647 , n700 );
and ( n1649 , n875 , n1055 );
and ( n1650 , n959 , n970 );
nor ( n1651 , n1649 , n1650 );
xnor ( n1652 , n1651 , n1036 );
xor ( n1653 , n1648 , n1652 );
buf ( n1654 , n492 );
buf ( n1655 , n1654 );
xor ( n1656 , n1655 , n1469 );
and ( n1657 , n682 , n1656 );
xor ( n1658 , n1653 , n1657 );
xor ( n1659 , n1644 , n1658 );
xor ( n1660 , n1623 , n1659 );
xor ( n1661 , n1607 , n1660 );
and ( n1662 , n1515 , n1519 );
and ( n1663 , n1520 , n1523 );
or ( n1664 , n1662 , n1663 );
xor ( n1665 , n1661 , n1664 );
buf ( n1666 , n1665 );
and ( n1667 , n1578 , n1582 );
and ( n1668 , n1582 , n1587 );
and ( n1669 , n1578 , n1587 );
or ( n1670 , n1667 , n1668 , n1669 );
and ( n1671 , n1575 , n777 );
not ( n1672 , n456 );
and ( n1673 , n1672 , n476 );
and ( n1674 , n460 , n456 );
or ( n1675 , n1673 , n1674 );
buf ( n1676 , n1675 );
buf ( n1677 , n1676 );
and ( n1678 , n1677 , n774 );
nor ( n1679 , n1671 , n1678 );
xnor ( n1680 , n1679 , n750 );
and ( n1681 , n1087 , n935 );
and ( n1682 , n1189 , n855 );
nor ( n1683 , n1681 , n1682 );
xnor ( n1684 , n1683 , n925 );
xor ( n1685 , n1680 , n1684 );
and ( n1686 , n784 , n1322 );
and ( n1687 , n844 , n1199 );
nor ( n1688 , n1686 , n1687 );
xnor ( n1689 , n1688 , n1296 );
xor ( n1690 , n1685 , n1689 );
xor ( n1691 , n1670 , n1690 );
and ( n1692 , n1537 , n1549 );
and ( n1693 , n1549 , n1557 );
and ( n1694 , n1537 , n1557 );
or ( n1695 , n1692 , n1693 , n1694 );
xor ( n1696 , n1691 , n1695 );
and ( n1697 , n1563 , n1567 );
and ( n1698 , n1567 , n1588 );
and ( n1699 , n1563 , n1588 );
or ( n1700 , n1697 , n1698 , n1699 );
and ( n1701 , n760 , n1542 );
and ( n1702 , n772 , n1442 );
nor ( n1703 , n1701 , n1702 );
xnor ( n1704 , n1703 , n1548 );
and ( n1705 , n1311 , n753 );
and ( n1706 , n1411 , n751 );
nor ( n1707 , n1705 , n1706 );
xnor ( n1708 , n1707 , n765 );
and ( n1709 , n916 , n1110 );
and ( n1710 , n996 , n1007 );
nor ( n1711 , n1709 , n1710 );
xnor ( n1712 , n1711 , n1096 );
xor ( n1713 , n1708 , n1712 );
buf ( n1714 , n492 );
buf ( n1715 , n1714 );
xor ( n1716 , n1715 , n1539 );
and ( n1717 , n743 , n1716 );
xor ( n1718 , n1713 , n1717 );
xor ( n1719 , n1704 , n1718 );
and ( n1720 , n1554 , n1556 );
xor ( n1721 , n1719 , n1720 );
xor ( n1722 , n1700 , n1721 );
and ( n1723 , n1533 , n1558 );
and ( n1724 , n1558 , n1589 );
and ( n1725 , n1533 , n1589 );
or ( n1726 , n1723 , n1724 , n1725 );
xor ( n1727 , n1722 , n1726 );
xor ( n1728 , n1696 , n1727 );
and ( n1729 , n1529 , n1590 );
and ( n1730 , n1590 , n1595 );
and ( n1731 , n1529 , n1595 );
or ( n1732 , n1729 , n1730 , n1731 );
xor ( n1733 , n1728 , n1732 );
and ( n1734 , n1596 , n1597 );
xor ( n1735 , n1733 , n1734 );
buf ( n1736 , n1735 );
not ( n1737 , n455 );
and ( n1738 , n1737 , n1666 );
and ( n1739 , n1736 , n455 );
or ( n1740 , n1738 , n1739 );
and ( n1741 , n1627 , n1643 );
and ( n1742 , n1643 , n1658 );
and ( n1743 , n1627 , n1658 );
or ( n1744 , n1741 , n1742 , n1743 );
and ( n1745 , n1630 , n708 );
buf ( n1746 , n507 );
buf ( n1747 , n1746 );
and ( n1748 , n1747 , n705 );
nor ( n1749 , n1745 , n1748 );
xnor ( n1750 , n1749 , n689 );
not ( n1751 , n1657 );
buf ( n1752 , n491 );
buf ( n1753 , n1752 );
and ( n1754 , n1655 , n1469 );
not ( n1755 , n1754 );
and ( n1756 , n1753 , n1755 );
and ( n1757 , n1751 , n1756 );
xor ( n1758 , n1750 , n1757 );
and ( n1759 , n1633 , n1637 );
and ( n1760 , n1637 , n1642 );
and ( n1761 , n1633 , n1642 );
or ( n1762 , n1759 , n1760 , n1761 );
xor ( n1763 , n1758 , n1762 );
and ( n1764 , n1648 , n1652 );
and ( n1765 , n1652 , n1657 );
and ( n1766 , n1648 , n1657 );
or ( n1767 , n1764 , n1765 , n1766 );
xor ( n1768 , n1763 , n1767 );
xor ( n1769 , n1744 , n1768 );
and ( n1770 , n1615 , n1616 );
and ( n1771 , n1616 , n1621 );
and ( n1772 , n1615 , n1621 );
or ( n1773 , n1770 , n1771 , n1772 );
and ( n1774 , n1349 , n692 );
and ( n1775 , n1500 , n690 );
nor ( n1776 , n1774 , n1775 );
xnor ( n1777 , n1776 , n700 );
and ( n1778 , n959 , n1055 );
and ( n1779 , n1027 , n970 );
nor ( n1780 , n1778 , n1779 );
xnor ( n1781 , n1780 , n1036 );
xor ( n1782 , n1777 , n1781 );
and ( n1783 , n817 , n1241 );
and ( n1784 , n875 , n1148 );
nor ( n1785 , n1783 , n1784 );
xnor ( n1786 , n1785 , n1247 );
xor ( n1787 , n1782 , n1786 );
xor ( n1788 , n1773 , n1787 );
and ( n1789 , n1137 , n894 );
and ( n1790 , n1228 , n828 );
nor ( n1791 , n1789 , n1790 );
xnor ( n1792 , n1791 , n884 );
and ( n1793 , n703 , n1482 );
and ( n1794 , n711 , n1381 );
nor ( n1795 , n1793 , n1794 );
xnor ( n1796 , n1795 , n1472 );
xor ( n1797 , n1792 , n1796 );
xor ( n1798 , n1753 , n1655 );
not ( n1799 , n1656 );
and ( n1800 , n1798 , n1799 );
and ( n1801 , n682 , n1800 );
and ( n1802 , n695 , n1656 );
nor ( n1803 , n1801 , n1802 );
xnor ( n1804 , n1803 , n1756 );
xor ( n1805 , n1797 , n1804 );
xor ( n1806 , n1788 , n1805 );
xor ( n1807 , n1769 , n1806 );
and ( n1808 , n1611 , n1622 );
and ( n1809 , n1622 , n1659 );
and ( n1810 , n1611 , n1659 );
or ( n1811 , n1808 , n1809 , n1810 );
xor ( n1812 , n1807 , n1811 );
and ( n1813 , n1607 , n1660 );
and ( n1814 , n1661 , n1664 );
or ( n1815 , n1813 , n1814 );
xor ( n1816 , n1812 , n1815 );
buf ( n1817 , n1816 );
and ( n1818 , n1670 , n1690 );
and ( n1819 , n1690 , n1695 );
and ( n1820 , n1670 , n1695 );
or ( n1821 , n1818 , n1819 , n1820 );
and ( n1822 , n1704 , n1718 );
and ( n1823 , n1718 , n1720 );
and ( n1824 , n1704 , n1720 );
or ( n1825 , n1822 , n1823 , n1824 );
buf ( n1826 , n491 );
buf ( n1827 , n1826 );
xor ( n1828 , n1827 , n1715 );
not ( n1829 , n1716 );
and ( n1830 , n1828 , n1829 );
and ( n1831 , n743 , n1830 );
and ( n1832 , n760 , n1716 );
nor ( n1833 , n1831 , n1832 );
and ( n1834 , n1715 , n1539 );
not ( n1835 , n1834 );
and ( n1836 , n1827 , n1835 );
xnor ( n1837 , n1833 , n1836 );
not ( n1838 , n1717 );
and ( n1839 , n1838 , n1836 );
xor ( n1840 , n1837 , n1839 );
and ( n1841 , n1411 , n753 );
and ( n1842 , n1575 , n751 );
nor ( n1843 , n1841 , n1842 );
xnor ( n1844 , n1843 , n765 );
and ( n1845 , n996 , n1110 );
and ( n1846 , n1087 , n1007 );
nor ( n1847 , n1845 , n1846 );
xnor ( n1848 , n1847 , n1096 );
xor ( n1849 , n1844 , n1848 );
and ( n1850 , n844 , n1322 );
and ( n1851 , n916 , n1199 );
nor ( n1852 , n1850 , n1851 );
xnor ( n1853 , n1852 , n1296 );
xor ( n1854 , n1849 , n1853 );
xor ( n1855 , n1840 , n1854 );
xor ( n1856 , n1825 , n1855 );
and ( n1857 , n1708 , n1712 );
and ( n1858 , n1712 , n1717 );
and ( n1859 , n1708 , n1717 );
or ( n1860 , n1857 , n1858 , n1859 );
and ( n1861 , n1680 , n1684 );
and ( n1862 , n1684 , n1689 );
and ( n1863 , n1680 , n1689 );
or ( n1864 , n1861 , n1862 , n1863 );
xor ( n1865 , n1860 , n1864 );
and ( n1866 , n1677 , n777 );
not ( n1867 , n456 );
and ( n1868 , n1867 , n475 );
and ( n1869 , n459 , n456 );
or ( n1870 , n1868 , n1869 );
buf ( n1871 , n1870 );
buf ( n1872 , n1871 );
and ( n1873 , n1872 , n774 );
nor ( n1874 , n1866 , n1873 );
xnor ( n1875 , n1874 , n750 );
and ( n1876 , n1189 , n935 );
and ( n1877 , n1311 , n855 );
nor ( n1878 , n1876 , n1877 );
xnor ( n1879 , n1878 , n925 );
xor ( n1880 , n1875 , n1879 );
and ( n1881 , n772 , n1542 );
and ( n1882 , n784 , n1442 );
nor ( n1883 , n1881 , n1882 );
xnor ( n1884 , n1883 , n1548 );
xor ( n1885 , n1880 , n1884 );
xor ( n1886 , n1865 , n1885 );
xor ( n1887 , n1856 , n1886 );
xor ( n1888 , n1821 , n1887 );
and ( n1889 , n1700 , n1721 );
and ( n1890 , n1721 , n1726 );
and ( n1891 , n1700 , n1726 );
or ( n1892 , n1889 , n1890 , n1891 );
xor ( n1893 , n1888 , n1892 );
and ( n1894 , n1696 , n1727 );
and ( n1895 , n1727 , n1732 );
and ( n1896 , n1696 , n1732 );
or ( n1897 , n1894 , n1895 , n1896 );
xor ( n1898 , n1893 , n1897 );
and ( n1899 , n1733 , n1734 );
xor ( n1900 , n1898 , n1899 );
buf ( n1901 , n1900 );
not ( n1902 , n455 );
and ( n1903 , n1902 , n1817 );
and ( n1904 , n1901 , n455 );
or ( n1905 , n1903 , n1904 );
and ( n1906 , n1773 , n1787 );
and ( n1907 , n1787 , n1805 );
and ( n1908 , n1773 , n1805 );
or ( n1909 , n1906 , n1907 , n1908 );
and ( n1910 , n1777 , n1781 );
and ( n1911 , n1781 , n1786 );
and ( n1912 , n1777 , n1786 );
or ( n1913 , n1910 , n1911 , n1912 );
and ( n1914 , n1792 , n1796 );
and ( n1915 , n1796 , n1804 );
and ( n1916 , n1792 , n1804 );
or ( n1917 , n1914 , n1915 , n1916 );
xor ( n1918 , n1913 , n1917 );
and ( n1919 , n1747 , n708 );
buf ( n1920 , n506 );
buf ( n1921 , n1920 );
and ( n1922 , n1921 , n705 );
nor ( n1923 , n1919 , n1922 );
xnor ( n1924 , n1923 , n689 );
and ( n1925 , n1500 , n692 );
and ( n1926 , n1630 , n690 );
nor ( n1927 , n1925 , n1926 );
xnor ( n1928 , n1927 , n700 );
xor ( n1929 , n1924 , n1928 );
buf ( n1930 , n490 );
buf ( n1931 , n1930 );
xor ( n1932 , n1931 , n1753 );
and ( n1933 , n682 , n1932 );
xor ( n1934 , n1929 , n1933 );
xor ( n1935 , n1918 , n1934 );
xor ( n1936 , n1909 , n1935 );
and ( n1937 , n1758 , n1762 );
and ( n1938 , n1762 , n1767 );
and ( n1939 , n1758 , n1767 );
or ( n1940 , n1937 , n1938 , n1939 );
and ( n1941 , n1228 , n894 );
and ( n1942 , n1349 , n828 );
nor ( n1943 , n1941 , n1942 );
xnor ( n1944 , n1943 , n884 );
and ( n1945 , n1027 , n1055 );
and ( n1946 , n1137 , n970 );
nor ( n1947 , n1945 , n1946 );
xnor ( n1948 , n1947 , n1036 );
xor ( n1949 , n1944 , n1948 );
and ( n1950 , n875 , n1241 );
and ( n1951 , n959 , n1148 );
nor ( n1952 , n1950 , n1951 );
xnor ( n1953 , n1952 , n1247 );
xor ( n1954 , n1949 , n1953 );
xor ( n1955 , n1940 , n1954 );
and ( n1956 , n1750 , n1757 );
and ( n1957 , n711 , n1482 );
and ( n1958 , n817 , n1381 );
nor ( n1959 , n1957 , n1958 );
xnor ( n1960 , n1959 , n1472 );
xor ( n1961 , n1956 , n1960 );
and ( n1962 , n695 , n1800 );
and ( n1963 , n703 , n1656 );
nor ( n1964 , n1962 , n1963 );
xnor ( n1965 , n1964 , n1756 );
xor ( n1966 , n1961 , n1965 );
xor ( n1967 , n1955 , n1966 );
xor ( n1968 , n1936 , n1967 );
and ( n1969 , n1744 , n1768 );
and ( n1970 , n1768 , n1806 );
and ( n1971 , n1744 , n1806 );
or ( n1972 , n1969 , n1970 , n1971 );
xor ( n1973 , n1968 , n1972 );
and ( n1974 , n1807 , n1811 );
and ( n1975 , n1812 , n1815 );
or ( n1976 , n1974 , n1975 );
xor ( n1977 , n1973 , n1976 );
buf ( n1978 , n1977 );
and ( n1979 , n1875 , n1879 );
and ( n1980 , n1879 , n1884 );
and ( n1981 , n1875 , n1884 );
or ( n1982 , n1979 , n1980 , n1981 );
and ( n1983 , n1844 , n1848 );
and ( n1984 , n1848 , n1853 );
and ( n1985 , n1844 , n1853 );
or ( n1986 , n1983 , n1984 , n1985 );
and ( n1987 , n1872 , n777 );
not ( n1988 , n456 );
and ( n1989 , n1988 , n474 );
and ( n1990 , n458 , n456 );
or ( n1991 , n1989 , n1990 );
buf ( n1992 , n1991 );
buf ( n1993 , n1992 );
and ( n1994 , n1993 , n774 );
nor ( n1995 , n1987 , n1994 );
xnor ( n1996 , n1995 , n750 );
and ( n1997 , n1575 , n753 );
and ( n1998 , n1677 , n751 );
nor ( n1999 , n1997 , n1998 );
xnor ( n2000 , n1999 , n765 );
xor ( n2001 , n1996 , n2000 );
buf ( n2002 , n490 );
buf ( n2003 , n2002 );
xor ( n2004 , n2003 , n1827 );
and ( n2005 , n743 , n2004 );
xor ( n2006 , n2001 , n2005 );
xnor ( n2007 , n1986 , n2006 );
xor ( n2008 , n1982 , n2007 );
and ( n2009 , n1837 , n1839 );
and ( n2010 , n1839 , n1854 );
and ( n2011 , n1837 , n1854 );
or ( n2012 , n2009 , n2010 , n2011 );
xor ( n2013 , n2008 , n2012 );
and ( n2014 , n1860 , n1864 );
and ( n2015 , n1864 , n1885 );
and ( n2016 , n1860 , n1885 );
or ( n2017 , n2014 , n2015 , n2016 );
and ( n2018 , n784 , n1542 );
and ( n2019 , n844 , n1442 );
nor ( n2020 , n2018 , n2019 );
xnor ( n2021 , n2020 , n1548 );
and ( n2022 , n760 , n1830 );
and ( n2023 , n772 , n1716 );
nor ( n2024 , n2022 , n2023 );
xnor ( n2025 , n2024 , n1836 );
xor ( n2026 , n2021 , n2025 );
and ( n2027 , n1311 , n935 );
and ( n2028 , n1411 , n855 );
nor ( n2029 , n2027 , n2028 );
xnor ( n2030 , n2029 , n925 );
and ( n2031 , n1087 , n1110 );
and ( n2032 , n1189 , n1007 );
nor ( n2033 , n2031 , n2032 );
xnor ( n2034 , n2033 , n1096 );
xor ( n2035 , n2030 , n2034 );
and ( n2036 , n916 , n1322 );
and ( n2037 , n996 , n1199 );
nor ( n2038 , n2036 , n2037 );
xnor ( n2039 , n2038 , n1296 );
xor ( n2040 , n2035 , n2039 );
xor ( n2041 , n2026 , n2040 );
xor ( n2042 , n2017 , n2041 );
and ( n2043 , n1825 , n1855 );
and ( n2044 , n1855 , n1886 );
and ( n2045 , n1825 , n1886 );
or ( n2046 , n2043 , n2044 , n2045 );
xor ( n2047 , n2042 , n2046 );
xor ( n2048 , n2013 , n2047 );
and ( n2049 , n1821 , n1887 );
and ( n2050 , n1887 , n1892 );
and ( n2051 , n1821 , n1892 );
or ( n2052 , n2049 , n2050 , n2051 );
xor ( n2053 , n2048 , n2052 );
not ( n2054 , n2053 );
and ( n2055 , n1893 , n1897 );
and ( n2056 , n1898 , n1899 );
or ( n2057 , n2055 , n2056 );
xor ( n2058 , n2054 , n2057 );
buf ( n2059 , n2058 );
not ( n2060 , n455 );
and ( n2061 , n2060 , n1978 );
and ( n2062 , n2059 , n455 );
or ( n2063 , n2061 , n2062 );
and ( n2064 , n1940 , n1954 );
and ( n2065 , n1954 , n1966 );
and ( n2066 , n1940 , n1966 );
or ( n2067 , n2064 , n2065 , n2066 );
and ( n2068 , n1944 , n1948 );
and ( n2069 , n1948 , n1953 );
and ( n2070 , n1944 , n1953 );
or ( n2071 , n2068 , n2069 , n2070 );
and ( n2072 , n1349 , n894 );
and ( n2073 , n1500 , n828 );
nor ( n2074 , n2072 , n2073 );
xnor ( n2075 , n2074 , n884 );
and ( n2076 , n959 , n1241 );
and ( n2077 , n1027 , n1148 );
nor ( n2078 , n2076 , n2077 );
xnor ( n2079 , n2078 , n1247 );
xor ( n2080 , n2075 , n2079 );
and ( n2081 , n817 , n1482 );
and ( n2082 , n875 , n1381 );
nor ( n2083 , n2081 , n2082 );
xnor ( n2084 , n2083 , n1472 );
xor ( n2085 , n2080 , n2084 );
xor ( n2086 , n2071 , n2085 );
and ( n2087 , n1630 , n692 );
and ( n2088 , n1747 , n690 );
nor ( n2089 , n2087 , n2088 );
xnor ( n2090 , n2089 , n700 );
and ( n2091 , n1137 , n1055 );
and ( n2092 , n1228 , n970 );
nor ( n2093 , n2091 , n2092 );
xnor ( n2094 , n2093 , n1036 );
xor ( n2095 , n2090 , n2094 );
buf ( n2096 , n489 );
buf ( n2097 , n2096 );
xor ( n2098 , n2097 , n1931 );
not ( n2099 , n1932 );
and ( n2100 , n2098 , n2099 );
and ( n2101 , n682 , n2100 );
and ( n2102 , n695 , n1932 );
nor ( n2103 , n2101 , n2102 );
and ( n2104 , n1931 , n1753 );
not ( n2105 , n2104 );
and ( n2106 , n2097 , n2105 );
xnor ( n2107 , n2103 , n2106 );
xor ( n2108 , n2095 , n2107 );
xor ( n2109 , n2086 , n2108 );
xor ( n2110 , n2067 , n2109 );
and ( n2111 , n1956 , n1960 );
and ( n2112 , n1960 , n1965 );
and ( n2113 , n1956 , n1965 );
or ( n2114 , n2111 , n2112 , n2113 );
and ( n2115 , n1913 , n1917 );
and ( n2116 , n1917 , n1934 );
and ( n2117 , n1913 , n1934 );
or ( n2118 , n2115 , n2116 , n2117 );
xor ( n2119 , n2114 , n2118 );
and ( n2120 , n1921 , n708 );
buf ( n2121 , n505 );
buf ( n2122 , n2121 );
and ( n2123 , n2122 , n705 );
nor ( n2124 , n2120 , n2123 );
xnor ( n2125 , n2124 , n689 );
not ( n2126 , n1933 );
and ( n2127 , n2126 , n2106 );
xor ( n2128 , n2125 , n2127 );
and ( n2129 , n1924 , n1928 );
and ( n2130 , n1928 , n1933 );
and ( n2131 , n1924 , n1933 );
or ( n2132 , n2129 , n2130 , n2131 );
xor ( n2133 , n2128 , n2132 );
and ( n2134 , n703 , n1800 );
and ( n2135 , n711 , n1656 );
nor ( n2136 , n2134 , n2135 );
xnor ( n2137 , n2136 , n1756 );
xor ( n2138 , n2133 , n2137 );
xor ( n2139 , n2119 , n2138 );
xor ( n2140 , n2110 , n2139 );
and ( n2141 , n1909 , n1935 );
and ( n2142 , n1935 , n1967 );
and ( n2143 , n1909 , n1967 );
or ( n2144 , n2141 , n2142 , n2143 );
xor ( n2145 , n2140 , n2144 );
and ( n2146 , n1968 , n1972 );
and ( n2147 , n1973 , n1976 );
or ( n2148 , n2146 , n2147 );
xor ( n2149 , n2145 , n2148 );
buf ( n2150 , n2149 );
and ( n2151 , n2017 , n2041 );
and ( n2152 , n2041 , n2046 );
and ( n2153 , n2017 , n2046 );
or ( n2154 , n2151 , n2152 , n2153 );
and ( n2155 , n2030 , n2034 );
and ( n2156 , n2034 , n2039 );
and ( n2157 , n2030 , n2039 );
or ( n2158 , n2155 , n2156 , n2157 );
and ( n2159 , n1677 , n753 );
and ( n2160 , n1872 , n751 );
nor ( n2161 , n2159 , n2160 );
xnor ( n2162 , n2161 , n765 );
and ( n2163 , n1411 , n935 );
and ( n2164 , n1575 , n855 );
nor ( n2165 , n2163 , n2164 );
xnor ( n2166 , n2165 , n925 );
xor ( n2167 , n2162 , n2166 );
and ( n2168 , n1189 , n1110 );
and ( n2169 , n1311 , n1007 );
nor ( n2170 , n2168 , n2169 );
xnor ( n2171 , n2170 , n1096 );
xor ( n2172 , n2167 , n2171 );
xor ( n2173 , n2158 , n2172 );
and ( n2174 , n996 , n1322 );
and ( n2175 , n1087 , n1199 );
nor ( n2176 , n2174 , n2175 );
xnor ( n2177 , n2176 , n1296 );
and ( n2178 , n844 , n1542 );
and ( n2179 , n916 , n1442 );
nor ( n2180 , n2178 , n2179 );
xnor ( n2181 , n2180 , n1548 );
xor ( n2182 , n2177 , n2181 );
buf ( n2183 , n489 );
buf ( n2184 , n2183 );
xor ( n2185 , n2184 , n2003 );
not ( n2186 , n2004 );
and ( n2187 , n2185 , n2186 );
and ( n2188 , n743 , n2187 );
and ( n2189 , n760 , n2004 );
nor ( n2190 , n2188 , n2189 );
and ( n2191 , n2003 , n1827 );
not ( n2192 , n2191 );
and ( n2193 , n2184 , n2192 );
xnor ( n2194 , n2190 , n2193 );
xor ( n2195 , n2182 , n2194 );
xor ( n2196 , n2173 , n2195 );
and ( n2197 , n1982 , n2007 );
and ( n2198 , n2007 , n2012 );
and ( n2199 , n1982 , n2012 );
or ( n2200 , n2197 , n2198 , n2199 );
xor ( n2201 , n2196 , n2200 );
and ( n2202 , n1993 , n777 );
not ( n2203 , n456 );
and ( n2204 , n2203 , n473 );
and ( n2205 , n457 , n456 );
or ( n2206 , n2204 , n2205 );
buf ( n2207 , n2206 );
buf ( n2208 , n2207 );
and ( n2209 , n2208 , n774 );
nor ( n2210 , n2202 , n2209 );
xnor ( n2211 , n2210 , n750 );
not ( n2212 , n2005 );
and ( n2213 , n2212 , n2193 );
xor ( n2214 , n2211 , n2213 );
and ( n2215 , n1996 , n2000 );
and ( n2216 , n2000 , n2005 );
and ( n2217 , n1996 , n2005 );
or ( n2218 , n2215 , n2216 , n2217 );
xor ( n2219 , n2214 , n2218 );
and ( n2220 , n772 , n1830 );
and ( n2221 , n784 , n1716 );
nor ( n2222 , n2220 , n2221 );
xnor ( n2223 , n2222 , n1836 );
xor ( n2224 , n2219 , n2223 );
or ( n2225 , n1986 , n2006 );
xor ( n2226 , n2224 , n2225 );
and ( n2227 , n2021 , n2025 );
and ( n2228 , n2025 , n2040 );
and ( n2229 , n2021 , n2040 );
or ( n2230 , n2227 , n2228 , n2229 );
xor ( n2231 , n2226 , n2230 );
xor ( n2232 , n2201 , n2231 );
xor ( n2233 , n2154 , n2232 );
and ( n2234 , n2013 , n2047 );
and ( n2235 , n2047 , n2052 );
and ( n2236 , n2013 , n2052 );
or ( n2237 , n2234 , n2235 , n2236 );
xor ( n2238 , n2233 , n2237 );
not ( n2239 , n2238 );
and ( n2240 , n2054 , n2057 );
or ( n2241 , n2053 , n2240 );
xor ( n2242 , n2239 , n2241 );
buf ( n2243 , n2242 );
not ( n2244 , n455 );
and ( n2245 , n2244 , n2150 );
and ( n2246 , n2243 , n455 );
or ( n2247 , n2245 , n2246 );
and ( n2248 , n2114 , n2118 );
and ( n2249 , n2118 , n2138 );
and ( n2250 , n2114 , n2138 );
or ( n2251 , n2248 , n2249 , n2250 );
and ( n2252 , n2122 , n708 );
not ( n2253 , n2252 );
xnor ( n2254 , n2253 , n689 );
and ( n2255 , n1747 , n692 );
and ( n2256 , n1921 , n690 );
nor ( n2257 , n2255 , n2256 );
xnor ( n2258 , n2257 , n700 );
xor ( n2259 , n2254 , n2258 );
and ( n2260 , n682 , n2097 );
xor ( n2261 , n2259 , n2260 );
and ( n2262 , n1228 , n1055 );
and ( n2263 , n1349 , n970 );
nor ( n2264 , n2262 , n2263 );
xnor ( n2265 , n2264 , n1036 );
and ( n2266 , n1027 , n1241 );
and ( n2267 , n1137 , n1148 );
nor ( n2268 , n2266 , n2267 );
xnor ( n2269 , n2268 , n1247 );
xor ( n2270 , n2265 , n2269 );
and ( n2271 , n695 , n2100 );
and ( n2272 , n703 , n1932 );
nor ( n2273 , n2271 , n2272 );
xnor ( n2274 , n2273 , n2106 );
xor ( n2275 , n2270 , n2274 );
xor ( n2276 , n2261 , n2275 );
and ( n2277 , n1500 , n894 );
and ( n2278 , n1630 , n828 );
nor ( n2279 , n2277 , n2278 );
xnor ( n2280 , n2279 , n884 );
and ( n2281 , n875 , n1482 );
and ( n2282 , n959 , n1381 );
nor ( n2283 , n2281 , n2282 );
xnor ( n2284 , n2283 , n1472 );
xor ( n2285 , n2280 , n2284 );
and ( n2286 , n711 , n1800 );
and ( n2287 , n817 , n1656 );
nor ( n2288 , n2286 , n2287 );
xnor ( n2289 , n2288 , n1756 );
xor ( n2290 , n2285 , n2289 );
xor ( n2291 , n2276 , n2290 );
xor ( n2292 , n2251 , n2291 );
and ( n2293 , n2128 , n2132 );
and ( n2294 , n2132 , n2137 );
and ( n2295 , n2128 , n2137 );
or ( n2296 , n2293 , n2294 , n2295 );
and ( n2297 , n2071 , n2085 );
and ( n2298 , n2085 , n2108 );
and ( n2299 , n2071 , n2108 );
or ( n2300 , n2297 , n2298 , n2299 );
xor ( n2301 , n2296 , n2300 );
and ( n2302 , n2075 , n2079 );
and ( n2303 , n2079 , n2084 );
and ( n2304 , n2075 , n2084 );
or ( n2305 , n2302 , n2303 , n2304 );
and ( n2306 , n2090 , n2094 );
and ( n2307 , n2094 , n2107 );
and ( n2308 , n2090 , n2107 );
or ( n2309 , n2306 , n2307 , n2308 );
xor ( n2310 , n2305 , n2309 );
and ( n2311 , n2125 , n2127 );
xor ( n2312 , n2310 , n2311 );
xor ( n2313 , n2301 , n2312 );
xor ( n2314 , n2292 , n2313 );
and ( n2315 , n2067 , n2109 );
and ( n2316 , n2109 , n2139 );
and ( n2317 , n2067 , n2139 );
or ( n2318 , n2315 , n2316 , n2317 );
xor ( n2319 , n2314 , n2318 );
and ( n2320 , n2140 , n2144 );
and ( n2321 , n2145 , n2148 );
or ( n2322 , n2320 , n2321 );
xor ( n2323 , n2319 , n2322 );
buf ( n2324 , n2323 );
and ( n2325 , n1872 , n753 );
and ( n2326 , n1993 , n751 );
nor ( n2327 , n2325 , n2326 );
xnor ( n2328 , n2327 , n765 );
and ( n2329 , n1311 , n1110 );
and ( n2330 , n1411 , n1007 );
nor ( n2331 , n2329 , n2330 );
xnor ( n2332 , n2331 , n1096 );
xor ( n2333 , n2328 , n2332 );
and ( n2334 , n1087 , n1322 );
and ( n2335 , n1189 , n1199 );
nor ( n2336 , n2334 , n2335 );
xnor ( n2337 , n2336 , n1296 );
xor ( n2338 , n2333 , n2337 );
and ( n2339 , n2214 , n2218 );
and ( n2340 , n2218 , n2223 );
and ( n2341 , n2214 , n2223 );
or ( n2342 , n2339 , n2340 , n2341 );
xor ( n2343 , n2338 , n2342 );
and ( n2344 , n2158 , n2172 );
and ( n2345 , n2172 , n2195 );
and ( n2346 , n2158 , n2195 );
or ( n2347 , n2344 , n2345 , n2346 );
xor ( n2348 , n2343 , n2347 );
and ( n2349 , n2196 , n2200 );
and ( n2350 , n2200 , n2231 );
and ( n2351 , n2196 , n2231 );
or ( n2352 , n2349 , n2350 , n2351 );
xor ( n2353 , n2348 , n2352 );
and ( n2354 , n760 , n2187 );
and ( n2355 , n772 , n2004 );
nor ( n2356 , n2354 , n2355 );
xnor ( n2357 , n2356 , n2193 );
and ( n2358 , n1575 , n935 );
and ( n2359 , n1677 , n855 );
nor ( n2360 , n2358 , n2359 );
xnor ( n2361 , n2360 , n925 );
and ( n2362 , n916 , n1542 );
and ( n2363 , n996 , n1442 );
nor ( n2364 , n2362 , n2363 );
xnor ( n2365 , n2364 , n1548 );
xor ( n2366 , n2361 , n2365 );
and ( n2367 , n784 , n1830 );
and ( n2368 , n844 , n1716 );
nor ( n2369 , n2367 , n2368 );
xnor ( n2370 , n2369 , n1836 );
xor ( n2371 , n2366 , n2370 );
xor ( n2372 , n2357 , n2371 );
and ( n2373 , n2208 , n777 );
not ( n2374 , n2373 );
xnor ( n2375 , n2374 , n750 );
and ( n2376 , n743 , n2184 );
xor ( n2377 , n2375 , n2376 );
xor ( n2378 , n2372 , n2377 );
and ( n2379 , n2211 , n2213 );
and ( n2380 , n2162 , n2166 );
and ( n2381 , n2166 , n2171 );
and ( n2382 , n2162 , n2171 );
or ( n2383 , n2380 , n2381 , n2382 );
xor ( n2384 , n2379 , n2383 );
and ( n2385 , n2177 , n2181 );
and ( n2386 , n2181 , n2194 );
and ( n2387 , n2177 , n2194 );
or ( n2388 , n2385 , n2386 , n2387 );
xor ( n2389 , n2384 , n2388 );
xor ( n2390 , n2378 , n2389 );
and ( n2391 , n2224 , n2225 );
and ( n2392 , n2225 , n2230 );
and ( n2393 , n2224 , n2230 );
or ( n2394 , n2391 , n2392 , n2393 );
xor ( n2395 , n2390 , n2394 );
xor ( n2396 , n2353 , n2395 );
and ( n2397 , n2154 , n2232 );
and ( n2398 , n2232 , n2237 );
and ( n2399 , n2154 , n2237 );
or ( n2400 , n2397 , n2398 , n2399 );
xnor ( n2401 , n2396 , n2400 );
and ( n2402 , n2239 , n2241 );
or ( n2403 , n2238 , n2402 );
xor ( n2404 , n2401 , n2403 );
buf ( n2405 , n2404 );
not ( n2406 , n455 );
and ( n2407 , n2406 , n2324 );
and ( n2408 , n2405 , n455 );
or ( n2409 , n2407 , n2408 );
and ( n2410 , n2296 , n2300 );
and ( n2411 , n2300 , n2312 );
and ( n2412 , n2296 , n2312 );
or ( n2413 , n2410 , n2411 , n2412 );
and ( n2414 , n2305 , n2309 );
and ( n2415 , n2309 , n2311 );
and ( n2416 , n2305 , n2311 );
or ( n2417 , n2414 , n2415 , n2416 );
not ( n2418 , n689 );
and ( n2419 , n703 , n2100 );
and ( n2420 , n711 , n1932 );
nor ( n2421 , n2419 , n2420 );
xnor ( n2422 , n2421 , n2106 );
xor ( n2423 , n2418 , n2422 );
and ( n2424 , n695 , n2097 );
xor ( n2425 , n2423 , n2424 );
xor ( n2426 , n2417 , n2425 );
and ( n2427 , n1921 , n692 );
and ( n2428 , n2122 , n690 );
nor ( n2429 , n2427 , n2428 );
xnor ( n2430 , n2429 , n700 );
and ( n2431 , n1630 , n894 );
and ( n2432 , n1747 , n828 );
nor ( n2433 , n2431 , n2432 );
xnor ( n2434 , n2433 , n884 );
xor ( n2435 , n2430 , n2434 );
and ( n2436 , n1137 , n1241 );
and ( n2437 , n1228 , n1148 );
nor ( n2438 , n2436 , n2437 );
xnor ( n2439 , n2438 , n1247 );
xor ( n2440 , n2435 , n2439 );
xor ( n2441 , n2426 , n2440 );
xor ( n2442 , n2413 , n2441 );
and ( n2443 , n2261 , n2275 );
and ( n2444 , n2275 , n2290 );
and ( n2445 , n2261 , n2290 );
or ( n2446 , n2443 , n2444 , n2445 );
and ( n2447 , n2254 , n2258 );
and ( n2448 , n2258 , n2260 );
and ( n2449 , n2254 , n2260 );
or ( n2450 , n2447 , n2448 , n2449 );
and ( n2451 , n2265 , n2269 );
and ( n2452 , n2269 , n2274 );
and ( n2453 , n2265 , n2274 );
or ( n2454 , n2451 , n2452 , n2453 );
xor ( n2455 , n2450 , n2454 );
and ( n2456 , n2280 , n2284 );
and ( n2457 , n2284 , n2289 );
and ( n2458 , n2280 , n2289 );
or ( n2459 , n2456 , n2457 , n2458 );
xor ( n2460 , n2455 , n2459 );
xor ( n2461 , n2446 , n2460 );
and ( n2462 , n1349 , n1055 );
and ( n2463 , n1500 , n970 );
nor ( n2464 , n2462 , n2463 );
xnor ( n2465 , n2464 , n1036 );
not ( n2466 , n2465 );
and ( n2467 , n959 , n1482 );
and ( n2468 , n1027 , n1381 );
nor ( n2469 , n2467 , n2468 );
xnor ( n2470 , n2469 , n1472 );
xor ( n2471 , n2466 , n2470 );
and ( n2472 , n817 , n1800 );
and ( n2473 , n875 , n1656 );
nor ( n2474 , n2472 , n2473 );
xnor ( n2475 , n2474 , n1756 );
xor ( n2476 , n2471 , n2475 );
xor ( n2477 , n2461 , n2476 );
xor ( n2478 , n2442 , n2477 );
and ( n2479 , n2251 , n2291 );
and ( n2480 , n2291 , n2313 );
and ( n2481 , n2251 , n2313 );
or ( n2482 , n2479 , n2480 , n2481 );
xor ( n2483 , n2478 , n2482 );
and ( n2484 , n2314 , n2318 );
and ( n2485 , n2319 , n2322 );
or ( n2486 , n2484 , n2485 );
xor ( n2487 , n2483 , n2486 );
buf ( n2488 , n2487 );
and ( n2489 , n2378 , n2389 );
and ( n2490 , n2389 , n2394 );
and ( n2491 , n2378 , n2394 );
or ( n2492 , n2489 , n2490 , n2491 );
and ( n2493 , n2375 , n2376 );
and ( n2494 , n2328 , n2332 );
and ( n2495 , n2332 , n2337 );
and ( n2496 , n2328 , n2337 );
or ( n2497 , n2494 , n2495 , n2496 );
xor ( n2498 , n2493 , n2497 );
and ( n2499 , n1993 , n753 );
and ( n2500 , n2208 , n751 );
nor ( n2501 , n2499 , n2500 );
xnor ( n2502 , n2501 , n765 );
and ( n2503 , n1677 , n935 );
and ( n2504 , n1872 , n855 );
nor ( n2505 , n2503 , n2504 );
xnor ( n2506 , n2505 , n925 );
xor ( n2507 , n2502 , n2506 );
and ( n2508 , n1189 , n1322 );
and ( n2509 , n1311 , n1199 );
nor ( n2510 , n2508 , n2509 );
xnor ( n2511 , n2510 , n1296 );
xor ( n2512 , n2507 , n2511 );
xor ( n2513 , n2498 , n2512 );
and ( n2514 , n2338 , n2342 );
and ( n2515 , n2342 , n2347 );
and ( n2516 , n2338 , n2347 );
or ( n2517 , n2514 , n2515 , n2516 );
xor ( n2518 , n2513 , n2517 );
and ( n2519 , n2357 , n2371 );
and ( n2520 , n2371 , n2377 );
and ( n2521 , n2357 , n2377 );
or ( n2522 , n2519 , n2520 , n2521 );
and ( n2523 , n2379 , n2383 );
and ( n2524 , n2383 , n2388 );
and ( n2525 , n2379 , n2388 );
or ( n2526 , n2523 , n2524 , n2525 );
xor ( n2527 , n2522 , n2526 );
not ( n2528 , n750 );
and ( n2529 , n772 , n2187 );
and ( n2530 , n784 , n2004 );
nor ( n2531 , n2529 , n2530 );
xnor ( n2532 , n2531 , n2193 );
xor ( n2533 , n2528 , n2532 );
and ( n2534 , n760 , n2184 );
xor ( n2535 , n2533 , n2534 );
and ( n2536 , n1411 , n1110 );
and ( n2537 , n1575 , n1007 );
nor ( n2538 , n2536 , n2537 );
xnor ( n2539 , n2538 , n1096 );
not ( n2540 , n2539 );
and ( n2541 , n996 , n1542 );
and ( n2542 , n1087 , n1442 );
nor ( n2543 , n2541 , n2542 );
xnor ( n2544 , n2543 , n1548 );
xor ( n2545 , n2540 , n2544 );
and ( n2546 , n844 , n1830 );
and ( n2547 , n916 , n1716 );
nor ( n2548 , n2546 , n2547 );
xnor ( n2549 , n2548 , n1836 );
xor ( n2550 , n2545 , n2549 );
xor ( n2551 , n2535 , n2550 );
and ( n2552 , n2361 , n2365 );
and ( n2553 , n2365 , n2370 );
and ( n2554 , n2361 , n2370 );
or ( n2555 , n2552 , n2553 , n2554 );
xor ( n2556 , n2551 , n2555 );
xor ( n2557 , n2527 , n2556 );
xor ( n2558 , n2518 , n2557 );
xor ( n2559 , n2492 , n2558 );
and ( n2560 , n2348 , n2352 );
and ( n2561 , n2352 , n2395 );
and ( n2562 , n2348 , n2395 );
or ( n2563 , n2560 , n2561 , n2562 );
xor ( n2564 , n2559 , n2563 );
or ( n2565 , n2396 , n2400 );
xnor ( n2566 , n2564 , n2565 );
and ( n2567 , n2401 , n2403 );
xor ( n2568 , n2566 , n2567 );
buf ( n2569 , n2568 );
not ( n2570 , n455 );
and ( n2571 , n2570 , n2488 );
and ( n2572 , n2569 , n455 );
or ( n2573 , n2571 , n2572 );
and ( n2574 , n2413 , n2441 );
and ( n2575 , n2441 , n2477 );
and ( n2576 , n2413 , n2477 );
or ( n2577 , n2574 , n2575 , n2576 );
and ( n2578 , n2446 , n2460 );
and ( n2579 , n2460 , n2476 );
and ( n2580 , n2446 , n2476 );
or ( n2581 , n2578 , n2579 , n2580 );
and ( n2582 , n2450 , n2454 );
and ( n2583 , n2454 , n2459 );
and ( n2584 , n2450 , n2459 );
or ( n2585 , n2582 , n2583 , n2584 );
and ( n2586 , n1747 , n894 );
and ( n2587 , n1921 , n828 );
nor ( n2588 , n2586 , n2587 );
xnor ( n2589 , n2588 , n884 );
and ( n2590 , n1228 , n1241 );
and ( n2591 , n1349 , n1148 );
nor ( n2592 , n2590 , n2591 );
xnor ( n2593 , n2592 , n1247 );
xor ( n2594 , n2589 , n2593 );
and ( n2595 , n703 , n2097 );
xor ( n2596 , n2594 , n2595 );
xor ( n2597 , n2585 , n2596 );
buf ( n2598 , n2465 );
and ( n2599 , n2122 , n692 );
not ( n2600 , n2599 );
xnor ( n2601 , n2600 , n700 );
not ( n2602 , n2601 );
xor ( n2603 , n2598 , n2602 );
and ( n2604 , n711 , n2100 );
and ( n2605 , n817 , n1932 );
nor ( n2606 , n2604 , n2605 );
xnor ( n2607 , n2606 , n2106 );
xor ( n2608 , n2603 , n2607 );
xor ( n2609 , n2597 , n2608 );
xor ( n2610 , n2581 , n2609 );
and ( n2611 , n2466 , n2470 );
and ( n2612 , n2470 , n2475 );
and ( n2613 , n2466 , n2475 );
or ( n2614 , n2611 , n2612 , n2613 );
and ( n2615 , n2417 , n2425 );
and ( n2616 , n2425 , n2440 );
and ( n2617 , n2417 , n2440 );
or ( n2618 , n2615 , n2616 , n2617 );
xor ( n2619 , n2614 , n2618 );
and ( n2620 , n2418 , n2422 );
and ( n2621 , n2422 , n2424 );
and ( n2622 , n2418 , n2424 );
or ( n2623 , n2620 , n2621 , n2622 );
and ( n2624 , n2430 , n2434 );
and ( n2625 , n2434 , n2439 );
and ( n2626 , n2430 , n2439 );
or ( n2627 , n2624 , n2625 , n2626 );
xor ( n2628 , n2623 , n2627 );
and ( n2629 , n1500 , n1055 );
and ( n2630 , n1630 , n970 );
nor ( n2631 , n2629 , n2630 );
xnor ( n2632 , n2631 , n1036 );
and ( n2633 , n1027 , n1482 );
and ( n2634 , n1137 , n1381 );
nor ( n2635 , n2633 , n2634 );
xnor ( n2636 , n2635 , n1472 );
xor ( n2637 , n2632 , n2636 );
and ( n2638 , n875 , n1800 );
and ( n2639 , n959 , n1656 );
nor ( n2640 , n2638 , n2639 );
xnor ( n2641 , n2640 , n1756 );
xor ( n2642 , n2637 , n2641 );
xor ( n2643 , n2628 , n2642 );
xor ( n2644 , n2619 , n2643 );
xor ( n2645 , n2610 , n2644 );
xor ( n2646 , n2577 , n2645 );
and ( n2647 , n2478 , n2482 );
and ( n2648 , n2483 , n2486 );
or ( n2649 , n2647 , n2648 );
xor ( n2650 , n2646 , n2649 );
buf ( n2651 , n2650 );
and ( n2652 , n2513 , n2517 );
and ( n2653 , n2517 , n2557 );
and ( n2654 , n2513 , n2557 );
or ( n2655 , n2652 , n2653 , n2654 );
and ( n2656 , n2522 , n2526 );
and ( n2657 , n2526 , n2556 );
and ( n2658 , n2522 , n2556 );
or ( n2659 , n2656 , n2657 , n2658 );
and ( n2660 , n2502 , n2506 );
and ( n2661 , n2506 , n2511 );
and ( n2662 , n2502 , n2511 );
or ( n2663 , n2660 , n2661 , n2662 );
and ( n2664 , n2208 , n753 );
not ( n2665 , n2664 );
xnor ( n2666 , n2665 , n765 );
and ( n2667 , n1872 , n935 );
and ( n2668 , n1993 , n855 );
nor ( n2669 , n2667 , n2668 );
xnor ( n2670 , n2669 , n925 );
xor ( n2671 , n2666 , n2670 );
and ( n2672 , n1311 , n1322 );
and ( n2673 , n1411 , n1199 );
nor ( n2674 , n2672 , n2673 );
xnor ( n2675 , n2674 , n1296 );
xor ( n2676 , n2671 , n2675 );
xor ( n2677 , n2663 , n2676 );
and ( n2678 , n2535 , n2550 );
and ( n2679 , n2550 , n2555 );
and ( n2680 , n2535 , n2555 );
or ( n2681 , n2678 , n2679 , n2680 );
xor ( n2682 , n2677 , n2681 );
xor ( n2683 , n2659 , n2682 );
and ( n2684 , n2493 , n2497 );
and ( n2685 , n2497 , n2512 );
and ( n2686 , n2493 , n2512 );
or ( n2687 , n2684 , n2685 , n2686 );
and ( n2688 , n784 , n2187 );
and ( n2689 , n844 , n2004 );
nor ( n2690 , n2688 , n2689 );
xnor ( n2691 , n2690 , n2193 );
and ( n2692 , n772 , n2184 );
xor ( n2693 , n2691 , n2692 );
and ( n2694 , n1575 , n1110 );
and ( n2695 , n1677 , n1007 );
nor ( n2696 , n2694 , n2695 );
xnor ( n2697 , n2696 , n1096 );
and ( n2698 , n1087 , n1542 );
and ( n2699 , n1189 , n1442 );
nor ( n2700 , n2698 , n2699 );
xnor ( n2701 , n2700 , n1548 );
xor ( n2702 , n2697 , n2701 );
and ( n2703 , n916 , n1830 );
and ( n2704 , n996 , n1716 );
nor ( n2705 , n2703 , n2704 );
xnor ( n2706 , n2705 , n1836 );
xor ( n2707 , n2702 , n2706 );
xor ( n2708 , n2693 , n2707 );
xor ( n2709 , n2687 , n2708 );
and ( n2710 , n2528 , n2532 );
and ( n2711 , n2532 , n2534 );
and ( n2712 , n2528 , n2534 );
or ( n2713 , n2710 , n2711 , n2712 );
and ( n2714 , n2540 , n2544 );
and ( n2715 , n2544 , n2549 );
and ( n2716 , n2540 , n2549 );
or ( n2717 , n2714 , n2715 , n2716 );
xor ( n2718 , n2713 , n2717 );
buf ( n2719 , n2539 );
xor ( n2720 , n2718 , n2719 );
xor ( n2721 , n2709 , n2720 );
xor ( n2722 , n2683 , n2721 );
xor ( n2723 , n2655 , n2722 );
and ( n2724 , n2492 , n2558 );
and ( n2725 , n2558 , n2563 );
and ( n2726 , n2492 , n2563 );
or ( n2727 , n2724 , n2725 , n2726 );
xor ( n2728 , n2723 , n2727 );
or ( n2729 , n2564 , n2565 );
xor ( n2730 , n2728 , n2729 );
and ( n2731 , n2566 , n2567 );
xor ( n2732 , n2730 , n2731 );
buf ( n2733 , n2732 );
not ( n2734 , n455 );
and ( n2735 , n2734 , n2651 );
and ( n2736 , n2733 , n455 );
or ( n2737 , n2735 , n2736 );
and ( n2738 , n2614 , n2618 );
and ( n2739 , n2618 , n2643 );
and ( n2740 , n2614 , n2643 );
or ( n2741 , n2738 , n2739 , n2740 );
and ( n2742 , n2598 , n2602 );
and ( n2743 , n2602 , n2607 );
and ( n2744 , n2598 , n2607 );
or ( n2745 , n2742 , n2743 , n2744 );
and ( n2746 , n1630 , n1055 );
and ( n2747 , n1747 , n970 );
nor ( n2748 , n2746 , n2747 );
xnor ( n2749 , n2748 , n1036 );
and ( n2750 , n1137 , n1482 );
and ( n2751 , n1228 , n1381 );
nor ( n2752 , n2750 , n2751 );
xnor ( n2753 , n2752 , n1472 );
xor ( n2754 , n2749 , n2753 );
and ( n2755 , n711 , n2097 );
xor ( n2756 , n2754 , n2755 );
xor ( n2757 , n2745 , n2756 );
buf ( n2758 , n2601 );
and ( n2759 , n959 , n1800 );
and ( n2760 , n1027 , n1656 );
nor ( n2761 , n2759 , n2760 );
xnor ( n2762 , n2761 , n1756 );
xor ( n2763 , n2758 , n2762 );
and ( n2764 , n817 , n2100 );
and ( n2765 , n875 , n1932 );
nor ( n2766 , n2764 , n2765 );
xnor ( n2767 , n2766 , n2106 );
xor ( n2768 , n2763 , n2767 );
xor ( n2769 , n2757 , n2768 );
xor ( n2770 , n2741 , n2769 );
and ( n2771 , n2623 , n2627 );
and ( n2772 , n2627 , n2642 );
and ( n2773 , n2623 , n2642 );
or ( n2774 , n2771 , n2772 , n2773 );
and ( n2775 , n2585 , n2596 );
and ( n2776 , n2596 , n2608 );
and ( n2777 , n2585 , n2608 );
or ( n2778 , n2775 , n2776 , n2777 );
xor ( n2779 , n2774 , n2778 );
and ( n2780 , n2589 , n2593 );
and ( n2781 , n2593 , n2595 );
and ( n2782 , n2589 , n2595 );
or ( n2783 , n2780 , n2781 , n2782 );
and ( n2784 , n2632 , n2636 );
and ( n2785 , n2636 , n2641 );
and ( n2786 , n2632 , n2641 );
or ( n2787 , n2784 , n2785 , n2786 );
xor ( n2788 , n2783 , n2787 );
not ( n2789 , n700 );
and ( n2790 , n1921 , n894 );
and ( n2791 , n2122 , n828 );
nor ( n2792 , n2790 , n2791 );
xnor ( n2793 , n2792 , n884 );
xor ( n2794 , n2789 , n2793 );
and ( n2795 , n1349 , n1241 );
and ( n2796 , n1500 , n1148 );
nor ( n2797 , n2795 , n2796 );
xnor ( n2798 , n2797 , n1247 );
xor ( n2799 , n2794 , n2798 );
xor ( n2800 , n2788 , n2799 );
xor ( n2801 , n2779 , n2800 );
xor ( n2802 , n2770 , n2801 );
and ( n2803 , n2581 , n2609 );
and ( n2804 , n2609 , n2644 );
and ( n2805 , n2581 , n2644 );
or ( n2806 , n2803 , n2804 , n2805 );
xor ( n2807 , n2802 , n2806 );
and ( n2808 , n2577 , n2645 );
and ( n2809 , n2646 , n2649 );
or ( n2810 , n2808 , n2809 );
xor ( n2811 , n2807 , n2810 );
buf ( n2812 , n2811 );
and ( n2813 , n2713 , n2717 );
and ( n2814 , n2717 , n2719 );
and ( n2815 , n2713 , n2719 );
or ( n2816 , n2813 , n2814 , n2815 );
not ( n2817 , n765 );
and ( n2818 , n1411 , n1322 );
and ( n2819 , n1575 , n1199 );
nor ( n2820 , n2818 , n2819 );
xnor ( n2821 , n2820 , n1296 );
xor ( n2822 , n2817 , n2821 );
and ( n2823 , n2697 , n2701 );
and ( n2824 , n2701 , n2706 );
and ( n2825 , n2697 , n2706 );
or ( n2826 , n2823 , n2824 , n2825 );
xor ( n2827 , n2822 , n2826 );
and ( n2828 , n2666 , n2670 );
and ( n2829 , n2670 , n2675 );
and ( n2830 , n2666 , n2675 );
or ( n2831 , n2828 , n2829 , n2830 );
xor ( n2832 , n2827 , n2831 );
xor ( n2833 , n2816 , n2832 );
and ( n2834 , n2663 , n2676 );
and ( n2835 , n2676 , n2681 );
and ( n2836 , n2663 , n2681 );
or ( n2837 , n2834 , n2835 , n2836 );
xor ( n2838 , n2833 , n2837 );
and ( n2839 , n2687 , n2708 );
and ( n2840 , n2708 , n2720 );
and ( n2841 , n2687 , n2720 );
or ( n2842 , n2839 , n2840 , n2841 );
and ( n2843 , n1993 , n935 );
and ( n2844 , n2208 , n855 );
nor ( n2845 , n2843 , n2844 );
xnor ( n2846 , n2845 , n925 );
and ( n2847 , n1677 , n1110 );
and ( n2848 , n1872 , n1007 );
nor ( n2849 , n2847 , n2848 );
xnor ( n2850 , n2849 , n1096 );
xor ( n2851 , n2846 , n2850 );
and ( n2852 , n1189 , n1542 );
and ( n2853 , n1311 , n1442 );
nor ( n2854 , n2852 , n2853 );
xnor ( n2855 , n2854 , n1548 );
xor ( n2856 , n2851 , n2855 );
and ( n2857 , n996 , n1830 );
and ( n2858 , n1087 , n1716 );
nor ( n2859 , n2857 , n2858 );
xnor ( n2860 , n2859 , n1836 );
and ( n2861 , n844 , n2187 );
and ( n2862 , n916 , n2004 );
nor ( n2863 , n2861 , n2862 );
xnor ( n2864 , n2863 , n2193 );
xor ( n2865 , n2860 , n2864 );
and ( n2866 , n784 , n2184 );
xor ( n2867 , n2865 , n2866 );
xor ( n2868 , n2856 , n2867 );
and ( n2869 , n2691 , n2692 );
and ( n2870 , n2692 , n2707 );
and ( n2871 , n2691 , n2707 );
or ( n2872 , n2869 , n2870 , n2871 );
xor ( n2873 , n2868 , n2872 );
xor ( n2874 , n2842 , n2873 );
and ( n2875 , n2659 , n2682 );
and ( n2876 , n2682 , n2721 );
and ( n2877 , n2659 , n2721 );
or ( n2878 , n2875 , n2876 , n2877 );
xor ( n2879 , n2874 , n2878 );
xor ( n2880 , n2838 , n2879 );
and ( n2881 , n2655 , n2722 );
and ( n2882 , n2722 , n2727 );
and ( n2883 , n2655 , n2727 );
or ( n2884 , n2881 , n2882 , n2883 );
xor ( n2885 , n2880 , n2884 );
and ( n2886 , n2728 , n2729 );
and ( n2887 , n2730 , n2731 );
or ( n2888 , n2886 , n2887 );
xor ( n2889 , n2885 , n2888 );
buf ( n2890 , n2889 );
not ( n2891 , n455 );
and ( n2892 , n2891 , n2812 );
and ( n2893 , n2890 , n455 );
or ( n2894 , n2892 , n2893 );
and ( n2895 , n2741 , n2769 );
and ( n2896 , n2769 , n2801 );
and ( n2897 , n2741 , n2801 );
or ( n2898 , n2895 , n2896 , n2897 );
and ( n2899 , n2745 , n2756 );
and ( n2900 , n2756 , n2768 );
and ( n2901 , n2745 , n2768 );
or ( n2902 , n2899 , n2900 , n2901 );
and ( n2903 , n2774 , n2778 );
and ( n2904 , n2778 , n2800 );
and ( n2905 , n2774 , n2800 );
or ( n2906 , n2903 , n2904 , n2905 );
xor ( n2907 , n2902 , n2906 );
and ( n2908 , n2783 , n2787 );
and ( n2909 , n2787 , n2799 );
and ( n2910 , n2783 , n2799 );
or ( n2911 , n2908 , n2909 , n2910 );
and ( n2912 , n2749 , n2753 );
and ( n2913 , n2753 , n2755 );
and ( n2914 , n2749 , n2755 );
or ( n2915 , n2912 , n2913 , n2914 );
and ( n2916 , n2789 , n2793 );
and ( n2917 , n2793 , n2798 );
and ( n2918 , n2789 , n2798 );
or ( n2919 , n2916 , n2917 , n2918 );
xor ( n2920 , n2915 , n2919 );
and ( n2921 , n2122 , n894 );
not ( n2922 , n2921 );
xnor ( n2923 , n2922 , n884 );
not ( n2924 , n2923 );
xor ( n2925 , n2920 , n2924 );
xor ( n2926 , n2911 , n2925 );
and ( n2927 , n2758 , n2762 );
and ( n2928 , n2762 , n2767 );
and ( n2929 , n2758 , n2767 );
or ( n2930 , n2927 , n2928 , n2929 );
and ( n2931 , n1747 , n1055 );
and ( n2932 , n1921 , n970 );
nor ( n2933 , n2931 , n2932 );
xnor ( n2934 , n2933 , n1036 );
and ( n2935 , n1228 , n1482 );
and ( n2936 , n1349 , n1381 );
nor ( n2937 , n2935 , n2936 );
xnor ( n2938 , n2937 , n1472 );
xor ( n2939 , n2934 , n2938 );
and ( n2940 , n1027 , n1800 );
and ( n2941 , n1137 , n1656 );
nor ( n2942 , n2940 , n2941 );
xnor ( n2943 , n2942 , n1756 );
xor ( n2944 , n2939 , n2943 );
xor ( n2945 , n2930 , n2944 );
and ( n2946 , n1500 , n1241 );
and ( n2947 , n1630 , n1148 );
nor ( n2948 , n2946 , n2947 );
xnor ( n2949 , n2948 , n1247 );
and ( n2950 , n875 , n2100 );
and ( n2951 , n959 , n1932 );
nor ( n2952 , n2950 , n2951 );
xnor ( n2953 , n2952 , n2106 );
xor ( n2954 , n2949 , n2953 );
and ( n2955 , n817 , n2097 );
xor ( n2956 , n2954 , n2955 );
xor ( n2957 , n2945 , n2956 );
xor ( n2958 , n2926 , n2957 );
xor ( n2959 , n2907 , n2958 );
xor ( n2960 , n2898 , n2959 );
and ( n2961 , n2802 , n2806 );
and ( n2962 , n2807 , n2810 );
or ( n2963 , n2961 , n2962 );
xor ( n2964 , n2960 , n2963 );
buf ( n2965 , n2964 );
and ( n2966 , n2842 , n2873 );
and ( n2967 , n2873 , n2878 );
and ( n2968 , n2842 , n2878 );
or ( n2969 , n2966 , n2967 , n2968 );
and ( n2970 , n2856 , n2867 );
and ( n2971 , n2867 , n2872 );
and ( n2972 , n2856 , n2872 );
or ( n2973 , n2970 , n2971 , n2972 );
and ( n2974 , n2822 , n2826 );
and ( n2975 , n2826 , n2831 );
and ( n2976 , n2822 , n2831 );
or ( n2977 , n2974 , n2975 , n2976 );
and ( n2978 , n1087 , n1830 );
and ( n2979 , n1189 , n1716 );
nor ( n2980 , n2978 , n2979 );
xnor ( n2981 , n2980 , n1836 );
and ( n2982 , n1575 , n1322 );
and ( n2983 , n1677 , n1199 );
nor ( n2984 , n2982 , n2983 );
xnor ( n2985 , n2984 , n1296 );
and ( n2986 , n916 , n2187 );
and ( n2987 , n996 , n2004 );
nor ( n2988 , n2986 , n2987 );
xnor ( n2989 , n2988 , n2193 );
xor ( n2990 , n2985 , n2989 );
and ( n2991 , n844 , n2184 );
xor ( n2992 , n2990 , n2991 );
xor ( n2993 , n2981 , n2992 );
and ( n2994 , n2817 , n2821 );
xor ( n2995 , n2993 , n2994 );
xor ( n2996 , n2977 , n2995 );
and ( n2997 , n2846 , n2850 );
and ( n2998 , n2850 , n2855 );
and ( n2999 , n2846 , n2855 );
or ( n3000 , n2997 , n2998 , n2999 );
and ( n3001 , n2860 , n2864 );
and ( n3002 , n2864 , n2866 );
and ( n3003 , n2860 , n2866 );
or ( n3004 , n3001 , n3002 , n3003 );
xor ( n3005 , n3000 , n3004 );
and ( n3006 , n2208 , n935 );
not ( n3007 , n3006 );
xnor ( n3008 , n3007 , n925 );
and ( n3009 , n1872 , n1110 );
and ( n3010 , n1993 , n1007 );
nor ( n3011 , n3009 , n3010 );
xnor ( n3012 , n3011 , n1096 );
xor ( n3013 , n3008 , n3012 );
and ( n3014 , n1311 , n1542 );
and ( n3015 , n1411 , n1442 );
nor ( n3016 , n3014 , n3015 );
xnor ( n3017 , n3016 , n1548 );
xor ( n3018 , n3013 , n3017 );
xor ( n3019 , n3005 , n3018 );
xor ( n3020 , n2996 , n3019 );
xor ( n3021 , n2973 , n3020 );
and ( n3022 , n2816 , n2832 );
and ( n3023 , n2832 , n2837 );
and ( n3024 , n2816 , n2837 );
or ( n3025 , n3022 , n3023 , n3024 );
xor ( n3026 , n3021 , n3025 );
xor ( n3027 , n2969 , n3026 );
and ( n3028 , n2838 , n2879 );
and ( n3029 , n2879 , n2884 );
and ( n3030 , n2838 , n2884 );
or ( n3031 , n3028 , n3029 , n3030 );
xor ( n3032 , n3027 , n3031 );
not ( n3033 , n3032 );
and ( n3034 , n2885 , n2888 );
xor ( n3035 , n3033 , n3034 );
buf ( n3036 , n3035 );
not ( n3037 , n455 );
and ( n3038 , n3037 , n2965 );
and ( n3039 , n3036 , n455 );
or ( n3040 , n3038 , n3039 );
and ( n3041 , n2911 , n2925 );
and ( n3042 , n2925 , n2957 );
and ( n3043 , n2911 , n2957 );
or ( n3044 , n3041 , n3042 , n3043 );
and ( n3045 , n2949 , n2953 );
and ( n3046 , n2953 , n2955 );
and ( n3047 , n2949 , n2955 );
or ( n3048 , n3045 , n3046 , n3047 );
not ( n3049 , n884 );
and ( n3050 , n1921 , n1055 );
and ( n3051 , n2122 , n970 );
nor ( n3052 , n3050 , n3051 );
xnor ( n3053 , n3052 , n1036 );
xor ( n3054 , n3049 , n3053 );
and ( n3055 , n1349 , n1482 );
and ( n3056 , n1500 , n1381 );
nor ( n3057 , n3055 , n3056 );
xnor ( n3058 , n3057 , n1472 );
xor ( n3059 , n3054 , n3058 );
xor ( n3060 , n3048 , n3059 );
and ( n3061 , n1630 , n1241 );
and ( n3062 , n1747 , n1148 );
nor ( n3063 , n3061 , n3062 );
xnor ( n3064 , n3063 , n1247 );
and ( n3065 , n1137 , n1800 );
and ( n3066 , n1228 , n1656 );
nor ( n3067 , n3065 , n3066 );
xnor ( n3068 , n3067 , n1756 );
xor ( n3069 , n3064 , n3068 );
and ( n3070 , n959 , n2100 );
and ( n3071 , n1027 , n1932 );
nor ( n3072 , n3070 , n3071 );
xnor ( n3073 , n3072 , n2106 );
xor ( n3074 , n3069 , n3073 );
xor ( n3075 , n3060 , n3074 );
xor ( n3076 , n3044 , n3075 );
and ( n3077 , n2915 , n2919 );
and ( n3078 , n2919 , n2924 );
and ( n3079 , n2915 , n2924 );
or ( n3080 , n3077 , n3078 , n3079 );
and ( n3081 , n2930 , n2944 );
and ( n3082 , n2944 , n2956 );
and ( n3083 , n2930 , n2956 );
or ( n3084 , n3081 , n3082 , n3083 );
xor ( n3085 , n3080 , n3084 );
and ( n3086 , n2934 , n2938 );
and ( n3087 , n2938 , n2943 );
and ( n3088 , n2934 , n2943 );
or ( n3089 , n3086 , n3087 , n3088 );
buf ( n3090 , n2923 );
xor ( n3091 , n3089 , n3090 );
and ( n3092 , n875 , n2097 );
xor ( n3093 , n3091 , n3092 );
xor ( n3094 , n3085 , n3093 );
xor ( n3095 , n3076 , n3094 );
and ( n3096 , n2902 , n2906 );
and ( n3097 , n2906 , n2958 );
and ( n3098 , n2902 , n2958 );
or ( n3099 , n3096 , n3097 , n3098 );
xor ( n3100 , n3095 , n3099 );
and ( n3101 , n2898 , n2959 );
and ( n3102 , n2960 , n2963 );
or ( n3103 , n3101 , n3102 );
xor ( n3104 , n3100 , n3103 );
buf ( n3105 , n3104 );
and ( n3106 , n916 , n2184 );
and ( n3107 , n3008 , n3012 );
and ( n3108 , n3012 , n3017 );
and ( n3109 , n3008 , n3017 );
or ( n3110 , n3107 , n3108 , n3109 );
xor ( n3111 , n3106 , n3110 );
and ( n3112 , n2985 , n2989 );
and ( n3113 , n2989 , n2991 );
and ( n3114 , n2985 , n2991 );
or ( n3115 , n3112 , n3113 , n3114 );
not ( n3116 , n925 );
and ( n3117 , n1993 , n1110 );
and ( n3118 , n2208 , n1007 );
nor ( n3119 , n3117 , n3118 );
xnor ( n3120 , n3119 , n1096 );
xor ( n3121 , n3116 , n3120 );
and ( n3122 , n1411 , n1542 );
and ( n3123 , n1575 , n1442 );
nor ( n3124 , n3122 , n3123 );
xnor ( n3125 , n3124 , n1548 );
xor ( n3126 , n3121 , n3125 );
xor ( n3127 , n3115 , n3126 );
and ( n3128 , n1677 , n1322 );
and ( n3129 , n1872 , n1199 );
nor ( n3130 , n3128 , n3129 );
xnor ( n3131 , n3130 , n1296 );
and ( n3132 , n1189 , n1830 );
and ( n3133 , n1311 , n1716 );
nor ( n3134 , n3132 , n3133 );
xnor ( n3135 , n3134 , n1836 );
xor ( n3136 , n3131 , n3135 );
and ( n3137 , n996 , n2187 );
and ( n3138 , n1087 , n2004 );
nor ( n3139 , n3137 , n3138 );
xnor ( n3140 , n3139 , n2193 );
xor ( n3141 , n3136 , n3140 );
xor ( n3142 , n3127 , n3141 );
xor ( n3143 , n3111 , n3142 );
and ( n3144 , n2981 , n2992 );
and ( n3145 , n2992 , n2994 );
and ( n3146 , n2981 , n2994 );
or ( n3147 , n3144 , n3145 , n3146 );
and ( n3148 , n3000 , n3004 );
and ( n3149 , n3004 , n3018 );
and ( n3150 , n3000 , n3018 );
or ( n3151 , n3148 , n3149 , n3150 );
xor ( n3152 , n3147 , n3151 );
and ( n3153 , n2977 , n2995 );
and ( n3154 , n2995 , n3019 );
and ( n3155 , n2977 , n3019 );
or ( n3156 , n3153 , n3154 , n3155 );
xor ( n3157 , n3152 , n3156 );
xor ( n3158 , n3143 , n3157 );
and ( n3159 , n2973 , n3020 );
and ( n3160 , n3020 , n3025 );
and ( n3161 , n2973 , n3025 );
or ( n3162 , n3159 , n3160 , n3161 );
xor ( n3163 , n3158 , n3162 );
and ( n3164 , n2969 , n3026 );
and ( n3165 , n3026 , n3031 );
and ( n3166 , n2969 , n3031 );
or ( n3167 , n3164 , n3165 , n3166 );
xor ( n3168 , n3163 , n3167 );
and ( n3169 , n3033 , n3034 );
or ( n3170 , n3032 , n3169 );
xor ( n3171 , n3168 , n3170 );
buf ( n3172 , n3171 );
not ( n3173 , n455 );
and ( n3174 , n3173 , n3105 );
and ( n3175 , n3172 , n455 );
or ( n3176 , n3174 , n3175 );
and ( n3177 , n3080 , n3084 );
and ( n3178 , n3084 , n3093 );
and ( n3179 , n3080 , n3093 );
or ( n3180 , n3177 , n3178 , n3179 );
and ( n3181 , n3049 , n3053 );
and ( n3182 , n3053 , n3058 );
and ( n3183 , n3049 , n3058 );
or ( n3184 , n3181 , n3182 , n3183 );
and ( n3185 , n3064 , n3068 );
and ( n3186 , n3068 , n3073 );
and ( n3187 , n3064 , n3073 );
or ( n3188 , n3185 , n3186 , n3187 );
xor ( n3189 , n3184 , n3188 );
and ( n3190 , n2122 , n1055 );
not ( n3191 , n3190 );
xnor ( n3192 , n3191 , n1036 );
and ( n3193 , n1228 , n1800 );
and ( n3194 , n1349 , n1656 );
nor ( n3195 , n3193 , n3194 );
xnor ( n3196 , n3195 , n1756 );
xor ( n3197 , n3192 , n3196 );
and ( n3198 , n1027 , n2100 );
and ( n3199 , n1137 , n1932 );
nor ( n3200 , n3198 , n3199 );
xnor ( n3201 , n3200 , n2106 );
xor ( n3202 , n3197 , n3201 );
xor ( n3203 , n3189 , n3202 );
xor ( n3204 , n3180 , n3203 );
and ( n3205 , n3089 , n3090 );
and ( n3206 , n3090 , n3092 );
and ( n3207 , n3089 , n3092 );
or ( n3208 , n3205 , n3206 , n3207 );
and ( n3209 , n3048 , n3059 );
and ( n3210 , n3059 , n3074 );
and ( n3211 , n3048 , n3074 );
or ( n3212 , n3209 , n3210 , n3211 );
xor ( n3213 , n3208 , n3212 );
and ( n3214 , n1747 , n1241 );
and ( n3215 , n1921 , n1148 );
nor ( n3216 , n3214 , n3215 );
xnor ( n3217 , n3216 , n1247 );
not ( n3218 , n3217 );
and ( n3219 , n1500 , n1482 );
and ( n3220 , n1630 , n1381 );
nor ( n3221 , n3219 , n3220 );
xnor ( n3222 , n3221 , n1472 );
xor ( n3223 , n3218 , n3222 );
and ( n3224 , n959 , n2097 );
xor ( n3225 , n3223 , n3224 );
xor ( n3226 , n3213 , n3225 );
xor ( n3227 , n3204 , n3226 );
and ( n3228 , n3044 , n3075 );
and ( n3229 , n3075 , n3094 );
and ( n3230 , n3044 , n3094 );
or ( n3231 , n3228 , n3229 , n3230 );
xor ( n3232 , n3227 , n3231 );
and ( n3233 , n3095 , n3099 );
and ( n3234 , n3100 , n3103 );
or ( n3235 , n3233 , n3234 );
xor ( n3236 , n3232 , n3235 );
buf ( n3237 , n3236 );
and ( n3238 , n3106 , n3110 );
and ( n3239 , n3110 , n3142 );
and ( n3240 , n3106 , n3142 );
or ( n3241 , n3238 , n3239 , n3240 );
and ( n3242 , n1872 , n1322 );
and ( n3243 , n1993 , n1199 );
nor ( n3244 , n3242 , n3243 );
xnor ( n3245 , n3244 , n1296 );
not ( n3246 , n3245 );
and ( n3247 , n1575 , n1542 );
and ( n3248 , n1677 , n1442 );
nor ( n3249 , n3247 , n3248 );
xnor ( n3250 , n3249 , n1548 );
xor ( n3251 , n3246 , n3250 );
and ( n3252 , n996 , n2184 );
xor ( n3253 , n3251 , n3252 );
and ( n3254 , n3116 , n3120 );
and ( n3255 , n3120 , n3125 );
and ( n3256 , n3116 , n3125 );
or ( n3257 , n3254 , n3255 , n3256 );
and ( n3258 , n3131 , n3135 );
and ( n3259 , n3135 , n3140 );
and ( n3260 , n3131 , n3140 );
or ( n3261 , n3258 , n3259 , n3260 );
xor ( n3262 , n3257 , n3261 );
and ( n3263 , n2208 , n1110 );
not ( n3264 , n3263 );
xnor ( n3265 , n3264 , n1096 );
and ( n3266 , n1311 , n1830 );
and ( n3267 , n1411 , n1716 );
nor ( n3268 , n3266 , n3267 );
xnor ( n3269 , n3268 , n1836 );
xor ( n3270 , n3265 , n3269 );
and ( n3271 , n1087 , n2187 );
and ( n3272 , n1189 , n2004 );
nor ( n3273 , n3271 , n3272 );
xnor ( n3274 , n3273 , n2193 );
xor ( n3275 , n3270 , n3274 );
xor ( n3276 , n3262 , n3275 );
xor ( n3277 , n3253 , n3276 );
and ( n3278 , n3115 , n3126 );
and ( n3279 , n3126 , n3141 );
and ( n3280 , n3115 , n3141 );
or ( n3281 , n3278 , n3279 , n3280 );
xor ( n3282 , n3277 , n3281 );
xor ( n3283 , n3241 , n3282 );
and ( n3284 , n3147 , n3151 );
and ( n3285 , n3151 , n3156 );
and ( n3286 , n3147 , n3156 );
or ( n3287 , n3284 , n3285 , n3286 );
xor ( n3288 , n3283 , n3287 );
and ( n3289 , n3143 , n3157 );
and ( n3290 , n3157 , n3162 );
and ( n3291 , n3143 , n3162 );
or ( n3292 , n3289 , n3290 , n3291 );
xor ( n3293 , n3288 , n3292 );
and ( n3294 , n3163 , n3167 );
and ( n3295 , n3168 , n3170 );
or ( n3296 , n3294 , n3295 );
xor ( n3297 , n3293 , n3296 );
buf ( n3298 , n3297 );
not ( n3299 , n455 );
and ( n3300 , n3299 , n3237 );
and ( n3301 , n3298 , n455 );
or ( n3302 , n3300 , n3301 );
and ( n3303 , n3184 , n3188 );
and ( n3304 , n3188 , n3202 );
and ( n3305 , n3184 , n3202 );
or ( n3306 , n3303 , n3304 , n3305 );
and ( n3307 , n3208 , n3212 );
and ( n3308 , n3212 , n3225 );
and ( n3309 , n3208 , n3225 );
or ( n3310 , n3307 , n3308 , n3309 );
xor ( n3311 , n3306 , n3310 );
and ( n3312 , n3218 , n3222 );
and ( n3313 , n3222 , n3224 );
and ( n3314 , n3218 , n3224 );
or ( n3315 , n3312 , n3313 , n3314 );
not ( n3316 , n1036 );
and ( n3317 , n1921 , n1241 );
and ( n3318 , n2122 , n1148 );
nor ( n3319 , n3317 , n3318 );
xnor ( n3320 , n3319 , n1247 );
xor ( n3321 , n3316 , n3320 );
and ( n3322 , n1349 , n1800 );
and ( n3323 , n1500 , n1656 );
nor ( n3324 , n3322 , n3323 );
xnor ( n3325 , n3324 , n1756 );
xor ( n3326 , n3321 , n3325 );
xor ( n3327 , n3315 , n3326 );
and ( n3328 , n3192 , n3196 );
and ( n3329 , n3196 , n3201 );
and ( n3330 , n3192 , n3201 );
or ( n3331 , n3328 , n3329 , n3330 );
buf ( n3332 , n3217 );
xor ( n3333 , n3331 , n3332 );
and ( n3334 , n1630 , n1482 );
and ( n3335 , n1747 , n1381 );
nor ( n3336 , n3334 , n3335 );
xnor ( n3337 , n3336 , n1472 );
and ( n3338 , n1137 , n2100 );
and ( n3339 , n1228 , n1932 );
nor ( n3340 , n3338 , n3339 );
xnor ( n3341 , n3340 , n2106 );
xor ( n3342 , n3337 , n3341 );
and ( n3343 , n1027 , n2097 );
xor ( n3344 , n3342 , n3343 );
xor ( n3345 , n3333 , n3344 );
xor ( n3346 , n3327 , n3345 );
xor ( n3347 , n3311 , n3346 );
and ( n3348 , n3180 , n3203 );
and ( n3349 , n3203 , n3226 );
and ( n3350 , n3180 , n3226 );
or ( n3351 , n3348 , n3349 , n3350 );
xor ( n3352 , n3347 , n3351 );
and ( n3353 , n3227 , n3231 );
and ( n3354 , n3232 , n3235 );
or ( n3355 , n3353 , n3354 );
xor ( n3356 , n3352 , n3355 );
buf ( n3357 , n3356 );
and ( n3358 , n3257 , n3261 );
and ( n3359 , n3261 , n3275 );
and ( n3360 , n3257 , n3275 );
or ( n3361 , n3358 , n3359 , n3360 );
and ( n3362 , n3246 , n3250 );
and ( n3363 , n3250 , n3252 );
and ( n3364 , n3246 , n3252 );
or ( n3365 , n3362 , n3363 , n3364 );
not ( n3366 , n1096 );
and ( n3367 , n1993 , n1322 );
and ( n3368 , n2208 , n1199 );
nor ( n3369 , n3367 , n3368 );
xnor ( n3370 , n3369 , n1296 );
xor ( n3371 , n3366 , n3370 );
and ( n3372 , n1411 , n1830 );
and ( n3373 , n1575 , n1716 );
nor ( n3374 , n3372 , n3373 );
xnor ( n3375 , n3374 , n1836 );
xor ( n3376 , n3371 , n3375 );
xor ( n3377 , n3365 , n3376 );
and ( n3378 , n3265 , n3269 );
and ( n3379 , n3269 , n3274 );
and ( n3380 , n3265 , n3274 );
or ( n3381 , n3378 , n3379 , n3380 );
buf ( n3382 , n3245 );
xor ( n3383 , n3381 , n3382 );
and ( n3384 , n1677 , n1542 );
and ( n3385 , n1872 , n1442 );
nor ( n3386 , n3384 , n3385 );
xnor ( n3387 , n3386 , n1548 );
and ( n3388 , n1189 , n2187 );
and ( n3389 , n1311 , n2004 );
nor ( n3390 , n3388 , n3389 );
xnor ( n3391 , n3390 , n2193 );
xor ( n3392 , n3387 , n3391 );
and ( n3393 , n1087 , n2184 );
xor ( n3394 , n3392 , n3393 );
xor ( n3395 , n3383 , n3394 );
xor ( n3396 , n3377 , n3395 );
xor ( n3397 , n3361 , n3396 );
and ( n3398 , n3253 , n3276 );
and ( n3399 , n3276 , n3281 );
and ( n3400 , n3253 , n3281 );
or ( n3401 , n3398 , n3399 , n3400 );
xor ( n3402 , n3397 , n3401 );
and ( n3403 , n3241 , n3282 );
and ( n3404 , n3282 , n3287 );
and ( n3405 , n3241 , n3287 );
or ( n3406 , n3403 , n3404 , n3405 );
xor ( n3407 , n3402 , n3406 );
and ( n3408 , n3288 , n3292 );
and ( n3409 , n3293 , n3296 );
or ( n3410 , n3408 , n3409 );
xor ( n3411 , n3407 , n3410 );
buf ( n3412 , n3411 );
not ( n3413 , n455 );
and ( n3414 , n3413 , n3357 );
and ( n3415 , n3412 , n455 );
or ( n3416 , n3414 , n3415 );
and ( n3417 , n3331 , n3332 );
and ( n3418 , n3332 , n3344 );
and ( n3419 , n3331 , n3344 );
or ( n3420 , n3417 , n3418 , n3419 );
and ( n3421 , n3315 , n3326 );
and ( n3422 , n3326 , n3345 );
and ( n3423 , n3315 , n3345 );
or ( n3424 , n3421 , n3422 , n3423 );
xor ( n3425 , n3420 , n3424 );
and ( n3426 , n3316 , n3320 );
and ( n3427 , n3320 , n3325 );
and ( n3428 , n3316 , n3325 );
or ( n3429 , n3426 , n3427 , n3428 );
and ( n3430 , n2122 , n1241 );
not ( n3431 , n3430 );
xnor ( n3432 , n3431 , n1247 );
and ( n3433 , n1228 , n2100 );
and ( n3434 , n1349 , n1932 );
nor ( n3435 , n3433 , n3434 );
xnor ( n3436 , n3435 , n2106 );
xor ( n3437 , n3432 , n3436 );
and ( n3438 , n1137 , n2097 );
xor ( n3439 , n3437 , n3438 );
xor ( n3440 , n3429 , n3439 );
and ( n3441 , n3337 , n3341 );
and ( n3442 , n3341 , n3343 );
and ( n3443 , n3337 , n3343 );
or ( n3444 , n3441 , n3442 , n3443 );
and ( n3445 , n1747 , n1482 );
and ( n3446 , n1921 , n1381 );
nor ( n3447 , n3445 , n3446 );
xnor ( n3448 , n3447 , n1472 );
not ( n3449 , n3448 );
xor ( n3450 , n3444 , n3449 );
and ( n3451 , n1500 , n1800 );
and ( n3452 , n1630 , n1656 );
nor ( n3453 , n3451 , n3452 );
xnor ( n3454 , n3453 , n1756 );
xor ( n3455 , n3450 , n3454 );
xor ( n3456 , n3440 , n3455 );
xor ( n3457 , n3425 , n3456 );
and ( n3458 , n3306 , n3310 );
and ( n3459 , n3310 , n3346 );
and ( n3460 , n3306 , n3346 );
or ( n3461 , n3458 , n3459 , n3460 );
xor ( n3462 , n3457 , n3461 );
and ( n3463 , n3347 , n3351 );
and ( n3464 , n3352 , n3355 );
or ( n3465 , n3463 , n3464 );
xor ( n3466 , n3462 , n3465 );
buf ( n3467 , n3466 );
and ( n3468 , n3381 , n3382 );
and ( n3469 , n3382 , n3394 );
and ( n3470 , n3381 , n3394 );
or ( n3471 , n3468 , n3469 , n3470 );
and ( n3472 , n3365 , n3376 );
and ( n3473 , n3376 , n3395 );
and ( n3474 , n3365 , n3395 );
or ( n3475 , n3472 , n3473 , n3474 );
xor ( n3476 , n3471 , n3475 );
and ( n3477 , n3366 , n3370 );
and ( n3478 , n3370 , n3375 );
and ( n3479 , n3366 , n3375 );
or ( n3480 , n3477 , n3478 , n3479 );
and ( n3481 , n2208 , n1322 );
not ( n3482 , n3481 );
xnor ( n3483 , n3482 , n1296 );
and ( n3484 , n1311 , n2187 );
and ( n3485 , n1411 , n2004 );
nor ( n3486 , n3484 , n3485 );
xnor ( n3487 , n3486 , n2193 );
xor ( n3488 , n3483 , n3487 );
and ( n3489 , n1189 , n2184 );
xor ( n3490 , n3488 , n3489 );
xor ( n3491 , n3480 , n3490 );
and ( n3492 , n3387 , n3391 );
and ( n3493 , n3391 , n3393 );
and ( n3494 , n3387 , n3393 );
or ( n3495 , n3492 , n3493 , n3494 );
and ( n3496 , n1872 , n1542 );
and ( n3497 , n1993 , n1442 );
nor ( n3498 , n3496 , n3497 );
xnor ( n3499 , n3498 , n1548 );
not ( n3500 , n3499 );
xor ( n3501 , n3495 , n3500 );
and ( n3502 , n1575 , n1830 );
and ( n3503 , n1677 , n1716 );
nor ( n3504 , n3502 , n3503 );
xnor ( n3505 , n3504 , n1836 );
xor ( n3506 , n3501 , n3505 );
xor ( n3507 , n3491 , n3506 );
xor ( n3508 , n3476 , n3507 );
and ( n3509 , n3361 , n3396 );
and ( n3510 , n3396 , n3401 );
and ( n3511 , n3361 , n3401 );
or ( n3512 , n3509 , n3510 , n3511 );
xor ( n3513 , n3508 , n3512 );
and ( n3514 , n3402 , n3406 );
and ( n3515 , n3407 , n3410 );
or ( n3516 , n3514 , n3515 );
xor ( n3517 , n3513 , n3516 );
buf ( n3518 , n3517 );
not ( n3519 , n455 );
and ( n3520 , n3519 , n3467 );
and ( n3521 , n3518 , n455 );
or ( n3522 , n3520 , n3521 );
and ( n3523 , n3420 , n3424 );
and ( n3524 , n3424 , n3456 );
and ( n3525 , n3420 , n3456 );
or ( n3526 , n3523 , n3524 , n3525 );
and ( n3527 , n3444 , n3449 );
and ( n3528 , n3449 , n3454 );
and ( n3529 , n3444 , n3454 );
or ( n3530 , n3527 , n3528 , n3529 );
and ( n3531 , n3429 , n3439 );
and ( n3532 , n3439 , n3455 );
and ( n3533 , n3429 , n3455 );
or ( n3534 , n3531 , n3532 , n3533 );
xor ( n3535 , n3530 , n3534 );
and ( n3536 , n3432 , n3436 );
and ( n3537 , n3436 , n3438 );
and ( n3538 , n3432 , n3438 );
or ( n3539 , n3536 , n3537 , n3538 );
not ( n3540 , n1247 );
and ( n3541 , n1921 , n1482 );
and ( n3542 , n2122 , n1381 );
nor ( n3543 , n3541 , n3542 );
xnor ( n3544 , n3543 , n1472 );
xor ( n3545 , n3540 , n3544 );
and ( n3546 , n1349 , n2100 );
and ( n3547 , n1500 , n1932 );
nor ( n3548 , n3546 , n3547 );
xnor ( n3549 , n3548 , n2106 );
xor ( n3550 , n3545 , n3549 );
xor ( n3551 , n3539 , n3550 );
buf ( n3552 , n3448 );
and ( n3553 , n1630 , n1800 );
and ( n3554 , n1747 , n1656 );
nor ( n3555 , n3553 , n3554 );
xnor ( n3556 , n3555 , n1756 );
xor ( n3557 , n3552 , n3556 );
and ( n3558 , n1228 , n2097 );
xor ( n3559 , n3557 , n3558 );
xor ( n3560 , n3551 , n3559 );
xor ( n3561 , n3535 , n3560 );
xor ( n3562 , n3526 , n3561 );
and ( n3563 , n3457 , n3461 );
and ( n3564 , n3462 , n3465 );
or ( n3565 , n3563 , n3564 );
xor ( n3566 , n3562 , n3565 );
buf ( n3567 , n3566 );
and ( n3568 , n3471 , n3475 );
and ( n3569 , n3475 , n3507 );
and ( n3570 , n3471 , n3507 );
or ( n3571 , n3568 , n3569 , n3570 );
and ( n3572 , n3495 , n3500 );
and ( n3573 , n3500 , n3505 );
and ( n3574 , n3495 , n3505 );
or ( n3575 , n3572 , n3573 , n3574 );
and ( n3576 , n3480 , n3490 );
and ( n3577 , n3490 , n3506 );
and ( n3578 , n3480 , n3506 );
or ( n3579 , n3576 , n3577 , n3578 );
xor ( n3580 , n3575 , n3579 );
and ( n3581 , n3483 , n3487 );
and ( n3582 , n3487 , n3489 );
and ( n3583 , n3483 , n3489 );
or ( n3584 , n3581 , n3582 , n3583 );
not ( n3585 , n1296 );
and ( n3586 , n1993 , n1542 );
and ( n3587 , n2208 , n1442 );
nor ( n3588 , n3586 , n3587 );
xnor ( n3589 , n3588 , n1548 );
xor ( n3590 , n3585 , n3589 );
and ( n3591 , n1411 , n2187 );
and ( n3592 , n1575 , n2004 );
nor ( n3593 , n3591 , n3592 );
xnor ( n3594 , n3593 , n2193 );
xor ( n3595 , n3590 , n3594 );
xor ( n3596 , n3584 , n3595 );
buf ( n3597 , n3499 );
and ( n3598 , n1677 , n1830 );
and ( n3599 , n1872 , n1716 );
nor ( n3600 , n3598 , n3599 );
xnor ( n3601 , n3600 , n1836 );
xor ( n3602 , n3597 , n3601 );
and ( n3603 , n1311 , n2184 );
xor ( n3604 , n3602 , n3603 );
xor ( n3605 , n3596 , n3604 );
xor ( n3606 , n3580 , n3605 );
xor ( n3607 , n3571 , n3606 );
and ( n3608 , n3508 , n3512 );
and ( n3609 , n3513 , n3516 );
or ( n3610 , n3608 , n3609 );
xor ( n3611 , n3607 , n3610 );
buf ( n3612 , n3611 );
not ( n3613 , n455 );
and ( n3614 , n3613 , n3567 );
and ( n3615 , n3612 , n455 );
or ( n3616 , n3614 , n3615 );
and ( n3617 , n3552 , n3556 );
and ( n3618 , n3556 , n3558 );
and ( n3619 , n3552 , n3558 );
or ( n3620 , n3617 , n3618 , n3619 );
and ( n3621 , n3539 , n3550 );
and ( n3622 , n3550 , n3559 );
and ( n3623 , n3539 , n3559 );
or ( n3624 , n3621 , n3622 , n3623 );
xor ( n3625 , n3620 , n3624 );
and ( n3626 , n3540 , n3544 );
and ( n3627 , n3544 , n3549 );
and ( n3628 , n3540 , n3549 );
or ( n3629 , n3626 , n3627 , n3628 );
and ( n3630 , n2122 , n1482 );
not ( n3631 , n3630 );
xnor ( n3632 , n3631 , n1472 );
not ( n3633 , n3632 );
xor ( n3634 , n3629 , n3633 );
and ( n3635 , n1747 , n1800 );
and ( n3636 , n1921 , n1656 );
nor ( n3637 , n3635 , n3636 );
xnor ( n3638 , n3637 , n1756 );
and ( n3639 , n1500 , n2100 );
and ( n3640 , n1630 , n1932 );
nor ( n3641 , n3639 , n3640 );
xnor ( n3642 , n3641 , n2106 );
xor ( n3643 , n3638 , n3642 );
and ( n3644 , n1349 , n2097 );
xor ( n3645 , n3643 , n3644 );
xor ( n3646 , n3634 , n3645 );
xor ( n3647 , n3625 , n3646 );
and ( n3648 , n3530 , n3534 );
and ( n3649 , n3534 , n3560 );
and ( n3650 , n3530 , n3560 );
or ( n3651 , n3648 , n3649 , n3650 );
xor ( n3652 , n3647 , n3651 );
and ( n3653 , n3526 , n3561 );
and ( n3654 , n3562 , n3565 );
or ( n3655 , n3653 , n3654 );
xor ( n3656 , n3652 , n3655 );
buf ( n3657 , n3656 );
and ( n3658 , n3597 , n3601 );
and ( n3659 , n3601 , n3603 );
and ( n3660 , n3597 , n3603 );
or ( n3661 , n3658 , n3659 , n3660 );
and ( n3662 , n3584 , n3595 );
and ( n3663 , n3595 , n3604 );
and ( n3664 , n3584 , n3604 );
or ( n3665 , n3662 , n3663 , n3664 );
xor ( n3666 , n3661 , n3665 );
and ( n3667 , n3585 , n3589 );
and ( n3668 , n3589 , n3594 );
and ( n3669 , n3585 , n3594 );
or ( n3670 , n3667 , n3668 , n3669 );
and ( n3671 , n2208 , n1542 );
not ( n3672 , n3671 );
xnor ( n3673 , n3672 , n1548 );
not ( n3674 , n3673 );
xor ( n3675 , n3670 , n3674 );
and ( n3676 , n1872 , n1830 );
and ( n3677 , n1993 , n1716 );
nor ( n3678 , n3676 , n3677 );
xnor ( n3679 , n3678 , n1836 );
and ( n3680 , n1575 , n2187 );
and ( n3681 , n1677 , n2004 );
nor ( n3682 , n3680 , n3681 );
xnor ( n3683 , n3682 , n2193 );
xor ( n3684 , n3679 , n3683 );
and ( n3685 , n1411 , n2184 );
xor ( n3686 , n3684 , n3685 );
xor ( n3687 , n3675 , n3686 );
xor ( n3688 , n3666 , n3687 );
and ( n3689 , n3575 , n3579 );
and ( n3690 , n3579 , n3605 );
and ( n3691 , n3575 , n3605 );
or ( n3692 , n3689 , n3690 , n3691 );
xor ( n3693 , n3688 , n3692 );
and ( n3694 , n3571 , n3606 );
and ( n3695 , n3607 , n3610 );
or ( n3696 , n3694 , n3695 );
xor ( n3697 , n3693 , n3696 );
buf ( n3698 , n3697 );
not ( n3699 , n455 );
and ( n3700 , n3699 , n3657 );
and ( n3701 , n3698 , n455 );
or ( n3702 , n3700 , n3701 );
and ( n3703 , n3629 , n3633 );
and ( n3704 , n3633 , n3645 );
and ( n3705 , n3629 , n3645 );
or ( n3706 , n3703 , n3704 , n3705 );
not ( n3707 , n1472 );
and ( n3708 , n1921 , n1800 );
and ( n3709 , n2122 , n1656 );
nor ( n3710 , n3708 , n3709 );
xnor ( n3711 , n3710 , n1756 );
xor ( n3712 , n3707 , n3711 );
and ( n3713 , n1500 , n2097 );
xor ( n3714 , n3712 , n3713 );
xor ( n3715 , n3706 , n3714 );
and ( n3716 , n3638 , n3642 );
and ( n3717 , n3642 , n3644 );
and ( n3718 , n3638 , n3644 );
or ( n3719 , n3716 , n3717 , n3718 );
buf ( n3720 , n3632 );
xor ( n3721 , n3719 , n3720 );
and ( n3722 , n1630 , n2100 );
and ( n3723 , n1747 , n1932 );
nor ( n3724 , n3722 , n3723 );
xnor ( n3725 , n3724 , n2106 );
xor ( n3726 , n3721 , n3725 );
xor ( n3727 , n3715 , n3726 );
and ( n3728 , n3620 , n3624 );
and ( n3729 , n3624 , n3646 );
and ( n3730 , n3620 , n3646 );
or ( n3731 , n3728 , n3729 , n3730 );
xor ( n3732 , n3727 , n3731 );
and ( n3733 , n3647 , n3651 );
and ( n3734 , n3652 , n3655 );
or ( n3735 , n3733 , n3734 );
xor ( n3736 , n3732 , n3735 );
buf ( n3737 , n3736 );
and ( n3738 , n3670 , n3674 );
and ( n3739 , n3674 , n3686 );
and ( n3740 , n3670 , n3686 );
or ( n3741 , n3738 , n3739 , n3740 );
not ( n3742 , n1548 );
and ( n3743 , n1993 , n1830 );
and ( n3744 , n2208 , n1716 );
nor ( n3745 , n3743 , n3744 );
xnor ( n3746 , n3745 , n1836 );
xor ( n3747 , n3742 , n3746 );
and ( n3748 , n1575 , n2184 );
xor ( n3749 , n3747 , n3748 );
xor ( n3750 , n3741 , n3749 );
and ( n3751 , n3679 , n3683 );
and ( n3752 , n3683 , n3685 );
and ( n3753 , n3679 , n3685 );
or ( n3754 , n3751 , n3752 , n3753 );
buf ( n3755 , n3673 );
xor ( n3756 , n3754 , n3755 );
and ( n3757 , n1677 , n2187 );
and ( n3758 , n1872 , n2004 );
nor ( n3759 , n3757 , n3758 );
xnor ( n3760 , n3759 , n2193 );
xor ( n3761 , n3756 , n3760 );
xor ( n3762 , n3750 , n3761 );
and ( n3763 , n3661 , n3665 );
and ( n3764 , n3665 , n3687 );
and ( n3765 , n3661 , n3687 );
or ( n3766 , n3763 , n3764 , n3765 );
xor ( n3767 , n3762 , n3766 );
and ( n3768 , n3688 , n3692 );
and ( n3769 , n3693 , n3696 );
or ( n3770 , n3768 , n3769 );
xor ( n3771 , n3767 , n3770 );
buf ( n3772 , n3771 );
not ( n3773 , n455 );
and ( n3774 , n3773 , n3737 );
and ( n3775 , n3772 , n455 );
or ( n3776 , n3774 , n3775 );
and ( n3777 , n3706 , n3714 );
and ( n3778 , n3714 , n3726 );
and ( n3779 , n3706 , n3726 );
or ( n3780 , n3777 , n3778 , n3779 );
and ( n3781 , n2122 , n1800 );
not ( n3782 , n3781 );
xnor ( n3783 , n3782 , n1756 );
not ( n3784 , n3783 );
and ( n3785 , n1747 , n2100 );
and ( n3786 , n1921 , n1932 );
nor ( n3787 , n3785 , n3786 );
xnor ( n3788 , n3787 , n2106 );
xor ( n3789 , n3784 , n3788 );
and ( n3790 , n1630 , n2097 );
xor ( n3791 , n3789 , n3790 );
and ( n3792 , n3707 , n3711 );
and ( n3793 , n3711 , n3713 );
and ( n3794 , n3707 , n3713 );
or ( n3795 , n3792 , n3793 , n3794 );
xor ( n3796 , n3791 , n3795 );
and ( n3797 , n3719 , n3720 );
and ( n3798 , n3720 , n3725 );
and ( n3799 , n3719 , n3725 );
or ( n3800 , n3797 , n3798 , n3799 );
xor ( n3801 , n3796 , n3800 );
xor ( n3802 , n3780 , n3801 );
and ( n3803 , n3727 , n3731 );
and ( n3804 , n3732 , n3735 );
or ( n3805 , n3803 , n3804 );
xor ( n3806 , n3802 , n3805 );
buf ( n3807 , n3806 );
and ( n3808 , n3742 , n3746 );
and ( n3809 , n3746 , n3748 );
and ( n3810 , n3742 , n3748 );
or ( n3811 , n3808 , n3809 , n3810 );
and ( n3812 , n3754 , n3755 );
and ( n3813 , n3755 , n3760 );
and ( n3814 , n3754 , n3760 );
or ( n3815 , n3812 , n3813 , n3814 );
xor ( n3816 , n3811 , n3815 );
and ( n3817 , n2208 , n1830 );
not ( n3818 , n3817 );
xnor ( n3819 , n3818 , n1836 );
not ( n3820 , n3819 );
and ( n3821 , n1872 , n2187 );
and ( n3822 , n1993 , n2004 );
nor ( n3823 , n3821 , n3822 );
xnor ( n3824 , n3823 , n2193 );
xor ( n3825 , n3820 , n3824 );
and ( n3826 , n1677 , n2184 );
xor ( n3827 , n3825 , n3826 );
xor ( n3828 , n3816 , n3827 );
and ( n3829 , n3741 , n3749 );
and ( n3830 , n3749 , n3761 );
and ( n3831 , n3741 , n3761 );
or ( n3832 , n3829 , n3830 , n3831 );
xor ( n3833 , n3828 , n3832 );
and ( n3834 , n3762 , n3766 );
and ( n3835 , n3767 , n3770 );
or ( n3836 , n3834 , n3835 );
xor ( n3837 , n3833 , n3836 );
buf ( n3838 , n3837 );
not ( n3839 , n455 );
and ( n3840 , n3839 , n3807 );
and ( n3841 , n3838 , n455 );
or ( n3842 , n3840 , n3841 );
and ( n3843 , n3784 , n3788 );
and ( n3844 , n3788 , n3790 );
and ( n3845 , n3784 , n3790 );
or ( n3846 , n3843 , n3844 , n3845 );
buf ( n3847 , n3783 );
xor ( n3848 , n3846 , n3847 );
not ( n3849 , n1756 );
and ( n3850 , n1921 , n2100 );
and ( n3851 , n2122 , n1932 );
nor ( n3852 , n3850 , n3851 );
xnor ( n3853 , n3852 , n2106 );
xor ( n3854 , n3849 , n3853 );
and ( n3855 , n1747 , n2097 );
xor ( n3856 , n3854 , n3855 );
xor ( n3857 , n3848 , n3856 );
and ( n3858 , n3791 , n3795 );
and ( n3859 , n3795 , n3800 );
and ( n3860 , n3791 , n3800 );
or ( n3861 , n3858 , n3859 , n3860 );
xor ( n3862 , n3857 , n3861 );
and ( n3863 , n3780 , n3801 );
and ( n3864 , n3802 , n3805 );
or ( n3865 , n3863 , n3864 );
xor ( n3866 , n3862 , n3865 );
buf ( n3867 , n3866 );
and ( n3868 , n3820 , n3824 );
and ( n3869 , n3824 , n3826 );
and ( n3870 , n3820 , n3826 );
or ( n3871 , n3868 , n3869 , n3870 );
buf ( n3872 , n3819 );
xor ( n3873 , n3871 , n3872 );
not ( n3874 , n1836 );
and ( n3875 , n1993 , n2187 );
and ( n3876 , n2208 , n2004 );
nor ( n3877 , n3875 , n3876 );
xnor ( n3878 , n3877 , n2193 );
xor ( n3879 , n3874 , n3878 );
and ( n3880 , n1872 , n2184 );
xor ( n3881 , n3879 , n3880 );
xor ( n3882 , n3873 , n3881 );
and ( n3883 , n3811 , n3815 );
and ( n3884 , n3815 , n3827 );
and ( n3885 , n3811 , n3827 );
or ( n3886 , n3883 , n3884 , n3885 );
xor ( n3887 , n3882 , n3886 );
and ( n3888 , n3828 , n3832 );
and ( n3889 , n3833 , n3836 );
or ( n3890 , n3888 , n3889 );
xor ( n3891 , n3887 , n3890 );
buf ( n3892 , n3891 );
not ( n3893 , n455 );
and ( n3894 , n3893 , n3867 );
and ( n3895 , n3892 , n455 );
or ( n3896 , n3894 , n3895 );
and ( n3897 , n3849 , n3853 );
and ( n3898 , n3853 , n3855 );
and ( n3899 , n3849 , n3855 );
or ( n3900 , n3897 , n3898 , n3899 );
and ( n3901 , n2122 , n2100 );
not ( n3902 , n3901 );
xnor ( n3903 , n3902 , n2106 );
xor ( n3904 , n3900 , n3903 );
and ( n3905 , n1921 , n2097 );
not ( n3906 , n3905 );
xor ( n3907 , n3904 , n3906 );
and ( n3908 , n3846 , n3847 );
and ( n3909 , n3847 , n3856 );
and ( n3910 , n3846 , n3856 );
or ( n3911 , n3908 , n3909 , n3910 );
xor ( n3912 , n3907 , n3911 );
and ( n3913 , n3857 , n3861 );
and ( n3914 , n3862 , n3865 );
or ( n3915 , n3913 , n3914 );
xor ( n3916 , n3912 , n3915 );
buf ( n3917 , n3916 );
and ( n3918 , n3874 , n3878 );
and ( n3919 , n3878 , n3880 );
and ( n3920 , n3874 , n3880 );
or ( n3921 , n3918 , n3919 , n3920 );
and ( n3922 , n2208 , n2187 );
not ( n3923 , n3922 );
xnor ( n3924 , n3923 , n2193 );
xor ( n3925 , n3921 , n3924 );
and ( n3926 , n1993 , n2184 );
not ( n3927 , n3926 );
xor ( n3928 , n3925 , n3927 );
and ( n3929 , n3871 , n3872 );
and ( n3930 , n3872 , n3881 );
and ( n3931 , n3871 , n3881 );
or ( n3932 , n3929 , n3930 , n3931 );
xor ( n3933 , n3928 , n3932 );
and ( n3934 , n3882 , n3886 );
and ( n3935 , n3887 , n3890 );
or ( n3936 , n3934 , n3935 );
xor ( n3937 , n3933 , n3936 );
buf ( n3938 , n3937 );
not ( n3939 , n455 );
and ( n3940 , n3939 , n3917 );
and ( n3941 , n3938 , n455 );
or ( n3942 , n3940 , n3941 );
and ( n3943 , n3900 , n3903 );
and ( n3944 , n3903 , n3906 );
and ( n3945 , n3900 , n3906 );
or ( n3946 , n3943 , n3944 , n3945 );
buf ( n3947 , n3905 );
not ( n3948 , n2106 );
xor ( n3949 , n3947 , n3948 );
and ( n3950 , n2122 , n2097 );
xor ( n3951 , n3949 , n3950 );
xor ( n3952 , n3946 , n3951 );
and ( n3953 , n3907 , n3911 );
and ( n3954 , n3912 , n3915 );
or ( n3955 , n3953 , n3954 );
xor ( n3956 , n3952 , n3955 );
buf ( n3957 , n3956 );
and ( n3958 , n3921 , n3924 );
and ( n3959 , n3924 , n3927 );
and ( n3960 , n3921 , n3927 );
or ( n3961 , n3958 , n3959 , n3960 );
buf ( n3962 , n3926 );
not ( n3963 , n2193 );
xor ( n3964 , n3962 , n3963 );
and ( n3965 , n2208 , n2184 );
xor ( n3966 , n3964 , n3965 );
xor ( n3967 , n3961 , n3966 );
and ( n3968 , n3928 , n3932 );
and ( n3969 , n3933 , n3936 );
or ( n3970 , n3968 , n3969 );
xor ( n3971 , n3967 , n3970 );
buf ( n3972 , n3971 );
not ( n3973 , n455 );
and ( n3974 , n3973 , n3957 );
and ( n3975 , n3972 , n455 );
or ( n3976 , n3974 , n3975 );
buf ( n3977 , n504 );
buf ( n3978 , n3977 );
buf ( n3979 , n770 );
buf ( n3980 , n3979 );
and ( n3981 , n3978 , n3980 );
buf ( n3982 , n3981 );
buf ( n3983 , n3982 );
buf ( n3984 , n536 );
buf ( n3985 , n3984 );
buf ( n3986 , n550 );
buf ( n3987 , n3986 );
buf ( n3988 , n551 );
buf ( n3989 , n3988 );
xor ( n3990 , n3987 , n3989 );
and ( n3991 , n3985 , n3990 );
not ( n3992 , n3991 );
buf ( n3993 , n549 );
buf ( n3994 , n3993 );
and ( n3995 , n3987 , n3989 );
not ( n3996 , n3995 );
and ( n3997 , n3994 , n3996 );
and ( n3998 , n3992 , n3997 );
buf ( n3999 , n469 );
buf ( n4000 , n3999 );
and ( n4001 , n3998 , n4000 );
buf ( n4002 , n548 );
buf ( n4003 , n4002 );
xor ( n4004 , n4003 , n3994 );
and ( n4005 , n3985 , n4004 );
and ( n4006 , n4001 , n4005 );
buf ( n4007 , n468 );
buf ( n4008 , n4007 );
and ( n4009 , n4005 , n4008 );
and ( n4010 , n4001 , n4008 );
or ( n4011 , n4006 , n4009 , n4010 );
buf ( n4012 , n534 );
buf ( n4013 , n4012 );
xor ( n4014 , n3994 , n3987 );
not ( n4015 , n3990 );
and ( n4016 , n4014 , n4015 );
and ( n4017 , n4013 , n4016 );
buf ( n4018 , n533 );
buf ( n4019 , n4018 );
and ( n4020 , n4019 , n3990 );
nor ( n4021 , n4017 , n4020 );
xnor ( n4022 , n4021 , n3997 );
xor ( n4023 , n4011 , n4022 );
not ( n4024 , n4005 );
buf ( n4025 , n547 );
buf ( n4026 , n4025 );
and ( n4027 , n4003 , n3994 );
not ( n4028 , n4027 );
and ( n4029 , n4026 , n4028 );
and ( n4030 , n4024 , n4029 );
buf ( n4031 , n467 );
buf ( n4032 , n4031 );
xor ( n4033 , n4030 , n4032 );
buf ( n4034 , n532 );
buf ( n4035 , n4034 );
buf ( n4036 , n552 );
buf ( n4037 , n4036 );
xor ( n4038 , n3989 , n4037 );
not ( n4039 , n4037 );
and ( n4040 , n4038 , n4039 );
and ( n4041 , n4035 , n4040 );
buf ( n4042 , n531 );
buf ( n4043 , n4042 );
and ( n4044 , n4043 , n4037 );
nor ( n4045 , n4041 , n4044 );
xnor ( n4046 , n4045 , n3989 );
xor ( n4047 , n4033 , n4046 );
xor ( n4048 , n4026 , n4003 );
not ( n4049 , n4004 );
and ( n4050 , n4048 , n4049 );
and ( n4051 , n3985 , n4050 );
buf ( n4052 , n535 );
buf ( n4053 , n4052 );
and ( n4054 , n4053 , n4004 );
nor ( n4055 , n4051 , n4054 );
xnor ( n4056 , n4055 , n4029 );
xor ( n4057 , n4047 , n4056 );
xor ( n4058 , n4023 , n4057 );
and ( n4059 , n4019 , n4040 );
and ( n4060 , n4035 , n4037 );
nor ( n4061 , n4059 , n4060 );
xnor ( n4062 , n4061 , n3989 );
and ( n4063 , n4053 , n4016 );
and ( n4064 , n4013 , n3990 );
nor ( n4065 , n4063 , n4064 );
xnor ( n4066 , n4065 , n3997 );
and ( n4067 , n4062 , n4066 );
xor ( n4068 , n4001 , n4005 );
xor ( n4069 , n4068 , n4008 );
and ( n4070 , n4066 , n4069 );
and ( n4071 , n4062 , n4069 );
or ( n4072 , n4067 , n4070 , n4071 );
xor ( n4073 , n4058 , n4072 );
xor ( n4074 , n3998 , n4000 );
and ( n4075 , n4013 , n4040 );
and ( n4076 , n4019 , n4037 );
nor ( n4077 , n4075 , n4076 );
xnor ( n4078 , n4077 , n3989 );
and ( n4079 , n4074 , n4078 );
and ( n4080 , n3985 , n4016 );
and ( n4081 , n4053 , n3990 );
nor ( n4082 , n4080 , n4081 );
xnor ( n4083 , n4082 , n3997 );
and ( n4084 , n4078 , n4083 );
and ( n4085 , n4074 , n4083 );
or ( n4086 , n4079 , n4084 , n4085 );
xor ( n4087 , n4062 , n4066 );
xor ( n4088 , n4087 , n4069 );
and ( n4089 , n4086 , n4088 );
xor ( n4090 , n4086 , n4088 );
xor ( n4091 , n4074 , n4078 );
xor ( n4092 , n4091 , n4083 );
and ( n4093 , n3985 , n4037 );
not ( n4094 , n4093 );
and ( n4095 , n4094 , n3989 );
buf ( n4096 , n471 );
buf ( n4097 , n4096 );
and ( n4098 , n4095 , n4097 );
and ( n4099 , n4098 , n3991 );
buf ( n4100 , n470 );
buf ( n4101 , n4100 );
and ( n4102 , n3991 , n4101 );
and ( n4103 , n4098 , n4101 );
or ( n4104 , n4099 , n4102 , n4103 );
and ( n4105 , n4092 , n4104 );
xor ( n4106 , n4092 , n4104 );
and ( n4107 , n4053 , n4040 );
and ( n4108 , n4013 , n4037 );
nor ( n4109 , n4107 , n4108 );
xnor ( n4110 , n4109 , n3989 );
xor ( n4111 , n4098 , n3991 );
xor ( n4112 , n4111 , n4101 );
and ( n4113 , n4110 , n4112 );
xor ( n4114 , n4110 , n4112 );
and ( n4115 , n3985 , n4040 );
and ( n4116 , n4053 , n4037 );
nor ( n4117 , n4115 , n4116 );
xnor ( n4118 , n4117 , n3989 );
xor ( n4119 , n4095 , n4097 );
and ( n4120 , n4118 , n4119 );
xor ( n4121 , n4118 , n4119 );
buf ( n4122 , n472 );
buf ( n4123 , n4122 );
and ( n4124 , n4093 , n4123 );
and ( n4125 , n4121 , n4124 );
or ( n4126 , n4120 , n4125 );
and ( n4127 , n4114 , n4126 );
or ( n4128 , n4113 , n4127 );
and ( n4129 , n4106 , n4128 );
or ( n4130 , n4105 , n4129 );
and ( n4131 , n4090 , n4130 );
or ( n4132 , n4089 , n4131 );
xor ( n4133 , n4073 , n4132 );
buf ( n4134 , n4133 );
buf ( n4135 , n1221 );
buf ( n4136 , n547 );
xor ( n4137 , n4135 , n4136 );
buf ( n4138 , n1126 );
buf ( n4139 , n548 );
and ( n4140 , n4138 , n4139 );
buf ( n4141 , n1024 );
buf ( n4142 , n549 );
and ( n4143 , n4141 , n4142 );
buf ( n4144 , n950 );
buf ( n4145 , n550 );
and ( n4146 , n4144 , n4145 );
buf ( n4147 , n868 );
buf ( n4148 , n551 );
and ( n4149 , n4147 , n4148 );
buf ( n4150 , n814 );
buf ( n4151 , n552 );
and ( n4152 , n4150 , n4151 );
and ( n4153 , n4148 , n4152 );
and ( n4154 , n4147 , n4152 );
or ( n4155 , n4149 , n4153 , n4154 );
and ( n4156 , n4145 , n4155 );
and ( n4157 , n4144 , n4155 );
or ( n4158 , n4146 , n4156 , n4157 );
and ( n4159 , n4142 , n4158 );
and ( n4160 , n4141 , n4158 );
or ( n4161 , n4143 , n4159 , n4160 );
and ( n4162 , n4139 , n4161 );
and ( n4163 , n4138 , n4161 );
or ( n4164 , n4140 , n4162 , n4163 );
xor ( n4165 , n4137 , n4164 );
buf ( n4166 , n4165 );
not ( n4167 , n454 );
and ( n4168 , n4167 , n4134 );
and ( n4169 , n4166 , n454 );
or ( n4170 , n4168 , n4169 );
buf ( n4171 , n4170 );
buf ( n4172 , n472 );
xor ( n4173 , n4171 , n4172 );
buf ( n4174 , n4173 );
xor ( n4175 , n454 , n455 );
xor ( n4176 , n4175 , n456 );
not ( n4177 , n4176 );
and ( n4178 , n4177 , n3983 );
and ( n4179 , n4174 , n4176 );
or ( n4180 , n4178 , n4179 );
buf ( n4181 , n782 );
buf ( n4182 , n4181 );
xor ( n4183 , n4182 , n3980 );
not ( n4184 , n3980 );
and ( n4185 , n4183 , n4184 );
and ( n4186 , n3978 , n4185 );
buf ( n4187 , n503 );
buf ( n4188 , n4187 );
and ( n4189 , n4188 , n3980 );
nor ( n4190 , n4186 , n4189 );
xnor ( n4191 , n4190 , n4182 );
not ( n4192 , n3981 );
and ( n4193 , n4192 , n4182 );
xor ( n4194 , n4191 , n4193 );
buf ( n4195 , n4194 );
and ( n4196 , n4033 , n4046 );
and ( n4197 , n4046 , n4056 );
and ( n4198 , n4033 , n4056 );
or ( n4199 , n4196 , n4197 , n4198 );
and ( n4200 , n4053 , n4050 );
and ( n4201 , n4013 , n4004 );
nor ( n4202 , n4200 , n4201 );
xnor ( n4203 , n4202 , n4029 );
buf ( n4204 , n546 );
buf ( n4205 , n4204 );
xor ( n4206 , n4205 , n4026 );
and ( n4207 , n3985 , n4206 );
xor ( n4208 , n4203 , n4207 );
buf ( n4209 , n466 );
buf ( n4210 , n4209 );
xor ( n4211 , n4208 , n4210 );
xor ( n4212 , n4199 , n4211 );
and ( n4213 , n4030 , n4032 );
and ( n4214 , n4043 , n4040 );
buf ( n4215 , n530 );
buf ( n4216 , n4215 );
and ( n4217 , n4216 , n4037 );
nor ( n4218 , n4214 , n4217 );
xnor ( n4219 , n4218 , n3989 );
xor ( n4220 , n4213 , n4219 );
and ( n4221 , n4019 , n4016 );
and ( n4222 , n4035 , n3990 );
nor ( n4223 , n4221 , n4222 );
xnor ( n4224 , n4223 , n3997 );
xor ( n4225 , n4220 , n4224 );
xor ( n4226 , n4212 , n4225 );
and ( n4227 , n4011 , n4022 );
and ( n4228 , n4022 , n4057 );
and ( n4229 , n4011 , n4057 );
or ( n4230 , n4227 , n4228 , n4229 );
xor ( n4231 , n4226 , n4230 );
and ( n4232 , n4058 , n4072 );
and ( n4233 , n4073 , n4132 );
or ( n4234 , n4232 , n4233 );
xor ( n4235 , n4231 , n4234 );
buf ( n4236 , n4235 );
buf ( n4237 , n1342 );
buf ( n4238 , n546 );
xor ( n4239 , n4237 , n4238 );
and ( n4240 , n4135 , n4136 );
and ( n4241 , n4136 , n4164 );
and ( n4242 , n4135 , n4164 );
or ( n4243 , n4240 , n4241 , n4242 );
xor ( n4244 , n4239 , n4243 );
buf ( n4245 , n4244 );
not ( n4246 , n454 );
and ( n4247 , n4246 , n4236 );
and ( n4248 , n4245 , n454 );
or ( n4249 , n4247 , n4248 );
buf ( n4250 , n4249 );
buf ( n4251 , n471 );
xor ( n4252 , n4250 , n4251 );
and ( n4253 , n4171 , n4172 );
xor ( n4254 , n4252 , n4253 );
buf ( n4255 , n4254 );
not ( n4256 , n4176 );
and ( n4257 , n4256 , n4195 );
and ( n4258 , n4255 , n4176 );
or ( n4259 , n4257 , n4258 );
and ( n4260 , n4188 , n4185 );
buf ( n4261 , n502 );
buf ( n4262 , n4261 );
and ( n4263 , n4262 , n3980 );
nor ( n4264 , n4260 , n4263 );
xnor ( n4265 , n4264 , n4182 );
buf ( n4266 , n842 );
buf ( n4267 , n4266 );
xor ( n4268 , n4267 , n4182 );
and ( n4269 , n3978 , n4268 );
xor ( n4270 , n4265 , n4269 );
and ( n4271 , n4191 , n4193 );
xor ( n4272 , n4270 , n4271 );
buf ( n4273 , n4272 );
and ( n4274 , n4213 , n4219 );
and ( n4275 , n4219 , n4224 );
and ( n4276 , n4213 , n4224 );
or ( n4277 , n4274 , n4275 , n4276 );
and ( n4278 , n4203 , n4207 );
and ( n4279 , n4207 , n4210 );
and ( n4280 , n4203 , n4210 );
or ( n4281 , n4278 , n4279 , n4280 );
and ( n4282 , n4035 , n4016 );
and ( n4283 , n4043 , n3990 );
nor ( n4284 , n4282 , n4283 );
xnor ( n4285 , n4284 , n3997 );
xor ( n4286 , n4281 , n4285 );
buf ( n4287 , n545 );
buf ( n4288 , n4287 );
xor ( n4289 , n4288 , n4205 );
not ( n4290 , n4206 );
and ( n4291 , n4289 , n4290 );
and ( n4292 , n3985 , n4291 );
and ( n4293 , n4053 , n4206 );
nor ( n4294 , n4292 , n4293 );
and ( n4295 , n4205 , n4026 );
not ( n4296 , n4295 );
and ( n4297 , n4288 , n4296 );
xnor ( n4298 , n4294 , n4297 );
xor ( n4299 , n4286 , n4298 );
xor ( n4300 , n4277 , n4299 );
not ( n4301 , n4207 );
and ( n4302 , n4301 , n4297 );
buf ( n4303 , n465 );
buf ( n4304 , n4303 );
xor ( n4305 , n4302 , n4304 );
and ( n4306 , n4216 , n4040 );
buf ( n4307 , n529 );
buf ( n4308 , n4307 );
and ( n4309 , n4308 , n4037 );
nor ( n4310 , n4306 , n4309 );
xnor ( n4311 , n4310 , n3989 );
xor ( n4312 , n4305 , n4311 );
and ( n4313 , n4013 , n4050 );
and ( n4314 , n4019 , n4004 );
nor ( n4315 , n4313 , n4314 );
xnor ( n4316 , n4315 , n4029 );
xor ( n4317 , n4312 , n4316 );
xor ( n4318 , n4300 , n4317 );
and ( n4319 , n4199 , n4211 );
and ( n4320 , n4211 , n4225 );
and ( n4321 , n4199 , n4225 );
or ( n4322 , n4319 , n4320 , n4321 );
xor ( n4323 , n4318 , n4322 );
and ( n4324 , n4226 , n4230 );
and ( n4325 , n4231 , n4234 );
or ( n4326 , n4324 , n4325 );
xor ( n4327 , n4323 , n4326 );
buf ( n4328 , n4327 );
buf ( n4329 , n1458 );
buf ( n4330 , n545 );
xor ( n4331 , n4329 , n4330 );
and ( n4332 , n4237 , n4238 );
and ( n4333 , n4238 , n4243 );
and ( n4334 , n4237 , n4243 );
or ( n4335 , n4332 , n4333 , n4334 );
xor ( n4336 , n4331 , n4335 );
buf ( n4337 , n4336 );
not ( n4338 , n454 );
and ( n4339 , n4338 , n4328 );
and ( n4340 , n4337 , n454 );
or ( n4341 , n4339 , n4340 );
buf ( n4342 , n4341 );
buf ( n4343 , n470 );
xor ( n4344 , n4342 , n4343 );
and ( n4345 , n4250 , n4251 );
and ( n4346 , n4251 , n4253 );
and ( n4347 , n4250 , n4253 );
or ( n4348 , n4345 , n4346 , n4347 );
xor ( n4349 , n4344 , n4348 );
buf ( n4350 , n4349 );
not ( n4351 , n4176 );
and ( n4352 , n4351 , n4273 );
and ( n4353 , n4350 , n4176 );
or ( n4354 , n4352 , n4353 );
buf ( n4355 , n914 );
buf ( n4356 , n4355 );
xor ( n4357 , n4356 , n4267 );
not ( n4358 , n4268 );
and ( n4359 , n4357 , n4358 );
and ( n4360 , n3978 , n4359 );
and ( n4361 , n4188 , n4268 );
nor ( n4362 , n4360 , n4361 );
and ( n4363 , n4267 , n4182 );
not ( n4364 , n4363 );
and ( n4365 , n4356 , n4364 );
xnor ( n4366 , n4362 , n4365 );
and ( n4367 , n4262 , n4185 );
buf ( n4368 , n501 );
buf ( n4369 , n4368 );
and ( n4370 , n4369 , n3980 );
nor ( n4371 , n4367 , n4370 );
xnor ( n4372 , n4371 , n4182 );
not ( n4373 , n4269 );
and ( n4374 , n4373 , n4365 );
xor ( n4375 , n4372 , n4374 );
xor ( n4376 , n4366 , n4375 );
and ( n4377 , n4265 , n4269 );
and ( n4378 , n4270 , n4271 );
or ( n4379 , n4377 , n4378 );
xor ( n4380 , n4376 , n4379 );
buf ( n4381 , n4380 );
and ( n4382 , n4277 , n4299 );
and ( n4383 , n4299 , n4317 );
and ( n4384 , n4277 , n4317 );
or ( n4385 , n4382 , n4383 , n4384 );
and ( n4386 , n4281 , n4285 );
and ( n4387 , n4285 , n4298 );
and ( n4388 , n4281 , n4298 );
or ( n4389 , n4386 , n4387 , n4388 );
and ( n4390 , n4302 , n4304 );
and ( n4391 , n4019 , n4050 );
and ( n4392 , n4035 , n4004 );
nor ( n4393 , n4391 , n4392 );
xnor ( n4394 , n4393 , n4029 );
xor ( n4395 , n4390 , n4394 );
and ( n4396 , n4053 , n4291 );
and ( n4397 , n4013 , n4206 );
nor ( n4398 , n4396 , n4397 );
xnor ( n4399 , n4398 , n4297 );
xor ( n4400 , n4395 , n4399 );
xor ( n4401 , n4389 , n4400 );
and ( n4402 , n4305 , n4311 );
and ( n4403 , n4311 , n4316 );
and ( n4404 , n4305 , n4316 );
or ( n4405 , n4402 , n4403 , n4404 );
and ( n4406 , n4043 , n4016 );
and ( n4407 , n4216 , n3990 );
nor ( n4408 , n4406 , n4407 );
xnor ( n4409 , n4408 , n3997 );
xor ( n4410 , n4405 , n4409 );
and ( n4411 , n4308 , n4040 );
buf ( n4412 , n528 );
buf ( n4413 , n4412 );
and ( n4414 , n4413 , n4037 );
nor ( n4415 , n4411 , n4414 );
xnor ( n4416 , n4415 , n3989 );
buf ( n4417 , n544 );
buf ( n4418 , n4417 );
xor ( n4419 , n4418 , n4288 );
and ( n4420 , n3985 , n4419 );
xor ( n4421 , n4416 , n4420 );
buf ( n4422 , n464 );
buf ( n4423 , n4422 );
xor ( n4424 , n4421 , n4423 );
xor ( n4425 , n4410 , n4424 );
xor ( n4426 , n4401 , n4425 );
xor ( n4427 , n4385 , n4426 );
and ( n4428 , n4318 , n4322 );
and ( n4429 , n4323 , n4326 );
or ( n4430 , n4428 , n4429 );
xor ( n4431 , n4427 , n4430 );
buf ( n4432 , n4431 );
buf ( n4433 , n1603 );
buf ( n4434 , n544 );
xor ( n4435 , n4433 , n4434 );
and ( n4436 , n4329 , n4330 );
and ( n4437 , n4330 , n4335 );
and ( n4438 , n4329 , n4335 );
or ( n4439 , n4436 , n4437 , n4438 );
xor ( n4440 , n4435 , n4439 );
buf ( n4441 , n4440 );
not ( n4442 , n454 );
and ( n4443 , n4442 , n4432 );
and ( n4444 , n4441 , n454 );
or ( n4445 , n4443 , n4444 );
buf ( n4446 , n4445 );
buf ( n4447 , n469 );
xor ( n4448 , n4446 , n4447 );
and ( n4449 , n4342 , n4343 );
and ( n4450 , n4343 , n4348 );
and ( n4451 , n4342 , n4348 );
or ( n4452 , n4449 , n4450 , n4451 );
xor ( n4453 , n4448 , n4452 );
buf ( n4454 , n4453 );
not ( n4455 , n4176 );
and ( n4456 , n4455 , n4381 );
and ( n4457 , n4454 , n4176 );
or ( n4458 , n4456 , n4457 );
and ( n4459 , n4369 , n4185 );
buf ( n4460 , n500 );
buf ( n4461 , n4460 );
and ( n4462 , n4461 , n3980 );
nor ( n4463 , n4459 , n4462 );
xnor ( n4464 , n4463 , n4182 );
and ( n4465 , n4188 , n4359 );
and ( n4466 , n4262 , n4268 );
nor ( n4467 , n4465 , n4466 );
xnor ( n4468 , n4467 , n4365 );
xor ( n4469 , n4464 , n4468 );
buf ( n4470 , n994 );
buf ( n4471 , n4470 );
xor ( n4472 , n4471 , n4356 );
and ( n4473 , n3978 , n4472 );
xor ( n4474 , n4469 , n4473 );
and ( n4475 , n4372 , n4374 );
xor ( n4476 , n4474 , n4475 );
and ( n4477 , n4366 , n4375 );
and ( n4478 , n4376 , n4379 );
or ( n4479 , n4477 , n4478 );
xor ( n4480 , n4476 , n4479 );
buf ( n4481 , n4480 );
and ( n4482 , n4405 , n4409 );
and ( n4483 , n4409 , n4424 );
and ( n4484 , n4405 , n4424 );
or ( n4485 , n4482 , n4483 , n4484 );
and ( n4486 , n4216 , n4016 );
and ( n4487 , n4308 , n3990 );
nor ( n4488 , n4486 , n4487 );
xnor ( n4489 , n4488 , n3997 );
and ( n4490 , n4013 , n4291 );
and ( n4491 , n4019 , n4206 );
nor ( n4492 , n4490 , n4491 );
xnor ( n4493 , n4492 , n4297 );
xor ( n4494 , n4489 , n4493 );
buf ( n4495 , n543 );
buf ( n4496 , n4495 );
xor ( n4497 , n4496 , n4418 );
not ( n4498 , n4419 );
and ( n4499 , n4497 , n4498 );
and ( n4500 , n3985 , n4499 );
and ( n4501 , n4053 , n4419 );
nor ( n4502 , n4500 , n4501 );
and ( n4503 , n4418 , n4288 );
not ( n4504 , n4503 );
and ( n4505 , n4496 , n4504 );
xnor ( n4506 , n4502 , n4505 );
xor ( n4507 , n4494 , n4506 );
xor ( n4508 , n4485 , n4507 );
and ( n4509 , n4390 , n4394 );
and ( n4510 , n4394 , n4399 );
and ( n4511 , n4390 , n4399 );
or ( n4512 , n4509 , n4510 , n4511 );
and ( n4513 , n4416 , n4420 );
and ( n4514 , n4420 , n4423 );
and ( n4515 , n4416 , n4423 );
or ( n4516 , n4513 , n4514 , n4515 );
xor ( n4517 , n4512 , n4516 );
not ( n4518 , n4420 );
and ( n4519 , n4518 , n4505 );
buf ( n4520 , n463 );
buf ( n4521 , n4520 );
xor ( n4522 , n4519 , n4521 );
and ( n4523 , n4413 , n4040 );
buf ( n4524 , n527 );
buf ( n4525 , n4524 );
and ( n4526 , n4525 , n4037 );
nor ( n4527 , n4523 , n4526 );
xnor ( n4528 , n4527 , n3989 );
xor ( n4529 , n4522 , n4528 );
and ( n4530 , n4035 , n4050 );
and ( n4531 , n4043 , n4004 );
nor ( n4532 , n4530 , n4531 );
xnor ( n4533 , n4532 , n4029 );
xor ( n4534 , n4529 , n4533 );
xor ( n4535 , n4517 , n4534 );
xor ( n4536 , n4508 , n4535 );
and ( n4537 , n4389 , n4400 );
and ( n4538 , n4400 , n4425 );
and ( n4539 , n4389 , n4425 );
or ( n4540 , n4537 , n4538 , n4539 );
xor ( n4541 , n4536 , n4540 );
and ( n4542 , n4385 , n4426 );
and ( n4543 , n4427 , n4430 );
or ( n4544 , n4542 , n4543 );
xor ( n4545 , n4541 , n4544 );
buf ( n4546 , n4545 );
buf ( n4547 , n1740 );
buf ( n4548 , n543 );
xor ( n4549 , n4547 , n4548 );
and ( n4550 , n4433 , n4434 );
and ( n4551 , n4434 , n4439 );
and ( n4552 , n4433 , n4439 );
or ( n4553 , n4550 , n4551 , n4552 );
xor ( n4554 , n4549 , n4553 );
buf ( n4555 , n4554 );
not ( n4556 , n454 );
and ( n4557 , n4556 , n4546 );
and ( n4558 , n4555 , n454 );
or ( n4559 , n4557 , n4558 );
buf ( n4560 , n4559 );
and ( n4561 , n4446 , n4447 );
and ( n4562 , n4447 , n4452 );
and ( n4563 , n4446 , n4452 );
or ( n4564 , n4561 , n4562 , n4563 );
xor ( n4565 , n4560 , n4564 );
buf ( n4566 , n4565 );
not ( n4567 , n4176 );
and ( n4568 , n4567 , n4481 );
and ( n4569 , n4566 , n4176 );
or ( n4570 , n4568 , n4569 );
and ( n4571 , n4464 , n4468 );
and ( n4572 , n4468 , n4473 );
and ( n4573 , n4464 , n4473 );
or ( n4574 , n4571 , n4572 , n4573 );
and ( n4575 , n4461 , n4185 );
buf ( n4576 , n499 );
buf ( n4577 , n4576 );
and ( n4578 , n4577 , n3980 );
nor ( n4579 , n4575 , n4578 );
xnor ( n4580 , n4579 , n4182 );
not ( n4581 , n4473 );
buf ( n4582 , n1085 );
buf ( n4583 , n4582 );
and ( n4584 , n4471 , n4356 );
not ( n4585 , n4584 );
and ( n4586 , n4583 , n4585 );
and ( n4587 , n4581 , n4586 );
xor ( n4588 , n4580 , n4587 );
and ( n4589 , n4262 , n4359 );
and ( n4590 , n4369 , n4268 );
nor ( n4591 , n4589 , n4590 );
xnor ( n4592 , n4591 , n4365 );
xor ( n4593 , n4588 , n4592 );
xor ( n4594 , n4583 , n4471 );
not ( n4595 , n4472 );
and ( n4596 , n4594 , n4595 );
and ( n4597 , n3978 , n4596 );
and ( n4598 , n4188 , n4472 );
nor ( n4599 , n4597 , n4598 );
xnor ( n4600 , n4599 , n4586 );
xor ( n4601 , n4593 , n4600 );
xor ( n4602 , n4574 , n4601 );
and ( n4603 , n4474 , n4475 );
and ( n4604 , n4476 , n4479 );
or ( n4605 , n4603 , n4604 );
xor ( n4606 , n4602 , n4605 );
buf ( n4607 , n4606 );
and ( n4608 , n4512 , n4516 );
and ( n4609 , n4516 , n4534 );
and ( n4610 , n4512 , n4534 );
or ( n4611 , n4608 , n4609 , n4610 );
and ( n4612 , n4522 , n4528 );
and ( n4613 , n4528 , n4533 );
and ( n4614 , n4522 , n4533 );
or ( n4615 , n4612 , n4613 , n4614 );
and ( n4616 , n4308 , n4016 );
and ( n4617 , n4413 , n3990 );
nor ( n4618 , n4616 , n4617 );
xnor ( n4619 , n4618 , n3997 );
xor ( n4620 , n4615 , n4619 );
and ( n4621 , n4053 , n4499 );
and ( n4622 , n4013 , n4419 );
nor ( n4623 , n4621 , n4622 );
xnor ( n4624 , n4623 , n4505 );
xor ( n4625 , n4620 , n4624 );
xor ( n4626 , n4611 , n4625 );
and ( n4627 , n4489 , n4493 );
and ( n4628 , n4493 , n4506 );
and ( n4629 , n4489 , n4506 );
or ( n4630 , n4627 , n4628 , n4629 );
and ( n4631 , n4519 , n4521 );
and ( n4632 , n4043 , n4050 );
and ( n4633 , n4216 , n4004 );
nor ( n4634 , n4632 , n4633 );
xnor ( n4635 , n4634 , n4029 );
xor ( n4636 , n4631 , n4635 );
and ( n4637 , n4019 , n4291 );
and ( n4638 , n4035 , n4206 );
nor ( n4639 , n4637 , n4638 );
xnor ( n4640 , n4639 , n4297 );
xor ( n4641 , n4636 , n4640 );
xor ( n4642 , n4630 , n4641 );
and ( n4643 , n4525 , n4040 );
buf ( n4644 , n526 );
buf ( n4645 , n4644 );
and ( n4646 , n4645 , n4037 );
nor ( n4647 , n4643 , n4646 );
xnor ( n4648 , n4647 , n3989 );
buf ( n4649 , n542 );
buf ( n4650 , n4649 );
xor ( n4651 , n4650 , n4496 );
and ( n4652 , n3985 , n4651 );
xor ( n4653 , n4648 , n4652 );
buf ( n4654 , n462 );
buf ( n4655 , n4654 );
xor ( n4656 , n4653 , n4655 );
xor ( n4657 , n4642 , n4656 );
xor ( n4658 , n4626 , n4657 );
and ( n4659 , n4485 , n4507 );
and ( n4660 , n4507 , n4535 );
and ( n4661 , n4485 , n4535 );
or ( n4662 , n4659 , n4660 , n4661 );
xor ( n4663 , n4658 , n4662 );
and ( n4664 , n4536 , n4540 );
and ( n4665 , n4541 , n4544 );
or ( n4666 , n4664 , n4665 );
xor ( n4667 , n4663 , n4666 );
buf ( n4668 , n4667 );
buf ( n4669 , n1905 );
buf ( n4670 , n542 );
xor ( n4671 , n4669 , n4670 );
and ( n4672 , n4547 , n4548 );
and ( n4673 , n4548 , n4553 );
and ( n4674 , n4547 , n4553 );
or ( n4675 , n4672 , n4673 , n4674 );
xor ( n4676 , n4671 , n4675 );
buf ( n4677 , n4676 );
not ( n4678 , n454 );
and ( n4679 , n4678 , n4668 );
and ( n4680 , n4677 , n454 );
or ( n4681 , n4679 , n4680 );
buf ( n4682 , n4681 );
and ( n4683 , n4560 , n4564 );
xor ( n4684 , n4682 , n4683 );
buf ( n4685 , n4684 );
not ( n4686 , n4176 );
and ( n4687 , n4686 , n4607 );
and ( n4688 , n4685 , n4176 );
or ( n4689 , n4687 , n4688 );
and ( n4690 , n4580 , n4587 );
and ( n4691 , n4188 , n4596 );
and ( n4692 , n4262 , n4472 );
nor ( n4693 , n4691 , n4692 );
xnor ( n4694 , n4693 , n4586 );
xor ( n4695 , n4690 , n4694 );
and ( n4696 , n4577 , n4185 );
buf ( n4697 , n498 );
buf ( n4698 , n4697 );
and ( n4699 , n4698 , n3980 );
nor ( n4700 , n4696 , n4699 );
xnor ( n4701 , n4700 , n4182 );
and ( n4702 , n4369 , n4359 );
and ( n4703 , n4461 , n4268 );
nor ( n4704 , n4702 , n4703 );
xnor ( n4705 , n4704 , n4365 );
xor ( n4706 , n4701 , n4705 );
buf ( n4707 , n1187 );
buf ( n4708 , n4707 );
xor ( n4709 , n4708 , n4583 );
and ( n4710 , n3978 , n4709 );
xor ( n4711 , n4706 , n4710 );
xor ( n4712 , n4695 , n4711 );
and ( n4713 , n4588 , n4592 );
and ( n4714 , n4592 , n4600 );
and ( n4715 , n4588 , n4600 );
or ( n4716 , n4713 , n4714 , n4715 );
xor ( n4717 , n4712 , n4716 );
and ( n4718 , n4574 , n4601 );
and ( n4719 , n4602 , n4605 );
or ( n4720 , n4718 , n4719 );
xor ( n4721 , n4717 , n4720 );
buf ( n4722 , n4721 );
and ( n4723 , n4611 , n4625 );
and ( n4724 , n4625 , n4657 );
and ( n4725 , n4611 , n4657 );
or ( n4726 , n4723 , n4724 , n4725 );
and ( n4727 , n4630 , n4641 );
and ( n4728 , n4641 , n4656 );
and ( n4729 , n4630 , n4656 );
or ( n4730 , n4727 , n4728 , n4729 );
and ( n4731 , n4631 , n4635 );
and ( n4732 , n4635 , n4640 );
and ( n4733 , n4631 , n4640 );
or ( n4734 , n4731 , n4732 , n4733 );
and ( n4735 , n4648 , n4652 );
and ( n4736 , n4652 , n4655 );
and ( n4737 , n4648 , n4655 );
or ( n4738 , n4735 , n4736 , n4737 );
xor ( n4739 , n4734 , n4738 );
buf ( n4740 , n541 );
buf ( n4741 , n4740 );
xor ( n4742 , n4741 , n4650 );
not ( n4743 , n4651 );
and ( n4744 , n4742 , n4743 );
and ( n4745 , n3985 , n4744 );
and ( n4746 , n4053 , n4651 );
nor ( n4747 , n4745 , n4746 );
and ( n4748 , n4650 , n4496 );
not ( n4749 , n4748 );
and ( n4750 , n4741 , n4749 );
xnor ( n4751 , n4747 , n4750 );
xor ( n4752 , n4739 , n4751 );
xor ( n4753 , n4730 , n4752 );
and ( n4754 , n4615 , n4619 );
and ( n4755 , n4619 , n4624 );
and ( n4756 , n4615 , n4624 );
or ( n4757 , n4754 , n4755 , n4756 );
and ( n4758 , n4413 , n4016 );
and ( n4759 , n4525 , n3990 );
nor ( n4760 , n4758 , n4759 );
xnor ( n4761 , n4760 , n3997 );
and ( n4762 , n4035 , n4291 );
and ( n4763 , n4043 , n4206 );
nor ( n4764 , n4762 , n4763 );
xnor ( n4765 , n4764 , n4297 );
xor ( n4766 , n4761 , n4765 );
and ( n4767 , n4013 , n4499 );
and ( n4768 , n4019 , n4419 );
nor ( n4769 , n4767 , n4768 );
xnor ( n4770 , n4769 , n4505 );
xor ( n4771 , n4766 , n4770 );
xor ( n4772 , n4757 , n4771 );
not ( n4773 , n4652 );
and ( n4774 , n4773 , n4750 );
buf ( n4775 , n461 );
buf ( n4776 , n4775 );
xor ( n4777 , n4774 , n4776 );
and ( n4778 , n4645 , n4040 );
buf ( n4779 , n525 );
buf ( n4780 , n4779 );
and ( n4781 , n4780 , n4037 );
nor ( n4782 , n4778 , n4781 );
xnor ( n4783 , n4782 , n3989 );
xor ( n4784 , n4777 , n4783 );
and ( n4785 , n4216 , n4050 );
and ( n4786 , n4308 , n4004 );
nor ( n4787 , n4785 , n4786 );
xnor ( n4788 , n4787 , n4029 );
xor ( n4789 , n4784 , n4788 );
xor ( n4790 , n4772 , n4789 );
xor ( n4791 , n4753 , n4790 );
xor ( n4792 , n4726 , n4791 );
and ( n4793 , n4658 , n4662 );
and ( n4794 , n4663 , n4666 );
or ( n4795 , n4793 , n4794 );
xor ( n4796 , n4792 , n4795 );
buf ( n4797 , n4796 );
buf ( n4798 , n2063 );
buf ( n4799 , n541 );
xor ( n4800 , n4798 , n4799 );
and ( n4801 , n4669 , n4670 );
and ( n4802 , n4670 , n4675 );
and ( n4803 , n4669 , n4675 );
or ( n4804 , n4801 , n4802 , n4803 );
xor ( n4805 , n4800 , n4804 );
buf ( n4806 , n4805 );
not ( n4807 , n454 );
and ( n4808 , n4807 , n4797 );
and ( n4809 , n4806 , n454 );
or ( n4810 , n4808 , n4809 );
buf ( n4811 , n4810 );
and ( n4812 , n4682 , n4683 );
xor ( n4813 , n4811 , n4812 );
buf ( n4814 , n4813 );
not ( n4815 , n4176 );
and ( n4816 , n4815 , n4722 );
and ( n4817 , n4814 , n4176 );
or ( n4818 , n4816 , n4817 );
and ( n4819 , n4698 , n4185 );
buf ( n4820 , n497 );
buf ( n4821 , n4820 );
and ( n4822 , n4821 , n3980 );
nor ( n4823 , n4819 , n4822 );
xnor ( n4824 , n4823 , n4182 );
not ( n4825 , n4710 );
buf ( n4826 , n1309 );
buf ( n4827 , n4826 );
and ( n4828 , n4708 , n4583 );
not ( n4829 , n4828 );
and ( n4830 , n4827 , n4829 );
and ( n4831 , n4825 , n4830 );
xor ( n4832 , n4824 , n4831 );
and ( n4833 , n4701 , n4705 );
and ( n4834 , n4705 , n4710 );
and ( n4835 , n4701 , n4710 );
or ( n4836 , n4833 , n4834 , n4835 );
xor ( n4837 , n4832 , n4836 );
and ( n4838 , n4461 , n4359 );
and ( n4839 , n4577 , n4268 );
nor ( n4840 , n4838 , n4839 );
xnor ( n4841 , n4840 , n4365 );
and ( n4842 , n4262 , n4596 );
and ( n4843 , n4369 , n4472 );
nor ( n4844 , n4842 , n4843 );
xnor ( n4845 , n4844 , n4586 );
xor ( n4846 , n4841 , n4845 );
xor ( n4847 , n4827 , n4708 );
not ( n4848 , n4709 );
and ( n4849 , n4847 , n4848 );
and ( n4850 , n3978 , n4849 );
and ( n4851 , n4188 , n4709 );
nor ( n4852 , n4850 , n4851 );
xnor ( n4853 , n4852 , n4830 );
xor ( n4854 , n4846 , n4853 );
xor ( n4855 , n4837 , n4854 );
and ( n4856 , n4690 , n4694 );
and ( n4857 , n4694 , n4711 );
and ( n4858 , n4690 , n4711 );
or ( n4859 , n4856 , n4857 , n4858 );
xor ( n4860 , n4855 , n4859 );
and ( n4861 , n4712 , n4716 );
and ( n4862 , n4717 , n4720 );
or ( n4863 , n4861 , n4862 );
xor ( n4864 , n4860 , n4863 );
buf ( n4865 , n4864 );
and ( n4866 , n4757 , n4771 );
and ( n4867 , n4771 , n4789 );
and ( n4868 , n4757 , n4789 );
or ( n4869 , n4866 , n4867 , n4868 );
and ( n4870 , n4761 , n4765 );
and ( n4871 , n4765 , n4770 );
and ( n4872 , n4761 , n4770 );
or ( n4873 , n4870 , n4871 , n4872 );
and ( n4874 , n4777 , n4783 );
and ( n4875 , n4783 , n4788 );
and ( n4876 , n4777 , n4788 );
or ( n4877 , n4874 , n4875 , n4876 );
xor ( n4878 , n4873 , n4877 );
and ( n4879 , n4780 , n4040 );
buf ( n4880 , n524 );
buf ( n4881 , n4880 );
and ( n4882 , n4881 , n4037 );
nor ( n4883 , n4879 , n4882 );
xnor ( n4884 , n4883 , n3989 );
buf ( n4885 , n540 );
buf ( n4886 , n4885 );
xor ( n4887 , n4886 , n4741 );
and ( n4888 , n3985 , n4887 );
xor ( n4889 , n4884 , n4888 );
buf ( n4890 , n460 );
buf ( n4891 , n4890 );
xor ( n4892 , n4889 , n4891 );
xor ( n4893 , n4878 , n4892 );
xor ( n4894 , n4869 , n4893 );
and ( n4895 , n4734 , n4738 );
and ( n4896 , n4738 , n4751 );
and ( n4897 , n4734 , n4751 );
or ( n4898 , n4895 , n4896 , n4897 );
and ( n4899 , n4525 , n4016 );
and ( n4900 , n4645 , n3990 );
nor ( n4901 , n4899 , n4900 );
xnor ( n4902 , n4901 , n3997 );
and ( n4903 , n4019 , n4499 );
and ( n4904 , n4035 , n4419 );
nor ( n4905 , n4903 , n4904 );
xnor ( n4906 , n4905 , n4505 );
xor ( n4907 , n4902 , n4906 );
and ( n4908 , n4053 , n4744 );
and ( n4909 , n4013 , n4651 );
nor ( n4910 , n4908 , n4909 );
xnor ( n4911 , n4910 , n4750 );
xor ( n4912 , n4907 , n4911 );
xor ( n4913 , n4898 , n4912 );
and ( n4914 , n4774 , n4776 );
and ( n4915 , n4308 , n4050 );
and ( n4916 , n4413 , n4004 );
nor ( n4917 , n4915 , n4916 );
xnor ( n4918 , n4917 , n4029 );
xor ( n4919 , n4914 , n4918 );
and ( n4920 , n4043 , n4291 );
and ( n4921 , n4216 , n4206 );
nor ( n4922 , n4920 , n4921 );
xnor ( n4923 , n4922 , n4297 );
xor ( n4924 , n4919 , n4923 );
xor ( n4925 , n4913 , n4924 );
xor ( n4926 , n4894 , n4925 );
and ( n4927 , n4730 , n4752 );
and ( n4928 , n4752 , n4790 );
and ( n4929 , n4730 , n4790 );
or ( n4930 , n4927 , n4928 , n4929 );
xor ( n4931 , n4926 , n4930 );
and ( n4932 , n4726 , n4791 );
and ( n4933 , n4792 , n4795 );
or ( n4934 , n4932 , n4933 );
xor ( n4935 , n4931 , n4934 );
buf ( n4936 , n4935 );
buf ( n4937 , n2247 );
buf ( n4938 , n540 );
xor ( n4939 , n4937 , n4938 );
and ( n4940 , n4798 , n4799 );
and ( n4941 , n4799 , n4804 );
and ( n4942 , n4798 , n4804 );
or ( n4943 , n4940 , n4941 , n4942 );
xor ( n4944 , n4939 , n4943 );
buf ( n4945 , n4944 );
not ( n4946 , n454 );
and ( n4947 , n4946 , n4936 );
and ( n4948 , n4945 , n454 );
or ( n4949 , n4947 , n4948 );
buf ( n4950 , n4949 );
and ( n4951 , n4811 , n4812 );
xor ( n4952 , n4950 , n4951 );
buf ( n4953 , n4952 );
not ( n4954 , n4176 );
and ( n4955 , n4954 , n4865 );
and ( n4956 , n4953 , n4176 );
or ( n4957 , n4955 , n4956 );
and ( n4958 , n4832 , n4836 );
and ( n4959 , n4836 , n4854 );
and ( n4960 , n4832 , n4854 );
or ( n4961 , n4958 , n4959 , n4960 );
and ( n4962 , n4841 , n4845 );
and ( n4963 , n4845 , n4853 );
and ( n4964 , n4841 , n4853 );
or ( n4965 , n4962 , n4963 , n4964 );
and ( n4966 , n4821 , n4185 );
buf ( n4967 , n496 );
buf ( n4968 , n4967 );
and ( n4969 , n4968 , n3980 );
nor ( n4970 , n4966 , n4969 );
xnor ( n4971 , n4970 , n4182 );
and ( n4972 , n4188 , n4849 );
and ( n4973 , n4262 , n4709 );
nor ( n4974 , n4972 , n4973 );
xnor ( n4975 , n4974 , n4830 );
xor ( n4976 , n4971 , n4975 );
buf ( n4977 , n1409 );
buf ( n4978 , n4977 );
xor ( n4979 , n4978 , n4827 );
and ( n4980 , n3978 , n4979 );
xor ( n4981 , n4976 , n4980 );
xor ( n4982 , n4965 , n4981 );
and ( n4983 , n4824 , n4831 );
and ( n4984 , n4577 , n4359 );
and ( n4985 , n4698 , n4268 );
nor ( n4986 , n4984 , n4985 );
xnor ( n4987 , n4986 , n4365 );
xor ( n4988 , n4983 , n4987 );
and ( n4989 , n4369 , n4596 );
and ( n4990 , n4461 , n4472 );
nor ( n4991 , n4989 , n4990 );
xnor ( n4992 , n4991 , n4586 );
xor ( n4993 , n4988 , n4992 );
xor ( n4994 , n4982 , n4993 );
xor ( n4995 , n4961 , n4994 );
and ( n4996 , n4855 , n4859 );
and ( n4997 , n4860 , n4863 );
or ( n4998 , n4996 , n4997 );
xor ( n4999 , n4995 , n4998 );
buf ( n5000 , n4999 );
and ( n5001 , n4898 , n4912 );
and ( n5002 , n4912 , n4924 );
and ( n5003 , n4898 , n4924 );
or ( n5004 , n5001 , n5002 , n5003 );
and ( n5005 , n4884 , n4888 );
and ( n5006 , n4888 , n4891 );
and ( n5007 , n4884 , n4891 );
or ( n5008 , n5005 , n5006 , n5007 );
and ( n5009 , n4914 , n4918 );
and ( n5010 , n4918 , n4923 );
and ( n5011 , n4914 , n4923 );
or ( n5012 , n5009 , n5010 , n5011 );
xor ( n5013 , n5008 , n5012 );
not ( n5014 , n4888 );
buf ( n5015 , n539 );
buf ( n5016 , n5015 );
and ( n5017 , n4886 , n4741 );
not ( n5018 , n5017 );
and ( n5019 , n5016 , n5018 );
and ( n5020 , n5014 , n5019 );
buf ( n5021 , n459 );
buf ( n5022 , n5021 );
xor ( n5023 , n5020 , n5022 );
and ( n5024 , n4881 , n4040 );
buf ( n5025 , n523 );
buf ( n5026 , n5025 );
and ( n5027 , n5026 , n4037 );
nor ( n5028 , n5024 , n5027 );
xnor ( n5029 , n5028 , n3989 );
xor ( n5030 , n5023 , n5029 );
xor ( n5031 , n5016 , n4886 );
not ( n5032 , n4887 );
and ( n5033 , n5031 , n5032 );
and ( n5034 , n3985 , n5033 );
and ( n5035 , n4053 , n4887 );
nor ( n5036 , n5034 , n5035 );
xnor ( n5037 , n5036 , n5019 );
xor ( n5038 , n5030 , n5037 );
xor ( n5039 , n5013 , n5038 );
xor ( n5040 , n5004 , n5039 );
and ( n5041 , n4873 , n4877 );
and ( n5042 , n4877 , n4892 );
and ( n5043 , n4873 , n4892 );
or ( n5044 , n5041 , n5042 , n5043 );
and ( n5045 , n4645 , n4016 );
and ( n5046 , n4780 , n3990 );
nor ( n5047 , n5045 , n5046 );
xnor ( n5048 , n5047 , n3997 );
and ( n5049 , n4413 , n4050 );
and ( n5050 , n4525 , n4004 );
nor ( n5051 , n5049 , n5050 );
xnor ( n5052 , n5051 , n4029 );
xor ( n5053 , n5048 , n5052 );
and ( n5054 , n4216 , n4291 );
and ( n5055 , n4308 , n4206 );
nor ( n5056 , n5054 , n5055 );
xnor ( n5057 , n5056 , n4297 );
xor ( n5058 , n5053 , n5057 );
xor ( n5059 , n5044 , n5058 );
and ( n5060 , n4902 , n4906 );
and ( n5061 , n4906 , n4911 );
and ( n5062 , n4902 , n4911 );
or ( n5063 , n5060 , n5061 , n5062 );
and ( n5064 , n4035 , n4499 );
and ( n5065 , n4043 , n4419 );
nor ( n5066 , n5064 , n5065 );
xnor ( n5067 , n5066 , n4505 );
xor ( n5068 , n5063 , n5067 );
and ( n5069 , n4013 , n4744 );
and ( n5070 , n4019 , n4651 );
nor ( n5071 , n5069 , n5070 );
xnor ( n5072 , n5071 , n4750 );
xor ( n5073 , n5068 , n5072 );
xor ( n5074 , n5059 , n5073 );
xor ( n5075 , n5040 , n5074 );
and ( n5076 , n4869 , n4893 );
and ( n5077 , n4893 , n4925 );
and ( n5078 , n4869 , n4925 );
or ( n5079 , n5076 , n5077 , n5078 );
xor ( n5080 , n5075 , n5079 );
and ( n5081 , n4926 , n4930 );
and ( n5082 , n4931 , n4934 );
or ( n5083 , n5081 , n5082 );
xor ( n5084 , n5080 , n5083 );
buf ( n5085 , n5084 );
buf ( n5086 , n2409 );
buf ( n5087 , n539 );
xor ( n5088 , n5086 , n5087 );
and ( n5089 , n4937 , n4938 );
and ( n5090 , n4938 , n4943 );
and ( n5091 , n4937 , n4943 );
or ( n5092 , n5089 , n5090 , n5091 );
xor ( n5093 , n5088 , n5092 );
buf ( n5094 , n5093 );
not ( n5095 , n454 );
and ( n5096 , n5095 , n5085 );
and ( n5097 , n5094 , n454 );
or ( n5098 , n5096 , n5097 );
buf ( n5099 , n5098 );
and ( n5100 , n4950 , n4951 );
xor ( n5101 , n5099 , n5100 );
buf ( n5102 , n5101 );
not ( n5103 , n4176 );
and ( n5104 , n5103 , n5000 );
and ( n5105 , n5102 , n4176 );
or ( n5106 , n5104 , n5105 );
and ( n5107 , n4983 , n4987 );
and ( n5108 , n4987 , n4992 );
and ( n5109 , n4983 , n4992 );
or ( n5110 , n5107 , n5108 , n5109 );
and ( n5111 , n4968 , n4185 );
buf ( n5112 , n495 );
buf ( n5113 , n5112 );
and ( n5114 , n5113 , n3980 );
nor ( n5115 , n5111 , n5114 );
xnor ( n5116 , n5115 , n4182 );
and ( n5117 , n4262 , n4849 );
and ( n5118 , n4369 , n4709 );
nor ( n5119 , n5117 , n5118 );
xnor ( n5120 , n5119 , n4830 );
xor ( n5121 , n5116 , n5120 );
buf ( n5122 , n1573 );
buf ( n5123 , n5122 );
xor ( n5124 , n5123 , n4978 );
not ( n5125 , n4979 );
and ( n5126 , n5124 , n5125 );
and ( n5127 , n3978 , n5126 );
and ( n5128 , n4188 , n4979 );
nor ( n5129 , n5127 , n5128 );
and ( n5130 , n4978 , n4827 );
not ( n5131 , n5130 );
and ( n5132 , n5123 , n5131 );
xnor ( n5133 , n5129 , n5132 );
xor ( n5134 , n5121 , n5133 );
xor ( n5135 , n5110 , n5134 );
and ( n5136 , n4698 , n4359 );
and ( n5137 , n4821 , n4268 );
nor ( n5138 , n5136 , n5137 );
xnor ( n5139 , n5138 , n4365 );
not ( n5140 , n4980 );
and ( n5141 , n5140 , n5132 );
xor ( n5142 , n5139 , n5141 );
and ( n5143 , n4971 , n4975 );
and ( n5144 , n4975 , n4980 );
and ( n5145 , n4971 , n4980 );
or ( n5146 , n5143 , n5144 , n5145 );
xor ( n5147 , n5142 , n5146 );
and ( n5148 , n4461 , n4596 );
and ( n5149 , n4577 , n4472 );
nor ( n5150 , n5148 , n5149 );
xnor ( n5151 , n5150 , n4586 );
xor ( n5152 , n5147 , n5151 );
xor ( n5153 , n5135 , n5152 );
and ( n5154 , n4965 , n4981 );
and ( n5155 , n4981 , n4993 );
and ( n5156 , n4965 , n4993 );
or ( n5157 , n5154 , n5155 , n5156 );
xor ( n5158 , n5153 , n5157 );
and ( n5159 , n4961 , n4994 );
and ( n5160 , n4995 , n4998 );
or ( n5161 , n5159 , n5160 );
xor ( n5162 , n5158 , n5161 );
buf ( n5163 , n5162 );
and ( n5164 , n5044 , n5058 );
and ( n5165 , n5058 , n5073 );
and ( n5166 , n5044 , n5073 );
or ( n5167 , n5164 , n5165 , n5166 );
and ( n5168 , n5023 , n5029 );
and ( n5169 , n5029 , n5037 );
and ( n5170 , n5023 , n5037 );
or ( n5171 , n5168 , n5169 , n5170 );
and ( n5172 , n4525 , n4050 );
and ( n5173 , n4645 , n4004 );
nor ( n5174 , n5172 , n5173 );
xnor ( n5175 , n5174 , n4029 );
and ( n5176 , n4308 , n4291 );
and ( n5177 , n4413 , n4206 );
nor ( n5178 , n5176 , n5177 );
xnor ( n5179 , n5178 , n4297 );
xor ( n5180 , n5175 , n5179 );
and ( n5181 , n4053 , n5033 );
and ( n5182 , n4013 , n4887 );
nor ( n5183 , n5181 , n5182 );
xnor ( n5184 , n5183 , n5019 );
xor ( n5185 , n5180 , n5184 );
xor ( n5186 , n5171 , n5185 );
and ( n5187 , n5020 , n5022 );
and ( n5188 , n4780 , n4016 );
and ( n5189 , n4881 , n3990 );
nor ( n5190 , n5188 , n5189 );
xnor ( n5191 , n5190 , n3997 );
xor ( n5192 , n5187 , n5191 );
and ( n5193 , n4043 , n4499 );
and ( n5194 , n4216 , n4419 );
nor ( n5195 , n5193 , n5194 );
xnor ( n5196 , n5195 , n4505 );
xor ( n5197 , n5192 , n5196 );
xor ( n5198 , n5186 , n5197 );
xor ( n5199 , n5167 , n5198 );
and ( n5200 , n5063 , n5067 );
and ( n5201 , n5067 , n5072 );
and ( n5202 , n5063 , n5072 );
or ( n5203 , n5200 , n5201 , n5202 );
and ( n5204 , n5008 , n5012 );
and ( n5205 , n5012 , n5038 );
and ( n5206 , n5008 , n5038 );
or ( n5207 , n5204 , n5205 , n5206 );
xor ( n5208 , n5203 , n5207 );
and ( n5209 , n5048 , n5052 );
and ( n5210 , n5052 , n5057 );
and ( n5211 , n5048 , n5057 );
or ( n5212 , n5209 , n5210 , n5211 );
and ( n5213 , n4019 , n4744 );
and ( n5214 , n4035 , n4651 );
nor ( n5215 , n5213 , n5214 );
xnor ( n5216 , n5215 , n4750 );
xor ( n5217 , n5212 , n5216 );
and ( n5218 , n5026 , n4040 );
buf ( n5219 , n522 );
buf ( n5220 , n5219 );
and ( n5221 , n5220 , n4037 );
nor ( n5222 , n5218 , n5221 );
xnor ( n5223 , n5222 , n3989 );
buf ( n5224 , n538 );
buf ( n5225 , n5224 );
xor ( n5226 , n5225 , n5016 );
and ( n5227 , n3985 , n5226 );
xor ( n5228 , n5223 , n5227 );
buf ( n5229 , n458 );
buf ( n5230 , n5229 );
xor ( n5231 , n5228 , n5230 );
xor ( n5232 , n5217 , n5231 );
xor ( n5233 , n5208 , n5232 );
xor ( n5234 , n5199 , n5233 );
and ( n5235 , n5004 , n5039 );
and ( n5236 , n5039 , n5074 );
and ( n5237 , n5004 , n5074 );
or ( n5238 , n5235 , n5236 , n5237 );
xor ( n5239 , n5234 , n5238 );
and ( n5240 , n5075 , n5079 );
and ( n5241 , n5080 , n5083 );
or ( n5242 , n5240 , n5241 );
xor ( n5243 , n5239 , n5242 );
buf ( n5244 , n5243 );
buf ( n5245 , n2573 );
buf ( n5246 , n538 );
xor ( n5247 , n5245 , n5246 );
and ( n5248 , n5086 , n5087 );
and ( n5249 , n5087 , n5092 );
and ( n5250 , n5086 , n5092 );
or ( n5251 , n5248 , n5249 , n5250 );
xor ( n5252 , n5247 , n5251 );
buf ( n5253 , n5252 );
not ( n5254 , n454 );
and ( n5255 , n5254 , n5244 );
and ( n5256 , n5253 , n454 );
or ( n5257 , n5255 , n5256 );
buf ( n5258 , n5257 );
and ( n5259 , n5099 , n5100 );
xor ( n5260 , n5258 , n5259 );
buf ( n5261 , n5260 );
not ( n5262 , n4176 );
and ( n5263 , n5262 , n5163 );
and ( n5264 , n5261 , n4176 );
or ( n5265 , n5263 , n5264 );
and ( n5266 , n5142 , n5146 );
and ( n5267 , n5146 , n5151 );
and ( n5268 , n5142 , n5151 );
or ( n5269 , n5266 , n5267 , n5268 );
and ( n5270 , n5113 , n4185 );
buf ( n5271 , n494 );
buf ( n5272 , n5271 );
and ( n5273 , n5272 , n3980 );
nor ( n5274 , n5270 , n5273 );
xnor ( n5275 , n5274 , n4182 );
and ( n5276 , n4577 , n4596 );
and ( n5277 , n4698 , n4472 );
nor ( n5278 , n5276 , n5277 );
xnor ( n5279 , n5278 , n4586 );
xor ( n5280 , n5275 , n5279 );
and ( n5281 , n4188 , n5126 );
and ( n5282 , n4262 , n4979 );
nor ( n5283 , n5281 , n5282 );
xnor ( n5284 , n5283 , n5132 );
xor ( n5285 , n5280 , n5284 );
xor ( n5286 , n5269 , n5285 );
and ( n5287 , n5116 , n5120 );
and ( n5288 , n5120 , n5133 );
and ( n5289 , n5116 , n5133 );
or ( n5290 , n5287 , n5288 , n5289 );
and ( n5291 , n5139 , n5141 );
xor ( n5292 , n5290 , n5291 );
and ( n5293 , n4821 , n4359 );
and ( n5294 , n4968 , n4268 );
nor ( n5295 , n5293 , n5294 );
xnor ( n5296 , n5295 , n4365 );
and ( n5297 , n4369 , n4849 );
and ( n5298 , n4461 , n4709 );
nor ( n5299 , n5297 , n5298 );
xnor ( n5300 , n5299 , n4830 );
xor ( n5301 , n5296 , n5300 );
buf ( n5302 , n1675 );
buf ( n5303 , n5302 );
xor ( n5304 , n5303 , n5123 );
and ( n5305 , n3978 , n5304 );
xor ( n5306 , n5301 , n5305 );
xor ( n5307 , n5292 , n5306 );
xor ( n5308 , n5286 , n5307 );
and ( n5309 , n5110 , n5134 );
and ( n5310 , n5134 , n5152 );
and ( n5311 , n5110 , n5152 );
or ( n5312 , n5309 , n5310 , n5311 );
xor ( n5313 , n5308 , n5312 );
and ( n5314 , n5153 , n5157 );
and ( n5315 , n5158 , n5161 );
or ( n5316 , n5314 , n5315 );
xor ( n5317 , n5313 , n5316 );
buf ( n5318 , n5317 );
and ( n5319 , n5203 , n5207 );
and ( n5320 , n5207 , n5232 );
and ( n5321 , n5203 , n5232 );
or ( n5322 , n5319 , n5320 , n5321 );
and ( n5323 , n4881 , n4016 );
and ( n5324 , n5026 , n3990 );
nor ( n5325 , n5323 , n5324 );
xnor ( n5326 , n5325 , n3997 );
and ( n5327 , n4216 , n4499 );
and ( n5328 , n4308 , n4419 );
nor ( n5329 , n5327 , n5328 );
xnor ( n5330 , n5329 , n4505 );
xor ( n5331 , n5326 , n5330 );
and ( n5332 , n4035 , n4744 );
and ( n5333 , n4043 , n4651 );
nor ( n5334 , n5332 , n5333 );
xnor ( n5335 , n5334 , n4750 );
xor ( n5336 , n5331 , n5335 );
and ( n5337 , n4645 , n4050 );
and ( n5338 , n4780 , n4004 );
nor ( n5339 , n5337 , n5338 );
xnor ( n5340 , n5339 , n4029 );
and ( n5341 , n4013 , n5033 );
and ( n5342 , n4019 , n4887 );
nor ( n5343 , n5341 , n5342 );
xnor ( n5344 , n5343 , n5019 );
xor ( n5345 , n5340 , n5344 );
buf ( n5346 , n537 );
buf ( n5347 , n5346 );
xor ( n5348 , n5347 , n5225 );
not ( n5349 , n5226 );
and ( n5350 , n5348 , n5349 );
and ( n5351 , n3985 , n5350 );
and ( n5352 , n4053 , n5226 );
nor ( n5353 , n5351 , n5352 );
and ( n5354 , n5225 , n5016 );
not ( n5355 , n5354 );
and ( n5356 , n5347 , n5355 );
xnor ( n5357 , n5353 , n5356 );
xor ( n5358 , n5345 , n5357 );
xor ( n5359 , n5336 , n5358 );
not ( n5360 , n5227 );
and ( n5361 , n5360 , n5356 );
buf ( n5362 , n457 );
buf ( n5363 , n5362 );
xor ( n5364 , n5361 , n5363 );
and ( n5365 , n5220 , n4040 );
buf ( n5366 , n521 );
buf ( n5367 , n5366 );
and ( n5368 , n5367 , n4037 );
nor ( n5369 , n5365 , n5368 );
xnor ( n5370 , n5369 , n3989 );
xor ( n5371 , n5364 , n5370 );
and ( n5372 , n4413 , n4291 );
and ( n5373 , n4525 , n4206 );
nor ( n5374 , n5372 , n5373 );
xnor ( n5375 , n5374 , n4297 );
xor ( n5376 , n5371 , n5375 );
xor ( n5377 , n5359 , n5376 );
xor ( n5378 , n5322 , n5377 );
and ( n5379 , n5212 , n5216 );
and ( n5380 , n5216 , n5231 );
and ( n5381 , n5212 , n5231 );
or ( n5382 , n5379 , n5380 , n5381 );
and ( n5383 , n5171 , n5185 );
and ( n5384 , n5185 , n5197 );
and ( n5385 , n5171 , n5197 );
or ( n5386 , n5383 , n5384 , n5385 );
xor ( n5387 , n5382 , n5386 );
and ( n5388 , n5175 , n5179 );
and ( n5389 , n5179 , n5184 );
and ( n5390 , n5175 , n5184 );
or ( n5391 , n5388 , n5389 , n5390 );
and ( n5392 , n5187 , n5191 );
and ( n5393 , n5191 , n5196 );
and ( n5394 , n5187 , n5196 );
or ( n5395 , n5392 , n5393 , n5394 );
xor ( n5396 , n5391 , n5395 );
and ( n5397 , n5223 , n5227 );
and ( n5398 , n5227 , n5230 );
and ( n5399 , n5223 , n5230 );
or ( n5400 , n5397 , n5398 , n5399 );
xor ( n5401 , n5396 , n5400 );
xor ( n5402 , n5387 , n5401 );
xor ( n5403 , n5378 , n5402 );
and ( n5404 , n5167 , n5198 );
and ( n5405 , n5198 , n5233 );
and ( n5406 , n5167 , n5233 );
or ( n5407 , n5404 , n5405 , n5406 );
xor ( n5408 , n5403 , n5407 );
and ( n5409 , n5234 , n5238 );
and ( n5410 , n5239 , n5242 );
or ( n5411 , n5409 , n5410 );
xor ( n5412 , n5408 , n5411 );
buf ( n5413 , n5412 );
buf ( n5414 , n2737 );
buf ( n5415 , n537 );
xor ( n5416 , n5414 , n5415 );
and ( n5417 , n5245 , n5246 );
and ( n5418 , n5246 , n5251 );
and ( n5419 , n5245 , n5251 );
or ( n5420 , n5417 , n5418 , n5419 );
xor ( n5421 , n5416 , n5420 );
buf ( n5422 , n5421 );
not ( n5423 , n454 );
and ( n5424 , n5423 , n5413 );
and ( n5425 , n5422 , n454 );
or ( n5426 , n5424 , n5425 );
buf ( n5427 , n5426 );
and ( n5428 , n5258 , n5259 );
xor ( n5429 , n5427 , n5428 );
buf ( n5430 , n5429 );
not ( n5431 , n4176 );
and ( n5432 , n5431 , n5318 );
and ( n5433 , n5430 , n4176 );
or ( n5434 , n5432 , n5433 );
and ( n5435 , n5290 , n5291 );
and ( n5436 , n5291 , n5306 );
and ( n5437 , n5290 , n5306 );
or ( n5438 , n5435 , n5436 , n5437 );
and ( n5439 , n4968 , n4359 );
and ( n5440 , n5113 , n4268 );
nor ( n5441 , n5439 , n5440 );
xnor ( n5442 , n5441 , n4365 );
not ( n5443 , n5305 );
buf ( n5444 , n1870 );
buf ( n5445 , n5444 );
and ( n5446 , n5303 , n5123 );
not ( n5447 , n5446 );
and ( n5448 , n5445 , n5447 );
and ( n5449 , n5443 , n5448 );
xor ( n5450 , n5442 , n5449 );
and ( n5451 , n4698 , n4596 );
and ( n5452 , n4821 , n4472 );
nor ( n5453 , n5451 , n5452 );
xnor ( n5454 , n5453 , n4586 );
xor ( n5455 , n5450 , n5454 );
xor ( n5456 , n5445 , n5303 );
not ( n5457 , n5304 );
and ( n5458 , n5456 , n5457 );
and ( n5459 , n3978 , n5458 );
and ( n5460 , n4188 , n5304 );
nor ( n5461 , n5459 , n5460 );
xnor ( n5462 , n5461 , n5448 );
xor ( n5463 , n5455 , n5462 );
xor ( n5464 , n5438 , n5463 );
and ( n5465 , n5275 , n5279 );
and ( n5466 , n5279 , n5284 );
and ( n5467 , n5275 , n5284 );
or ( n5468 , n5465 , n5466 , n5467 );
and ( n5469 , n5296 , n5300 );
and ( n5470 , n5300 , n5305 );
and ( n5471 , n5296 , n5305 );
or ( n5472 , n5469 , n5470 , n5471 );
xor ( n5473 , n5468 , n5472 );
and ( n5474 , n5272 , n4185 );
buf ( n5475 , n493 );
buf ( n5476 , n5475 );
and ( n5477 , n5476 , n3980 );
nor ( n5478 , n5474 , n5477 );
xnor ( n5479 , n5478 , n4182 );
and ( n5480 , n4461 , n4849 );
and ( n5481 , n4577 , n4709 );
nor ( n5482 , n5480 , n5481 );
xnor ( n5483 , n5482 , n4830 );
xor ( n5484 , n5479 , n5483 );
and ( n5485 , n4262 , n5126 );
and ( n5486 , n4369 , n4979 );
nor ( n5487 , n5485 , n5486 );
xnor ( n5488 , n5487 , n5132 );
xor ( n5489 , n5484 , n5488 );
xor ( n5490 , n5473 , n5489 );
xor ( n5491 , n5464 , n5490 );
and ( n5492 , n5269 , n5285 );
and ( n5493 , n5285 , n5307 );
and ( n5494 , n5269 , n5307 );
or ( n5495 , n5492 , n5493 , n5494 );
xor ( n5496 , n5491 , n5495 );
and ( n5497 , n5308 , n5312 );
and ( n5498 , n5313 , n5316 );
or ( n5499 , n5497 , n5498 );
xor ( n5500 , n5496 , n5499 );
buf ( n5501 , n5500 );
and ( n5502 , n5382 , n5386 );
and ( n5503 , n5386 , n5401 );
and ( n5504 , n5382 , n5401 );
or ( n5505 , n5502 , n5503 , n5504 );
and ( n5506 , n5026 , n4016 );
and ( n5507 , n5220 , n3990 );
nor ( n5508 , n5506 , n5507 );
xnor ( n5509 , n5508 , n3997 );
and ( n5510 , n4525 , n4291 );
and ( n5511 , n4645 , n4206 );
nor ( n5512 , n5510 , n5511 );
xnor ( n5513 , n5512 , n4297 );
xor ( n5514 , n5509 , n5513 );
and ( n5515 , n4053 , n5350 );
and ( n5516 , n4013 , n5226 );
nor ( n5517 , n5515 , n5516 );
xnor ( n5518 , n5517 , n5356 );
xor ( n5519 , n5514 , n5518 );
and ( n5520 , n5361 , n5363 );
and ( n5521 , n4780 , n4050 );
and ( n5522 , n4881 , n4004 );
nor ( n5523 , n5521 , n5522 );
xnor ( n5524 , n5523 , n4029 );
xor ( n5525 , n5520 , n5524 );
and ( n5526 , n4308 , n4499 );
and ( n5527 , n4413 , n4419 );
nor ( n5528 , n5526 , n5527 );
xnor ( n5529 , n5528 , n4505 );
xor ( n5530 , n5525 , n5529 );
xor ( n5531 , n5519 , n5530 );
and ( n5532 , n5367 , n4040 );
not ( n5533 , n5532 );
xnor ( n5534 , n5533 , n3989 );
and ( n5535 , n3985 , n5347 );
xor ( n5536 , n5534 , n5535 );
and ( n5537 , n4043 , n4744 );
and ( n5538 , n4216 , n4651 );
nor ( n5539 , n5537 , n5538 );
xnor ( n5540 , n5539 , n4750 );
xor ( n5541 , n5536 , n5540 );
and ( n5542 , n4019 , n5033 );
and ( n5543 , n4035 , n4887 );
nor ( n5544 , n5542 , n5543 );
xnor ( n5545 , n5544 , n5019 );
xor ( n5546 , n5541 , n5545 );
xor ( n5547 , n5531 , n5546 );
xor ( n5548 , n5505 , n5547 );
and ( n5549 , n5391 , n5395 );
and ( n5550 , n5395 , n5400 );
and ( n5551 , n5391 , n5400 );
or ( n5552 , n5549 , n5550 , n5551 );
and ( n5553 , n5336 , n5358 );
and ( n5554 , n5358 , n5376 );
and ( n5555 , n5336 , n5376 );
or ( n5556 , n5553 , n5554 , n5555 );
xor ( n5557 , n5552 , n5556 );
and ( n5558 , n5326 , n5330 );
and ( n5559 , n5330 , n5335 );
and ( n5560 , n5326 , n5335 );
or ( n5561 , n5558 , n5559 , n5560 );
and ( n5562 , n5340 , n5344 );
and ( n5563 , n5344 , n5357 );
and ( n5564 , n5340 , n5357 );
or ( n5565 , n5562 , n5563 , n5564 );
xor ( n5566 , n5561 , n5565 );
and ( n5567 , n5364 , n5370 );
and ( n5568 , n5370 , n5375 );
and ( n5569 , n5364 , n5375 );
or ( n5570 , n5567 , n5568 , n5569 );
xor ( n5571 , n5566 , n5570 );
xor ( n5572 , n5557 , n5571 );
xor ( n5573 , n5548 , n5572 );
and ( n5574 , n5322 , n5377 );
and ( n5575 , n5377 , n5402 );
and ( n5576 , n5322 , n5402 );
or ( n5577 , n5574 , n5575 , n5576 );
xor ( n5578 , n5573 , n5577 );
and ( n5579 , n5403 , n5407 );
and ( n5580 , n5408 , n5411 );
or ( n5581 , n5579 , n5580 );
xor ( n5582 , n5578 , n5581 );
buf ( n5583 , n5582 );
buf ( n5584 , n2894 );
and ( n5585 , n5414 , n5415 );
and ( n5586 , n5415 , n5420 );
and ( n5587 , n5414 , n5420 );
or ( n5588 , n5585 , n5586 , n5587 );
xor ( n5589 , n5584 , n5588 );
buf ( n5590 , n5589 );
not ( n5591 , n454 );
and ( n5592 , n5591 , n5583 );
and ( n5593 , n5590 , n454 );
or ( n5594 , n5592 , n5593 );
buf ( n5595 , n5594 );
and ( n5596 , n5427 , n5428 );
xor ( n5597 , n5595 , n5596 );
buf ( n5598 , n5597 );
not ( n5599 , n4176 );
and ( n5600 , n5599 , n5501 );
and ( n5601 , n5598 , n4176 );
or ( n5602 , n5600 , n5601 );
and ( n5603 , n5438 , n5463 );
and ( n5604 , n5463 , n5490 );
and ( n5605 , n5438 , n5490 );
or ( n5606 , n5603 , n5604 , n5605 );
and ( n5607 , n5468 , n5472 );
and ( n5608 , n5472 , n5489 );
and ( n5609 , n5468 , n5489 );
or ( n5610 , n5607 , n5608 , n5609 );
and ( n5611 , n5479 , n5483 );
and ( n5612 , n5483 , n5488 );
and ( n5613 , n5479 , n5488 );
or ( n5614 , n5611 , n5612 , n5613 );
and ( n5615 , n5442 , n5449 );
xor ( n5616 , n5614 , n5615 );
and ( n5617 , n4821 , n4596 );
and ( n5618 , n4968 , n4472 );
nor ( n5619 , n5617 , n5618 );
xnor ( n5620 , n5619 , n4586 );
xor ( n5621 , n5616 , n5620 );
xor ( n5622 , n5610 , n5621 );
and ( n5623 , n5450 , n5454 );
and ( n5624 , n5454 , n5462 );
and ( n5625 , n5450 , n5462 );
or ( n5626 , n5623 , n5624 , n5625 );
and ( n5627 , n5476 , n4185 );
buf ( n5628 , n492 );
buf ( n5629 , n5628 );
and ( n5630 , n5629 , n3980 );
nor ( n5631 , n5627 , n5630 );
xnor ( n5632 , n5631 , n4182 );
and ( n5633 , n4369 , n5126 );
and ( n5634 , n4461 , n4979 );
nor ( n5635 , n5633 , n5634 );
xnor ( n5636 , n5635 , n5132 );
xor ( n5637 , n5632 , n5636 );
and ( n5638 , n4188 , n5458 );
and ( n5639 , n4262 , n5304 );
nor ( n5640 , n5638 , n5639 );
xnor ( n5641 , n5640 , n5448 );
xor ( n5642 , n5637 , n5641 );
xor ( n5643 , n5626 , n5642 );
and ( n5644 , n5113 , n4359 );
and ( n5645 , n5272 , n4268 );
nor ( n5646 , n5644 , n5645 );
xnor ( n5647 , n5646 , n4365 );
and ( n5648 , n4577 , n4849 );
and ( n5649 , n4698 , n4709 );
nor ( n5650 , n5648 , n5649 );
xnor ( n5651 , n5650 , n4830 );
xor ( n5652 , n5647 , n5651 );
buf ( n5653 , n1991 );
buf ( n5654 , n5653 );
xor ( n5655 , n5654 , n5445 );
and ( n5656 , n3978 , n5655 );
xor ( n5657 , n5652 , n5656 );
xor ( n5658 , n5643 , n5657 );
xor ( n5659 , n5622 , n5658 );
xor ( n5660 , n5606 , n5659 );
and ( n5661 , n5491 , n5495 );
and ( n5662 , n5496 , n5499 );
or ( n5663 , n5661 , n5662 );
xor ( n5664 , n5660 , n5663 );
buf ( n5665 , n5664 );
and ( n5666 , n5573 , n5577 );
and ( n5667 , n5552 , n5556 );
and ( n5668 , n5556 , n5571 );
and ( n5669 , n5552 , n5571 );
or ( n5670 , n5667 , n5668 , n5669 );
and ( n5671 , n5561 , n5565 );
and ( n5672 , n5565 , n5570 );
and ( n5673 , n5561 , n5570 );
or ( n5674 , n5671 , n5672 , n5673 );
and ( n5675 , n5536 , n5540 );
and ( n5676 , n5540 , n5545 );
and ( n5677 , n5536 , n5545 );
or ( n5678 , n5675 , n5676 , n5677 );
xor ( n5679 , n5674 , n5678 );
and ( n5680 , n5220 , n4016 );
and ( n5681 , n5367 , n3990 );
nor ( n5682 , n5680 , n5681 );
xnor ( n5683 , n5682 , n3997 );
and ( n5684 , n4881 , n4050 );
and ( n5685 , n5026 , n4004 );
nor ( n5686 , n5684 , n5685 );
xnor ( n5687 , n5686 , n4029 );
xor ( n5688 , n5683 , n5687 );
and ( n5689 , n4216 , n4744 );
and ( n5690 , n4308 , n4651 );
nor ( n5691 , n5689 , n5690 );
xnor ( n5692 , n5691 , n4750 );
xor ( n5693 , n5688 , n5692 );
xor ( n5694 , n5679 , n5693 );
xor ( n5695 , n5670 , n5694 );
and ( n5696 , n5519 , n5530 );
and ( n5697 , n5530 , n5546 );
and ( n5698 , n5519 , n5546 );
or ( n5699 , n5696 , n5697 , n5698 );
and ( n5700 , n5520 , n5524 );
and ( n5701 , n5524 , n5529 );
and ( n5702 , n5520 , n5529 );
or ( n5703 , n5700 , n5701 , n5702 );
and ( n5704 , n5534 , n5535 );
xor ( n5705 , n5703 , n5704 );
and ( n5706 , n4035 , n5033 );
and ( n5707 , n4043 , n4887 );
nor ( n5708 , n5706 , n5707 );
xnor ( n5709 , n5708 , n5019 );
xor ( n5710 , n5705 , n5709 );
xor ( n5711 , n5699 , n5710 );
not ( n5712 , n3989 );
and ( n5713 , n4413 , n4499 );
and ( n5714 , n4525 , n4419 );
nor ( n5715 , n5713 , n5714 );
xnor ( n5716 , n5715 , n4505 );
xnor ( n5717 , n5712 , n5716 );
and ( n5718 , n5509 , n5513 );
and ( n5719 , n5513 , n5518 );
and ( n5720 , n5509 , n5518 );
or ( n5721 , n5718 , n5719 , n5720 );
xor ( n5722 , n5717 , n5721 );
and ( n5723 , n4645 , n4291 );
and ( n5724 , n4780 , n4206 );
nor ( n5725 , n5723 , n5724 );
xnor ( n5726 , n5725 , n4297 );
and ( n5727 , n4013 , n5350 );
and ( n5728 , n4019 , n5226 );
nor ( n5729 , n5727 , n5728 );
xnor ( n5730 , n5729 , n5356 );
xor ( n5731 , n5726 , n5730 );
and ( n5732 , n4053 , n5347 );
xor ( n5733 , n5731 , n5732 );
xor ( n5734 , n5722 , n5733 );
xor ( n5735 , n5711 , n5734 );
xor ( n5736 , n5695 , n5735 );
and ( n5737 , n5505 , n5547 );
and ( n5738 , n5547 , n5572 );
and ( n5739 , n5505 , n5572 );
or ( n5740 , n5737 , n5738 , n5739 );
xor ( n5741 , n5736 , n5740 );
xor ( n5742 , n5666 , n5741 );
and ( n5743 , n5578 , n5581 );
xor ( n5744 , n5742 , n5743 );
buf ( n5745 , n5744 );
buf ( n5746 , n3040 );
and ( n5747 , n5584 , n5588 );
xor ( n5748 , n5746 , n5747 );
buf ( n5749 , n5748 );
not ( n5750 , n454 );
and ( n5751 , n5750 , n5745 );
and ( n5752 , n5749 , n454 );
or ( n5753 , n5751 , n5752 );
buf ( n5754 , n5753 );
and ( n5755 , n5595 , n5596 );
xor ( n5756 , n5754 , n5755 );
buf ( n5757 , n5756 );
not ( n5758 , n4176 );
and ( n5759 , n5758 , n5665 );
and ( n5760 , n5757 , n4176 );
or ( n5761 , n5759 , n5760 );
and ( n5762 , n5626 , n5642 );
and ( n5763 , n5642 , n5657 );
and ( n5764 , n5626 , n5657 );
or ( n5765 , n5762 , n5763 , n5764 );
and ( n5766 , n5629 , n4185 );
buf ( n5767 , n491 );
buf ( n5768 , n5767 );
and ( n5769 , n5768 , n3980 );
nor ( n5770 , n5766 , n5769 );
xnor ( n5771 , n5770 , n4182 );
not ( n5772 , n5656 );
buf ( n5773 , n2206 );
buf ( n5774 , n5773 );
and ( n5775 , n5654 , n5445 );
not ( n5776 , n5775 );
and ( n5777 , n5774 , n5776 );
and ( n5778 , n5772 , n5777 );
xor ( n5779 , n5771 , n5778 );
and ( n5780 , n5632 , n5636 );
and ( n5781 , n5636 , n5641 );
and ( n5782 , n5632 , n5641 );
or ( n5783 , n5780 , n5781 , n5782 );
xor ( n5784 , n5779 , n5783 );
and ( n5785 , n5647 , n5651 );
and ( n5786 , n5651 , n5656 );
and ( n5787 , n5647 , n5656 );
or ( n5788 , n5785 , n5786 , n5787 );
xor ( n5789 , n5784 , n5788 );
xor ( n5790 , n5765 , n5789 );
and ( n5791 , n5614 , n5615 );
and ( n5792 , n5615 , n5620 );
and ( n5793 , n5614 , n5620 );
or ( n5794 , n5791 , n5792 , n5793 );
and ( n5795 , n4968 , n4596 );
and ( n5796 , n5113 , n4472 );
nor ( n5797 , n5795 , n5796 );
xnor ( n5798 , n5797 , n4586 );
and ( n5799 , n4262 , n5458 );
and ( n5800 , n4369 , n5304 );
nor ( n5801 , n5799 , n5800 );
xnor ( n5802 , n5801 , n5448 );
xor ( n5803 , n5798 , n5802 );
xor ( n5804 , n5774 , n5654 );
not ( n5805 , n5655 );
and ( n5806 , n5804 , n5805 );
and ( n5807 , n3978 , n5806 );
and ( n5808 , n4188 , n5655 );
nor ( n5809 , n5807 , n5808 );
xnor ( n5810 , n5809 , n5777 );
xor ( n5811 , n5803 , n5810 );
xor ( n5812 , n5794 , n5811 );
and ( n5813 , n5272 , n4359 );
and ( n5814 , n5476 , n4268 );
nor ( n5815 , n5813 , n5814 );
xnor ( n5816 , n5815 , n4365 );
and ( n5817 , n4698 , n4849 );
and ( n5818 , n4821 , n4709 );
nor ( n5819 , n5817 , n5818 );
xnor ( n5820 , n5819 , n4830 );
xor ( n5821 , n5816 , n5820 );
and ( n5822 , n4461 , n5126 );
and ( n5823 , n4577 , n4979 );
nor ( n5824 , n5822 , n5823 );
xnor ( n5825 , n5824 , n5132 );
xor ( n5826 , n5821 , n5825 );
xor ( n5827 , n5812 , n5826 );
xor ( n5828 , n5790 , n5827 );
and ( n5829 , n5610 , n5621 );
and ( n5830 , n5621 , n5658 );
and ( n5831 , n5610 , n5658 );
or ( n5832 , n5829 , n5830 , n5831 );
xor ( n5833 , n5828 , n5832 );
and ( n5834 , n5606 , n5659 );
and ( n5835 , n5660 , n5663 );
or ( n5836 , n5834 , n5835 );
xor ( n5837 , n5833 , n5836 );
buf ( n5838 , n5837 );
and ( n5839 , n5736 , n5740 );
and ( n5840 , n5670 , n5694 );
and ( n5841 , n5694 , n5735 );
and ( n5842 , n5670 , n5735 );
or ( n5843 , n5840 , n5841 , n5842 );
and ( n5844 , n5699 , n5710 );
and ( n5845 , n5710 , n5734 );
and ( n5846 , n5699 , n5734 );
or ( n5847 , n5844 , n5845 , n5846 );
and ( n5848 , n5703 , n5704 );
and ( n5849 , n5704 , n5709 );
and ( n5850 , n5703 , n5709 );
or ( n5851 , n5848 , n5849 , n5850 );
and ( n5852 , n4525 , n4499 );
and ( n5853 , n4645 , n4419 );
nor ( n5854 , n5852 , n5853 );
xnor ( n5855 , n5854 , n4505 );
and ( n5856 , n4308 , n4744 );
and ( n5857 , n4413 , n4651 );
nor ( n5858 , n5856 , n5857 );
xnor ( n5859 , n5858 , n4750 );
xor ( n5860 , n5855 , n5859 );
and ( n5861 , n4013 , n5347 );
xor ( n5862 , n5860 , n5861 );
xor ( n5863 , n5851 , n5862 );
and ( n5864 , n5726 , n5730 );
and ( n5865 , n5730 , n5732 );
and ( n5866 , n5726 , n5732 );
or ( n5867 , n5864 , n5865 , n5866 );
or ( n5868 , n5712 , n5716 );
xor ( n5869 , n5867 , n5868 );
and ( n5870 , n4019 , n5350 );
and ( n5871 , n4035 , n5226 );
nor ( n5872 , n5870 , n5871 );
xnor ( n5873 , n5872 , n5356 );
xor ( n5874 , n5869 , n5873 );
xor ( n5875 , n5863 , n5874 );
xor ( n5876 , n5847 , n5875 );
and ( n5877 , n5674 , n5678 );
and ( n5878 , n5678 , n5693 );
and ( n5879 , n5674 , n5693 );
or ( n5880 , n5877 , n5878 , n5879 );
and ( n5881 , n5717 , n5721 );
and ( n5882 , n5721 , n5733 );
and ( n5883 , n5717 , n5733 );
or ( n5884 , n5881 , n5882 , n5883 );
xor ( n5885 , n5880 , n5884 );
and ( n5886 , n4780 , n4291 );
and ( n5887 , n4881 , n4206 );
nor ( n5888 , n5886 , n5887 );
xnor ( n5889 , n5888 , n4297 );
and ( n5890 , n4043 , n5033 );
and ( n5891 , n4216 , n4887 );
nor ( n5892 , n5890 , n5891 );
xnor ( n5893 , n5892 , n5019 );
xor ( n5894 , n5889 , n5893 );
and ( n5895 , n5683 , n5687 );
and ( n5896 , n5687 , n5692 );
and ( n5897 , n5683 , n5692 );
or ( n5898 , n5895 , n5896 , n5897 );
xor ( n5899 , n5894 , n5898 );
and ( n5900 , n5367 , n4016 );
not ( n5901 , n5900 );
xnor ( n5902 , n5901 , n3997 );
and ( n5903 , n5026 , n4050 );
and ( n5904 , n5220 , n4004 );
nor ( n5905 , n5903 , n5904 );
xnor ( n5906 , n5905 , n4029 );
xnor ( n5907 , n5902 , n5906 );
xor ( n5908 , n5899 , n5907 );
xor ( n5909 , n5885 , n5908 );
xor ( n5910 , n5876 , n5909 );
xor ( n5911 , n5843 , n5910 );
xor ( n5912 , n5839 , n5911 );
and ( n5913 , n5666 , n5741 );
and ( n5914 , n5742 , n5743 );
or ( n5915 , n5913 , n5914 );
xor ( n5916 , n5912 , n5915 );
buf ( n5917 , n5916 );
buf ( n5918 , n3176 );
and ( n5919 , n5746 , n5747 );
xor ( n5920 , n5918 , n5919 );
buf ( n5921 , n5920 );
not ( n5922 , n454 );
and ( n5923 , n5922 , n5917 );
and ( n5924 , n5921 , n454 );
or ( n5925 , n5923 , n5924 );
buf ( n5926 , n5925 );
and ( n5927 , n5754 , n5755 );
xor ( n5928 , n5926 , n5927 );
buf ( n5929 , n5928 );
not ( n5930 , n4176 );
and ( n5931 , n5930 , n5838 );
and ( n5932 , n5929 , n4176 );
or ( n5933 , n5931 , n5932 );
and ( n5934 , n5794 , n5811 );
and ( n5935 , n5811 , n5826 );
and ( n5936 , n5794 , n5826 );
or ( n5937 , n5934 , n5935 , n5936 );
and ( n5938 , n5798 , n5802 );
and ( n5939 , n5802 , n5810 );
and ( n5940 , n5798 , n5810 );
or ( n5941 , n5938 , n5939 , n5940 );
and ( n5942 , n5816 , n5820 );
and ( n5943 , n5820 , n5825 );
and ( n5944 , n5816 , n5825 );
or ( n5945 , n5942 , n5943 , n5944 );
xor ( n5946 , n5941 , n5945 );
and ( n5947 , n5768 , n4185 );
buf ( n5948 , n490 );
buf ( n5949 , n5948 );
and ( n5950 , n5949 , n3980 );
nor ( n5951 , n5947 , n5950 );
xnor ( n5952 , n5951 , n4182 );
and ( n5953 , n5476 , n4359 );
and ( n5954 , n5629 , n4268 );
nor ( n5955 , n5953 , n5954 );
xnor ( n5956 , n5955 , n4365 );
xor ( n5957 , n5952 , n5956 );
and ( n5958 , n3978 , n5774 );
xor ( n5959 , n5957 , n5958 );
xor ( n5960 , n5946 , n5959 );
xor ( n5961 , n5937 , n5960 );
and ( n5962 , n5779 , n5783 );
and ( n5963 , n5783 , n5788 );
and ( n5964 , n5779 , n5788 );
or ( n5965 , n5962 , n5963 , n5964 );
and ( n5966 , n5113 , n4596 );
and ( n5967 , n5272 , n4472 );
nor ( n5968 , n5966 , n5967 );
xnor ( n5969 , n5968 , n4586 );
and ( n5970 , n4821 , n4849 );
and ( n5971 , n4968 , n4709 );
nor ( n5972 , n5970 , n5971 );
xnor ( n5973 , n5972 , n4830 );
xor ( n5974 , n5969 , n5973 );
and ( n5975 , n4577 , n5126 );
and ( n5976 , n4698 , n4979 );
nor ( n5977 , n5975 , n5976 );
xnor ( n5978 , n5977 , n5132 );
xor ( n5979 , n5974 , n5978 );
xor ( n5980 , n5965 , n5979 );
and ( n5981 , n5771 , n5778 );
and ( n5982 , n4369 , n5458 );
and ( n5983 , n4461 , n5304 );
nor ( n5984 , n5982 , n5983 );
xnor ( n5985 , n5984 , n5448 );
xor ( n5986 , n5981 , n5985 );
and ( n5987 , n4188 , n5806 );
and ( n5988 , n4262 , n5655 );
nor ( n5989 , n5987 , n5988 );
xnor ( n5990 , n5989 , n5777 );
xor ( n5991 , n5986 , n5990 );
xor ( n5992 , n5980 , n5991 );
xor ( n5993 , n5961 , n5992 );
and ( n5994 , n5765 , n5789 );
and ( n5995 , n5789 , n5827 );
and ( n5996 , n5765 , n5827 );
or ( n5997 , n5994 , n5995 , n5996 );
xor ( n5998 , n5993 , n5997 );
and ( n5999 , n5828 , n5832 );
and ( n6000 , n5833 , n5836 );
or ( n6001 , n5999 , n6000 );
xor ( n6002 , n5998 , n6001 );
buf ( n6003 , n6002 );
and ( n6004 , n5843 , n5910 );
and ( n6005 , n5880 , n5884 );
and ( n6006 , n5884 , n5908 );
and ( n6007 , n5880 , n5908 );
or ( n6008 , n6005 , n6006 , n6007 );
and ( n6009 , n5867 , n5868 );
and ( n6010 , n5868 , n5873 );
and ( n6011 , n5867 , n5873 );
or ( n6012 , n6009 , n6010 , n6011 );
and ( n6013 , n4881 , n4291 );
and ( n6014 , n5026 , n4206 );
nor ( n6015 , n6013 , n6014 );
xnor ( n6016 , n6015 , n4297 );
and ( n6017 , n4413 , n4744 );
and ( n6018 , n4525 , n4651 );
nor ( n6019 , n6017 , n6018 );
xnor ( n6020 , n6019 , n4750 );
xor ( n6021 , n6016 , n6020 );
and ( n6022 , n4019 , n5347 );
xor ( n6023 , n6021 , n6022 );
xor ( n6024 , n6012 , n6023 );
and ( n6025 , n5889 , n5893 );
and ( n6026 , n4216 , n5033 );
and ( n6027 , n4308 , n4887 );
nor ( n6028 , n6026 , n6027 );
xnor ( n6029 , n6028 , n5019 );
xor ( n6030 , n6025 , n6029 );
and ( n6031 , n4035 , n5350 );
and ( n6032 , n4043 , n5226 );
nor ( n6033 , n6031 , n6032 );
xnor ( n6034 , n6033 , n5356 );
xor ( n6035 , n6030 , n6034 );
xor ( n6036 , n6024 , n6035 );
xor ( n6037 , n6008 , n6036 );
and ( n6038 , n5851 , n5862 );
and ( n6039 , n5862 , n5874 );
and ( n6040 , n5851 , n5874 );
or ( n6041 , n6038 , n6039 , n6040 );
and ( n6042 , n5894 , n5898 );
and ( n6043 , n5898 , n5907 );
and ( n6044 , n5894 , n5907 );
or ( n6045 , n6042 , n6043 , n6044 );
xor ( n6046 , n6041 , n6045 );
and ( n6047 , n5855 , n5859 );
and ( n6048 , n5859 , n5861 );
and ( n6049 , n5855 , n5861 );
or ( n6050 , n6047 , n6048 , n6049 );
or ( n6051 , n5902 , n5906 );
xor ( n6052 , n6050 , n6051 );
not ( n6053 , n3997 );
and ( n6054 , n5220 , n4050 );
and ( n6055 , n5367 , n4004 );
nor ( n6056 , n6054 , n6055 );
xnor ( n6057 , n6056 , n4029 );
xor ( n6058 , n6053 , n6057 );
and ( n6059 , n4645 , n4499 );
and ( n6060 , n4780 , n4419 );
nor ( n6061 , n6059 , n6060 );
xnor ( n6062 , n6061 , n4505 );
xor ( n6063 , n6058 , n6062 );
xor ( n6064 , n6052 , n6063 );
xor ( n6065 , n6046 , n6064 );
xor ( n6066 , n6037 , n6065 );
and ( n6067 , n5847 , n5875 );
and ( n6068 , n5875 , n5909 );
and ( n6069 , n5847 , n5909 );
or ( n6070 , n6067 , n6068 , n6069 );
xor ( n6071 , n6066 , n6070 );
xor ( n6072 , n6004 , n6071 );
and ( n6073 , n5839 , n5911 );
and ( n6074 , n5912 , n5915 );
or ( n6075 , n6073 , n6074 );
xor ( n6076 , n6072 , n6075 );
buf ( n6077 , n6076 );
buf ( n6078 , n3302 );
and ( n6079 , n5918 , n5919 );
xor ( n6080 , n6078 , n6079 );
buf ( n6081 , n6080 );
not ( n6082 , n454 );
and ( n6083 , n6082 , n6077 );
and ( n6084 , n6081 , n454 );
or ( n6085 , n6083 , n6084 );
buf ( n6086 , n6085 );
and ( n6087 , n5926 , n5927 );
xor ( n6088 , n6086 , n6087 );
buf ( n6089 , n6088 );
not ( n6090 , n4176 );
and ( n6091 , n6090 , n6003 );
and ( n6092 , n6089 , n4176 );
or ( n6093 , n6091 , n6092 );
and ( n6094 , n5965 , n5979 );
and ( n6095 , n5979 , n5991 );
and ( n6096 , n5965 , n5991 );
or ( n6097 , n6094 , n6095 , n6096 );
and ( n6098 , n5969 , n5973 );
and ( n6099 , n5973 , n5978 );
and ( n6100 , n5969 , n5978 );
or ( n6101 , n6098 , n6099 , n6100 );
and ( n6102 , n5272 , n4596 );
and ( n6103 , n5476 , n4472 );
nor ( n6104 , n6102 , n6103 );
xnor ( n6105 , n6104 , n4586 );
and ( n6106 , n4698 , n5126 );
and ( n6107 , n4821 , n4979 );
nor ( n6108 , n6106 , n6107 );
xnor ( n6109 , n6108 , n5132 );
xor ( n6110 , n6105 , n6109 );
and ( n6111 , n4461 , n5458 );
and ( n6112 , n4577 , n5304 );
nor ( n6113 , n6111 , n6112 );
xnor ( n6114 , n6113 , n5448 );
xor ( n6115 , n6110 , n6114 );
xor ( n6116 , n6101 , n6115 );
and ( n6117 , n5629 , n4359 );
and ( n6118 , n5768 , n4268 );
nor ( n6119 , n6117 , n6118 );
xnor ( n6120 , n6119 , n4365 );
and ( n6121 , n4968 , n4849 );
and ( n6122 , n5113 , n4709 );
nor ( n6123 , n6121 , n6122 );
xnor ( n6124 , n6123 , n4830 );
xor ( n6125 , n6120 , n6124 );
and ( n6126 , n4188 , n5774 );
xor ( n6127 , n6125 , n6126 );
xor ( n6128 , n6116 , n6127 );
xor ( n6129 , n6097 , n6128 );
and ( n6130 , n5981 , n5985 );
and ( n6131 , n5985 , n5990 );
and ( n6132 , n5981 , n5990 );
or ( n6133 , n6130 , n6131 , n6132 );
and ( n6134 , n5941 , n5945 );
and ( n6135 , n5945 , n5959 );
and ( n6136 , n5941 , n5959 );
or ( n6137 , n6134 , n6135 , n6136 );
xor ( n6138 , n6133 , n6137 );
and ( n6139 , n5952 , n5956 );
and ( n6140 , n5956 , n5958 );
and ( n6141 , n5952 , n5958 );
or ( n6142 , n6139 , n6140 , n6141 );
and ( n6143 , n5949 , n4185 );
buf ( n6144 , n489 );
buf ( n6145 , n6144 );
and ( n6146 , n6145 , n3980 );
nor ( n6147 , n6143 , n6146 );
xnor ( n6148 , n6147 , n4182 );
xor ( n6149 , n6142 , n6148 );
and ( n6150 , n4262 , n5806 );
and ( n6151 , n4369 , n5655 );
nor ( n6152 , n6150 , n6151 );
xnor ( n6153 , n6152 , n5777 );
xor ( n6154 , n6149 , n6153 );
xor ( n6155 , n6138 , n6154 );
xor ( n6156 , n6129 , n6155 );
and ( n6157 , n5937 , n5960 );
and ( n6158 , n5960 , n5992 );
and ( n6159 , n5937 , n5992 );
or ( n6160 , n6157 , n6158 , n6159 );
xor ( n6161 , n6156 , n6160 );
and ( n6162 , n5993 , n5997 );
and ( n6163 , n5998 , n6001 );
or ( n6164 , n6162 , n6163 );
xor ( n6165 , n6161 , n6164 );
buf ( n6166 , n6165 );
and ( n6167 , n6066 , n6070 );
and ( n6168 , n6041 , n6045 );
and ( n6169 , n6045 , n6064 );
and ( n6170 , n6041 , n6064 );
or ( n6171 , n6168 , n6169 , n6170 );
and ( n6172 , n6025 , n6029 );
and ( n6173 , n6029 , n6034 );
and ( n6174 , n6025 , n6034 );
or ( n6175 , n6172 , n6173 , n6174 );
and ( n6176 , n5026 , n4291 );
and ( n6177 , n5220 , n4206 );
nor ( n6178 , n6176 , n6177 );
xnor ( n6179 , n6178 , n4297 );
and ( n6180 , n4525 , n4744 );
and ( n6181 , n4645 , n4651 );
nor ( n6182 , n6180 , n6181 );
xnor ( n6183 , n6182 , n4750 );
xor ( n6184 , n6179 , n6183 );
and ( n6185 , n4308 , n5033 );
and ( n6186 , n4413 , n4887 );
nor ( n6187 , n6185 , n6186 );
xnor ( n6188 , n6187 , n5019 );
xor ( n6189 , n6184 , n6188 );
xor ( n6190 , n6175 , n6189 );
and ( n6191 , n4780 , n4499 );
and ( n6192 , n4881 , n4419 );
nor ( n6193 , n6191 , n6192 );
xnor ( n6194 , n6193 , n4505 );
and ( n6195 , n4043 , n5350 );
and ( n6196 , n4216 , n5226 );
nor ( n6197 , n6195 , n6196 );
xnor ( n6198 , n6197 , n5356 );
xor ( n6199 , n6194 , n6198 );
and ( n6200 , n4035 , n5347 );
xor ( n6201 , n6199 , n6200 );
xor ( n6202 , n6190 , n6201 );
xor ( n6203 , n6171 , n6202 );
and ( n6204 , n6050 , n6051 );
and ( n6205 , n6051 , n6063 );
and ( n6206 , n6050 , n6063 );
or ( n6207 , n6204 , n6205 , n6206 );
and ( n6208 , n6012 , n6023 );
and ( n6209 , n6023 , n6035 );
and ( n6210 , n6012 , n6035 );
or ( n6211 , n6208 , n6209 , n6210 );
xor ( n6212 , n6207 , n6211 );
and ( n6213 , n6016 , n6020 );
and ( n6214 , n6020 , n6022 );
and ( n6215 , n6016 , n6022 );
or ( n6216 , n6213 , n6214 , n6215 );
and ( n6217 , n6053 , n6057 );
and ( n6218 , n6057 , n6062 );
and ( n6219 , n6053 , n6062 );
or ( n6220 , n6217 , n6218 , n6219 );
xor ( n6221 , n6216 , n6220 );
and ( n6222 , n5367 , n4050 );
not ( n6223 , n6222 );
xnor ( n6224 , n6223 , n4029 );
not ( n6225 , n6224 );
xor ( n6226 , n6221 , n6225 );
xor ( n6227 , n6212 , n6226 );
xor ( n6228 , n6203 , n6227 );
and ( n6229 , n6008 , n6036 );
and ( n6230 , n6036 , n6065 );
and ( n6231 , n6008 , n6065 );
or ( n6232 , n6229 , n6230 , n6231 );
xor ( n6233 , n6228 , n6232 );
xor ( n6234 , n6167 , n6233 );
and ( n6235 , n6004 , n6071 );
and ( n6236 , n6072 , n6075 );
or ( n6237 , n6235 , n6236 );
xor ( n6238 , n6234 , n6237 );
buf ( n6239 , n6238 );
buf ( n6240 , n3416 );
and ( n6241 , n6078 , n6079 );
xor ( n6242 , n6240 , n6241 );
buf ( n6243 , n6242 );
not ( n6244 , n454 );
and ( n6245 , n6244 , n6239 );
and ( n6246 , n6243 , n454 );
or ( n6247 , n6245 , n6246 );
buf ( n6248 , n6247 );
and ( n6249 , n6086 , n6087 );
xor ( n6250 , n6248 , n6249 );
buf ( n6251 , n6250 );
not ( n6252 , n4176 );
and ( n6253 , n6252 , n6166 );
and ( n6254 , n6251 , n4176 );
or ( n6255 , n6253 , n6254 );
and ( n6256 , n6133 , n6137 );
and ( n6257 , n6137 , n6154 );
and ( n6258 , n6133 , n6154 );
or ( n6259 , n6256 , n6257 , n6258 );
and ( n6260 , n6105 , n6109 );
and ( n6261 , n6109 , n6114 );
and ( n6262 , n6105 , n6114 );
or ( n6263 , n6260 , n6261 , n6262 );
and ( n6264 , n5476 , n4596 );
and ( n6265 , n5629 , n4472 );
nor ( n6266 , n6264 , n6265 );
xnor ( n6267 , n6266 , n4586 );
and ( n6268 , n4577 , n5458 );
and ( n6269 , n4698 , n5304 );
nor ( n6270 , n6268 , n6269 );
xnor ( n6271 , n6270 , n5448 );
xor ( n6272 , n6267 , n6271 );
and ( n6273 , n4369 , n5806 );
and ( n6274 , n4461 , n5655 );
nor ( n6275 , n6273 , n6274 );
xnor ( n6276 , n6275 , n5777 );
xor ( n6277 , n6272 , n6276 );
xor ( n6278 , n6263 , n6277 );
and ( n6279 , n5113 , n4849 );
and ( n6280 , n5272 , n4709 );
nor ( n6281 , n6279 , n6280 );
xnor ( n6282 , n6281 , n4830 );
and ( n6283 , n4821 , n5126 );
and ( n6284 , n4968 , n4979 );
nor ( n6285 , n6283 , n6284 );
xnor ( n6286 , n6285 , n5132 );
xor ( n6287 , n6282 , n6286 );
and ( n6288 , n4262 , n5774 );
xor ( n6289 , n6287 , n6288 );
xor ( n6290 , n6278 , n6289 );
xor ( n6291 , n6259 , n6290 );
and ( n6292 , n6120 , n6124 );
and ( n6293 , n6124 , n6126 );
and ( n6294 , n6120 , n6126 );
or ( n6295 , n6292 , n6293 , n6294 );
and ( n6296 , n6145 , n4185 );
not ( n6297 , n6296 );
xnor ( n6298 , n6297 , n4182 );
and ( n6299 , n5768 , n4359 );
and ( n6300 , n5949 , n4268 );
nor ( n6301 , n6299 , n6300 );
xnor ( n6302 , n6301 , n4365 );
xor ( n6303 , n6298 , n6302 );
xor ( n6304 , n6295 , n6303 );
and ( n6305 , n6142 , n6148 );
and ( n6306 , n6148 , n6153 );
and ( n6307 , n6142 , n6153 );
or ( n6308 , n6305 , n6306 , n6307 );
xor ( n6309 , n6304 , n6308 );
and ( n6310 , n6101 , n6115 );
and ( n6311 , n6115 , n6127 );
and ( n6312 , n6101 , n6127 );
or ( n6313 , n6310 , n6311 , n6312 );
xor ( n6314 , n6309 , n6313 );
xor ( n6315 , n6291 , n6314 );
and ( n6316 , n6097 , n6128 );
and ( n6317 , n6128 , n6155 );
and ( n6318 , n6097 , n6155 );
or ( n6319 , n6316 , n6317 , n6318 );
xor ( n6320 , n6315 , n6319 );
and ( n6321 , n6156 , n6160 );
and ( n6322 , n6161 , n6164 );
or ( n6323 , n6321 , n6322 );
xor ( n6324 , n6320 , n6323 );
buf ( n6325 , n6324 );
and ( n6326 , n6171 , n6202 );
and ( n6327 , n6202 , n6227 );
and ( n6328 , n6171 , n6227 );
or ( n6329 , n6326 , n6327 , n6328 );
and ( n6330 , n6207 , n6211 );
and ( n6331 , n6211 , n6226 );
and ( n6332 , n6207 , n6226 );
or ( n6333 , n6330 , n6331 , n6332 );
and ( n6334 , n6175 , n6189 );
and ( n6335 , n6189 , n6201 );
and ( n6336 , n6175 , n6201 );
or ( n6337 , n6334 , n6335 , n6336 );
and ( n6338 , n6216 , n6220 );
and ( n6339 , n6220 , n6225 );
and ( n6340 , n6216 , n6225 );
or ( n6341 , n6338 , n6339 , n6340 );
and ( n6342 , n6179 , n6183 );
and ( n6343 , n6183 , n6188 );
and ( n6344 , n6179 , n6188 );
or ( n6345 , n6342 , n6343 , n6344 );
buf ( n6346 , n6224 );
xor ( n6347 , n6345 , n6346 );
and ( n6348 , n4043 , n5347 );
xor ( n6349 , n6347 , n6348 );
xor ( n6350 , n6341 , n6349 );
and ( n6351 , n6194 , n6198 );
and ( n6352 , n6198 , n6200 );
and ( n6353 , n6194 , n6200 );
or ( n6354 , n6351 , n6352 , n6353 );
and ( n6355 , n4881 , n4499 );
and ( n6356 , n5026 , n4419 );
nor ( n6357 , n6355 , n6356 );
xnor ( n6358 , n6357 , n4505 );
and ( n6359 , n4413 , n5033 );
and ( n6360 , n4525 , n4887 );
nor ( n6361 , n6359 , n6360 );
xnor ( n6362 , n6361 , n5019 );
xor ( n6363 , n6358 , n6362 );
and ( n6364 , n4216 , n5350 );
and ( n6365 , n4308 , n5226 );
nor ( n6366 , n6364 , n6365 );
xnor ( n6367 , n6366 , n5356 );
xor ( n6368 , n6363 , n6367 );
xor ( n6369 , n6354 , n6368 );
not ( n6370 , n4029 );
and ( n6371 , n5220 , n4291 );
and ( n6372 , n5367 , n4206 );
nor ( n6373 , n6371 , n6372 );
xnor ( n6374 , n6373 , n4297 );
xor ( n6375 , n6370 , n6374 );
and ( n6376 , n4645 , n4744 );
and ( n6377 , n4780 , n4651 );
nor ( n6378 , n6376 , n6377 );
xnor ( n6379 , n6378 , n4750 );
xor ( n6380 , n6375 , n6379 );
xor ( n6381 , n6369 , n6380 );
xor ( n6382 , n6350 , n6381 );
xor ( n6383 , n6337 , n6382 );
xor ( n6384 , n6333 , n6383 );
xor ( n6385 , n6329 , n6384 );
and ( n6386 , n6228 , n6232 );
xor ( n6387 , n6385 , n6386 );
and ( n6388 , n6167 , n6233 );
and ( n6389 , n6234 , n6237 );
or ( n6390 , n6388 , n6389 );
xor ( n6391 , n6387 , n6390 );
buf ( n6392 , n6391 );
buf ( n6393 , n3522 );
and ( n6394 , n6240 , n6241 );
xor ( n6395 , n6393 , n6394 );
buf ( n6396 , n6395 );
not ( n6397 , n454 );
and ( n6398 , n6397 , n6392 );
and ( n6399 , n6396 , n454 );
or ( n6400 , n6398 , n6399 );
buf ( n6401 , n6400 );
and ( n6402 , n6248 , n6249 );
xor ( n6403 , n6401 , n6402 );
buf ( n6404 , n6403 );
not ( n6405 , n4176 );
and ( n6406 , n6405 , n6325 );
and ( n6407 , n6404 , n4176 );
or ( n6408 , n6406 , n6407 );
and ( n6409 , n6304 , n6308 );
and ( n6410 , n6308 , n6313 );
and ( n6411 , n6304 , n6313 );
or ( n6412 , n6409 , n6410 , n6411 );
and ( n6413 , n6263 , n6277 );
and ( n6414 , n6277 , n6289 );
and ( n6415 , n6263 , n6289 );
or ( n6416 , n6413 , n6414 , n6415 );
and ( n6417 , n6295 , n6303 );
xor ( n6418 , n6416 , n6417 );
and ( n6419 , n6267 , n6271 );
and ( n6420 , n6271 , n6276 );
and ( n6421 , n6267 , n6276 );
or ( n6422 , n6419 , n6420 , n6421 );
and ( n6423 , n6282 , n6286 );
and ( n6424 , n6286 , n6288 );
and ( n6425 , n6282 , n6288 );
or ( n6426 , n6423 , n6424 , n6425 );
xor ( n6427 , n6422 , n6426 );
and ( n6428 , n6298 , n6302 );
xor ( n6429 , n6427 , n6428 );
xor ( n6430 , n6418 , n6429 );
xor ( n6431 , n6412 , n6430 );
not ( n6432 , n4182 );
and ( n6433 , n5949 , n4359 );
and ( n6434 , n6145 , n4268 );
nor ( n6435 , n6433 , n6434 );
xnor ( n6436 , n6435 , n4365 );
xnor ( n6437 , n6432 , n6436 );
and ( n6438 , n5629 , n4596 );
and ( n6439 , n5768 , n4472 );
nor ( n6440 , n6438 , n6439 );
xnor ( n6441 , n6440 , n4586 );
and ( n6442 , n4698 , n5458 );
and ( n6443 , n4821 , n5304 );
nor ( n6444 , n6442 , n6443 );
xnor ( n6445 , n6444 , n5448 );
xor ( n6446 , n6441 , n6445 );
and ( n6447 , n4461 , n5806 );
and ( n6448 , n4577 , n5655 );
nor ( n6449 , n6447 , n6448 );
xnor ( n6450 , n6449 , n5777 );
xor ( n6451 , n6446 , n6450 );
xor ( n6452 , n6437 , n6451 );
and ( n6453 , n5272 , n4849 );
and ( n6454 , n5476 , n4709 );
nor ( n6455 , n6453 , n6454 );
xnor ( n6456 , n6455 , n4830 );
and ( n6457 , n4968 , n5126 );
and ( n6458 , n5113 , n4979 );
nor ( n6459 , n6457 , n6458 );
xnor ( n6460 , n6459 , n5132 );
xor ( n6461 , n6456 , n6460 );
and ( n6462 , n4369 , n5774 );
xor ( n6463 , n6461 , n6462 );
xor ( n6464 , n6452 , n6463 );
xor ( n6465 , n6431 , n6464 );
and ( n6466 , n6259 , n6290 );
and ( n6467 , n6290 , n6314 );
and ( n6468 , n6259 , n6314 );
or ( n6469 , n6466 , n6467 , n6468 );
xor ( n6470 , n6465 , n6469 );
and ( n6471 , n6315 , n6319 );
and ( n6472 , n6320 , n6323 );
or ( n6473 , n6471 , n6472 );
xor ( n6474 , n6470 , n6473 );
buf ( n6475 , n6474 );
and ( n6476 , n6333 , n6383 );
and ( n6477 , n6341 , n6349 );
and ( n6478 , n6349 , n6381 );
and ( n6479 , n6341 , n6381 );
or ( n6480 , n6477 , n6478 , n6479 );
and ( n6481 , n6358 , n6362 );
and ( n6482 , n6362 , n6367 );
and ( n6483 , n6358 , n6367 );
or ( n6484 , n6481 , n6482 , n6483 );
and ( n6485 , n6370 , n6374 );
and ( n6486 , n6374 , n6379 );
and ( n6487 , n6370 , n6379 );
or ( n6488 , n6485 , n6486 , n6487 );
xor ( n6489 , n6484 , n6488 );
and ( n6490 , n5367 , n4291 );
not ( n6491 , n6490 );
xnor ( n6492 , n6491 , n4297 );
and ( n6493 , n4525 , n5033 );
and ( n6494 , n4645 , n4887 );
nor ( n6495 , n6493 , n6494 );
xnor ( n6496 , n6495 , n5019 );
xor ( n6497 , n6492 , n6496 );
and ( n6498 , n4308 , n5350 );
and ( n6499 , n4413 , n5226 );
nor ( n6500 , n6498 , n6499 );
xnor ( n6501 , n6500 , n5356 );
xor ( n6502 , n6497 , n6501 );
xor ( n6503 , n6489 , n6502 );
xor ( n6504 , n6480 , n6503 );
and ( n6505 , n6345 , n6346 );
and ( n6506 , n6346 , n6348 );
and ( n6507 , n6345 , n6348 );
or ( n6508 , n6505 , n6506 , n6507 );
and ( n6509 , n6354 , n6368 );
and ( n6510 , n6368 , n6380 );
and ( n6511 , n6354 , n6380 );
or ( n6512 , n6509 , n6510 , n6511 );
xor ( n6513 , n6508 , n6512 );
and ( n6514 , n5026 , n4499 );
and ( n6515 , n5220 , n4419 );
nor ( n6516 , n6514 , n6515 );
xnor ( n6517 , n6516 , n4505 );
not ( n6518 , n6517 );
and ( n6519 , n4780 , n4744 );
and ( n6520 , n4881 , n4651 );
nor ( n6521 , n6519 , n6520 );
xnor ( n6522 , n6521 , n4750 );
xor ( n6523 , n6518 , n6522 );
and ( n6524 , n4216 , n5347 );
xor ( n6525 , n6523 , n6524 );
xor ( n6526 , n6513 , n6525 );
xor ( n6527 , n6504 , n6526 );
and ( n6528 , n6337 , n6382 );
xor ( n6529 , n6527 , n6528 );
xor ( n6530 , n6476 , n6529 );
and ( n6531 , n6329 , n6384 );
and ( n6532 , n6384 , n6386 );
and ( n6533 , n6329 , n6386 );
or ( n6534 , n6531 , n6532 , n6533 );
xor ( n6535 , n6530 , n6534 );
and ( n6536 , n6387 , n6390 );
xor ( n6537 , n6535 , n6536 );
buf ( n6538 , n6537 );
buf ( n6539 , n3616 );
and ( n6540 , n6393 , n6394 );
xor ( n6541 , n6539 , n6540 );
buf ( n6542 , n6541 );
not ( n6543 , n454 );
and ( n6544 , n6543 , n6538 );
and ( n6545 , n6542 , n454 );
or ( n6546 , n6544 , n6545 );
buf ( n6547 , n6546 );
and ( n6548 , n6401 , n6402 );
xor ( n6549 , n6547 , n6548 );
buf ( n6550 , n6549 );
not ( n6551 , n4176 );
and ( n6552 , n6551 , n6475 );
and ( n6553 , n6550 , n4176 );
or ( n6554 , n6552 , n6553 );
and ( n6555 , n6416 , n6417 );
and ( n6556 , n6417 , n6429 );
and ( n6557 , n6416 , n6429 );
or ( n6558 , n6555 , n6556 , n6557 );
and ( n6559 , n6441 , n6445 );
and ( n6560 , n6445 , n6450 );
and ( n6561 , n6441 , n6450 );
or ( n6562 , n6559 , n6560 , n6561 );
and ( n6563 , n5476 , n4849 );
and ( n6564 , n5629 , n4709 );
nor ( n6565 , n6563 , n6564 );
xnor ( n6566 , n6565 , n4830 );
and ( n6567 , n4577 , n5806 );
and ( n6568 , n4698 , n5655 );
nor ( n6569 , n6567 , n6568 );
xnor ( n6570 , n6569 , n5777 );
xor ( n6571 , n6566 , n6570 );
and ( n6572 , n4461 , n5774 );
xor ( n6573 , n6571 , n6572 );
xor ( n6574 , n6562 , n6573 );
and ( n6575 , n5768 , n4596 );
and ( n6576 , n5949 , n4472 );
nor ( n6577 , n6575 , n6576 );
xnor ( n6578 , n6577 , n4586 );
and ( n6579 , n5113 , n5126 );
and ( n6580 , n5272 , n4979 );
nor ( n6581 , n6579 , n6580 );
xnor ( n6582 , n6581 , n5132 );
xor ( n6583 , n6578 , n6582 );
and ( n6584 , n4821 , n5458 );
and ( n6585 , n4968 , n5304 );
nor ( n6586 , n6584 , n6585 );
xnor ( n6587 , n6586 , n5448 );
xor ( n6588 , n6583 , n6587 );
xor ( n6589 , n6574 , n6588 );
xor ( n6590 , n6558 , n6589 );
and ( n6591 , n6422 , n6426 );
and ( n6592 , n6426 , n6428 );
and ( n6593 , n6422 , n6428 );
or ( n6594 , n6591 , n6592 , n6593 );
and ( n6595 , n6437 , n6451 );
and ( n6596 , n6451 , n6463 );
and ( n6597 , n6437 , n6463 );
or ( n6598 , n6595 , n6596 , n6597 );
xor ( n6599 , n6594 , n6598 );
and ( n6600 , n6456 , n6460 );
and ( n6601 , n6460 , n6462 );
and ( n6602 , n6456 , n6462 );
or ( n6603 , n6600 , n6601 , n6602 );
or ( n6604 , n6432 , n6436 );
xor ( n6605 , n6603 , n6604 );
and ( n6606 , n6145 , n4359 );
not ( n6607 , n6606 );
xnor ( n6608 , n6607 , n4365 );
not ( n6609 , n6608 );
xor ( n6610 , n6605 , n6609 );
xor ( n6611 , n6599 , n6610 );
xor ( n6612 , n6590 , n6611 );
and ( n6613 , n6412 , n6430 );
and ( n6614 , n6430 , n6464 );
and ( n6615 , n6412 , n6464 );
or ( n6616 , n6613 , n6614 , n6615 );
xor ( n6617 , n6612 , n6616 );
and ( n6618 , n6465 , n6469 );
and ( n6619 , n6470 , n6473 );
or ( n6620 , n6618 , n6619 );
xor ( n6621 , n6617 , n6620 );
buf ( n6622 , n6621 );
and ( n6623 , n6527 , n6528 );
and ( n6624 , n6484 , n6488 );
and ( n6625 , n6488 , n6502 );
and ( n6626 , n6484 , n6502 );
or ( n6627 , n6624 , n6625 , n6626 );
and ( n6628 , n6508 , n6512 );
and ( n6629 , n6512 , n6525 );
and ( n6630 , n6508 , n6525 );
or ( n6631 , n6628 , n6629 , n6630 );
xor ( n6632 , n6627 , n6631 );
and ( n6633 , n6518 , n6522 );
and ( n6634 , n6522 , n6524 );
and ( n6635 , n6518 , n6524 );
or ( n6636 , n6633 , n6634 , n6635 );
not ( n6637 , n4297 );
and ( n6638 , n5220 , n4499 );
and ( n6639 , n5367 , n4419 );
nor ( n6640 , n6638 , n6639 );
xnor ( n6641 , n6640 , n4505 );
xor ( n6642 , n6637 , n6641 );
and ( n6643 , n4645 , n5033 );
and ( n6644 , n4780 , n4887 );
nor ( n6645 , n6643 , n6644 );
xnor ( n6646 , n6645 , n5019 );
xor ( n6647 , n6642 , n6646 );
xor ( n6648 , n6636 , n6647 );
and ( n6649 , n6492 , n6496 );
and ( n6650 , n6496 , n6501 );
and ( n6651 , n6492 , n6501 );
or ( n6652 , n6649 , n6650 , n6651 );
buf ( n6653 , n6517 );
xor ( n6654 , n6652 , n6653 );
and ( n6655 , n4881 , n4744 );
and ( n6656 , n5026 , n4651 );
nor ( n6657 , n6655 , n6656 );
xnor ( n6658 , n6657 , n4750 );
and ( n6659 , n4413 , n5350 );
and ( n6660 , n4525 , n5226 );
nor ( n6661 , n6659 , n6660 );
xnor ( n6662 , n6661 , n5356 );
xor ( n6663 , n6658 , n6662 );
and ( n6664 , n4308 , n5347 );
xor ( n6665 , n6663 , n6664 );
xor ( n6666 , n6654 , n6665 );
xor ( n6667 , n6648 , n6666 );
xor ( n6668 , n6632 , n6667 );
and ( n6669 , n6480 , n6503 );
and ( n6670 , n6503 , n6526 );
and ( n6671 , n6480 , n6526 );
or ( n6672 , n6669 , n6670 , n6671 );
xor ( n6673 , n6668 , n6672 );
xor ( n6674 , n6623 , n6673 );
and ( n6675 , n6476 , n6529 );
and ( n6676 , n6529 , n6534 );
and ( n6677 , n6476 , n6534 );
or ( n6678 , n6675 , n6676 , n6677 );
xor ( n6679 , n6674 , n6678 );
and ( n6680 , n6535 , n6536 );
xor ( n6681 , n6679 , n6680 );
buf ( n6682 , n6681 );
buf ( n6683 , n3702 );
and ( n6684 , n6539 , n6540 );
xor ( n6685 , n6683 , n6684 );
buf ( n6686 , n6685 );
not ( n6687 , n454 );
and ( n6688 , n6687 , n6682 );
and ( n6689 , n6686 , n454 );
or ( n6690 , n6688 , n6689 );
buf ( n6691 , n6690 );
and ( n6692 , n6547 , n6548 );
xor ( n6693 , n6691 , n6692 );
buf ( n6694 , n6693 );
not ( n6695 , n4176 );
and ( n6696 , n6695 , n6622 );
and ( n6697 , n6694 , n4176 );
or ( n6698 , n6696 , n6697 );
and ( n6699 , n6558 , n6589 );
and ( n6700 , n6589 , n6611 );
and ( n6701 , n6558 , n6611 );
or ( n6702 , n6699 , n6700 , n6701 );
and ( n6703 , n6594 , n6598 );
and ( n6704 , n6598 , n6610 );
and ( n6705 , n6594 , n6610 );
or ( n6706 , n6703 , n6704 , n6705 );
and ( n6707 , n6566 , n6570 );
and ( n6708 , n6570 , n6572 );
and ( n6709 , n6566 , n6572 );
or ( n6710 , n6707 , n6708 , n6709 );
and ( n6711 , n5629 , n4849 );
and ( n6712 , n5768 , n4709 );
nor ( n6713 , n6711 , n6712 );
xnor ( n6714 , n6713 , n4830 );
and ( n6715 , n4968 , n5458 );
and ( n6716 , n5113 , n5304 );
nor ( n6717 , n6715 , n6716 );
xnor ( n6718 , n6717 , n5448 );
xor ( n6719 , n6714 , n6718 );
and ( n6720 , n4698 , n5806 );
and ( n6721 , n4821 , n5655 );
nor ( n6722 , n6720 , n6721 );
xnor ( n6723 , n6722 , n5777 );
xor ( n6724 , n6719 , n6723 );
xor ( n6725 , n6710 , n6724 );
not ( n6726 , n4365 );
and ( n6727 , n5949 , n4596 );
and ( n6728 , n6145 , n4472 );
nor ( n6729 , n6727 , n6728 );
xnor ( n6730 , n6729 , n4586 );
xor ( n6731 , n6726 , n6730 );
and ( n6732 , n5272 , n5126 );
and ( n6733 , n5476 , n4979 );
nor ( n6734 , n6732 , n6733 );
xnor ( n6735 , n6734 , n5132 );
xor ( n6736 , n6731 , n6735 );
xor ( n6737 , n6725 , n6736 );
xor ( n6738 , n6706 , n6737 );
and ( n6739 , n6603 , n6604 );
and ( n6740 , n6604 , n6609 );
and ( n6741 , n6603 , n6609 );
or ( n6742 , n6739 , n6740 , n6741 );
and ( n6743 , n6562 , n6573 );
and ( n6744 , n6573 , n6588 );
and ( n6745 , n6562 , n6588 );
or ( n6746 , n6743 , n6744 , n6745 );
xor ( n6747 , n6742 , n6746 );
and ( n6748 , n6578 , n6582 );
and ( n6749 , n6582 , n6587 );
and ( n6750 , n6578 , n6587 );
or ( n6751 , n6748 , n6749 , n6750 );
buf ( n6752 , n6608 );
xor ( n6753 , n6751 , n6752 );
and ( n6754 , n4577 , n5774 );
xor ( n6755 , n6753 , n6754 );
xor ( n6756 , n6747 , n6755 );
xor ( n6757 , n6738 , n6756 );
xor ( n6758 , n6702 , n6757 );
and ( n6759 , n6612 , n6616 );
and ( n6760 , n6617 , n6620 );
or ( n6761 , n6759 , n6760 );
xor ( n6762 , n6758 , n6761 );
buf ( n6763 , n6762 );
and ( n6764 , n6668 , n6672 );
and ( n6765 , n6652 , n6653 );
and ( n6766 , n6653 , n6665 );
and ( n6767 , n6652 , n6665 );
or ( n6768 , n6765 , n6766 , n6767 );
and ( n6769 , n6636 , n6647 );
and ( n6770 , n6647 , n6666 );
and ( n6771 , n6636 , n6666 );
or ( n6772 , n6769 , n6770 , n6771 );
xor ( n6773 , n6768 , n6772 );
and ( n6774 , n6637 , n6641 );
and ( n6775 , n6641 , n6646 );
and ( n6776 , n6637 , n6646 );
or ( n6777 , n6774 , n6775 , n6776 );
and ( n6778 , n5367 , n4499 );
not ( n6779 , n6778 );
xnor ( n6780 , n6779 , n4505 );
and ( n6781 , n4525 , n5350 );
and ( n6782 , n4645 , n5226 );
nor ( n6783 , n6781 , n6782 );
xnor ( n6784 , n6783 , n5356 );
xor ( n6785 , n6780 , n6784 );
and ( n6786 , n4413 , n5347 );
xor ( n6787 , n6785 , n6786 );
xor ( n6788 , n6777 , n6787 );
and ( n6789 , n6658 , n6662 );
and ( n6790 , n6662 , n6664 );
and ( n6791 , n6658 , n6664 );
or ( n6792 , n6789 , n6790 , n6791 );
and ( n6793 , n5026 , n4744 );
and ( n6794 , n5220 , n4651 );
nor ( n6795 , n6793 , n6794 );
xnor ( n6796 , n6795 , n4750 );
not ( n6797 , n6796 );
xor ( n6798 , n6792 , n6797 );
and ( n6799 , n4780 , n5033 );
and ( n6800 , n4881 , n4887 );
nor ( n6801 , n6799 , n6800 );
xnor ( n6802 , n6801 , n5019 );
xor ( n6803 , n6798 , n6802 );
xor ( n6804 , n6788 , n6803 );
xor ( n6805 , n6773 , n6804 );
and ( n6806 , n6627 , n6631 );
and ( n6807 , n6631 , n6667 );
and ( n6808 , n6627 , n6667 );
or ( n6809 , n6806 , n6807 , n6808 );
xor ( n6810 , n6805 , n6809 );
xor ( n6811 , n6764 , n6810 );
and ( n6812 , n6623 , n6673 );
and ( n6813 , n6673 , n6678 );
and ( n6814 , n6623 , n6678 );
or ( n6815 , n6812 , n6813 , n6814 );
xor ( n6816 , n6811 , n6815 );
and ( n6817 , n6679 , n6680 );
xor ( n6818 , n6816 , n6817 );
buf ( n6819 , n6818 );
buf ( n6820 , n3776 );
and ( n6821 , n6683 , n6684 );
xor ( n6822 , n6820 , n6821 );
buf ( n6823 , n6822 );
not ( n6824 , n454 );
and ( n6825 , n6824 , n6819 );
and ( n6826 , n6823 , n454 );
or ( n6827 , n6825 , n6826 );
buf ( n6828 , n6827 );
and ( n6829 , n6691 , n6692 );
xor ( n6830 , n6828 , n6829 );
buf ( n6831 , n6830 );
not ( n6832 , n4176 );
and ( n6833 , n6832 , n6763 );
and ( n6834 , n6831 , n4176 );
or ( n6835 , n6833 , n6834 );
and ( n6836 , n6742 , n6746 );
and ( n6837 , n6746 , n6755 );
and ( n6838 , n6742 , n6755 );
or ( n6839 , n6836 , n6837 , n6838 );
and ( n6840 , n6714 , n6718 );
and ( n6841 , n6718 , n6723 );
and ( n6842 , n6714 , n6723 );
or ( n6843 , n6840 , n6841 , n6842 );
and ( n6844 , n6726 , n6730 );
and ( n6845 , n6730 , n6735 );
and ( n6846 , n6726 , n6735 );
or ( n6847 , n6844 , n6845 , n6846 );
xor ( n6848 , n6843 , n6847 );
and ( n6849 , n6145 , n4596 );
not ( n6850 , n6849 );
xnor ( n6851 , n6850 , n4586 );
and ( n6852 , n5113 , n5458 );
and ( n6853 , n5272 , n5304 );
nor ( n6854 , n6852 , n6853 );
xnor ( n6855 , n6854 , n5448 );
xor ( n6856 , n6851 , n6855 );
and ( n6857 , n4821 , n5806 );
and ( n6858 , n4968 , n5655 );
nor ( n6859 , n6857 , n6858 );
xnor ( n6860 , n6859 , n5777 );
xor ( n6861 , n6856 , n6860 );
xor ( n6862 , n6848 , n6861 );
xor ( n6863 , n6839 , n6862 );
and ( n6864 , n6751 , n6752 );
and ( n6865 , n6752 , n6754 );
and ( n6866 , n6751 , n6754 );
or ( n6867 , n6864 , n6865 , n6866 );
and ( n6868 , n6710 , n6724 );
and ( n6869 , n6724 , n6736 );
and ( n6870 , n6710 , n6736 );
or ( n6871 , n6868 , n6869 , n6870 );
xor ( n6872 , n6867 , n6871 );
and ( n6873 , n5768 , n4849 );
and ( n6874 , n5949 , n4709 );
nor ( n6875 , n6873 , n6874 );
xnor ( n6876 , n6875 , n4830 );
not ( n6877 , n6876 );
and ( n6878 , n5476 , n5126 );
and ( n6879 , n5629 , n4979 );
nor ( n6880 , n6878 , n6879 );
xnor ( n6881 , n6880 , n5132 );
xor ( n6882 , n6877 , n6881 );
and ( n6883 , n4698 , n5774 );
xor ( n6884 , n6882 , n6883 );
xor ( n6885 , n6872 , n6884 );
xor ( n6886 , n6863 , n6885 );
and ( n6887 , n6706 , n6737 );
and ( n6888 , n6737 , n6756 );
and ( n6889 , n6706 , n6756 );
or ( n6890 , n6887 , n6888 , n6889 );
xor ( n6891 , n6886 , n6890 );
and ( n6892 , n6702 , n6757 );
and ( n6893 , n6758 , n6761 );
or ( n6894 , n6892 , n6893 );
xor ( n6895 , n6891 , n6894 );
buf ( n6896 , n6895 );
and ( n6897 , n6805 , n6809 );
and ( n6898 , n6768 , n6772 );
and ( n6899 , n6772 , n6804 );
and ( n6900 , n6768 , n6804 );
or ( n6901 , n6898 , n6899 , n6900 );
and ( n6902 , n6792 , n6797 );
and ( n6903 , n6797 , n6802 );
and ( n6904 , n6792 , n6802 );
or ( n6905 , n6902 , n6903 , n6904 );
and ( n6906 , n6777 , n6787 );
and ( n6907 , n6787 , n6803 );
and ( n6908 , n6777 , n6803 );
or ( n6909 , n6906 , n6907 , n6908 );
xor ( n6910 , n6905 , n6909 );
and ( n6911 , n6780 , n6784 );
and ( n6912 , n6784 , n6786 );
and ( n6913 , n6780 , n6786 );
or ( n6914 , n6911 , n6912 , n6913 );
not ( n6915 , n4505 );
and ( n6916 , n5220 , n4744 );
and ( n6917 , n5367 , n4651 );
nor ( n6918 , n6916 , n6917 );
xnor ( n6919 , n6918 , n4750 );
xor ( n6920 , n6915 , n6919 );
and ( n6921 , n4645 , n5350 );
and ( n6922 , n4780 , n5226 );
nor ( n6923 , n6921 , n6922 );
xnor ( n6924 , n6923 , n5356 );
xor ( n6925 , n6920 , n6924 );
xor ( n6926 , n6914 , n6925 );
buf ( n6927 , n6796 );
and ( n6928 , n4881 , n5033 );
and ( n6929 , n5026 , n4887 );
nor ( n6930 , n6928 , n6929 );
xnor ( n6931 , n6930 , n5019 );
xor ( n6932 , n6927 , n6931 );
and ( n6933 , n4525 , n5347 );
xor ( n6934 , n6932 , n6933 );
xor ( n6935 , n6926 , n6934 );
xor ( n6936 , n6910 , n6935 );
xor ( n6937 , n6901 , n6936 );
xor ( n6938 , n6897 , n6937 );
and ( n6939 , n6764 , n6810 );
and ( n6940 , n6810 , n6815 );
and ( n6941 , n6764 , n6815 );
or ( n6942 , n6939 , n6940 , n6941 );
xor ( n6943 , n6938 , n6942 );
and ( n6944 , n6816 , n6817 );
xor ( n6945 , n6943 , n6944 );
buf ( n6946 , n6945 );
buf ( n6947 , n3842 );
and ( n6948 , n6820 , n6821 );
xor ( n6949 , n6947 , n6948 );
buf ( n6950 , n6949 );
not ( n6951 , n454 );
and ( n6952 , n6951 , n6946 );
and ( n6953 , n6950 , n454 );
or ( n6954 , n6952 , n6953 );
buf ( n6955 , n6954 );
and ( n6956 , n6828 , n6829 );
xor ( n6957 , n6955 , n6956 );
buf ( n6958 , n6957 );
not ( n6959 , n4176 );
and ( n6960 , n6959 , n6896 );
and ( n6961 , n6958 , n4176 );
or ( n6962 , n6960 , n6961 );
and ( n6963 , n6843 , n6847 );
and ( n6964 , n6847 , n6861 );
and ( n6965 , n6843 , n6861 );
or ( n6966 , n6963 , n6964 , n6965 );
and ( n6967 , n6867 , n6871 );
and ( n6968 , n6871 , n6884 );
and ( n6969 , n6867 , n6884 );
or ( n6970 , n6967 , n6968 , n6969 );
xor ( n6971 , n6966 , n6970 );
and ( n6972 , n6877 , n6881 );
and ( n6973 , n6881 , n6883 );
and ( n6974 , n6877 , n6883 );
or ( n6975 , n6972 , n6973 , n6974 );
not ( n6976 , n4586 );
and ( n6977 , n5949 , n4849 );
and ( n6978 , n6145 , n4709 );
nor ( n6979 , n6977 , n6978 );
xnor ( n6980 , n6979 , n4830 );
xor ( n6981 , n6976 , n6980 );
and ( n6982 , n5272 , n5458 );
and ( n6983 , n5476 , n5304 );
nor ( n6984 , n6982 , n6983 );
xnor ( n6985 , n6984 , n5448 );
xor ( n6986 , n6981 , n6985 );
xor ( n6987 , n6975 , n6986 );
and ( n6988 , n6851 , n6855 );
and ( n6989 , n6855 , n6860 );
and ( n6990 , n6851 , n6860 );
or ( n6991 , n6988 , n6989 , n6990 );
buf ( n6992 , n6876 );
xor ( n6993 , n6991 , n6992 );
and ( n6994 , n5629 , n5126 );
and ( n6995 , n5768 , n4979 );
nor ( n6996 , n6994 , n6995 );
xnor ( n6997 , n6996 , n5132 );
and ( n6998 , n4968 , n5806 );
and ( n6999 , n5113 , n5655 );
nor ( n7000 , n6998 , n6999 );
xnor ( n7001 , n7000 , n5777 );
xor ( n7002 , n6997 , n7001 );
and ( n7003 , n4821 , n5774 );
xor ( n7004 , n7002 , n7003 );
xor ( n7005 , n6993 , n7004 );
xor ( n7006 , n6987 , n7005 );
xor ( n7007 , n6971 , n7006 );
and ( n7008 , n6839 , n6862 );
and ( n7009 , n6862 , n6885 );
and ( n7010 , n6839 , n6885 );
or ( n7011 , n7008 , n7009 , n7010 );
xor ( n7012 , n7007 , n7011 );
and ( n7013 , n6886 , n6890 );
and ( n7014 , n6891 , n6894 );
or ( n7015 , n7013 , n7014 );
xor ( n7016 , n7012 , n7015 );
buf ( n7017 , n7016 );
and ( n7018 , n6901 , n6936 );
and ( n7019 , n6927 , n6931 );
and ( n7020 , n6931 , n6933 );
and ( n7021 , n6927 , n6933 );
or ( n7022 , n7019 , n7020 , n7021 );
and ( n7023 , n6914 , n6925 );
and ( n7024 , n6925 , n6934 );
and ( n7025 , n6914 , n6934 );
or ( n7026 , n7023 , n7024 , n7025 );
xor ( n7027 , n7022 , n7026 );
and ( n7028 , n6915 , n6919 );
and ( n7029 , n6919 , n6924 );
and ( n7030 , n6915 , n6924 );
or ( n7031 , n7028 , n7029 , n7030 );
and ( n7032 , n5367 , n4744 );
not ( n7033 , n7032 );
xnor ( n7034 , n7033 , n4750 );
not ( n7035 , n7034 );
xor ( n7036 , n7031 , n7035 );
and ( n7037 , n5026 , n5033 );
and ( n7038 , n5220 , n4887 );
nor ( n7039 , n7037 , n7038 );
xnor ( n7040 , n7039 , n5019 );
and ( n7041 , n4780 , n5350 );
and ( n7042 , n4881 , n5226 );
nor ( n7043 , n7041 , n7042 );
xnor ( n7044 , n7043 , n5356 );
xor ( n7045 , n7040 , n7044 );
and ( n7046 , n4645 , n5347 );
xor ( n7047 , n7045 , n7046 );
xor ( n7048 , n7036 , n7047 );
xor ( n7049 , n7027 , n7048 );
and ( n7050 , n6905 , n6909 );
and ( n7051 , n6909 , n6935 );
and ( n7052 , n6905 , n6935 );
or ( n7053 , n7050 , n7051 , n7052 );
xor ( n7054 , n7049 , n7053 );
xor ( n7055 , n7018 , n7054 );
and ( n7056 , n6897 , n6937 );
and ( n7057 , n6937 , n6942 );
and ( n7058 , n6897 , n6942 );
or ( n7059 , n7056 , n7057 , n7058 );
xor ( n7060 , n7055 , n7059 );
and ( n7061 , n6943 , n6944 );
xor ( n7062 , n7060 , n7061 );
buf ( n7063 , n7062 );
buf ( n7064 , n3896 );
and ( n7065 , n6947 , n6948 );
xor ( n7066 , n7064 , n7065 );
buf ( n7067 , n7066 );
not ( n7068 , n454 );
and ( n7069 , n7068 , n7063 );
and ( n7070 , n7067 , n454 );
or ( n7071 , n7069 , n7070 );
buf ( n7072 , n7071 );
and ( n7073 , n6955 , n6956 );
xor ( n7074 , n7072 , n7073 );
buf ( n7075 , n7074 );
not ( n7076 , n4176 );
and ( n7077 , n7076 , n7017 );
and ( n7078 , n7075 , n4176 );
or ( n7079 , n7077 , n7078 );
and ( n7080 , n6991 , n6992 );
and ( n7081 , n6992 , n7004 );
and ( n7082 , n6991 , n7004 );
or ( n7083 , n7080 , n7081 , n7082 );
and ( n7084 , n6975 , n6986 );
and ( n7085 , n6986 , n7005 );
and ( n7086 , n6975 , n7005 );
or ( n7087 , n7084 , n7085 , n7086 );
xor ( n7088 , n7083 , n7087 );
and ( n7089 , n6976 , n6980 );
and ( n7090 , n6980 , n6985 );
and ( n7091 , n6976 , n6985 );
or ( n7092 , n7089 , n7090 , n7091 );
and ( n7093 , n6145 , n4849 );
not ( n7094 , n7093 );
xnor ( n7095 , n7094 , n4830 );
and ( n7096 , n5113 , n5806 );
and ( n7097 , n5272 , n5655 );
nor ( n7098 , n7096 , n7097 );
xnor ( n7099 , n7098 , n5777 );
xor ( n7100 , n7095 , n7099 );
and ( n7101 , n4968 , n5774 );
xor ( n7102 , n7100 , n7101 );
xor ( n7103 , n7092 , n7102 );
and ( n7104 , n6997 , n7001 );
and ( n7105 , n7001 , n7003 );
and ( n7106 , n6997 , n7003 );
or ( n7107 , n7104 , n7105 , n7106 );
and ( n7108 , n5768 , n5126 );
and ( n7109 , n5949 , n4979 );
nor ( n7110 , n7108 , n7109 );
xnor ( n7111 , n7110 , n5132 );
not ( n7112 , n7111 );
xor ( n7113 , n7107 , n7112 );
and ( n7114 , n5476 , n5458 );
and ( n7115 , n5629 , n5304 );
nor ( n7116 , n7114 , n7115 );
xnor ( n7117 , n7116 , n5448 );
xor ( n7118 , n7113 , n7117 );
xor ( n7119 , n7103 , n7118 );
xor ( n7120 , n7088 , n7119 );
and ( n7121 , n6966 , n6970 );
and ( n7122 , n6970 , n7006 );
and ( n7123 , n6966 , n7006 );
or ( n7124 , n7121 , n7122 , n7123 );
xor ( n7125 , n7120 , n7124 );
and ( n7126 , n7007 , n7011 );
and ( n7127 , n7012 , n7015 );
or ( n7128 , n7126 , n7127 );
xor ( n7129 , n7125 , n7128 );
buf ( n7130 , n7129 );
and ( n7131 , n7049 , n7053 );
and ( n7132 , n7031 , n7035 );
and ( n7133 , n7035 , n7047 );
and ( n7134 , n7031 , n7047 );
or ( n7135 , n7132 , n7133 , n7134 );
not ( n7136 , n4750 );
and ( n7137 , n5220 , n5033 );
and ( n7138 , n5367 , n4887 );
nor ( n7139 , n7137 , n7138 );
xnor ( n7140 , n7139 , n5019 );
xor ( n7141 , n7136 , n7140 );
and ( n7142 , n4780 , n5347 );
xor ( n7143 , n7141 , n7142 );
xor ( n7144 , n7135 , n7143 );
and ( n7145 , n7040 , n7044 );
and ( n7146 , n7044 , n7046 );
and ( n7147 , n7040 , n7046 );
or ( n7148 , n7145 , n7146 , n7147 );
buf ( n7149 , n7034 );
xor ( n7150 , n7148 , n7149 );
and ( n7151 , n4881 , n5350 );
and ( n7152 , n5026 , n5226 );
nor ( n7153 , n7151 , n7152 );
xnor ( n7154 , n7153 , n5356 );
xor ( n7155 , n7150 , n7154 );
xor ( n7156 , n7144 , n7155 );
and ( n7157 , n7022 , n7026 );
and ( n7158 , n7026 , n7048 );
and ( n7159 , n7022 , n7048 );
or ( n7160 , n7157 , n7158 , n7159 );
xor ( n7161 , n7156 , n7160 );
xor ( n7162 , n7131 , n7161 );
and ( n7163 , n7018 , n7054 );
and ( n7164 , n7054 , n7059 );
and ( n7165 , n7018 , n7059 );
or ( n7166 , n7163 , n7164 , n7165 );
xor ( n7167 , n7162 , n7166 );
and ( n7168 , n7060 , n7061 );
xor ( n7169 , n7167 , n7168 );
buf ( n7170 , n7169 );
buf ( n7171 , n3942 );
and ( n7172 , n7064 , n7065 );
xor ( n7173 , n7171 , n7172 );
buf ( n7174 , n7173 );
not ( n7175 , n454 );
and ( n7176 , n7175 , n7170 );
and ( n7177 , n7174 , n454 );
or ( n7178 , n7176 , n7177 );
buf ( n7179 , n7178 );
and ( n7180 , n7072 , n7073 );
xor ( n7181 , n7179 , n7180 );
buf ( n7182 , n7181 );
not ( n7183 , n4176 );
and ( n7184 , n7183 , n7130 );
and ( n7185 , n7182 , n4176 );
or ( n7186 , n7184 , n7185 );
and ( n7187 , n7083 , n7087 );
and ( n7188 , n7087 , n7119 );
and ( n7189 , n7083 , n7119 );
or ( n7190 , n7187 , n7188 , n7189 );
and ( n7191 , n7107 , n7112 );
and ( n7192 , n7112 , n7117 );
and ( n7193 , n7107 , n7117 );
or ( n7194 , n7191 , n7192 , n7193 );
and ( n7195 , n7092 , n7102 );
and ( n7196 , n7102 , n7118 );
and ( n7197 , n7092 , n7118 );
or ( n7198 , n7195 , n7196 , n7197 );
xor ( n7199 , n7194 , n7198 );
and ( n7200 , n7095 , n7099 );
and ( n7201 , n7099 , n7101 );
and ( n7202 , n7095 , n7101 );
or ( n7203 , n7200 , n7201 , n7202 );
not ( n7204 , n4830 );
and ( n7205 , n5949 , n5126 );
and ( n7206 , n6145 , n4979 );
nor ( n7207 , n7205 , n7206 );
xnor ( n7208 , n7207 , n5132 );
xor ( n7209 , n7204 , n7208 );
and ( n7210 , n5272 , n5806 );
and ( n7211 , n5476 , n5655 );
nor ( n7212 , n7210 , n7211 );
xnor ( n7213 , n7212 , n5777 );
xor ( n7214 , n7209 , n7213 );
xor ( n7215 , n7203 , n7214 );
buf ( n7216 , n7111 );
and ( n7217 , n5629 , n5458 );
and ( n7218 , n5768 , n5304 );
nor ( n7219 , n7217 , n7218 );
xnor ( n7220 , n7219 , n5448 );
xor ( n7221 , n7216 , n7220 );
and ( n7222 , n5113 , n5774 );
xor ( n7223 , n7221 , n7222 );
xor ( n7224 , n7215 , n7223 );
xor ( n7225 , n7199 , n7224 );
xor ( n7226 , n7190 , n7225 );
and ( n7227 , n7120 , n7124 );
and ( n7228 , n7125 , n7128 );
or ( n7229 , n7227 , n7228 );
xor ( n7230 , n7226 , n7229 );
buf ( n7231 , n7230 );
and ( n7232 , n7136 , n7140 );
and ( n7233 , n7140 , n7142 );
and ( n7234 , n7136 , n7142 );
or ( n7235 , n7232 , n7233 , n7234 );
and ( n7236 , n7148 , n7149 );
and ( n7237 , n7149 , n7154 );
and ( n7238 , n7148 , n7154 );
or ( n7239 , n7236 , n7237 , n7238 );
xor ( n7240 , n7235 , n7239 );
and ( n7241 , n5367 , n5033 );
not ( n7242 , n7241 );
xnor ( n7243 , n7242 , n5019 );
not ( n7244 , n7243 );
and ( n7245 , n5026 , n5350 );
and ( n7246 , n5220 , n5226 );
nor ( n7247 , n7245 , n7246 );
xnor ( n7248 , n7247 , n5356 );
xor ( n7249 , n7244 , n7248 );
and ( n7250 , n4881 , n5347 );
xor ( n7251 , n7249 , n7250 );
xor ( n7252 , n7240 , n7251 );
and ( n7253 , n7135 , n7143 );
and ( n7254 , n7143 , n7155 );
and ( n7255 , n7135 , n7155 );
or ( n7256 , n7253 , n7254 , n7255 );
xor ( n7257 , n7252 , n7256 );
and ( n7258 , n7156 , n7160 );
xor ( n7259 , n7257 , n7258 );
and ( n7260 , n7131 , n7161 );
and ( n7261 , n7161 , n7166 );
and ( n7262 , n7131 , n7166 );
or ( n7263 , n7260 , n7261 , n7262 );
xor ( n7264 , n7259 , n7263 );
and ( n7265 , n7167 , n7168 );
xor ( n7266 , n7264 , n7265 );
buf ( n7267 , n7266 );
buf ( n7268 , n3976 );
and ( n7269 , n7171 , n7172 );
xor ( n7270 , n7268 , n7269 );
buf ( n7271 , n7270 );
not ( n7272 , n454 );
and ( n7273 , n7272 , n7267 );
and ( n7274 , n7271 , n454 );
or ( n7275 , n7273 , n7274 );
buf ( n7276 , n7275 );
and ( n7277 , n7179 , n7180 );
xor ( n7278 , n7276 , n7277 );
buf ( n7279 , n7278 );
not ( n7280 , n4176 );
and ( n7281 , n7280 , n7231 );
and ( n7282 , n7279 , n4176 );
or ( n7283 , n7281 , n7282 );
and ( n7284 , n7216 , n7220 );
and ( n7285 , n7220 , n7222 );
and ( n7286 , n7216 , n7222 );
or ( n7287 , n7284 , n7285 , n7286 );
and ( n7288 , n7203 , n7214 );
and ( n7289 , n7214 , n7223 );
and ( n7290 , n7203 , n7223 );
or ( n7291 , n7288 , n7289 , n7290 );
xor ( n7292 , n7287 , n7291 );
and ( n7293 , n7204 , n7208 );
and ( n7294 , n7208 , n7213 );
and ( n7295 , n7204 , n7213 );
or ( n7296 , n7293 , n7294 , n7295 );
and ( n7297 , n6145 , n5126 );
not ( n7298 , n7297 );
xnor ( n7299 , n7298 , n5132 );
not ( n7300 , n7299 );
xor ( n7301 , n7296 , n7300 );
and ( n7302 , n5768 , n5458 );
and ( n7303 , n5949 , n5304 );
nor ( n7304 , n7302 , n7303 );
xnor ( n7305 , n7304 , n5448 );
and ( n7306 , n5476 , n5806 );
and ( n7307 , n5629 , n5655 );
nor ( n7308 , n7306 , n7307 );
xnor ( n7309 , n7308 , n5777 );
xor ( n7310 , n7305 , n7309 );
and ( n7311 , n5272 , n5774 );
xor ( n7312 , n7310 , n7311 );
xor ( n7313 , n7301 , n7312 );
xor ( n7314 , n7292 , n7313 );
and ( n7315 , n7194 , n7198 );
and ( n7316 , n7198 , n7224 );
and ( n7317 , n7194 , n7224 );
or ( n7318 , n7315 , n7316 , n7317 );
xor ( n7319 , n7314 , n7318 );
and ( n7320 , n7190 , n7225 );
and ( n7321 , n7226 , n7229 );
or ( n7322 , n7320 , n7321 );
xor ( n7323 , n7319 , n7322 );
buf ( n7324 , n7323 );
and ( n7325 , n7252 , n7256 );
and ( n7326 , n7244 , n7248 );
and ( n7327 , n7248 , n7250 );
and ( n7328 , n7244 , n7250 );
or ( n7329 , n7326 , n7327 , n7328 );
buf ( n7330 , n7243 );
xor ( n7331 , n7329 , n7330 );
not ( n7332 , n5019 );
and ( n7333 , n5220 , n5350 );
and ( n7334 , n5367 , n5226 );
nor ( n7335 , n7333 , n7334 );
xnor ( n7336 , n7335 , n5356 );
xor ( n7337 , n7332 , n7336 );
and ( n7338 , n5026 , n5347 );
xor ( n7339 , n7337 , n7338 );
xor ( n7340 , n7331 , n7339 );
and ( n7341 , n7235 , n7239 );
and ( n7342 , n7239 , n7251 );
and ( n7343 , n7235 , n7251 );
or ( n7344 , n7341 , n7342 , n7343 );
xor ( n7345 , n7340 , n7344 );
xor ( n7346 , n7325 , n7345 );
and ( n7347 , n7257 , n7258 );
and ( n7348 , n7258 , n7263 );
and ( n7349 , n7257 , n7263 );
or ( n7350 , n7347 , n7348 , n7349 );
xor ( n7351 , n7346 , n7350 );
and ( n7352 , n7264 , n7265 );
xor ( n7353 , n7351 , n7352 );
buf ( n7354 , n7353 );
and ( n7355 , n7268 , n7269 );
buf ( n7356 , n7355 );
not ( n7357 , n454 );
and ( n7358 , n7357 , n7354 );
and ( n7359 , n7356 , n454 );
or ( n7360 , n7358 , n7359 );
buf ( n7361 , n7360 );
and ( n7362 , n7276 , n7277 );
xor ( n7363 , n7361 , n7362 );
buf ( n7364 , n7363 );
not ( n7365 , n4176 );
and ( n7366 , n7365 , n7324 );
and ( n7367 , n7364 , n4176 );
or ( n7368 , n7366 , n7367 );
and ( n7369 , n7296 , n7300 );
and ( n7370 , n7300 , n7312 );
and ( n7371 , n7296 , n7312 );
or ( n7372 , n7369 , n7370 , n7371 );
not ( n7373 , n5132 );
and ( n7374 , n5949 , n5458 );
and ( n7375 , n6145 , n5304 );
nor ( n7376 , n7374 , n7375 );
xnor ( n7377 , n7376 , n5448 );
xor ( n7378 , n7373 , n7377 );
and ( n7379 , n5476 , n5774 );
xor ( n7380 , n7378 , n7379 );
xor ( n7381 , n7372 , n7380 );
and ( n7382 , n7305 , n7309 );
and ( n7383 , n7309 , n7311 );
and ( n7384 , n7305 , n7311 );
or ( n7385 , n7382 , n7383 , n7384 );
buf ( n7386 , n7299 );
xor ( n7387 , n7385 , n7386 );
and ( n7388 , n5629 , n5806 );
and ( n7389 , n5768 , n5655 );
nor ( n7390 , n7388 , n7389 );
xnor ( n7391 , n7390 , n5777 );
xor ( n7392 , n7387 , n7391 );
xor ( n7393 , n7381 , n7392 );
and ( n7394 , n7287 , n7291 );
and ( n7395 , n7291 , n7313 );
and ( n7396 , n7287 , n7313 );
or ( n7397 , n7394 , n7395 , n7396 );
xor ( n7398 , n7393 , n7397 );
and ( n7399 , n7314 , n7318 );
and ( n7400 , n7319 , n7322 );
or ( n7401 , n7399 , n7400 );
xor ( n7402 , n7398 , n7401 );
buf ( n7403 , n7402 );
and ( n7404 , n7332 , n7336 );
and ( n7405 , n7336 , n7338 );
and ( n7406 , n7332 , n7338 );
or ( n7407 , n7404 , n7405 , n7406 );
and ( n7408 , n5367 , n5350 );
not ( n7409 , n7408 );
xnor ( n7410 , n7409 , n5356 );
xor ( n7411 , n7407 , n7410 );
and ( n7412 , n5220 , n5347 );
not ( n7413 , n7412 );
xor ( n7414 , n7411 , n7413 );
and ( n7415 , n7329 , n7330 );
and ( n7416 , n7330 , n7339 );
and ( n7417 , n7329 , n7339 );
or ( n7418 , n7415 , n7416 , n7417 );
xor ( n7419 , n7414 , n7418 );
and ( n7420 , n7340 , n7344 );
xor ( n7421 , n7419 , n7420 );
and ( n7422 , n7325 , n7345 );
and ( n7423 , n7345 , n7350 );
and ( n7424 , n7325 , n7350 );
or ( n7425 , n7422 , n7423 , n7424 );
xor ( n7426 , n7421 , n7425 );
and ( n7427 , n7351 , n7352 );
xor ( n7428 , n7426 , n7427 );
buf ( n7429 , n7428 );
not ( n7430 , n454 );
and ( n7431 , n7430 , n7429 );
and ( n7432 , C0 , n454 );
or ( n7433 , n7431 , n7432 );
buf ( n7434 , n7433 );
and ( n7435 , n7361 , n7362 );
xor ( n7436 , n7434 , n7435 );
buf ( n7437 , n7436 );
not ( n7438 , n4176 );
and ( n7439 , n7438 , n7403 );
and ( n7440 , n7437 , n4176 );
or ( n7441 , n7439 , n7440 );
and ( n7442 , n7373 , n7377 );
and ( n7443 , n7377 , n7379 );
and ( n7444 , n7373 , n7379 );
or ( n7445 , n7442 , n7443 , n7444 );
and ( n7446 , n7385 , n7386 );
and ( n7447 , n7386 , n7391 );
and ( n7448 , n7385 , n7391 );
or ( n7449 , n7446 , n7447 , n7448 );
xor ( n7450 , n7445 , n7449 );
and ( n7451 , n6145 , n5458 );
not ( n7452 , n7451 );
xnor ( n7453 , n7452 , n5448 );
not ( n7454 , n7453 );
and ( n7455 , n5768 , n5806 );
and ( n7456 , n5949 , n5655 );
nor ( n7457 , n7455 , n7456 );
xnor ( n7458 , n7457 , n5777 );
xor ( n7459 , n7454 , n7458 );
and ( n7460 , n5629 , n5774 );
xor ( n7461 , n7459 , n7460 );
xor ( n7462 , n7450 , n7461 );
and ( n7463 , n7372 , n7380 );
and ( n7464 , n7380 , n7392 );
and ( n7465 , n7372 , n7392 );
or ( n7466 , n7463 , n7464 , n7465 );
xor ( n7467 , n7462 , n7466 );
and ( n7468 , n7393 , n7397 );
and ( n7469 , n7398 , n7401 );
or ( n7470 , n7468 , n7469 );
xor ( n7471 , n7467 , n7470 );
buf ( n7472 , n7471 );
and ( n7473 , n7414 , n7418 );
and ( n7474 , n7407 , n7410 );
and ( n7475 , n7410 , n7413 );
and ( n7476 , n7407 , n7413 );
or ( n7477 , n7474 , n7475 , n7476 );
buf ( n7478 , n7412 );
not ( n7479 , n5356 );
xor ( n7480 , n7478 , n7479 );
and ( n7481 , n5367 , n5347 );
xor ( n7482 , n7480 , n7481 );
xor ( n7483 , n7477 , n7482 );
xor ( n7484 , n7473 , n7483 );
and ( n7485 , n7419 , n7420 );
and ( n7486 , n7420 , n7425 );
and ( n7487 , n7419 , n7425 );
or ( n7488 , n7485 , n7486 , n7487 );
xor ( n7489 , n7484 , n7488 );
and ( n7490 , n7426 , n7427 );
xor ( n7491 , n7489 , n7490 );
buf ( n7492 , n7491 );
not ( n7493 , n454 );
and ( n7494 , n7493 , n7492 );
and ( n7495 , C0 , n454 );
or ( n7496 , n7494 , n7495 );
buf ( n7497 , n7496 );
and ( n7498 , n7434 , n7435 );
xor ( n7499 , n7497 , n7498 );
buf ( n7500 , n7499 );
not ( n7501 , n4176 );
and ( n7502 , n7501 , n7472 );
and ( n7503 , n7500 , n4176 );
or ( n7504 , n7502 , n7503 );
and ( n7505 , n7454 , n7458 );
and ( n7506 , n7458 , n7460 );
and ( n7507 , n7454 , n7460 );
or ( n7508 , n7505 , n7506 , n7507 );
buf ( n7509 , n7453 );
xor ( n7510 , n7508 , n7509 );
not ( n7511 , n5448 );
and ( n7512 , n5949 , n5806 );
and ( n7513 , n6145 , n5655 );
nor ( n7514 , n7512 , n7513 );
xnor ( n7515 , n7514 , n5777 );
xor ( n7516 , n7511 , n7515 );
and ( n7517 , n5768 , n5774 );
xor ( n7518 , n7516 , n7517 );
xor ( n7519 , n7510 , n7518 );
and ( n7520 , n7445 , n7449 );
and ( n7521 , n7449 , n7461 );
and ( n7522 , n7445 , n7461 );
or ( n7523 , n7520 , n7521 , n7522 );
xor ( n7524 , n7519 , n7523 );
and ( n7525 , n7462 , n7466 );
and ( n7526 , n7467 , n7470 );
or ( n7527 , n7525 , n7526 );
xor ( n7528 , n7524 , n7527 );
buf ( n7529 , n7528 );
and ( n7530 , n7478 , n7479 );
and ( n7531 , n7479 , n7481 );
and ( n7532 , n7478 , n7481 );
or ( n7533 , n7530 , n7531 , n7532 );
and ( n7534 , n7477 , n7482 );
xor ( n7535 , n7533 , n7534 );
and ( n7536 , n7473 , n7483 );
and ( n7537 , n7483 , n7488 );
and ( n7538 , n7473 , n7488 );
or ( n7539 , n7536 , n7537 , n7538 );
xnor ( n7540 , n7535 , n7539 );
and ( n7541 , n7489 , n7490 );
xor ( n7542 , n7540 , n7541 );
buf ( n7543 , n7542 );
not ( n7544 , n454 );
and ( n7545 , n7544 , n7543 );
and ( n7546 , C0 , n454 );
or ( n7547 , n7545 , n7546 );
buf ( n7548 , n7547 );
and ( n7549 , n7497 , n7498 );
xor ( n7550 , n7548 , n7549 );
buf ( n7551 , n7550 );
not ( n7552 , n4176 );
and ( n7553 , n7552 , n7529 );
and ( n7554 , n7551 , n4176 );
or ( n7555 , n7553 , n7554 );
and ( n7556 , n7511 , n7515 );
and ( n7557 , n7515 , n7517 );
and ( n7558 , n7511 , n7517 );
or ( n7559 , n7556 , n7557 , n7558 );
and ( n7560 , n6145 , n5806 );
not ( n7561 , n7560 );
xnor ( n7562 , n7561 , n5777 );
xor ( n7563 , n7559 , n7562 );
and ( n7564 , n5949 , n5774 );
not ( n7565 , n7564 );
xor ( n7566 , n7563 , n7565 );
and ( n7567 , n7508 , n7509 );
and ( n7568 , n7509 , n7518 );
and ( n7569 , n7508 , n7518 );
or ( n7570 , n7567 , n7568 , n7569 );
xor ( n7571 , n7566 , n7570 );
and ( n7572 , n7519 , n7523 );
and ( n7573 , n7524 , n7527 );
or ( n7574 , n7572 , n7573 );
xor ( n7575 , n7571 , n7574 );
buf ( n7576 , n7575 );
and ( n7577 , n7548 , n7549 );
buf ( n7578 , n7577 );
buf ( n7579 , n7578 );
not ( n7580 , n4176 );
and ( n7581 , n7580 , n7576 );
and ( n7582 , n7579 , n4176 );
or ( n7583 , n7581 , n7582 );
and ( n7584 , n7559 , n7562 );
and ( n7585 , n7562 , n7565 );
and ( n7586 , n7559 , n7565 );
or ( n7587 , n7584 , n7585 , n7586 );
buf ( n7588 , n7564 );
not ( n7589 , n5777 );
xor ( n7590 , n7588 , n7589 );
and ( n7591 , n6145 , n5774 );
xor ( n7592 , n7590 , n7591 );
xor ( n7593 , n7587 , n7592 );
and ( n7594 , n7566 , n7570 );
and ( n7595 , n7571 , n7574 );
or ( n7596 , n7594 , n7595 );
xor ( n7597 , n7593 , n7596 );
buf ( n7598 , n7597 );
not ( n7599 , n4176 );
and ( n7600 , n7599 , n7598 );
and ( n7601 , C0 , n4176 );
or ( n7602 , n7600 , n7601 );
xor ( n7603 , n4093 , n4123 );
buf ( n7604 , n7603 );
xor ( n7605 , n4150 , n4151 );
buf ( n7606 , n7605 );
not ( n7607 , n454 );
and ( n7608 , n7607 , n7604 );
and ( n7609 , n7606 , n454 );
or ( n7610 , n7608 , n7609 );
xor ( n7611 , n4121 , n4124 );
buf ( n7612 , n7611 );
xor ( n7613 , n4147 , n4148 );
xor ( n7614 , n7613 , n4152 );
buf ( n7615 , n7614 );
not ( n7616 , n454 );
and ( n7617 , n7616 , n7612 );
and ( n7618 , n7615 , n454 );
or ( n7619 , n7617 , n7618 );
xor ( n7620 , n4114 , n4126 );
buf ( n7621 , n7620 );
xor ( n7622 , n4144 , n4145 );
xor ( n7623 , n7622 , n4155 );
buf ( n7624 , n7623 );
not ( n7625 , n454 );
and ( n7626 , n7625 , n7621 );
and ( n7627 , n7624 , n454 );
or ( n7628 , n7626 , n7627 );
xor ( n7629 , n4106 , n4128 );
buf ( n7630 , n7629 );
xor ( n7631 , n4141 , n4142 );
xor ( n7632 , n7631 , n4158 );
buf ( n7633 , n7632 );
not ( n7634 , n454 );
and ( n7635 , n7634 , n7630 );
and ( n7636 , n7633 , n454 );
or ( n7637 , n7635 , n7636 );
xor ( n7638 , n4090 , n4130 );
buf ( n7639 , n7638 );
xor ( n7640 , n4138 , n4139 );
xor ( n7641 , n7640 , n4161 );
buf ( n7642 , n7641 );
not ( n7643 , n454 );
and ( n7644 , n7643 , n7639 );
and ( n7645 , n7642 , n454 );
or ( n7646 , n7644 , n7645 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
endmodule
