// IWLS benchmark module "MultiplierA_16" printed on Wed May 29 22:12:32 2002
module MultiplierA_16(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \36 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ;
output
  \36 ;
reg
  \2 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ;
wire
  \164 ,
  \166 ,
  \168 ,
  \170 ,
  \172 ,
  \174 ,
  \176 ,
  \178 ,
  \180 ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ,
  \96 ,
  \97 ,
  \98 ,
  \99 ,
  \[30] ,
  \[31] ,
  \[32] ,
  \100 ,
  \101 ,
  \102 ,
  \103 ,
  \104 ,
  \105 ,
  \106 ,
  \107 ,
  \111 ,
  \113 ,
  \115 ,
  \117 ,
  \119 ,
  \121 ,
  \123 ,
  \125 ,
  \127 ,
  \129 ,
  \131 ,
  \133 ,
  \[17] ,
  \135 ,
  \137 ,
  \140 ,
  \141 ,
  \[18] ,
  \144 ,
  \146 ,
  \147 ,
  \148 ,
  \149 ,
  \150 ,
  \152 ,
  \[19] ,
  \154 ,
  \156 ,
  \158 ,
  \160 ,
  \162 ;
assign
  \164  = \11  & \1 ,
  \166  = \10  & \1 ,
  \168  = \9  & \1 ,
  \170  = \8  & \1 ,
  \172  = \7  & \1 ,
  \174  = \6  & \1 ,
  \176  = \5  & \1 ,
  \178  = \4  & \1 ,
  \180  = \3  & \1 ,
  \[20]  = \90 ,
  \[21]  = \91 ,
  \[22]  = \92 ,
  \[23]  = \93 ,
  \[24]  = \94 ,
  \[25]  = \95 ,
  \[26]  = \96 ,
  \36  = \87 ,
  \[27]  = \97 ,
  \[28]  = \98 ,
  \[29]  = \99 ,
  \86  = (\152  & \137 ) | ((\152  & \34 ) | (\137  & \34 )),
  \87  = (~\180  & \20 ) | (\180  & ~\20 ),
  \88  = (~\178  & (~\111  & \21 )) | ((~\178  & (\111  & ~\21 )) | ((\178  & (~\111  & ~\21 )) | (\178  & (\111  & \21 )))),
  \89  = (~\176  & (~\113  & \22 )) | ((~\176  & (\113  & ~\22 )) | ((\176  & (~\113  & ~\22 )) | (\176  & (\113  & \22 )))),
  \90  = (~\174  & (~\115  & \23 )) | ((~\174  & (\115  & ~\23 )) | ((\174  & (~\115  & ~\23 )) | (\174  & (\115  & \23 )))),
  \91  = (~\172  & (~\117  & \24 )) | ((~\172  & (\117  & ~\24 )) | ((\172  & (~\117  & ~\24 )) | (\172  & (\117  & \24 )))),
  \92  = (~\170  & (~\119  & \25 )) | ((~\170  & (\119  & ~\25 )) | ((\170  & (~\119  & ~\25 )) | (\170  & (\119  & \25 )))),
  \93  = (~\168  & (~\121  & \26 )) | ((~\168  & (\121  & ~\26 )) | ((\168  & (~\121  & ~\26 )) | (\168  & (\121  & \26 )))),
  \94  = (~\166  & (~\123  & \27 )) | ((~\166  & (\123  & ~\27 )) | ((\166  & (~\123  & ~\27 )) | (\166  & (\123  & \27 )))),
  \95  = (~\164  & (~\125  & \28 )) | ((~\164  & (\125  & ~\28 )) | ((\164  & (~\125  & ~\28 )) | (\164  & (\125  & \28 )))),
  \96  = (~\162  & (~\127  & \29 )) | ((~\162  & (\127  & ~\29 )) | ((\162  & (~\127  & ~\29 )) | (\162  & (\127  & \29 )))),
  \97  = (~\160  & (~\129  & \30 )) | ((~\160  & (\129  & ~\30 )) | ((\160  & (~\129  & ~\30 )) | (\160  & (\129  & \30 )))),
  \98  = (~\158  & (~\131  & \31 )) | ((~\158  & (\131  & ~\31 )) | ((\158  & (~\131  & ~\31 )) | (\158  & (\131  & \31 )))),
  \99  = (~\156  & (~\133  & \32 )) | ((~\156  & (\133  & ~\32 )) | ((\156  & (~\133  & ~\32 )) | (\156  & (\133  & \32 )))),
  \[30]  = \100 ,
  \[31]  = \101 ,
  \[32]  = \102 ,
  \100  = (~\154  & (~\135  & \33 )) | ((~\154  & (\135  & ~\33 )) | ((\154  & (~\135  & ~\33 )) | (\154  & (\135  & \33 )))),
  \101  = (~\152  & (~\137  & \34 )) | ((~\152  & (\137  & ~\34 )) | ((\152  & (~\137  & ~\34 )) | (\152  & (\137  & \34 )))),
  \102  = (~\140  & \2 ) | (\140  & ~\2 ),
  \103  = \141  & ~\86 ,
  \104  = \144  & \86 ,
  \105  = \146  & \86 ,
  \106  = \147  & \86 ,
  \107  = \149  | \148 ,
  \111  = \180  & \20 ,
  \113  = (\178  & \111 ) | ((\178  & \21 ) | (\111  & \21 )),
  \115  = (\176  & \113 ) | ((\176  & \22 ) | (\113  & \22 )),
  \117  = (\174  & \115 ) | ((\174  & \23 ) | (\115  & \23 )),
  \119  = (\172  & \117 ) | ((\172  & \24 ) | (\117  & \24 )),
  \121  = (\170  & \119 ) | ((\170  & \25 ) | (\119  & \25 )),
  \123  = (\168  & \121 ) | ((\168  & \26 ) | (\121  & \26 )),
  \125  = (\166  & \123 ) | ((\166  & \27 ) | (\123  & \27 )),
  \127  = (\164  & \125 ) | ((\164  & \28 ) | (\125  & \28 )),
  \129  = (\162  & \127 ) | ((\162  & \29 ) | (\127  & \29 )),
  \131  = (\160  & \129 ) | ((\160  & \30 ) | (\129  & \30 )),
  \133  = (\158  & \131 ) | ((\158  & \31 ) | (\131  & \31 )),
  \[17]  = \107 ,
  \135  = (\156  & \133 ) | ((\156  & \32 ) | (\133  & \32 )),
  \137  = (\154  & \135 ) | ((\154  & \33 ) | (\135  & \33 )),
  \140  = (~\150  & \86 ) | (\150  & ~\86 ),
  \141  = \150  & \2 ,
  \[18]  = \88 ,
  \144  = ~\150  & \2 ,
  \146  = \150  & ~\2 ,
  \147  = \150  & \2 ,
  \148  = \104  | \103 ,
  \149  = \106  | \105 ,
  \150  = \18  & \1 ,
  \152  = \17  & \1 ,
  \[19]  = \89 ,
  \154  = \16  & \1 ,
  \156  = \15  & \1 ,
  \158  = \14  & \1 ,
  \160  = \13  & \1 ,
  \162  = \12  & \1 ;
always begin
  \2  = \[17] ;
  \20  = \[18] ;
  \21  = \[19] ;
  \22  = \[20] ;
  \23  = \[21] ;
  \24  = \[22] ;
  \25  = \[23] ;
  \26  = \[24] ;
  \27  = \[25] ;
  \28  = \[26] ;
  \29  = \[27] ;
  \30  = \[28] ;
  \31  = \[29] ;
  \32  = \[30] ;
  \33  = \[31] ;
  \34  = \[32] ;
end
initial begin
  \2  = 0;
  \20  = 0;
  \21  = 0;
  \22  = 0;
  \23  = 0;
  \24  = 0;
  \25  = 0;
  \26  = 0;
  \27  = 0;
  \28  = 0;
  \29  = 0;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
end
endmodule

