//NOTE: no-implementation module stub

module REG16L (
    input wire DSPCLK,
    input wire CLKSIrenb,
    input wire GO_C,
    input wire [15:0] SSin,
    output reg [15:0] SIr
);

endmodule
