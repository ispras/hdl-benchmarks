module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 ;
output g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 ;
wire t_0 , t_1 , t_2 , t_3 , t_4 , t_5 , t_6 , t_7 , t_8 , t_9 , t_10 , t_11 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( g17 , n18 );
buf ( g18 , n19 );
buf ( g19 , n20 );
buf ( g20 , n21 );
buf ( g21 , n22 );
buf ( g22 , n23 );
buf ( g23 , n24 );
buf ( g24 , n25 );
buf ( g25 , n26 );
buf ( g26 , n27 );
buf ( g27 , n28 );
buf ( g28 , n29 );
buf ( g29 , n30 );
buf ( g30 , n31 );
buf ( g31 , n32 );
buf ( n18 , n1956 );
buf ( n19 , n1585 );
buf ( n20 , n1913 );
buf ( n21 , n1466 );
buf ( n22 , n1793 );
buf ( n23 , n466 );
buf ( n24 , n678 );
buf ( n25 , n1948 );
buf ( n26 , n1948 );
buf ( n27 , n1936 );
buf ( n28 , n1846 );
buf ( n29 , n1284 );
buf ( n30 , n1700 );
buf ( n31 , n908 );
buf ( n32 , n1091 );
nand ( n35 , n4 , n5 );
not ( n36 , n35 );
not ( n37 , n2 );
nand ( n38 , n37 , n3 );
not ( n39 , n38 );
not ( n40 , n1 );
nand ( n41 , n6 , n7 );
not ( n42 , n41 );
not ( n43 , n42 );
not ( n44 , n43 );
not ( n45 , n44 );
not ( n46 , n45 );
not ( n47 , n46 );
nor ( n48 , n40 , n47 );
not ( n49 , n6 );
not ( n50 , n1 );
not ( n51 , n3 );
not ( n52 , n12 );
nand ( n53 , n52 , n13 );
not ( n54 , n13 );
nand ( n55 , n54 , n12 );
nand ( n56 , n53 , n55 );
not ( n57 , n17 );
not ( n58 , n2 );
nor ( n59 , n58 , n4 );
and ( n60 , n57 , n59 );
and ( n61 , n56 , n60 );
not ( n62 , n13 );
nand ( n63 , n62 , n4 );
nor ( n64 , n63 , n2 );
and ( n65 , n64 , n12 );
nor ( n66 , n61 , n65 );
not ( n67 , n16 );
nand ( n68 , n67 , n15 );
not ( n69 , n68 );
not ( n70 , n69 );
not ( n71 , n70 );
not ( n72 , n71 );
or ( n73 , n66 , n72 );
not ( n74 , n17 );
not ( n75 , n15 );
nand ( n76 , n75 , n16 );
not ( n77 , n76 );
not ( n78 , n77 );
nor ( n79 , n74 , n78 );
not ( n80 , n63 );
not ( n81 , n2 );
nand ( n82 , n79 , n80 , n81 );
nand ( n83 , n73 , n82 );
not ( n84 , n10 );
not ( n85 , n11 );
nand ( n86 , n84 , n85 );
not ( n87 , n86 );
and ( n88 , n83 , n87 );
not ( n89 , n72 );
and ( n90 , n2 , n4 );
and ( n91 , n89 , n90 );
nor ( n92 , n88 , n91 );
not ( n93 , n5 );
or ( n94 , n92 , n93 );
not ( n95 , n5 );
nand ( n96 , n95 , n4 );
not ( n97 , n96 );
not ( n98 , n97 );
not ( n99 , n98 );
not ( n100 , n99 );
not ( n101 , n17 );
and ( n102 , n101 , n71 );
nand ( n103 , n2 , n102 );
or ( n104 , n100 , n103 );
nand ( n105 , n94 , n104 );
and ( n106 , n51 , n105 );
not ( n107 , n3 );
nand ( n108 , n107 , n2 );
not ( n109 , n108 );
nor ( n110 , n4 , n5 );
not ( n111 , n110 );
not ( n112 , n111 );
buf ( n113 , n112 );
nand ( n114 , n109 , n113 );
nor ( n115 , n53 , n86 );
or ( n116 , n3 , n115 );
not ( n117 , n4 );
nor ( n118 , n117 , n2 );
and ( n119 , n5 , n118 );
nand ( n120 , n116 , n119 );
and ( n121 , n114 , n120 );
nand ( n122 , n16 , n17 );
nor ( n123 , n15 , n122 );
not ( n124 , n123 );
nand ( n125 , n124 , n70 );
not ( n126 , n125 );
nor ( n127 , n121 , n126 );
nor ( n128 , n106 , n127 );
not ( n129 , n9 );
or ( n130 , n128 , n129 );
not ( n131 , n2 );
not ( n132 , n4 );
nand ( n133 , n132 , n5 );
nand ( n134 , n133 , n96 );
not ( n135 , n3 );
nand ( n136 , n78 , n70 );
not ( n137 , n136 );
nor ( n138 , n135 , n137 );
and ( n139 , n134 , n138 );
not ( n140 , n113 );
not ( n141 , n140 );
nor ( n142 , n17 , n76 );
not ( n143 , n142 );
nor ( n144 , n3 , n143 );
and ( n145 , n141 , n144 );
nor ( n146 , n139 , n145 );
or ( n147 , n131 , n146 );
nand ( n148 , n130 , n147 );
nand ( n149 , n49 , n50 , n148 );
and ( n150 , t_10 , n149 );
not ( n151 , n14 );
nor ( n152 , n150 , n151 );
not ( n153 , n3 );
or ( n154 , n1 , n2 );
nor ( n155 , n153 , n154 );
nand ( n156 , n9 , n155 , n125 );
nor ( n157 , n5 , n6 );
not ( n158 , n157 );
nor ( n159 , n156 , n4 , n158 );
or ( n160 , n152 , n159 );
nand ( n161 , n160 , n8 );
nand ( n162 , n1 , n2 );
nand ( n163 , n3 , n4 );
nor ( n164 , n162 , n163 );
or ( n165 , n4 , n154 );
nor ( n166 , n3 , n165 );
or ( n167 , n164 , n166 );
not ( n168 , n5 );
nand ( n169 , n167 , n168 );
not ( n170 , n2 );
not ( n171 , n16 );
nor ( n172 , n171 , n17 );
not ( n173 , n172 );
not ( n174 , n173 );
nor ( n175 , n12 , n15 );
and ( n176 , n4 , n10 );
not ( n177 , n176 );
not ( n178 , n9 );
nand ( n179 , n178 , n5 );
nor ( n180 , n177 , n179 );
nand ( n181 , n174 , n175 , n3 , n180 );
not ( n182 , n181 );
not ( n183 , n9 );
not ( n184 , n15 );
not ( n185 , n16 );
nand ( n186 , n184 , n185 );
not ( n187 , n186 );
not ( n188 , n187 );
not ( n189 , n188 );
not ( n190 , n3 );
nand ( n191 , n190 , n4 );
not ( n192 , n191 );
nand ( n193 , n10 , n192 );
not ( n194 , n193 );
not ( n195 , n194 );
or ( n196 , n189 , n195 );
not ( n197 , n10 );
nand ( n198 , n7 , n197 );
nor ( n199 , n198 , n12 );
not ( n200 , n3 );
nand ( n201 , n200 , n191 );
not ( n202 , n13 );
nor ( n203 , n15 , n16 );
and ( n204 , n17 , n203 );
nand ( n205 , n199 , n201 , n202 , n204 );
nand ( n206 , n196 , n205 );
nand ( n207 , n183 , n206 );
not ( n208 , n207 );
not ( n209 , n186 );
nor ( n210 , n209 , n197 );
nand ( n211 , n4 , n9 );
not ( n212 , n211 );
nand ( n213 , n210 , n212 );
not ( n214 , n213 );
not ( n215 , n3 );
nor ( n216 , n12 , n13 );
not ( n217 , n216 );
nand ( n218 , n215 , n217 );
nand ( n219 , n214 , n218 );
not ( n220 , n219 );
or ( n221 , n208 , n220 );
not ( n222 , n5 );
nand ( n223 , n221 , n222 );
not ( n224 , n223 );
or ( n225 , n182 , n224 );
not ( n226 , n11 );
nand ( n227 , n225 , n226 );
not ( n228 , n9 );
nor ( n229 , n3 , n5 );
nand ( n230 , n184 , n122 );
nand ( n231 , n197 , n229 , n230 );
not ( n232 , n3 );
nand ( n233 , n232 , n5 );
not ( n234 , n5 );
nand ( n235 , n234 , n3 );
nand ( n236 , n233 , n235 );
nor ( n237 , n203 , n13 );
nand ( n238 , n236 , n10 , n237 );
nand ( n239 , n231 , n238 );
not ( n240 , n239 );
or ( n241 , n228 , n240 );
not ( n242 , n9 );
and ( n243 , n7 , n242 );
and ( n244 , n197 , n243 );
nand ( n245 , n5 , n233 );
nand ( n246 , n244 , n202 , n245 , n204 );
nand ( n247 , n241 , n246 );
not ( n248 , n12 );
nand ( n249 , n247 , n248 );
not ( n250 , n10 );
nor ( n251 , n250 , n9 );
not ( n252 , n251 );
not ( n253 , n252 );
not ( n254 , n229 );
buf ( n255 , n203 );
or ( n256 , n254 , n255 );
nand ( n257 , n3 , n5 );
not ( n258 , n257 );
and ( n259 , n12 , n258 );
nor ( n260 , n13 , n15 );
nand ( n261 , n259 , n172 , n260 );
nand ( n262 , n256 , n261 );
nand ( n263 , n253 , n262 );
and ( n264 , n249 , n263 );
nor ( n265 , n264 , n11 );
nand ( n266 , n12 , n13 );
not ( n267 , n266 );
nor ( n268 , n9 , n257 );
nand ( n269 , n197 , n172 , n267 , n268 );
not ( n270 , n11 );
nor ( n271 , n269 , n270 , n15 );
or ( n272 , n265 , n271 );
not ( n273 , n4 );
nand ( n274 , n272 , n273 );
and ( n275 , n227 , n274 );
not ( n276 , n1 );
nor ( n277 , n275 , n276 );
not ( n278 , n9 );
nor ( n279 , n278 , n13 );
not ( n280 , n17 );
nand ( n281 , n184 , n280 );
not ( n282 , n281 );
not ( n283 , n282 );
not ( n284 , n4 );
and ( n285 , n284 , n3 );
nand ( n286 , n279 , n283 , n285 , n87 );
not ( n287 , n4 );
not ( n288 , n77 );
nor ( n289 , n287 , n288 );
not ( n290 , n11 );
nor ( n291 , n290 , n17 );
not ( n292 , n3 );
and ( n293 , n292 , n251 );
nand ( n294 , n289 , n13 , n291 , n293 );
nand ( n295 , n286 , n294 );
and ( n296 , n295 , n5 , n248 );
not ( n297 , n187 );
not ( n298 , n297 );
not ( n299 , n298 );
nand ( n300 , n3 , n253 );
not ( n301 , n12 );
nand ( n302 , n301 , n11 );
nor ( n303 , n13 , n302 );
and ( n304 , n97 , n303 );
not ( n305 , n11 );
not ( n306 , n133 );
and ( n307 , n305 , n306 );
nor ( n308 , n304 , n307 );
or ( n309 , n300 , n308 );
nand ( n310 , n5 , n192 );
not ( n311 , n11 );
and ( n312 , n311 , n251 );
nor ( n313 , n312 , n9 );
or ( n314 , n310 , n313 );
nand ( n315 , n309 , n314 );
and ( n316 , n299 , n315 );
nor ( n317 , n296 , n316 );
nor ( n318 , n1 , n317 );
not ( n319 , n9 );
nor ( n320 , n11 , n15 );
nor ( n321 , n10 , n12 );
nor ( n322 , n13 , n16 );
nand ( n323 , n17 , n321 , n322 );
not ( n324 , n3 );
not ( n325 , n7 );
or ( n326 , n323 , n324 , n325 );
not ( n327 , n16 );
nor ( n328 , n327 , n17 );
nand ( n329 , n10 , n328 );
or ( n330 , n3 , n329 );
nand ( n331 , n326 , n330 );
and ( n332 , n319 , n320 , n36 , n331 );
nor ( n333 , n277 , n318 , n332 );
or ( n334 , n333 , n8 );
nand ( n335 , n8 , n325 );
not ( n336 , n5 );
nor ( n337 , n6 , n15 );
nor ( n338 , n16 , n17 );
not ( n339 , n338 );
not ( n340 , n339 );
not ( n341 , n340 );
not ( n342 , n341 );
not ( n343 , n4 );
not ( n344 , n1 );
nor ( n345 , n344 , n3 );
and ( n346 , n343 , n345 );
nand ( n347 , n336 , n337 , n342 , n346 );
or ( n348 , n335 , n347 );
not ( n349 , n1 );
buf ( n350 , n255 );
buf ( n351 , n350 );
and ( n352 , n3 , n134 );
not ( n353 , n192 );
nor ( n354 , n353 , n179 );
nor ( n355 , n352 , n354 );
not ( n356 , n41 );
nand ( n357 , n356 , n8 );
or ( n358 , n355 , n357 );
nor ( n359 , n6 , n7 );
not ( n360 , n359 );
or ( n361 , n360 , n310 );
nand ( n362 , n358 , n361 );
and ( n363 , n351 , n362 );
not ( n364 , n285 );
nor ( n365 , n5 , n364 );
and ( n366 , n8 , n6 , n7 );
not ( n367 , n366 );
nand ( n368 , n360 , n367 );
and ( n369 , n365 , n368 );
nor ( n370 , n363 , n369 );
or ( n371 , n370 , n17 );
not ( n372 , n299 );
not ( n373 , n372 );
nor ( n374 , n367 , n310 );
and ( n375 , n9 , n374 );
not ( n376 , n3 );
not ( n377 , n306 );
or ( n378 , n376 , n377 );
not ( n379 , n4 );
nand ( n380 , n378 , n379 );
and ( n381 , n17 , n380 );
nor ( n382 , n375 , n381 );
or ( n383 , n373 , n382 );
nand ( n384 , n371 , n383 );
nand ( n385 , n349 , n384 );
nand ( n386 , n334 , n348 , n385 );
nand ( n387 , n170 , n386 );
not ( n388 , n1 );
not ( n389 , n253 );
not ( n390 , n389 );
not ( n391 , n302 );
not ( n392 , n237 );
not ( n393 , n392 );
not ( n394 , n393 );
not ( n395 , n394 );
and ( n396 , t_2 , n391 , n395 );
not ( n397 , n134 );
nor ( n398 , n3 , n11 );
nor ( n399 , n8 , n9 );
nor ( n400 , n12 , n13 );
not ( n401 , n400 );
not ( n402 , n401 );
nand ( n403 , n197 , n398 , n399 , n402 );
nand ( n404 , t_3 , n403 );
not ( n405 , n404 );
or ( n406 , n397 , n405 );
not ( n407 , n401 );
nor ( n408 , n8 , n9 );
nand ( n409 , n407 , n408 );
not ( n410 , n409 );
not ( n411 , n3 );
nand ( n412 , n410 , n87 , n112 , n411 );
nand ( n413 , n406 , n412 );
nor ( n414 , n6 , n17 );
and ( n415 , n413 , n414 );
not ( n416 , n13 );
nand ( n417 , n416 , n17 );
not ( n418 , n417 );
nand ( n419 , n418 , n87 , n408 , n248 );
nor ( n420 , n419 , n35 , n3 );
nor ( n421 , n415 , n420 );
not ( n422 , n372 );
or ( n423 , n421 , n422 );
not ( n424 , n3 );
not ( n425 , n5 );
nor ( n426 , n4 , n419 );
and ( n427 , n425 , n426 );
not ( n428 , n298 );
and ( n429 , n36 , n428 );
nor ( n430 , n427 , n429 );
or ( n431 , n424 , n430 );
nand ( n432 , n423 , n431 );
and ( n433 , n432 , n325 );
nor ( n434 , n396 , n433 );
not ( n435 , n2 );
or ( n436 , n434 , n435 );
buf ( n437 , n351 );
not ( n438 , n365 );
or ( n439 , n437 , n438 );
nand ( n440 , n436 , n439 );
nand ( n441 , n388 , n440 );
nor ( n442 , n11 , n12 );
not ( n443 , n442 );
not ( n444 , n443 );
not ( n445 , n444 );
not ( n446 , n445 );
not ( n447 , n16 );
nand ( n448 , n447 , n17 );
not ( n449 , n448 );
not ( n450 , n449 );
not ( n451 , n450 );
not ( n452 , n451 );
not ( n453 , n452 );
not ( n454 , n453 );
nor ( n455 , n10 , n454 );
nor ( n456 , n3 , n8 );
and ( n457 , n456 , n260 );
not ( n458 , n1 );
not ( n459 , n5 );
nand ( n460 , n459 , n2 );
not ( n461 , n243 );
nor ( n462 , n458 , n460 , n461 );
nand ( n463 , n446 , n455 , n457 , n462 );
nand ( n464 , n387 , n441 , n463 );
nand ( n465 , n464 , n151 );
nand ( n466 , n161 , n169 , n465 );
not ( n467 , n185 );
nand ( n468 , n5 , n426 );
not ( n469 , n17 );
not ( n470 , n469 );
not ( n471 , n6 );
nand ( n472 , n471 , n8 );
not ( n473 , n472 );
not ( n474 , n473 );
or ( n475 , n470 , n474 );
not ( n476 , n8 );
nor ( n477 , n9 , n10 );
and ( n478 , n476 , n477 );
not ( n479 , n417 );
and ( n480 , n479 , n442 );
nand ( n481 , n478 , n480 );
nand ( n482 , n475 , n481 );
nand ( n483 , n99 , n482 );
and ( n484 , n468 , n483 );
not ( n485 , n2 );
nor ( n486 , n484 , n485 );
not ( n487 , n5 );
nor ( n488 , n2 , n4 );
nand ( n489 , n488 , n414 );
nor ( n490 , n487 , n489 );
nor ( n491 , n486 , n490 );
or ( n492 , n491 , n7 );
not ( n493 , n357 );
or ( n494 , n17 , n112 );
nand ( n495 , n494 , n35 );
and ( n496 , n493 , n495 );
and ( n497 , n17 , n113 );
nor ( n498 , n496 , n497 );
or ( n499 , n2 , n498 );
nand ( n500 , n492 , n499 );
not ( n501 , n500 );
or ( n502 , n467 , n501 );
not ( n503 , n5 );
not ( n504 , n10 );
nor ( n505 , n504 , n12 );
not ( n506 , n9 );
nand ( n507 , t_4 , n506 );
not ( n508 , n17 );
not ( n509 , n118 );
nand ( n510 , n16 , n476 );
nor ( n511 , n509 , n510 );
nand ( n512 , n503 , n507 , n508 , n511 );
nand ( n513 , n502 , n512 );
and ( n514 , n184 , n513 );
or ( n515 , n7 , n35 );
nand ( n516 , n515 , n4 );
nand ( n517 , n2 , n516 );
not ( n518 , n11 );
nor ( n519 , n8 , n98 );
not ( n520 , n2 );
nand ( n521 , n9 , n266 );
not ( n522 , n12 );
nand ( n523 , n522 , n9 );
nor ( n524 , n13 , n523 );
not ( n525 , n524 );
nand ( n526 , t_5 , n525 );
nand ( n527 , n518 , n519 , n520 , n526 );
and ( n528 , n517 , n527 );
nor ( n529 , n528 , n437 );
nor ( n530 , n514 , n529 );
or ( n531 , n1 , n530 );
not ( n532 , n10 );
nor ( n533 , n532 , n11 );
not ( n534 , n533 );
and ( n535 , n186 , n9 );
not ( n536 , n4 );
not ( n537 , n401 );
not ( n538 , n537 );
nand ( n539 , n536 , n538 );
and ( n540 , n535 , n539 );
not ( n541 , n9 );
nand ( n542 , n4 , n142 );
not ( n543 , n542 );
and ( n544 , n541 , n543 );
nor ( n545 , n540 , n544 );
or ( n546 , n5 , n534 , n545 );
nor ( n547 , n11 , n13 );
nor ( n548 , n4 , n10 );
nand ( n549 , n11 , n548 , n267 , n174 );
and ( n550 , n451 , n199 );
nor ( n551 , t_8 , n550 );
not ( n552 , n551 );
not ( n553 , n4 );
nand ( n554 , n552 , n553 , n202 );
nand ( n555 , n248 , n176 , n172 );
nand ( n556 , n554 , n555 );
not ( n557 , n11 );
nand ( n558 , n556 , n557 );
and ( n559 , n549 , n558 );
nor ( n560 , n559 , n9 );
and ( n561 , n560 , n184 );
nor ( n562 , t_6 , n561 );
not ( n563 , n5 );
or ( n564 , n562 , n563 );
nand ( n565 , n546 , n564 );
nor ( n566 , n2 , n8 );
nand ( n567 , n565 , n1 , n566 );
nand ( n568 , n531 , n567 );
and ( n569 , n3 , n568 );
not ( n570 , n1 );
nand ( n571 , n570 , n437 );
not ( n572 , n4 );
not ( n573 , n1 );
and ( n574 , n2 , n573 );
nand ( n575 , n572 , n574 );
or ( n576 , n5 , n575 );
not ( n577 , n538 );
not ( n578 , n577 );
and ( n579 , n10 , n11 );
nand ( n580 , n579 , n188 );
not ( n581 , n580 );
not ( n582 , n581 );
or ( n583 , n9 , n576 , n578 , n582 );
not ( n584 , n9 );
not ( n585 , n2 );
nand ( n586 , n1 , n585 );
nor ( n587 , n584 , n586 );
or ( n588 , n11 , n587 );
not ( n589 , n574 );
or ( n590 , n9 , n589 );
nand ( n591 , n590 , n11 );
not ( n592 , n210 );
not ( n593 , n592 );
nand ( n594 , n588 , n591 , n593 );
nor ( n595 , n594 , n578 , n100 );
not ( n596 , n5 );
not ( n597 , n184 );
not ( n598 , n1 );
nor ( n599 , n598 , n4 );
not ( n600 , n599 );
nor ( n601 , n600 , n329 );
not ( n602 , n601 );
and ( n603 , n202 , n321 );
and ( n604 , n185 , n603 );
not ( n605 , n2 );
nor ( n606 , n605 , n1 );
and ( n607 , n4 , n606 );
and ( n608 , n325 , n607 );
nand ( n609 , n1 , n7 );
nor ( n610 , n609 , n488 );
nor ( n611 , n608 , n610 );
not ( n612 , n17 );
nor ( n613 , n611 , n612 );
nand ( n614 , n604 , n613 );
nand ( n615 , n602 , n614 );
not ( n616 , n615 );
or ( n617 , n597 , n616 );
not ( n618 , n586 );
nand ( n619 , n10 , n618 );
or ( n620 , n350 , n619 );
nand ( n621 , n617 , n620 );
not ( n622 , n9 );
nand ( n623 , n621 , n622 );
not ( n624 , n4 );
not ( n625 , n624 );
not ( n626 , n230 );
nor ( n627 , n10 , n626 );
not ( n628 , n627 );
or ( n629 , n625 , n628 );
nand ( n630 , n428 , n80 , n505 );
nand ( n631 , n629 , n630 );
nand ( n632 , n587 , n631 );
and ( n633 , n623 , n632 );
nor ( n634 , n633 , n11 );
not ( n635 , n9 );
and ( n636 , n635 , n607 , n577 , n581 );
nor ( n637 , n634 , n636 );
nor ( n638 , n596 , n637 );
or ( n639 , n595 , n638 );
not ( n640 , n3 );
nand ( n641 , n639 , n640 );
and ( n642 , n583 , n641 );
nor ( n643 , n642 , n8 );
nor ( n644 , n569 , t_11 , n643 );
or ( n645 , n644 , n14 );
not ( n646 , n1 );
and ( n647 , n9 , n49 );
not ( n648 , n89 );
not ( n649 , n648 );
not ( n650 , n649 );
not ( n651 , n650 );
nand ( n652 , n646 , n647 , n651 );
or ( n653 , n652 , n364 , n460 );
not ( n654 , n174 );
or ( n655 , n15 , n654 , n140 );
not ( n656 , n9 );
and ( n657 , n113 , n125 );
and ( n658 , n36 , n89 );
nor ( n659 , n657 , n658 );
or ( n660 , n656 , n659 );
nand ( n661 , n655 , n660 );
not ( n662 , n3 );
and ( n663 , n606 , n662 );
and ( n664 , n661 , n49 , n663 );
nand ( n665 , n46 , n618 , n134 );
not ( n666 , n158 );
not ( n667 , n1 );
nand ( n668 , n666 , n667 , n136 , n90 );
and ( n669 , n665 , n668 );
not ( n670 , n3 );
nor ( n671 , n669 , n670 );
nor ( n672 , n664 , n671 );
or ( n673 , n151 , n672 );
nand ( n674 , n653 , n673 );
and ( n675 , n8 , n674 );
and ( n676 , n5 , n164 );
nor ( n677 , n675 , n676 );
nand ( n678 , n645 , n677 );
not ( n679 , n2 );
not ( n680 , n1 );
not ( n681 , n3 );
nor ( n682 , n7 , n17 );
and ( n683 , n157 , n682 );
nor ( n684 , n683 , n17 );
or ( n685 , n681 , n684 );
not ( n686 , n9 );
and ( n687 , n686 , n493 );
nor ( n688 , n687 , n359 );
or ( n689 , n688 , n3 , n17 );
nand ( n690 , n3 , n366 );
nand ( n691 , n689 , n690 );
nand ( n692 , n5 , n691 );
not ( n693 , n3 );
nand ( n694 , n693 , n17 );
nand ( n695 , n685 , n692 , n694 );
and ( n696 , n695 , n185 );
not ( n697 , n235 );
and ( n698 , n697 , n174 , n476 , n507 );
nor ( n699 , n696 , n698 );
or ( n700 , n699 , n15 );
nand ( n701 , n10 , n697 );
not ( n702 , n9 );
and ( n703 , n702 , n303 );
not ( n704 , n11 );
and ( n705 , n704 , n521 );
nor ( n706 , n703 , n705 );
or ( n707 , n701 , n706 );
not ( n708 , n11 );
and ( n709 , n697 , n708 , n537 );
not ( n710 , n233 );
nor ( n711 , n709 , n710 );
not ( n712 , n9 );
or ( n713 , n711 , n712 );
nand ( n714 , n707 , n713 );
and ( n715 , n299 , n714 );
not ( n716 , n626 );
and ( n717 , n697 , n716 , n9 , n115 );
nor ( n718 , n715 , n717 );
or ( n719 , n718 , n8 );
nand ( n720 , n700 , n719 );
and ( n721 , n680 , n720 );
not ( n722 , n372 );
not ( n723 , n11 );
not ( n724 , n10 );
nor ( n725 , n724 , n8 );
and ( n726 , n723 , n725 );
and ( n727 , n9 , n525 );
or ( n728 , n254 , n727 );
or ( n729 , n257 , n525 );
nand ( n730 , n728 , n729 );
and ( n731 , n722 , n726 , n1 , n730 );
nor ( n732 , n721 , n731 );
not ( n733 , n4 );
or ( n734 , n732 , n733 );
not ( n735 , n408 );
not ( n736 , n735 );
nand ( n737 , n345 , n736 );
nand ( n738 , n5 , n533 , n373 );
or ( n739 , n737 , n738 );
not ( n740 , n9 );
not ( n741 , n5 );
not ( n742 , n345 );
not ( n743 , n230 );
or ( n744 , n742 , n743 );
nand ( n745 , n3 , n216 );
not ( n746 , n745 );
not ( n747 , n1 );
nand ( n748 , n746 , n281 , n747 );
nand ( n749 , n744 , n748 );
not ( n750 , n749 );
or ( n751 , n741 , n750 );
not ( n752 , n5 );
and ( n753 , n752 , n345 );
nand ( n754 , n716 , n248 , n753 );
nand ( n755 , n751 , n754 );
not ( n756 , n755 );
or ( n757 , n740 , n756 );
and ( n758 , n5 , n257 );
not ( n759 , n401 );
not ( n760 , n759 );
nor ( n761 , n758 , n760 , n609 );
not ( n762 , n9 );
nand ( n763 , n350 , n761 , n17 , n762 );
nand ( n764 , n757 , n763 );
and ( n765 , n197 , n764 );
not ( n766 , n55 );
not ( n767 , n1 );
nor ( n768 , n767 , n143 );
and ( n769 , n766 , n768 );
not ( n770 , n1 );
and ( n771 , n770 , n297 );
nor ( n772 , n769 , n771 );
not ( n773 , n268 );
nor ( n774 , n772 , n197 , n773 );
nor ( n775 , n765 , n774 );
or ( n776 , n775 , n11 );
nand ( n777 , n1 , n3 );
not ( n778 , n777 );
not ( n779 , n477 );
not ( n780 , n779 );
not ( n781 , n780 );
not ( n782 , n781 );
nand ( n783 , n11 , n142 );
nor ( n784 , n266 , n783 );
nand ( n785 , n778 , n782 , n5 , n784 );
nand ( n786 , n776 , n785 );
and ( n787 , n476 , n786 );
not ( n788 , n473 );
not ( n789 , n788 );
and ( n790 , n753 , n789 , n682 );
not ( n791 , n3 );
nor ( n792 , n791 , n1 );
and ( n793 , n17 , n5 , n792 );
nor ( n794 , n790 , n793 );
nor ( n795 , n373 , n794 );
nor ( n796 , n787 , n795 );
or ( n797 , n796 , n4 );
nand ( n798 , n734 , n739 , n797 );
nand ( n799 , n679 , n798 );
not ( n800 , n1 );
nand ( n801 , n4 , n800 );
not ( n802 , n17 );
and ( n803 , n8 , n802 );
not ( n804 , n803 );
or ( n805 , n6 , n235 , n804 );
and ( n806 , n710 , n736 );
nand ( n807 , n197 , n806 );
or ( n808 , n17 , n414 );
nand ( n809 , n202 , n444 , n808 );
or ( n810 , n807 , n809 );
nand ( n811 , n805 , n810 );
nor ( n812 , n7 , n16 );
and ( n813 , n811 , n184 , n812 );
buf ( n814 , n592 );
not ( n815 , n814 );
and ( n816 , n806 , n815 , n303 );
nor ( n817 , n813 , n816 );
or ( n818 , n801 , n817 );
not ( n819 , n204 );
not ( n820 , n819 );
and ( n821 , n710 , n820 );
and ( n822 , n697 , n373 );
nor ( n823 , n821 , n822 );
nor ( n824 , n1 , n4 );
not ( n825 , n824 );
or ( n826 , n823 , n825 );
not ( n827 , n11 );
not ( n828 , n452 );
not ( n829 , n781 );
nand ( n830 , n828 , n260 , n5 , n829 );
or ( n831 , n830 , n325 , n12 );
not ( n832 , n9 );
nor ( n833 , n832 , n96 );
not ( n834 , n833 );
or ( n835 , n834 , n814 );
nand ( n836 , n831 , n835 );
nand ( n837 , n1 , n456 , n827 , n836 );
nand ( n838 , n818 , n826 , n837 );
nand ( n839 , n2 , n838 );
not ( n840 , n198 );
not ( n841 , n538 );
nand ( n842 , n840 , n453 , n841 );
or ( n843 , n35 , n842 );
not ( n844 , n4 );
nand ( n845 , n844 , t_7 );
nand ( n846 , n843 , n845 );
nand ( n847 , n736 , n320 , n345 , n846 );
nand ( n848 , n799 , n839 , n847 );
nand ( n849 , n848 , n151 );
not ( n850 , n1 );
nand ( n851 , n647 , n850 , n125 );
not ( n852 , n851 );
or ( n853 , n48 , n852 );
nand ( n854 , n853 , n14 , n119 );
not ( n855 , n4 );
and ( n856 , n1 , n14 );
not ( n857 , n856 );
or ( n858 , n2 , n47 );
not ( n859 , n537 );
not ( n860 , n859 );
not ( n861 , n783 );
and ( n862 , n860 , n861 );
not ( n863 , n12 );
nand ( n864 , n184 , n13 , n328 );
nand ( n865 , n15 , n279 , n449 );
nand ( n866 , n864 , n865 );
not ( n867 , n866 );
or ( n868 , n863 , n867 );
and ( n869 , n288 , n202 );
and ( n870 , n13 , n68 );
nor ( n871 , n869 , n870 );
not ( n872 , n523 );
nand ( n873 , n871 , n17 , n872 );
nand ( n874 , n868 , n873 );
not ( n875 , n11 );
and ( n876 , n874 , n875 );
nor ( n877 , n862 , n876 );
or ( n878 , n10 , n877 );
not ( n879 , n9 );
nand ( n880 , n879 , n174 );
or ( n881 , n15 , n880 );
nand ( n882 , n878 , n881 );
not ( n883 , n5 );
nor ( n884 , n883 , n6 );
nand ( n885 , n882 , n2 , n884 );
nand ( n886 , n858 , n885 );
not ( n887 , n886 );
or ( n888 , n857 , n887 );
not ( n889 , n5 );
and ( n890 , n889 , n574 );
nand ( n891 , n651 , n647 , n890 );
nand ( n892 , n888 , n891 );
nand ( n893 , n855 , n892 );
and ( n894 , n854 , n893 );
not ( n895 , n3 );
nor ( n896 , n894 , n895 );
not ( n897 , n9 );
nor ( n898 , n897 , n10 );
not ( n899 , n60 );
nand ( n900 , n898 , n651 , n56 , t_9 );
not ( n901 , n11 );
nand ( n902 , n901 , n14 );
nor ( n903 , n1 , n3 );
nand ( n904 , n49 , n5 , n903 );
nor ( n905 , n900 , n902 , n904 );
or ( n906 , n896 , n905 );
nand ( n907 , n906 , n8 );
nand ( n908 , n849 , n169 , n907 );
nor ( n909 , n7 , n15 );
not ( n910 , n589 );
not ( n911 , n910 );
nand ( n912 , n4 , n17 );
not ( n913 , n4 );
nand ( n914 , n913 , n414 );
nand ( n915 , n912 , n914 );
and ( n916 , n915 , n456 , n577 );
not ( n917 , n9 );
and ( n918 , n916 , n917 , n87 );
and ( n919 , n49 , n285 , n803 );
nor ( n920 , n918 , n919 );
nor ( n921 , n911 , n920 );
nand ( n922 , n5 , n909 , n185 , n921 );
not ( n923 , n922 );
not ( n924 , n3 );
not ( n925 , n5 );
not ( n926 , n17 );
nand ( n927 , n926 , n255 );
not ( n928 , n927 );
and ( n929 , n4 , n359 , n928 );
or ( n930 , n16 , n357 );
not ( n931 , n11 );
nor ( n932 , n931 , n185 );
nor ( n933 , n202 , n12 );
nand ( n934 , n932 , n725 , n933 );
nand ( n935 , n930 , n934 );
not ( n936 , n4 );
nor ( n937 , n936 , n15 );
not ( n938 , n17 );
and ( n939 , n935 , n937 , n938 );
and ( n940 , n188 , n12 , n726 );
nor ( n941 , n939 , n940 );
nor ( n942 , n941 , n9 );
nor ( n943 , n929 , n942 );
nor ( n944 , n925 , n943 );
and ( n945 , n924 , n944 );
not ( n946 , n924 );
and ( n947 , n4 , n476 );
nand ( n948 , n11 , n537 );
or ( n949 , n948 , n252 , n255 );
not ( n950 , n187 );
and ( n951 , n950 , n526 );
and ( n952 , n230 , n898 , n933 );
nor ( n953 , n951 , n952 );
or ( n954 , n953 , n11 );
nand ( n955 , n949 , n954 );
and ( n956 , n947 , n955 );
not ( n957 , n17 );
not ( n958 , n4 );
not ( n959 , n958 );
not ( n960 , n368 );
or ( n961 , n959 , n960 );
not ( n962 , n78 );
not ( n963 , n962 );
not ( n964 , n963 );
nand ( n965 , n964 , n947 , n507 );
nand ( n966 , n961 , n965 );
and ( n967 , n957 , n966 );
nor ( n968 , n956 , n967 );
or ( n969 , n968 , n5 );
nand ( n970 , n937 , n453 );
nand ( n971 , n969 , n970 );
and ( n972 , n946 , n971 );
nor ( n973 , n945 , n972 );
not ( n974 , n973 );
not ( n975 , n1 );
nand ( n976 , n974 , n975 );
not ( n977 , n11 );
not ( n978 , n9 );
nand ( n979 , n12 , n978 );
or ( n980 , n281 , n979 );
not ( n981 , n5 );
nand ( n982 , n9 , n981 , n216 );
nand ( n983 , n980 , n982 );
nand ( n984 , n4 , n983 );
nor ( n985 , n5 , n9 );
nand ( n986 , n12 , n985 );
nand ( n987 , n306 , n524 );
and ( n988 , n984 , n986 , n987 );
or ( n989 , n988 , n3 );
nor ( n990 , n133 , n9 );
not ( n991 , n17 );
and ( n992 , n12 , n991 );
and ( n993 , n990 , n992 , n260 );
nor ( n994 , n993 , n833 );
not ( n995 , n3 );
or ( n996 , n994 , n995 );
nand ( n997 , n989 , n996 );
and ( n998 , n16 , n997 );
not ( n999 , n987 );
not ( n1000 , n3 );
nand ( n1001 , n999 , n1000 );
not ( n1002 , n212 );
not ( n1003 , n218 );
or ( n1004 , n1002 , n1003 );
nand ( n1005 , n1004 , n979 );
not ( n1006 , n5 );
nand ( n1007 , n3 , n211 );
nand ( n1008 , n1005 , n1006 , n1007 );
and ( n1009 , n1001 , n1008 );
nor ( n1010 , n1009 , n184 );
nor ( n1011 , n998 , n1010 );
or ( n1012 , n1011 , n197 );
not ( n1013 , n3 );
and ( n1014 , n1013 , n134 );
nor ( n1015 , n1014 , n113 );
nand ( n1016 , n244 , n260 , n248 , n451 );
or ( n1017 , n1015 , n1016 );
nand ( n1018 , n1012 , n1017 );
nand ( n1019 , n977 , n1018 );
and ( n1020 , n5 , n285 );
not ( n1021 , n964 );
not ( n1022 , n1021 );
and ( n1023 , n1020 , n267 , n1022 );
nand ( n1024 , n1023 , n291 , n782 );
and ( n1025 , n1019 , n1024 );
not ( n1026 , n1 );
nor ( n1027 , n1025 , n1026 );
nor ( n1028 , n15 , n16 );
not ( n1029 , n17 );
nor ( n1030 , n1029 , n11 );
not ( n1031 , n1030 );
not ( n1032 , n244 );
nor ( n1033 , n1031 , n163 , n1032 );
not ( n1034 , n578 );
and ( n1035 , n1028 , n1033 , n5 , n1034 );
or ( n1036 , n1027 , n1035 );
nand ( n1037 , n1036 , n476 );
and ( n1038 , n976 , n1037 );
nor ( n1039 , n1038 , n2 );
nand ( n1040 , n3 , n574 );
nor ( n1041 , n1040 , n4 , n7 );
nand ( n1042 , n17 , n1041 );
not ( n1043 , n1042 );
and ( n1044 , n87 , n410 , n1043 );
not ( n1045 , n162 );
nand ( n1046 , n1045 , n9 , n176 );
nor ( n1047 , n8 , n11 );
not ( n1048 , n1047 );
or ( n1049 , n1046 , n3 , n1048 );
not ( n1050 , n2 );
nor ( n1051 , n8 , n1050 , n252 );
and ( n1052 , n11 , n841 , n1051 );
nor ( n1053 , n1052 , n3 );
or ( n1054 , n825 , n1053 );
nand ( n1055 , n1049 , n1054 );
and ( n1056 , n373 , n1055 );
nor ( n1057 , n1044 , n1056 );
nor ( n1058 , n5 , n1057 );
nor ( n1059 , n923 , n1039 , n1058 );
or ( n1060 , n14 , n1059 );
not ( n1061 , n472 );
and ( n1062 , n9 , n1061 );
not ( n1063 , n79 );
nand ( n1064 , n12 , n69 );
and ( n1065 , n1063 , n1064 );
not ( n1066 , n2 );
nand ( n1067 , n1066 , n5 );
nor ( n1068 , n1065 , n1067 );
and ( n1069 , n1068 , n197 , n547 );
nor ( n1070 , n5 , n103 );
nor ( n1071 , n1069 , n1070 );
or ( n1072 , n151 , n353 , n1071 );
or ( n1073 , n151 , n108 );
nand ( n1074 , n1073 , n38 );
not ( n1075 , n5 );
and ( n1076 , n1074 , n1075 , n125 );
nor ( n1077 , n13 , n108 , n902 );
nand ( n1078 , n992 , n1077 , n5 , n197 );
nor ( n1079 , n650 , n1078 );
nor ( n1080 , n1076 , n1079 );
or ( n1081 , n4 , n1080 );
nand ( n1082 , n1072 , n1081 );
and ( n1083 , n1062 , n1082 );
not ( n1084 , n4 );
nor ( n1085 , n2 , n3 );
and ( n1086 , n1084 , n1085 );
nor ( n1087 , n1083 , n1086 );
or ( n1088 , n1 , n1087 );
not ( n1089 , n5 );
nand ( n1090 , n1089 , n164 );
nand ( n1091 , n1060 , n1088 , n1090 );
not ( n1092 , n11 );
not ( n1093 , n3 );
not ( n1094 , n17 );
and ( n1095 , n1094 , n359 );
not ( n1096 , n1 );
nand ( n1097 , n1095 , n90 , n1096 );
not ( n1098 , n613 );
nand ( n1099 , n1097 , n1098 );
and ( n1100 , n1099 , n604 );
nor ( n1101 , n1100 , n601 );
or ( n1102 , n1101 , n15 );
nand ( n1103 , n1102 , n620 );
and ( n1104 , n1093 , n1103 );
not ( n1105 , n4 );
not ( n1106 , n1 );
not ( n1107 , n260 );
or ( n1108 , n551 , n1106 , n1107 );
or ( n1109 , n592 , n1 );
nand ( n1110 , n1108 , n1109 );
and ( n1111 , n1105 , n39 , n1110 );
nor ( n1112 , n1104 , n1111 );
or ( n1113 , n1112 , n9 );
not ( n1114 , n9 );
nor ( n1115 , n1114 , n2 );
not ( n1116 , n1115 );
and ( n1117 , n346 , n627 );
nand ( n1118 , n176 , n188 );
and ( n1119 , n1 , n1118 );
and ( n1120 , n283 , n548 );
nor ( n1121 , n1120 , n1 );
nor ( n1122 , n1119 , n745 , n1121 );
nor ( n1123 , n1117 , n1122 );
or ( n1124 , n1116 , n1123 );
nand ( n1125 , n1113 , n1124 );
and ( n1126 , n1092 , n1125 );
and ( n1127 , n4 , n903 );
not ( n1128 , n1127 );
and ( n1129 , n2 , n390 , n303 );
nor ( n1130 , n1129 , n1115 );
or ( n1131 , n437 , n1130 );
not ( n1132 , n2 );
nor ( n1133 , n9 , n12 );
not ( n1134 , n864 );
nand ( n1135 , n1132 , n579 , n1133 , n1134 );
nand ( n1136 , n1131 , n1135 );
not ( n1137 , n1136 );
or ( n1138 , n1128 , n1137 );
nor ( n1139 , n10 , n38 );
not ( n1140 , n9 );
nand ( n1141 , n599 , n1139 , n1140 , n784 );
nand ( n1142 , n1138 , n1141 );
nor ( n1143 , n1126 , n1142 );
or ( n1144 , n1143 , n8 );
not ( n1145 , n2 );
and ( n1146 , n46 , n803 );
nor ( n1147 , n1146 , n17 );
or ( n1148 , n364 , n1147 );
not ( n1149 , n17 );
not ( n1150 , n1149 );
not ( n1151 , n690 );
or ( n1152 , n1150 , n1151 );
nand ( n1153 , n1152 , n4 );
nand ( n1154 , n1148 , n1153 );
and ( n1155 , n1145 , n1154 );
not ( n1156 , n3 );
nand ( n1157 , n9 , n118 );
or ( n1158 , n367 , n1157 );
not ( n1159 , n17 );
not ( n1160 , n59 );
not ( n1161 , n1160 );
not ( n1162 , n1161 );
not ( n1163 , n1162 );
not ( n1164 , n1163 );
or ( n1165 , n1159 , n1164 );
nand ( n1166 , n1158 , n1165 );
and ( n1167 , n1156 , n1166 );
nor ( n1168 , n1155 , n1167 );
or ( n1169 , n571 , n1168 );
nand ( n1170 , n1144 , n1169 );
and ( n1171 , n151 , n1170 );
and ( n1172 , n8 , n14 );
not ( n1173 , n1172 );
not ( n1174 , n4 );
nand ( n1175 , n3 , n618 );
or ( n1176 , n1174 , n47 , n1175 );
not ( n1177 , n1021 );
not ( n1178 , n17 );
nand ( n1179 , n1178 , n303 );
not ( n1180 , n1179 );
and ( n1181 , n1180 , n778 , n1161 );
not ( n1182 , n11 );
and ( n1183 , n872 , n479 );
not ( n1184 , n17 );
and ( n1185 , n1184 , n267 );
nor ( n1186 , n1183 , n1185 );
or ( n1187 , n364 , n162 , n1186 );
not ( n1188 , n9 );
nor ( n1189 , n1188 , n1 , n912 );
nand ( n1190 , n13 , n53 );
nand ( n1191 , n1189 , n1085 , n1190 );
nand ( n1192 , n1187 , n1191 );
and ( n1193 , n1182 , n1192 );
nor ( n1194 , n1181 , n1193 );
or ( n1195 , n1194 , n10 );
not ( n1196 , n3 );
not ( n1197 , n1 );
not ( n1198 , n17 );
or ( n1199 , n1198 , n1157 );
nand ( n1200 , n1199 , n1160 );
and ( n1201 , n1197 , n1200 );
nor ( n1202 , n9 , n17 );
nor ( n1203 , n4 , n162 );
and ( n1204 , n1202 , n1203 );
nor ( n1205 , n1201 , n1204 );
or ( n1206 , n1196 , n1205 );
nand ( n1207 , n1195 , n1206 );
and ( n1208 , n1177 , n1207 );
not ( n1209 , n3 );
nor ( n1210 , n648 , n1209 );
nor ( n1211 , n10 , n1031 );
nand ( n1212 , n1 , n9 );
not ( n1213 , n1212 );
and ( n1214 , n1211 , n1213 , n56 );
not ( n1215 , n1 );
nor ( n1216 , n1214 , n1215 );
or ( n1217 , n1162 , n1216 );
or ( n1218 , n211 , n154 );
nand ( n1219 , n1217 , n1218 );
and ( n1220 , n1210 , n1219 );
nor ( n1221 , n1208 , n1220 );
or ( n1222 , n1221 , n6 );
nand ( n1223 , n1176 , n1222 );
not ( n1224 , n1223 );
or ( n1225 , n1173 , n1224 );
not ( n1226 , n164 );
nand ( n1227 , n1225 , n1226 );
nor ( n1228 , n1171 , n1227 );
not ( n1229 , n5 );
or ( n1230 , n1228 , n1229 );
or ( n1231 , n151 , n47 , n1175 );
nand ( n1232 , n49 , n574 );
and ( n1233 , n14 , n144 );
and ( n1234 , n9 , n1210 );
nor ( n1235 , n1233 , n1234 );
or ( n1236 , n1232 , n1235 );
nand ( n1237 , n1231 , n1236 );
not ( n1238 , n4 );
and ( n1239 , n1237 , n8 , n1238 );
not ( n1240 , n581 );
not ( n1241 , n841 );
or ( n1242 , n9 , n1240 , n1241 , n575 );
not ( n1243 , n11 );
not ( n1244 , n2 );
or ( n1245 , n1118 , n1244 );
not ( n1246 , n2 );
nand ( n1247 , n248 , n548 , n1246 , n716 );
nand ( n1248 , n1245 , n1247 );
nand ( n1249 , n345 , n1248 );
and ( n1250 , n9 , n1249 );
not ( n1251 , n9 );
not ( n1252 , n350 );
not ( n1253 , n914 );
nand ( n1254 , n325 , n663 , n1253 );
not ( n1255 , n609 );
not ( n1256 , n2 );
or ( n1257 , n1256 , n191 );
not ( n1258 , n488 );
nand ( n1259 , n1257 , n1258 );
nand ( n1260 , n1255 , n17 , n1259 );
nand ( n1261 , n1254 , n1260 );
not ( n1262 , n1261 );
or ( n1263 , n1252 , n1262 );
nand ( n1264 , n1263 , n1042 );
and ( n1265 , n603 , n1264 );
nor ( n1266 , n592 , n586 , n353 );
nor ( n1267 , n1265 , n1266 );
and ( n1268 , n1251 , n1267 );
nor ( n1269 , n1250 , n1268 );
nand ( n1270 , n1243 , n1269 );
and ( n1271 , n1242 , n1270 );
nor ( n1272 , n1271 , n8 );
nor ( n1273 , n4 , n6 );
nand ( n1274 , n1 , n1085 , n1273 , n928 );
nor ( n1275 , n1274 , n476 , n7 );
or ( n1276 , n437 , n1164 );
nand ( n1277 , n49 , n118 , n909 , n342 );
nand ( n1278 , n1276 , n1277 );
and ( n1279 , n792 , n1278 );
nor ( n1280 , n1272 , n1275 , n1279 );
nor ( n1281 , n1280 , n14 );
nor ( n1282 , n1239 , n1281 );
or ( n1283 , n5 , n1282 );
nand ( n1284 , n1230 , n1283 );
not ( n1285 , n576 );
and ( n1286 , n151 , n188 );
nand ( n1287 , n1285 , n579 , n410 , n1286 );
not ( n1288 , n3 );
nor ( n1289 , n5 , n211 , n341 );
and ( n1290 , n14 , n15 );
and ( n1291 , n1289 , n1290 , n789 );
not ( n1292 , n4 );
not ( n1293 , n5 );
nor ( n1294 , n1293 , n86 );
nand ( n1295 , n1294 , n325 , n255 , n808 );
and ( n1296 , n580 , n1295 );
or ( n1297 , n1292 , n1296 );
not ( n1298 , n306 );
not ( n1299 , n339 );
nand ( n1300 , n197 , n320 , n359 , n1299 );
or ( n1301 , n1298 , n1300 );
nand ( n1302 , n1297 , n1301 );
and ( n1303 , n410 , n1302 );
not ( n1304 , n4 );
and ( n1305 , n184 , n451 );
and ( n1306 , n1304 , n1305 );
nor ( n1307 , n1303 , n1306 );
nor ( n1308 , n14 , n1307 );
nor ( n1309 , n1291 , n1308 );
or ( n1310 , n911 , n1309 );
and ( n1311 , n151 , n4 , n820 );
not ( n1312 , n1298 );
nor ( n1313 , n1311 , n1312 );
or ( n1314 , n154 , n1313 );
nor ( n1315 , n12 , n1048 );
or ( n1316 , n197 , n1157 , n394 );
not ( n1317 , n1067 );
or ( n1318 , n325 , n779 , n819 );
nand ( n1319 , n9 , n10 );
or ( n1320 , n1319 , n350 );
nand ( n1321 , n1318 , n1320 );
and ( n1322 , n202 , n1317 , n1321 );
not ( n1323 , n184 );
nor ( n1324 , n1323 , n389 , n173 , n460 );
nor ( n1325 , n1322 , n1324 );
or ( n1326 , n4 , n1325 );
nand ( n1327 , n1316 , n1326 );
nand ( n1328 , n1315 , n151 , n1 , n1327 );
nand ( n1329 , n1310 , n1314 , n1328 );
nand ( n1330 , n1288 , n1329 );
not ( n1331 , n140 );
not ( n1332 , n17 );
or ( n1333 , n1 , n14 );
not ( n1334 , n1333 );
and ( n1335 , n1332 , n1334 );
nor ( n1336 , n1335 , n856 );
or ( n1337 , n43 , n1336 );
nand ( n1338 , n1337 , n851 );
and ( n1339 , n8 , n1338 );
or ( n1340 , n820 , n1095 );
not ( n1341 , n1 );
nand ( n1342 , n1340 , n1341 );
nand ( n1343 , n1 , n476 );
not ( n1344 , n1343 );
nand ( n1345 , n1344 , n533 , n537 , n535 );
and ( n1346 , n1342 , n1345 );
nor ( n1347 , n1346 , n14 );
nor ( n1348 , n1339 , n1347 );
or ( n1349 , n2 , n1348 );
not ( n1350 , n1333 );
not ( n1351 , n2 );
or ( n1352 , n7 , n1351 , n419 );
nand ( n1353 , n1352 , n351 );
nand ( n1354 , n1350 , n1353 );
nand ( n1355 , n1349 , n1354 );
and ( n1356 , n1331 , n1355 );
not ( n1357 , n151 );
nor ( n1358 , n1 , n927 );
not ( n1359 , n1358 );
or ( n1360 , n1357 , n1359 );
not ( n1361 , n856 );
nand ( n1362 , n1360 , n1361 );
nand ( n1363 , n493 , n1362 );
not ( n1364 , n1343 );
and ( n1365 , n872 , n950 );
nor ( n1366 , n979 , n143 );
nor ( n1367 , n1365 , n1366 );
or ( n1368 , n1367 , n13 , n534 );
nand ( n1369 , n11 , n12 , n780 , n1134 );
nand ( n1370 , n1368 , n1369 );
nand ( n1371 , n1364 , n151 , n1370 );
and ( n1372 , n1363 , n1371 );
nor ( n1373 , n1372 , n2 , n1298 );
nor ( n1374 , n1356 , n1373 );
not ( n1375 , n2 );
not ( n1376 , n1312 );
nor ( n1377 , n1375 , n1376 );
not ( n1378 , n1333 );
nand ( n1379 , n1378 , n16 );
nand ( n1380 , n14 , n473 );
or ( n1381 , n16 , n1380 , n1216 );
nand ( n1382 , n1381 , n1333 );
nand ( n1383 , n15 , n1382 );
not ( n1384 , n1 );
nand ( n1385 , n151 , n44 , n340 );
nand ( n1386 , n14 , n16 );
not ( n1387 , n1386 );
not ( n1388 , n197 );
or ( n1389 , n11 , n1186 );
nand ( n1390 , n1389 , n1179 );
not ( n1391 , n1390 );
or ( n1392 , n1388 , n1391 );
not ( n1393 , n1202 );
nand ( n1394 , n1392 , n1393 );
nand ( n1395 , n49 , n1387 , n1394 );
and ( n1396 , n1385 , n1395 );
nor ( n1397 , n1396 , n476 );
or ( n1398 , n1384 , n1397 );
not ( n1399 , n1 );
nor ( n1400 , n7 , n14 );
nand ( n1401 , n1400 , n338 );
nand ( n1402 , n1386 , n1401 );
and ( n1403 , n473 , n1402 );
not ( n1404 , n448 );
nor ( n1405 , n7 , n8 );
nand ( n1406 , n1404 , n1405 , n477 );
or ( n1407 , n13 , n14 );
nor ( n1408 , n1406 , n443 , n1407 );
nor ( n1409 , n1403 , n1408 );
and ( n1410 , n1399 , n1409 );
nor ( n1411 , n1410 , n15 );
nand ( n1412 , n1398 , n1411 );
nand ( n1413 , n1379 , n1383 , n1412 );
nand ( n1414 , n1377 , n1413 );
not ( n1415 , n911 );
and ( n1416 , n185 , n1290 , n473 );
not ( n1417 , n1409 );
and ( n1418 , n184 , n1417 );
nor ( n1419 , n1416 , n1418 );
not ( n1420 , n1419 );
and ( n1421 , n1415 , n1420 );
not ( n1422 , n2 );
nor ( n1423 , n1 , n9 );
and ( n1424 , n11 , n1423 , n759 );
not ( n1425 , n11 );
and ( n1426 , n1425 , n1213 );
nor ( n1427 , n1424 , n1426 );
or ( n1428 , n255 , n1427 );
not ( n1429 , n11 );
not ( n1430 , n9 );
nand ( n1431 , n1429 , n1430 , n768 );
nand ( n1432 , n1428 , n1431 );
and ( n1433 , n725 , n1432 );
and ( n1434 , n359 , n1358 );
nor ( n1435 , n1433 , n1434 );
or ( n1436 , n14 , n1435 );
nand ( n1437 , n1436 , n1363 );
and ( n1438 , n1422 , n1437 );
nor ( n1439 , n1421 , n1438 );
or ( n1440 , n5 , n1439 );
not ( n1441 , n5 );
nor ( n1442 , n476 , n1232 );
and ( n1443 , n14 , n89 , n1442 );
not ( n1444 , n1442 );
not ( n1445 , n1402 );
or ( n1446 , n1444 , n1445 );
not ( n1447 , n9 );
and ( n1448 , n1447 , n566 );
or ( n1449 , n13 , n198 , n450 );
not ( n1450 , n1 );
or ( n1451 , n1450 , n329 );
nand ( n1452 , n1449 , n1451 );
nand ( n1453 , n1448 , n151 , n444 , n1452 );
nand ( n1454 , n1446 , n1453 );
and ( n1455 , n184 , n1454 );
nor ( n1456 , n1443 , n1455 );
or ( n1457 , n1441 , n1456 );
not ( n1458 , n2 );
nor ( n1459 , n1 , n819 );
and ( n1460 , n1458 , n1459 );
nand ( n1461 , n151 , n1460 );
nand ( n1462 , n1440 , n1457 , n1461 );
nand ( n1463 , n4 , n1462 );
nand ( n1464 , n1374 , n1414 , n1463 );
nand ( n1465 , n3 , n1464 );
nand ( n1466 , n1287 , n1330 , n1465 );
not ( n1467 , n2 );
not ( n1468 , n1467 );
nand ( n1469 , n1030 , n477 , n1405 , n759 );
nand ( n1470 , n255 , n1469 );
and ( n1471 , n792 , n1331 , n1470 );
not ( n1472 , n735 );
and ( n1473 , n229 , n1472 );
and ( n1474 , n197 , n480 , n1473 );
and ( n1475 , n6 , n803 , n1020 );
nor ( n1476 , n1474 , n1475 );
or ( n1477 , n609 , n1476 );
not ( n1478 , n1 );
or ( n1479 , n476 , n257 );
nand ( n1480 , n1473 , n321 , n547 );
nand ( n1481 , n1479 , n1480 );
nand ( n1482 , n1478 , n682 , n1273 , n1481 );
nand ( n1483 , n1477 , n1482 );
and ( n1484 , n437 , n1483 );
nor ( n1485 , n1471 , n1484 );
not ( n1486 , n1485 );
and ( n1487 , n1468 , n1486 );
not ( n1488 , n321 );
not ( n1489 , n716 );
or ( n1490 , n1488 , n1489 );
nand ( n1491 , n1490 , n9 );
not ( n1492 , n9 );
and ( n1493 , n1492 , n814 );
not ( n1494 , n5 );
nand ( n1495 , n476 , n1494 , n599 );
nor ( n1496 , n1493 , n11 , n1495 );
and ( n1497 , n1491 , n1496 );
nand ( n1498 , n10 , n399 );
nor ( n1499 , n11 , n17 );
not ( n1500 , n1499 );
or ( n1501 , n1021 , n1498 , n1500 );
not ( n1502 , n185 );
not ( n1503 , n49 );
not ( n1504 , n682 );
or ( n1505 , n1503 , n1504 );
or ( n1506 , n9 , n1202 );
nand ( n1507 , n1506 , n366 );
nand ( n1508 , n1505 , n1507 );
not ( n1509 , n1508 );
or ( n1510 , n1502 , n1509 );
not ( n1511 , n1498 );
nand ( n1512 , n1511 , n933 , n172 , n11 );
nand ( n1513 , n1510 , n1512 );
and ( n1514 , n1513 , n184 );
nor ( n1515 , n8 , n255 , n313 );
nor ( n1516 , n1514 , n1515 );
or ( n1517 , n1516 , n1 );
nand ( n1518 , n1501 , n1517 );
nand ( n1519 , n5 , n1518 );
not ( n1520 , n1 );
nor ( n1521 , n1520 , n5 );
or ( n1522 , n592 , n727 );
nand ( n1523 , n1522 , n1016 );
nand ( n1524 , n1047 , n1521 , n1523 );
and ( n1525 , n1519 , n1524 );
not ( n1526 , n4 );
nor ( n1527 , n1525 , n1526 );
nor ( n1528 , n1497 , n1527 );
or ( n1529 , n3 , n1528 );
not ( n1530 , n11 );
nand ( n1531 , n990 , n962 , n992 );
nand ( n1532 , n12 , n35 );
nand ( n1533 , n248 , n111 );
nand ( n1534 , n535 , n1532 , n1533 );
nand ( n1535 , n1531 , n1534 );
nand ( n1536 , n10 , n1535 );
not ( n1537 , n5 );
and ( n1538 , n1537 , n175 );
not ( n1539 , n779 );
nand ( n1540 , n1538 , n7 , n451 , n1539 );
and ( n1541 , n1536 , n1540 );
not ( n1542 , n3 );
nor ( n1543 , n1541 , n1542 );
not ( n1544 , n5 );
nand ( n1545 , n1544 , n548 , n175 );
nor ( n1546 , n1545 , n461 , n452 );
or ( n1547 , n1543 , n1546 );
nand ( n1548 , n1547 , n202 );
nand ( n1549 , n181 , n1548 );
and ( n1550 , n1530 , n1549 );
not ( n1551 , n1024 );
nor ( n1552 , n1550 , n1551 );
or ( n1553 , n1552 , n1343 );
nand ( n1554 , n36 , n1459 );
nand ( n1555 , n1529 , n1553 , n1554 );
not ( n1556 , n2 );
and ( n1557 , n1555 , n1556 );
nor ( n1558 , n1487 , n1557 );
or ( n1559 , n14 , n1558 );
not ( n1560 , n1 );
not ( n1561 , n1258 );
nand ( n1562 , n42 , n1172 );
not ( n1563 , n1562 );
and ( n1564 , n1561 , n1563 );
nor ( n1565 , n1564 , n90 );
or ( n1566 , n1560 , n1565 );
not ( n1567 , n1 );
not ( n1568 , n90 );
nor ( n1569 , n6 , n1568 );
nand ( n1570 , n14 , n136 );
not ( n1571 , n1570 );
nand ( n1572 , n8 , n1567 , n1569 , n1571 );
nand ( n1573 , n1566 , n1572 );
and ( n1574 , n3 , n1573 );
nor ( n1575 , n1574 , n166 );
or ( n1576 , n5 , n1575 );
not ( n1577 , n902 );
and ( n1578 , n118 , n1190 , n123 );
and ( n1579 , n509 , n899 );
not ( n1580 , n56 );
nor ( n1581 , n1579 , n650 , n1580 );
nor ( n1582 , n1578 , n1581 );
nor ( n1583 , n904 , n1582 );
nand ( n1584 , n898 , n1577 , n8 , n1583 );
nand ( n1585 , n1559 , n1576 , n1584 );
not ( n1586 , n3 );
and ( n1587 , n7 , n1521 , n1047 );
and ( n1588 , n1587 , n782 , n577 );
not ( n1589 , n1 );
nor ( n1590 , n1588 , n1589 );
or ( n1591 , n970 , n1590 );
not ( n1592 , n9 );
not ( n1593 , n1495 );
nand ( n1594 , n1592 , n533 , n422 , n1593 );
nand ( n1595 , n1591 , n1594 );
and ( n1596 , n151 , n1586 , n1595 );
not ( n1597 , n1 );
nor ( n1598 , n1597 , n111 , n1562 );
and ( n1599 , n3 , n1598 );
nor ( n1600 , n1596 , n1599 );
not ( n1601 , n1600 );
not ( n1602 , n5 );
not ( n1603 , n9 );
not ( n1604 , n1603 );
not ( n1605 , n1 );
nand ( n1606 , n1605 , n933 );
and ( n1607 , n11 , n1606 );
nor ( n1608 , n1607 , n193 );
not ( n1609 , n4 );
nand ( n1610 , n1609 , n778 );
not ( n1611 , n1610 );
not ( n1612 , n10 );
not ( n1613 , n547 );
or ( n1614 , n1612 , n1613 );
nand ( n1615 , n13 , n11 , n197 );
nand ( n1616 , n1614 , n1615 );
and ( n1617 , n12 , n1611 , n1616 );
nor ( n1618 , n1608 , n1617 );
or ( n1619 , n1618 , n510 );
nand ( n1620 , n366 , n1127 );
or ( n1621 , n16 , n1620 );
nand ( n1622 , n1619 , n1621 );
not ( n1623 , n1622 );
or ( n1624 , n1604 , n1623 );
or ( n1625 , n364 , n367 );
or ( n1626 , n353 , n360 );
nand ( n1627 , n1625 , n1626 );
not ( n1628 , n1 );
nand ( n1629 , n1627 , n1628 , n185 );
nand ( n1630 , n1624 , n1629 );
not ( n1631 , n17 );
and ( n1632 , n1630 , n1631 );
nor ( n1633 , n1 , n452 );
and ( n1634 , n4 , n1633 );
nor ( n1635 , n1632 , n1634 );
or ( n1636 , n1635 , n15 );
not ( n1637 , n9 );
not ( n1638 , n1637 );
not ( n1639 , n903 );
or ( n1640 , n1638 , n1639 );
nand ( n1641 , n12 , n778 , n279 );
nand ( n1642 , n1640 , n1641 );
nand ( n1643 , n947 , n533 , n722 , n1642 );
nand ( n1644 , n1636 , n1643 );
and ( n1645 , n151 , n1644 );
or ( n1646 , n45 , n1610 );
and ( n1647 , n898 , n1030 );
or ( n1648 , n137 , n53 );
not ( n1649 , n963 );
not ( n1650 , n1064 );
or ( n1651 , n1649 , n1650 );
nand ( n1652 , n1651 , n202 );
nand ( n1653 , n1648 , n1652 );
nand ( n1654 , n1647 , n49 , n1127 , n1653 );
nand ( n1655 , n1646 , n1654 );
and ( n1656 , n1172 , n1655 );
nor ( n1657 , n1645 , n1656 );
nor ( n1658 , n1602 , n1657 );
nor ( n1659 , n1601 , n1658 );
or ( n1660 , n2 , n1659 );
not ( n1661 , n4 );
and ( n1662 , n1661 , n1172 , n337 );
not ( n1663 , n654 );
and ( n1664 , n1662 , n1663 , n663 );
not ( n1665 , n17 );
and ( n1666 , n4 , n1568 );
nor ( n1667 , n1666 , n950 );
and ( n1668 , n1667 , n7 , n345 );
nor ( n1669 , n1668 , n1041 );
or ( n1670 , n1665 , n86 , n1669 );
not ( n1671 , n11 );
or ( n1672 , n814 , n1671 , n575 );
nand ( n1673 , n1670 , n1672 );
and ( n1674 , n410 , n1673 );
not ( n1675 , n1040 );
or ( n1676 , n4 , n351 );
nand ( n1677 , n4 , n337 , n803 , n812 );
nand ( n1678 , n1676 , n1677 );
and ( n1679 , n1675 , n1678 );
nor ( n1680 , n1674 , n1679 );
nor ( n1681 , n14 , n1680 );
nor ( n1682 , n1664 , n1681 );
or ( n1683 , n5 , n1682 );
not ( n1684 , n4 );
not ( n1685 , n17 );
nor ( n1686 , n1685 , n14 );
and ( n1687 , n184 , n1686 );
nor ( n1688 , n1 , n7 );
and ( n1689 , n1687 , n1688 , n398 );
and ( n1690 , n248 , n322 );
and ( n1691 , n1689 , n478 , n1690 );
nor ( n1692 , n1691 , n778 );
or ( n1693 , n1684 , n1692 );
not ( n1694 , n138 );
nand ( n1695 , n898 , n102 , n398 , n56 );
nand ( n1696 , n1694 , n1695 );
nand ( n1697 , n49 , n824 , n1172 , n1696 );
nand ( n1698 , n1693 , n1697 );
nand ( n1699 , n5 , n2 , n1698 );
nand ( n1700 , n1660 , n1683 , n1699 );
not ( n1701 , n14 );
not ( n1702 , n1405 );
nor ( n1703 , n1702 , n445 , n575 , n1107 );
not ( n1704 , n9 );
and ( n1705 , n1703 , n1704 , n455 );
or ( n1706 , n17 , n1095 );
nand ( n1707 , n1706 , n824 , n351 );
not ( n1708 , n4 );
not ( n1709 , n1708 );
not ( n1710 , n1426 );
or ( n1711 , n1709 , n1710 );
nand ( n1712 , n11 , n4 , n1423 );
nand ( n1713 , n1711 , n1712 );
nand ( n1714 , n248 , n725 , n393 , n1713 );
and ( n1715 , n1707 , n1714 );
nor ( n1716 , n1715 , n2 );
nor ( n1717 , n1705 , n1716 );
not ( n1718 , n1717 );
and ( n1719 , n1701 , n1718 );
not ( n1720 , n1 );
not ( n1721 , n184 );
not ( n1722 , n1401 );
not ( n1723 , n1722 );
or ( n1724 , n1721 , n1723 );
nand ( n1725 , n1724 , n1570 );
nand ( n1726 , n1720 , n1569 , n1725 );
or ( n1727 , n151 , n118 );
not ( n1728 , n1161 );
not ( n1729 , n928 );
or ( n1730 , n1728 , n1729 );
nand ( n1731 , n1730 , n151 );
nand ( n1732 , n1727 , n46 , n1731 );
not ( n1733 , n1732 );
nor ( n1734 , n151 , n6 );
nand ( n1735 , n1734 , n1163 , n882 );
not ( n1736 , n1735 );
or ( n1737 , n1733 , n1736 );
nand ( n1738 , n1737 , n1 );
nand ( n1739 , n1726 , n1738 );
and ( n1740 , n8 , n1739 );
nor ( n1741 , n1719 , n1740 );
or ( n1742 , n257 , n1741 );
and ( n1743 , n582 , n1300 );
not ( n1744 , n1407 );
nand ( n1745 , n1744 , n663 );
nor ( n1746 , n1743 , n1745 );
and ( n1747 , n1746 , n476 , n1133 );
not ( n1748 , n1 );
nor ( n1749 , n14 , n15 );
nand ( n1750 , n1748 , n342 , n1749 , n368 );
not ( n1751 , n1562 );
not ( n1752 , n1498 );
not ( n1753 , n11 );
nand ( n1754 , n1752 , n172 , n1749 , n1753 );
not ( n1755 , n1754 );
or ( n1756 , n1751 , n1755 );
nand ( n1757 , n1756 , n1 );
and ( n1758 , n1750 , n1757 );
nor ( n1759 , n1758 , n38 );
nor ( n1760 , n1747 , n1759 );
or ( n1761 , n100 , n1760 );
not ( n1762 , n1 );
not ( n1763 , n17 );
nor ( n1764 , n6 , n9 );
and ( n1765 , n1764 , n185 , n2 , n909 );
nand ( n1766 , n1762 , n1763 , n87 , n1765 );
and ( n1767 , n1766 , n594 );
not ( n1768 , n947 );
nor ( n1769 , n1767 , n1768 );
and ( n1770 , n1034 , n1769 );
and ( n1771 , n1163 , n1459 );
nor ( n1772 , n1770 , n1771 );
or ( n1773 , n14 , n1772 );
nand ( n1774 , n1773 , n165 );
and ( n1775 , n710 , n1774 );
not ( n1776 , n3 );
not ( n1777 , n1 );
and ( n1778 , n16 , n444 , n1051 );
nor ( n1779 , n2 , n6 );
and ( n1780 , n8 , n1779 , n812 );
nor ( n1781 , n1778 , n1780 );
or ( n1782 , n17 , n1777 , n1781 );
nand ( n1783 , n2 , n1633 );
nand ( n1784 , n1782 , n1783 );
and ( n1785 , n1776 , n1784 );
not ( n1786 , n454 );
and ( n1787 , n1786 , n155 );
nor ( n1788 , n1785 , n1787 );
not ( n1789 , n1331 );
not ( n1790 , n1749 );
nor ( n1791 , n1788 , n1789 , n1790 );
nor ( n1792 , n1775 , n1791 );
nand ( n1793 , n1742 , n1761 , n1792 );
not ( n1794 , n2 );
nand ( n1795 , n1047 , n1687 , n753 , n1690 );
not ( n1796 , n782 );
or ( n1797 , n1795 , n325 , n1796 );
not ( n1798 , n745 );
nand ( n1799 , n1798 , n1686 , n985 , n1405 );
and ( n1800 , n9 , n14 );
and ( n1801 , n1800 , n710 );
not ( n1802 , n788 );
nand ( n1803 , n1801 , n1802 , n102 , n56 );
nand ( n1804 , n1799 , n1803 );
and ( n1805 , n87 , n1804 );
and ( n1806 , n697 , n1286 );
nor ( n1807 , n1805 , n1806 );
or ( n1808 , n825 , n1807 );
nand ( n1809 , n1797 , n1808 );
not ( n1810 , n1809 );
or ( n1811 , n1794 , n1810 );
nand ( n1812 , n151 , n1177 , n1499 );
not ( n1813 , n293 );
or ( n1814 , n1812 , n8 , n1813 );
nand ( n1815 , n1286 , n1511 );
and ( n1816 , n197 , n1062 );
nand ( n1817 , n1816 , n14 , n56 , n125 );
nand ( n1818 , n1815 , n1817 );
and ( n1819 , n398 , n1818 );
not ( n1820 , n452 );
nand ( n1821 , n1820 , n1749 );
not ( n1822 , n1821 );
nor ( n1823 , n1819 , n1822 );
or ( n1824 , n1 , n1823 );
nand ( n1825 , n1814 , n1824 );
and ( n1826 , n36 , n1825 );
not ( n1827 , n1 );
nand ( n1828 , n533 , n229 );
nand ( n1829 , n259 , n282 , n1616 );
nand ( n1830 , n1828 , n1829 );
and ( n1831 , n16 , n1830 );
nor ( n1832 , t_0 , n1831 );
or ( n1833 , n4 , n1832 );
not ( n1834 , n11 );
not ( n1835 , n5 );
nand ( n1836 , n1834 , n1835 , n206 );
nand ( n1837 , n1833 , n1836 );
and ( n1838 , n1837 , n151 , n736 );
not ( n1839 , n3 );
not ( n1840 , n113 );
nor ( n1841 , n1839 , n1840 , n1562 );
nor ( n1842 , n1838 , n1841 );
nor ( n1843 , n1827 , n1842 );
nor ( n1844 , n1826 , n1843 );
or ( n1845 , n2 , n1844 );
nand ( n1846 , n1811 , n1845 );
not ( n1847 , n2 );
nand ( n1848 , n5 , n579 , n1286 );
or ( n1849 , n1848 , n1 , n409 );
not ( n1850 , n1 );
nand ( n1851 , n1850 , n1749 , n340 , n366 );
and ( n1852 , n1851 , n1757 );
or ( n1853 , n5 , n1852 );
nand ( n1854 , n1849 , n1853 );
and ( n1855 , n1847 , n1854 );
not ( n1856 , n911 );
nand ( n1857 , n1405 , n87 , n1133 , n1305 );
or ( n1858 , n1857 , n5 , n1407 );
not ( n1859 , n5 );
and ( n1860 , n789 , n1725 );
and ( n1861 , n299 , n1400 );
nor ( n1862 , n1860 , n1861 );
or ( n1863 , n1859 , n1862 );
nand ( n1864 , n1858 , n1863 );
and ( n1865 , n1856 , n1864 );
nor ( n1866 , n1855 , n1865 );
or ( n1867 , n163 , n1866 );
not ( n1868 , n481 );
and ( n1869 , n2 , n1868 );
not ( n1870 , n17 );
and ( n1871 , n1870 , n1779 );
nor ( n1872 , n1869 , n1871 );
not ( n1873 , n1688 );
not ( n1874 , n298 );
or ( n1875 , n1872 , n1873 , n1874 );
nor ( n1876 , n13 , n1319 , n443 );
and ( n1877 , n1876 , n476 , n618 );
nor ( n1878 , n1877 , n910 );
or ( n1879 , n351 , n1878 );
nand ( n1880 , n1875 , n1879 );
and ( n1881 , n5 , n1880 );
not ( n1882 , n5 );
and ( n1883 , n1882 , n1460 );
nor ( n1884 , n1881 , n1883 );
or ( n1885 , n364 , n1884 );
or ( n1886 , n14 , n1885 );
not ( n1887 , n5 );
not ( n1888 , n649 );
not ( n1889 , n607 );
nor ( n1890 , n1887 , n1888 , n1889 );
and ( n1891 , n1890 , n1800 , n789 );
nand ( n1892 , n890 , n87 , n1202 );
or ( n1893 , n1892 , n360 , n950 );
not ( n1894 , n9 );
and ( n1895 , n1894 , n11 , n890 );
nand ( n1896 , n5 , n9 );
nor ( n1897 , n11 , n1896 , n586 );
nor ( n1898 , n1895 , n1897 );
or ( n1899 , n814 , n1898 );
nand ( n1900 , n1893 , n1899 );
and ( n1901 , n80 , n1900 );
and ( n1902 , n172 , n1203 );
not ( n1903 , n5 );
and ( n1904 , n1902 , n1903 , n390 , n320 );
nor ( n1905 , n1901 , n1904 );
or ( n1906 , n12 , n8 , n1905 );
not ( n1907 , n576 );
nand ( n1908 , n1907 , n1305 );
nand ( n1909 , n1906 , n1908 );
and ( n1910 , n151 , n1909 );
nor ( n1911 , n1891 , n1910 );
or ( n1912 , n3 , n1911 );
nand ( n1913 , n1867 , n1886 , n1912 );
or ( n1914 , n1821 , n801 , n1067 );
not ( n1915 , n3 );
nor ( n1916 , n248 , n1896 , n392 );
and ( n1917 , n1916 , n176 , n618 );
nand ( n1918 , n325 , n910 , n112 );
not ( n1919 , n780 );
or ( n1920 , n1918 , n417 , n1919 );
not ( n1921 , n279 );
nor ( n1922 , n1921 , n255 , n111 );
nor ( n1923 , t_1 , n1922 );
or ( n1924 , n619 , n1923 );
nand ( n1925 , n1920 , n1924 );
and ( n1926 , n248 , n1925 );
nor ( n1927 , n1917 , n1926 );
or ( n1928 , n1048 , n1927 );
or ( n1929 , n437 , n576 );
nand ( n1930 , n1928 , n1929 );
and ( n1931 , n151 , n1930 );
not ( n1932 , n2 );
and ( n1933 , n1932 , n1598 );
nor ( n1934 , n1931 , n1933 );
or ( n1935 , n1915 , n1934 );
nand ( n1936 , n1914 , n1935 );
and ( n1937 , n185 , n1687 );
and ( n1938 , n1937 , n36 , n903 );
nor ( n1939 , n1938 , n1599 );
or ( n1940 , n2 , n1939 );
not ( n1941 , n5 );
not ( n1942 , n4 );
or ( n1943 , n1942 , n1380 , n137 );
not ( n1944 , n4 );
nand ( n1945 , n151 , n1944 , n1470 );
nand ( n1946 , n1943 , n1945 );
nand ( n1947 , n1941 , n1675 , n1946 );
nand ( n1948 , n1940 , n1947 );
not ( n1949 , n1 );
or ( n1950 , n1949 , n108 , n814 );
not ( n1951 , n1606 );
nand ( n1952 , n716 , n1139 , n1951 );
nand ( n1953 , n1950 , n1952 );
nand ( n1954 , n151 , n519 , n1953 );
not ( n1955 , n9 );
nor ( n1956 , n1954 , n1955 , n11 );
endmodule
