//NOTE: no-implementation module stub

module crp (
    output wire P,
    output wire R,
    input wire K_sub
);

endmodule
