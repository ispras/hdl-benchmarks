//NOTE: no-implementation module stub

module crp (
    output [31:0] P,
    input [31:0] R,
    input [31:0] K_sub
);
endmodule
