module OptKuznechikDecoder(
  input wire clk,
  input wire [127:0] encoded,
  input wire [255:0] key,
  output wire [127:0] out
);
  wire [7:0] literal_2043896[256] = '{8'hfc, 8'hee, 8'hdd, 8'h11, 8'hcf, 8'h6e, 8'h31, 8'h16, 8'hfb, 8'hc4, 8'hfa, 8'hda, 8'h23, 8'hc5, 8'h04, 8'h4d, 8'he9, 8'h77, 8'hf0, 8'hdb, 8'h93, 8'h2e, 8'h99, 8'hba, 8'h17, 8'h36, 8'hf1, 8'hbb, 8'h14, 8'hcd, 8'h5f, 8'hc1, 8'hf9, 8'h18, 8'h65, 8'h5a, 8'he2, 8'h5c, 8'hef, 8'h21, 8'h81, 8'h1c, 8'h3c, 8'h42, 8'h8b, 8'h01, 8'h8e, 8'h4f, 8'h05, 8'h84, 8'h02, 8'hae, 8'he3, 8'h6a, 8'h8f, 8'ha0, 8'h06, 8'h0b, 8'hed, 8'h98, 8'h7f, 8'hd4, 8'hd3, 8'h1f, 8'heb, 8'h34, 8'h2c, 8'h51, 8'hea, 8'hc8, 8'h48, 8'hab, 8'hf2, 8'h2a, 8'h68, 8'ha2, 8'hfd, 8'h3a, 8'hce, 8'hcc, 8'hb5, 8'h70, 8'h0e, 8'h56, 8'h08, 8'h0c, 8'h76, 8'h12, 8'hbf, 8'h72, 8'h13, 8'h47, 8'h9c, 8'hb7, 8'h5d, 8'h87, 8'h15, 8'ha1, 8'h96, 8'h29, 8'h10, 8'h7b, 8'h9a, 8'hc7, 8'hf3, 8'h91, 8'h78, 8'h6f, 8'h9d, 8'h9e, 8'hb2, 8'hb1, 8'h32, 8'h75, 8'h19, 8'h3d, 8'hff, 8'h35, 8'h8a, 8'h7e, 8'h6d, 8'h54, 8'hc6, 8'h80, 8'hc3, 8'hbd, 8'h0d, 8'h57, 8'hdf, 8'hf5, 8'h24, 8'ha9, 8'h3e, 8'ha8, 8'h43, 8'hc9, 8'hd7, 8'h79, 8'hd6, 8'hf6, 8'h7c, 8'h22, 8'hb9, 8'h03, 8'he0, 8'h0f, 8'hec, 8'hde, 8'h7a, 8'h94, 8'hb0, 8'hbc, 8'hdc, 8'he8, 8'h28, 8'h50, 8'h4e, 8'h33, 8'h0a, 8'h4a, 8'ha7, 8'h97, 8'h60, 8'h73, 8'h1e, 8'h00, 8'h62, 8'h44, 8'h1a, 8'hb8, 8'h38, 8'h82, 8'h64, 8'h9f, 8'h26, 8'h41, 8'had, 8'h45, 8'h46, 8'h92, 8'h27, 8'h5e, 8'h55, 8'h2f, 8'h8c, 8'ha3, 8'ha5, 8'h7d, 8'h69, 8'hd5, 8'h95, 8'h3b, 8'h07, 8'h58, 8'hb3, 8'h40, 8'h86, 8'hac, 8'h1d, 8'hf7, 8'h30, 8'h37, 8'h6b, 8'he4, 8'h88, 8'hd9, 8'he7, 8'h89, 8'he1, 8'h1b, 8'h83, 8'h49, 8'h4c, 8'h3f, 8'hf8, 8'hfe, 8'h8d, 8'h53, 8'haa, 8'h90, 8'hca, 8'hd8, 8'h85, 8'h61, 8'h20, 8'h71, 8'h67, 8'ha4, 8'h2d, 8'h2b, 8'h09, 8'h5b, 8'hcb, 8'h9b, 8'h25, 8'hd0, 8'hbe, 8'he5, 8'h6c, 8'h52, 8'h59, 8'ha6, 8'h74, 8'hd2, 8'he6, 8'hf4, 8'hb4, 8'hc0, 8'hd1, 8'h66, 8'haf, 8'hc2, 8'h39, 8'h4b, 8'h63, 8'hb6};
  wire [7:0] literal_2043910[256] = '{8'h00, 8'h94, 8'heb, 8'h7f, 8'h15, 8'h81, 8'hfe, 8'h6a, 8'h2a, 8'hbe, 8'hc1, 8'h55, 8'h3f, 8'hab, 8'hd4, 8'h40, 8'h54, 8'hc0, 8'hbf, 8'h2b, 8'h41, 8'hd5, 8'haa, 8'h3e, 8'h7e, 8'hea, 8'h95, 8'h01, 8'h6b, 8'hff, 8'h80, 8'h14, 8'ha8, 8'h3c, 8'h43, 8'hd7, 8'hbd, 8'h29, 8'h56, 8'hc2, 8'h82, 8'h16, 8'h69, 8'hfd, 8'h97, 8'h03, 8'h7c, 8'he8, 8'hfc, 8'h68, 8'h17, 8'h83, 8'he9, 8'h7d, 8'h02, 8'h96, 8'hd6, 8'h42, 8'h3d, 8'ha9, 8'hc3, 8'h57, 8'h28, 8'hbc, 8'h93, 8'h07, 8'h78, 8'hec, 8'h86, 8'h12, 8'h6d, 8'hf9, 8'hb9, 8'h2d, 8'h52, 8'hc6, 8'hac, 8'h38, 8'h47, 8'hd3, 8'hc7, 8'h53, 8'h2c, 8'hb8, 8'hd2, 8'h46, 8'h39, 8'had, 8'hed, 8'h79, 8'h06, 8'h92, 8'hf8, 8'h6c, 8'h13, 8'h87, 8'h3b, 8'haf, 8'hd0, 8'h44, 8'h2e, 8'hba, 8'hc5, 8'h51, 8'h11, 8'h85, 8'hfa, 8'h6e, 8'h04, 8'h90, 8'hef, 8'h7b, 8'h6f, 8'hfb, 8'h84, 8'h10, 8'h7a, 8'hee, 8'h91, 8'h05, 8'h45, 8'hd1, 8'hae, 8'h3a, 8'h50, 8'hc4, 8'hbb, 8'h2f, 8'he5, 8'h71, 8'h0e, 8'h9a, 8'hf0, 8'h64, 8'h1b, 8'h8f, 8'hcf, 8'h5b, 8'h24, 8'hb0, 8'hda, 8'h4e, 8'h31, 8'ha5, 8'hb1, 8'h25, 8'h5a, 8'hce, 8'ha4, 8'h30, 8'h4f, 8'hdb, 8'h9b, 8'h0f, 8'h70, 8'he4, 8'h8e, 8'h1a, 8'h65, 8'hf1, 8'h4d, 8'hd9, 8'ha6, 8'h32, 8'h58, 8'hcc, 8'hb3, 8'h27, 8'h67, 8'hf3, 8'h8c, 8'h18, 8'h72, 8'he6, 8'h99, 8'h0d, 8'h19, 8'h8d, 8'hf2, 8'h66, 8'h0c, 8'h98, 8'he7, 8'h73, 8'h33, 8'ha7, 8'hd8, 8'h4c, 8'h26, 8'hb2, 8'hcd, 8'h59, 8'h76, 8'he2, 8'h9d, 8'h09, 8'h63, 8'hf7, 8'h88, 8'h1c, 8'h5c, 8'hc8, 8'hb7, 8'h23, 8'h49, 8'hdd, 8'ha2, 8'h36, 8'h22, 8'hb6, 8'hc9, 8'h5d, 8'h37, 8'ha3, 8'hdc, 8'h48, 8'h08, 8'h9c, 8'he3, 8'h77, 8'h1d, 8'h89, 8'hf6, 8'h62, 8'hde, 8'h4a, 8'h35, 8'ha1, 8'hcb, 8'h5f, 8'h20, 8'hb4, 8'hf4, 8'h60, 8'h1f, 8'h8b, 8'he1, 8'h75, 8'h0a, 8'h9e, 8'h8a, 8'h1e, 8'h61, 8'hf5, 8'h9f, 8'h0b, 8'h74, 8'he0, 8'ha0, 8'h34, 8'h4b, 8'hdf, 8'hb5, 8'h21, 8'h5e, 8'hca};
  wire [7:0] literal_2043912[256] = '{8'h00, 8'h20, 8'h40, 8'h60, 8'h80, 8'ha0, 8'hc0, 8'he0, 8'hc3, 8'he3, 8'h83, 8'ha3, 8'h43, 8'h63, 8'h03, 8'h23, 8'h45, 8'h65, 8'h05, 8'h25, 8'hc5, 8'he5, 8'h85, 8'ha5, 8'h86, 8'ha6, 8'hc6, 8'he6, 8'h06, 8'h26, 8'h46, 8'h66, 8'h8a, 8'haa, 8'hca, 8'hea, 8'h0a, 8'h2a, 8'h4a, 8'h6a, 8'h49, 8'h69, 8'h09, 8'h29, 8'hc9, 8'he9, 8'h89, 8'ha9, 8'hcf, 8'hef, 8'h8f, 8'haf, 8'h4f, 8'h6f, 8'h0f, 8'h2f, 8'h0c, 8'h2c, 8'h4c, 8'h6c, 8'h8c, 8'hac, 8'hcc, 8'hec, 8'hd7, 8'hf7, 8'h97, 8'hb7, 8'h57, 8'h77, 8'h17, 8'h37, 8'h14, 8'h34, 8'h54, 8'h74, 8'h94, 8'hb4, 8'hd4, 8'hf4, 8'h92, 8'hb2, 8'hd2, 8'hf2, 8'h12, 8'h32, 8'h52, 8'h72, 8'h51, 8'h71, 8'h11, 8'h31, 8'hd1, 8'hf1, 8'h91, 8'hb1, 8'h5d, 8'h7d, 8'h1d, 8'h3d, 8'hdd, 8'hfd, 8'h9d, 8'hbd, 8'h9e, 8'hbe, 8'hde, 8'hfe, 8'h1e, 8'h3e, 8'h5e, 8'h7e, 8'h18, 8'h38, 8'h58, 8'h78, 8'h98, 8'hb8, 8'hd8, 8'hf8, 8'hdb, 8'hfb, 8'h9b, 8'hbb, 8'h5b, 8'h7b, 8'h1b, 8'h3b, 8'h6d, 8'h4d, 8'h2d, 8'h0d, 8'hed, 8'hcd, 8'had, 8'h8d, 8'hae, 8'h8e, 8'hee, 8'hce, 8'h2e, 8'h0e, 8'h6e, 8'h4e, 8'h28, 8'h08, 8'h68, 8'h48, 8'ha8, 8'h88, 8'he8, 8'hc8, 8'heb, 8'hcb, 8'hab, 8'h8b, 8'h6b, 8'h4b, 8'h2b, 8'h0b, 8'he7, 8'hc7, 8'ha7, 8'h87, 8'h67, 8'h47, 8'h27, 8'h07, 8'h24, 8'h04, 8'h64, 8'h44, 8'ha4, 8'h84, 8'he4, 8'hc4, 8'ha2, 8'h82, 8'he2, 8'hc2, 8'h22, 8'h02, 8'h62, 8'h42, 8'h61, 8'h41, 8'h21, 8'h01, 8'he1, 8'hc1, 8'ha1, 8'h81, 8'hba, 8'h9a, 8'hfa, 8'hda, 8'h3a, 8'h1a, 8'h7a, 8'h5a, 8'h79, 8'h59, 8'h39, 8'h19, 8'hf9, 8'hd9, 8'hb9, 8'h99, 8'hff, 8'hdf, 8'hbf, 8'h9f, 8'h7f, 8'h5f, 8'h3f, 8'h1f, 8'h3c, 8'h1c, 8'h7c, 8'h5c, 8'hbc, 8'h9c, 8'hfc, 8'hdc, 8'h30, 8'h10, 8'h70, 8'h50, 8'hb0, 8'h90, 8'hf0, 8'hd0, 8'hf3, 8'hd3, 8'hb3, 8'h93, 8'h73, 8'h53, 8'h33, 8'h13, 8'h75, 8'h55, 8'h35, 8'h15, 8'hf5, 8'hd5, 8'hb5, 8'h95, 8'hb6, 8'h96, 8'hf6, 8'hd6, 8'h36, 8'h16, 8'h76, 8'h56};
  wire [7:0] literal_2043914[256] = '{8'h00, 8'h85, 8'hc9, 8'h4c, 8'h51, 8'hd4, 8'h98, 8'h1d, 8'ha2, 8'h27, 8'h6b, 8'hee, 8'hf3, 8'h76, 8'h3a, 8'hbf, 8'h87, 8'h02, 8'h4e, 8'hcb, 8'hd6, 8'h53, 8'h1f, 8'h9a, 8'h25, 8'ha0, 8'hec, 8'h69, 8'h74, 8'hf1, 8'hbd, 8'h38, 8'hcd, 8'h48, 8'h04, 8'h81, 8'h9c, 8'h19, 8'h55, 8'hd0, 8'h6f, 8'hea, 8'ha6, 8'h23, 8'h3e, 8'hbb, 8'hf7, 8'h72, 8'h4a, 8'hcf, 8'h83, 8'h06, 8'h1b, 8'h9e, 8'hd2, 8'h57, 8'he8, 8'h6d, 8'h21, 8'ha4, 8'hb9, 8'h3c, 8'h70, 8'hf5, 8'h59, 8'hdc, 8'h90, 8'h15, 8'h08, 8'h8d, 8'hc1, 8'h44, 8'hfb, 8'h7e, 8'h32, 8'hb7, 8'haa, 8'h2f, 8'h63, 8'he6, 8'hde, 8'h5b, 8'h17, 8'h92, 8'h8f, 8'h0a, 8'h46, 8'hc3, 8'h7c, 8'hf9, 8'hb5, 8'h30, 8'h2d, 8'ha8, 8'he4, 8'h61, 8'h94, 8'h11, 8'h5d, 8'hd8, 8'hc5, 8'h40, 8'h0c, 8'h89, 8'h36, 8'hb3, 8'hff, 8'h7a, 8'h67, 8'he2, 8'hae, 8'h2b, 8'h13, 8'h96, 8'hda, 8'h5f, 8'h42, 8'hc7, 8'h8b, 8'h0e, 8'hb1, 8'h34, 8'h78, 8'hfd, 8'he0, 8'h65, 8'h29, 8'hac, 8'hb2, 8'h37, 8'h7b, 8'hfe, 8'he3, 8'h66, 8'h2a, 8'haf, 8'h10, 8'h95, 8'hd9, 8'h5c, 8'h41, 8'hc4, 8'h88, 8'h0d, 8'h35, 8'hb0, 8'hfc, 8'h79, 8'h64, 8'he1, 8'had, 8'h28, 8'h97, 8'h12, 8'h5e, 8'hdb, 8'hc6, 8'h43, 8'h0f, 8'h8a, 8'h7f, 8'hfa, 8'hb6, 8'h33, 8'h2e, 8'hab, 8'he7, 8'h62, 8'hdd, 8'h58, 8'h14, 8'h91, 8'h8c, 8'h09, 8'h45, 8'hc0, 8'hf8, 8'h7d, 8'h31, 8'hb4, 8'ha9, 8'h2c, 8'h60, 8'he5, 8'h5a, 8'hdf, 8'h93, 8'h16, 8'h0b, 8'h8e, 8'hc2, 8'h47, 8'heb, 8'h6e, 8'h22, 8'ha7, 8'hba, 8'h3f, 8'h73, 8'hf6, 8'h49, 8'hcc, 8'h80, 8'h05, 8'h18, 8'h9d, 8'hd1, 8'h54, 8'h6c, 8'he9, 8'ha5, 8'h20, 8'h3d, 8'hb8, 8'hf4, 8'h71, 8'hce, 8'h4b, 8'h07, 8'h82, 8'h9f, 8'h1a, 8'h56, 8'hd3, 8'h26, 8'ha3, 8'hef, 8'h6a, 8'h77, 8'hf2, 8'hbe, 8'h3b, 8'h84, 8'h01, 8'h4d, 8'hc8, 8'hd5, 8'h50, 8'h1c, 8'h99, 8'ha1, 8'h24, 8'h68, 8'hed, 8'hf0, 8'h75, 8'h39, 8'hbc, 8'h03, 8'h86, 8'hca, 8'h4f, 8'h52, 8'hd7, 8'h9b, 8'h1e};
  wire [7:0] literal_2043916[256] = '{8'h00, 8'h10, 8'h20, 8'h30, 8'h40, 8'h50, 8'h60, 8'h70, 8'h80, 8'h90, 8'ha0, 8'hb0, 8'hc0, 8'hd0, 8'he0, 8'hf0, 8'hc3, 8'hd3, 8'he3, 8'hf3, 8'h83, 8'h93, 8'ha3, 8'hb3, 8'h43, 8'h53, 8'h63, 8'h73, 8'h03, 8'h13, 8'h23, 8'h33, 8'h45, 8'h55, 8'h65, 8'h75, 8'h05, 8'h15, 8'h25, 8'h35, 8'hc5, 8'hd5, 8'he5, 8'hf5, 8'h85, 8'h95, 8'ha5, 8'hb5, 8'h86, 8'h96, 8'ha6, 8'hb6, 8'hc6, 8'hd6, 8'he6, 8'hf6, 8'h06, 8'h16, 8'h26, 8'h36, 8'h46, 8'h56, 8'h66, 8'h76, 8'h8a, 8'h9a, 8'haa, 8'hba, 8'hca, 8'hda, 8'hea, 8'hfa, 8'h0a, 8'h1a, 8'h2a, 8'h3a, 8'h4a, 8'h5a, 8'h6a, 8'h7a, 8'h49, 8'h59, 8'h69, 8'h79, 8'h09, 8'h19, 8'h29, 8'h39, 8'hc9, 8'hd9, 8'he9, 8'hf9, 8'h89, 8'h99, 8'ha9, 8'hb9, 8'hcf, 8'hdf, 8'hef, 8'hff, 8'h8f, 8'h9f, 8'haf, 8'hbf, 8'h4f, 8'h5f, 8'h6f, 8'h7f, 8'h0f, 8'h1f, 8'h2f, 8'h3f, 8'h0c, 8'h1c, 8'h2c, 8'h3c, 8'h4c, 8'h5c, 8'h6c, 8'h7c, 8'h8c, 8'h9c, 8'hac, 8'hbc, 8'hcc, 8'hdc, 8'hec, 8'hfc, 8'hd7, 8'hc7, 8'hf7, 8'he7, 8'h97, 8'h87, 8'hb7, 8'ha7, 8'h57, 8'h47, 8'h77, 8'h67, 8'h17, 8'h07, 8'h37, 8'h27, 8'h14, 8'h04, 8'h34, 8'h24, 8'h54, 8'h44, 8'h74, 8'h64, 8'h94, 8'h84, 8'hb4, 8'ha4, 8'hd4, 8'hc4, 8'hf4, 8'he4, 8'h92, 8'h82, 8'hb2, 8'ha2, 8'hd2, 8'hc2, 8'hf2, 8'he2, 8'h12, 8'h02, 8'h32, 8'h22, 8'h52, 8'h42, 8'h72, 8'h62, 8'h51, 8'h41, 8'h71, 8'h61, 8'h11, 8'h01, 8'h31, 8'h21, 8'hd1, 8'hc1, 8'hf1, 8'he1, 8'h91, 8'h81, 8'hb1, 8'ha1, 8'h5d, 8'h4d, 8'h7d, 8'h6d, 8'h1d, 8'h0d, 8'h3d, 8'h2d, 8'hdd, 8'hcd, 8'hfd, 8'hed, 8'h9d, 8'h8d, 8'hbd, 8'had, 8'h9e, 8'h8e, 8'hbe, 8'hae, 8'hde, 8'hce, 8'hfe, 8'hee, 8'h1e, 8'h0e, 8'h3e, 8'h2e, 8'h5e, 8'h4e, 8'h7e, 8'h6e, 8'h18, 8'h08, 8'h38, 8'h28, 8'h58, 8'h48, 8'h78, 8'h68, 8'h98, 8'h88, 8'hb8, 8'ha8, 8'hd8, 8'hc8, 8'hf8, 8'he8, 8'hdb, 8'hcb, 8'hfb, 8'heb, 8'h9b, 8'h8b, 8'hbb, 8'hab, 8'h5b, 8'h4b, 8'h7b, 8'h6b, 8'h1b, 8'h0b, 8'h3b, 8'h2b};
  wire [7:0] literal_2043918[256] = '{8'h00, 8'hc2, 8'h47, 8'h85, 8'h8e, 8'h4c, 8'hc9, 8'h0b, 8'hdf, 8'h1d, 8'h98, 8'h5a, 8'h51, 8'h93, 8'h16, 8'hd4, 8'h7d, 8'hbf, 8'h3a, 8'hf8, 8'hf3, 8'h31, 8'hb4, 8'h76, 8'ha2, 8'h60, 8'he5, 8'h27, 8'h2c, 8'hee, 8'h6b, 8'ha9, 8'hfa, 8'h38, 8'hbd, 8'h7f, 8'h74, 8'hb6, 8'h33, 8'hf1, 8'h25, 8'he7, 8'h62, 8'ha0, 8'hab, 8'h69, 8'hec, 8'h2e, 8'h87, 8'h45, 8'hc0, 8'h02, 8'h09, 8'hcb, 8'h4e, 8'h8c, 8'h58, 8'h9a, 8'h1f, 8'hdd, 8'hd6, 8'h14, 8'h91, 8'h53, 8'h37, 8'hf5, 8'h70, 8'hb2, 8'hb9, 8'h7b, 8'hfe, 8'h3c, 8'he8, 8'h2a, 8'haf, 8'h6d, 8'h66, 8'ha4, 8'h21, 8'he3, 8'h4a, 8'h88, 8'h0d, 8'hcf, 8'hc4, 8'h06, 8'h83, 8'h41, 8'h95, 8'h57, 8'hd2, 8'h10, 8'h1b, 8'hd9, 8'h5c, 8'h9e, 8'hcd, 8'h0f, 8'h8a, 8'h48, 8'h43, 8'h81, 8'h04, 8'hc6, 8'h12, 8'hd0, 8'h55, 8'h97, 8'h9c, 8'h5e, 8'hdb, 8'h19, 8'hb0, 8'h72, 8'hf7, 8'h35, 8'h3e, 8'hfc, 8'h79, 8'hbb, 8'h6f, 8'had, 8'h28, 8'hea, 8'he1, 8'h23, 8'ha6, 8'h64, 8'h6e, 8'hac, 8'h29, 8'heb, 8'he0, 8'h22, 8'ha7, 8'h65, 8'hb1, 8'h73, 8'hf6, 8'h34, 8'h3f, 8'hfd, 8'h78, 8'hba, 8'h13, 8'hd1, 8'h54, 8'h96, 8'h9d, 8'h5f, 8'hda, 8'h18, 8'hcc, 8'h0e, 8'h8b, 8'h49, 8'h42, 8'h80, 8'h05, 8'hc7, 8'h94, 8'h56, 8'hd3, 8'h11, 8'h1a, 8'hd8, 8'h5d, 8'h9f, 8'h4b, 8'h89, 8'h0c, 8'hce, 8'hc5, 8'h07, 8'h82, 8'h40, 8'he9, 8'h2b, 8'hae, 8'h6c, 8'h67, 8'ha5, 8'h20, 8'he2, 8'h36, 8'hf4, 8'h71, 8'hb3, 8'hb8, 8'h7a, 8'hff, 8'h3d, 8'h59, 8'h9b, 8'h1e, 8'hdc, 8'hd7, 8'h15, 8'h90, 8'h52, 8'h86, 8'h44, 8'hc1, 8'h03, 8'h08, 8'hca, 8'h4f, 8'h8d, 8'h24, 8'he6, 8'h63, 8'ha1, 8'haa, 8'h68, 8'hed, 8'h2f, 8'hfb, 8'h39, 8'hbc, 8'h7e, 8'h75, 8'hb7, 8'h32, 8'hf0, 8'ha3, 8'h61, 8'he4, 8'h26, 8'h2d, 8'hef, 8'h6a, 8'ha8, 8'h7c, 8'hbe, 8'h3b, 8'hf9, 8'hf2, 8'h30, 8'hb5, 8'h77, 8'hde, 8'h1c, 8'h99, 8'h5b, 8'h50, 8'h92, 8'h17, 8'hd5, 8'h01, 8'hc3, 8'h46, 8'h84, 8'h8f, 8'h4d, 8'hc8, 8'h0a};
  wire [7:0] literal_2043920[256] = '{8'h00, 8'hc0, 8'h43, 8'h83, 8'h86, 8'h46, 8'hc5, 8'h05, 8'hcf, 8'h0f, 8'h8c, 8'h4c, 8'h49, 8'h89, 8'h0a, 8'hca, 8'h5d, 8'h9d, 8'h1e, 8'hde, 8'hdb, 8'h1b, 8'h98, 8'h58, 8'h92, 8'h52, 8'hd1, 8'h11, 8'h14, 8'hd4, 8'h57, 8'h97, 8'hba, 8'h7a, 8'hf9, 8'h39, 8'h3c, 8'hfc, 8'h7f, 8'hbf, 8'h75, 8'hb5, 8'h36, 8'hf6, 8'hf3, 8'h33, 8'hb0, 8'h70, 8'he7, 8'h27, 8'ha4, 8'h64, 8'h61, 8'ha1, 8'h22, 8'he2, 8'h28, 8'he8, 8'h6b, 8'hab, 8'hae, 8'h6e, 8'hed, 8'h2d, 8'hb7, 8'h77, 8'hf4, 8'h34, 8'h31, 8'hf1, 8'h72, 8'hb2, 8'h78, 8'hb8, 8'h3b, 8'hfb, 8'hfe, 8'h3e, 8'hbd, 8'h7d, 8'hea, 8'h2a, 8'ha9, 8'h69, 8'h6c, 8'hac, 8'h2f, 8'hef, 8'h25, 8'he5, 8'h66, 8'ha6, 8'ha3, 8'h63, 8'he0, 8'h20, 8'h0d, 8'hcd, 8'h4e, 8'h8e, 8'h8b, 8'h4b, 8'hc8, 8'h08, 8'hc2, 8'h02, 8'h81, 8'h41, 8'h44, 8'h84, 8'h07, 8'hc7, 8'h50, 8'h90, 8'h13, 8'hd3, 8'hd6, 8'h16, 8'h95, 8'h55, 8'h9f, 8'h5f, 8'hdc, 8'h1c, 8'h19, 8'hd9, 8'h5a, 8'h9a, 8'had, 8'h6d, 8'hee, 8'h2e, 8'h2b, 8'heb, 8'h68, 8'ha8, 8'h62, 8'ha2, 8'h21, 8'he1, 8'he4, 8'h24, 8'ha7, 8'h67, 8'hf0, 8'h30, 8'hb3, 8'h73, 8'h76, 8'hb6, 8'h35, 8'hf5, 8'h3f, 8'hff, 8'h7c, 8'hbc, 8'hb9, 8'h79, 8'hfa, 8'h3a, 8'h17, 8'hd7, 8'h54, 8'h94, 8'h91, 8'h51, 8'hd2, 8'h12, 8'hd8, 8'h18, 8'h9b, 8'h5b, 8'h5e, 8'h9e, 8'h1d, 8'hdd, 8'h4a, 8'h8a, 8'h09, 8'hc9, 8'hcc, 8'h0c, 8'h8f, 8'h4f, 8'h85, 8'h45, 8'hc6, 8'h06, 8'h03, 8'hc3, 8'h40, 8'h80, 8'h1a, 8'hda, 8'h59, 8'h99, 8'h9c, 8'h5c, 8'hdf, 8'h1f, 8'hd5, 8'h15, 8'h96, 8'h56, 8'h53, 8'h93, 8'h10, 8'hd0, 8'h47, 8'h87, 8'h04, 8'hc4, 8'hc1, 8'h01, 8'h82, 8'h42, 8'h88, 8'h48, 8'hcb, 8'h0b, 8'h0e, 8'hce, 8'h4d, 8'h8d, 8'ha0, 8'h60, 8'he3, 8'h23, 8'h26, 8'he6, 8'h65, 8'ha5, 8'h6f, 8'haf, 8'h2c, 8'hec, 8'he9, 8'h29, 8'haa, 8'h6a, 8'hfd, 8'h3d, 8'hbe, 8'h7e, 8'h7b, 8'hbb, 8'h38, 8'hf8, 8'h32, 8'hf2, 8'h71, 8'hb1, 8'hb4, 8'h74, 8'hf7, 8'h37};
  wire [7:0] literal_2043923[256] = '{8'h00, 8'hfb, 8'h35, 8'hce, 8'h6a, 8'h91, 8'h5f, 8'ha4, 8'hd4, 8'h2f, 8'he1, 8'h1a, 8'hbe, 8'h45, 8'h8b, 8'h70, 8'h6b, 8'h90, 8'h5e, 8'ha5, 8'h01, 8'hfa, 8'h34, 8'hcf, 8'hbf, 8'h44, 8'h8a, 8'h71, 8'hd5, 8'h2e, 8'he0, 8'h1b, 8'hd6, 8'h2d, 8'he3, 8'h18, 8'hbc, 8'h47, 8'h89, 8'h72, 8'h02, 8'hf9, 8'h37, 8'hcc, 8'h68, 8'h93, 8'h5d, 8'ha6, 8'hbd, 8'h46, 8'h88, 8'h73, 8'hd7, 8'h2c, 8'he2, 8'h19, 8'h69, 8'h92, 8'h5c, 8'ha7, 8'h03, 8'hf8, 8'h36, 8'hcd, 8'h6f, 8'h94, 8'h5a, 8'ha1, 8'h05, 8'hfe, 8'h30, 8'hcb, 8'hbb, 8'h40, 8'h8e, 8'h75, 8'hd1, 8'h2a, 8'he4, 8'h1f, 8'h04, 8'hff, 8'h31, 8'hca, 8'h6e, 8'h95, 8'h5b, 8'ha0, 8'hd0, 8'h2b, 8'he5, 8'h1e, 8'hba, 8'h41, 8'h8f, 8'h74, 8'hb9, 8'h42, 8'h8c, 8'h77, 8'hd3, 8'h28, 8'he6, 8'h1d, 8'h6d, 8'h96, 8'h58, 8'ha3, 8'h07, 8'hfc, 8'h32, 8'hc9, 8'hd2, 8'h29, 8'he7, 8'h1c, 8'hb8, 8'h43, 8'h8d, 8'h76, 8'h06, 8'hfd, 8'h33, 8'hc8, 8'h6c, 8'h97, 8'h59, 8'ha2, 8'hde, 8'h25, 8'heb, 8'h10, 8'hb4, 8'h4f, 8'h81, 8'h7a, 8'h0a, 8'hf1, 8'h3f, 8'hc4, 8'h60, 8'h9b, 8'h55, 8'hae, 8'hb5, 8'h4e, 8'h80, 8'h7b, 8'hdf, 8'h24, 8'hea, 8'h11, 8'h61, 8'h9a, 8'h54, 8'haf, 8'h0b, 8'hf0, 8'h3e, 8'hc5, 8'h08, 8'hf3, 8'h3d, 8'hc6, 8'h62, 8'h99, 8'h57, 8'hac, 8'hdc, 8'h27, 8'he9, 8'h12, 8'hb6, 8'h4d, 8'h83, 8'h78, 8'h63, 8'h98, 8'h56, 8'had, 8'h09, 8'hf2, 8'h3c, 8'hc7, 8'hb7, 8'h4c, 8'h82, 8'h79, 8'hdd, 8'h26, 8'he8, 8'h13, 8'hb1, 8'h4a, 8'h84, 8'h7f, 8'hdb, 8'h20, 8'hee, 8'h15, 8'h65, 8'h9e, 8'h50, 8'hab, 8'h0f, 8'hf4, 8'h3a, 8'hc1, 8'hda, 8'h21, 8'hef, 8'h14, 8'hb0, 8'h4b, 8'h85, 8'h7e, 8'h0e, 8'hf5, 8'h3b, 8'hc0, 8'h64, 8'h9f, 8'h51, 8'haa, 8'h67, 8'h9c, 8'h52, 8'ha9, 8'h0d, 8'hf6, 8'h38, 8'hc3, 8'hb3, 8'h48, 8'h86, 8'h7d, 8'hd9, 8'h22, 8'hec, 8'h17, 8'h0c, 8'hf7, 8'h39, 8'hc2, 8'h66, 8'h9d, 8'h53, 8'ha8, 8'hd8, 8'h23, 8'hed, 8'h16, 8'hb2, 8'h49, 8'h87, 8'h7c};
  wire [7:0] literal_2051898[256] = '{8'ha5, 8'h2d, 8'h32, 8'h8f, 8'h0e, 8'h30, 8'h38, 8'hc0, 8'h54, 8'he6, 8'h9e, 8'h39, 8'h55, 8'h7e, 8'h52, 8'h91, 8'h64, 8'h03, 8'h57, 8'h5a, 8'h1c, 8'h60, 8'h07, 8'h18, 8'h21, 8'h72, 8'ha8, 8'hd1, 8'h29, 8'hc6, 8'ha4, 8'h3f, 8'he0, 8'h27, 8'h8d, 8'h0c, 8'h82, 8'hea, 8'hae, 8'hb4, 8'h9a, 8'h63, 8'h49, 8'he5, 8'h42, 8'he4, 8'h15, 8'hb7, 8'hc8, 8'h06, 8'h70, 8'h9d, 8'h41, 8'h75, 8'h19, 8'hc9, 8'haa, 8'hfc, 8'h4d, 8'hbf, 8'h2a, 8'h73, 8'h84, 8'hd5, 8'hc3, 8'haf, 8'h2b, 8'h86, 8'ha7, 8'hb1, 8'hb2, 8'h5b, 8'h46, 8'hd3, 8'h9f, 8'hfd, 8'hd4, 8'h0f, 8'h9c, 8'h2f, 8'h9b, 8'h43, 8'hef, 8'hd9, 8'h79, 8'hb6, 8'h53, 8'h7f, 8'hc1, 8'hf0, 8'h23, 8'he7, 8'h25, 8'h5e, 8'hb5, 8'h1e, 8'ha2, 8'hdf, 8'ha6, 8'hfe, 8'hac, 8'h22, 8'hf9, 8'he2, 8'h4a, 8'hbc, 8'h35, 8'hca, 8'hee, 8'h78, 8'h05, 8'h6b, 8'h51, 8'he1, 8'h59, 8'ha3, 8'hf2, 8'h71, 8'h56, 8'h11, 8'h6a, 8'h89, 8'h94, 8'h65, 8'h8c, 8'hbb, 8'h77, 8'h3c, 8'h7b, 8'h28, 8'hab, 8'hd2, 8'h31, 8'hde, 8'hc4, 8'h5f, 8'hcc, 8'hcf, 8'h76, 8'h2c, 8'hb8, 8'hd8, 8'h2e, 8'h36, 8'hdb, 8'h69, 8'hb3, 8'h14, 8'h95, 8'hbe, 8'h62, 8'ha1, 8'h3b, 8'h16, 8'h66, 8'he9, 8'h5c, 8'h6c, 8'h6d, 8'had, 8'h37, 8'h61, 8'h4b, 8'hb9, 8'he3, 8'hba, 8'hf1, 8'ha0, 8'h85, 8'h83, 8'hda, 8'h47, 8'hc5, 8'hb0, 8'h33, 8'hfa, 8'h96, 8'h6f, 8'h6e, 8'hc2, 8'hf6, 8'h50, 8'hff, 8'h5d, 8'ha9, 8'h8e, 8'h17, 8'h1b, 8'h97, 8'h7d, 8'hec, 8'h58, 8'hf7, 8'h1f, 8'hfb, 8'h7c, 8'h09, 8'h0d, 8'h7a, 8'h67, 8'h45, 8'h87, 8'hdc, 8'he8, 8'h4f, 8'h1d, 8'h4e, 8'h04, 8'heb, 8'hf8, 8'hf3, 8'h3e, 8'h3d, 8'hbd, 8'h8a, 8'h88, 8'hdd, 8'hcd, 8'h0b, 8'h13, 8'h98, 8'h02, 8'h93, 8'h80, 8'h90, 8'hd0, 8'h24, 8'h34, 8'hcb, 8'hed, 8'hf4, 8'hce, 8'h99, 8'h10, 8'h44, 8'h40, 8'h92, 8'h3a, 8'h01, 8'h26, 8'h12, 8'h1a, 8'h48, 8'h68, 8'hf5, 8'h81, 8'h8b, 8'hc7, 8'hd6, 8'h20, 8'h0a, 8'h08, 8'h00, 8'h4c, 8'hd7, 8'h74};

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [127:0] p0_encoded;
  reg [255:0] p0_key;
  reg [7:0] p1_literal_2043896[256];
  reg [7:0] p1_literal_2043910[256];
  reg [7:0] p1_literal_2043912[256];
  reg [7:0] p1_literal_2043914[256];
  reg [7:0] p1_literal_2043916[256];
  reg [7:0] p1_literal_2043918[256];
  reg [7:0] p1_literal_2043920[256];
  reg [7:0] p1_literal_2043923[256];
  reg [7:0] p8_literal_2051898[256];
  always_ff @ (posedge clk) begin
    p0_encoded <= encoded;
    p0_key <= key;
    p1_literal_2043896 <= literal_2043896;
    p1_literal_2043910 <= literal_2043910;
    p1_literal_2043912 <= literal_2043912;
    p1_literal_2043914 <= literal_2043914;
    p1_literal_2043916 <= literal_2043916;
    p1_literal_2043918 <= literal_2043918;
    p1_literal_2043920 <= literal_2043920;
    p1_literal_2043923 <= literal_2043923;
    p8_literal_2051898 <= literal_2051898;
  end

  // ===== Pipe stage 1:
  wire [127:0] p1_bit_slice_2043893_comb;
  wire [127:0] p1_addedKey__32_comb;
  wire [7:0] p1_array_index_2043911_comb;
  wire [7:0] p1_array_index_2043913_comb;
  wire [7:0] p1_array_index_2043915_comb;
  wire [7:0] p1_array_index_2043917_comb;
  wire [7:0] p1_array_index_2043919_comb;
  wire [7:0] p1_array_index_2043921_comb;
  wire [7:0] p1_array_index_2043924_comb;
  wire [7:0] p1_array_index_2043926_comb;
  wire [7:0] p1_array_index_2043927_comb;
  wire [7:0] p1_array_index_2043928_comb;
  wire [7:0] p1_array_index_2043929_comb;
  wire [7:0] p1_array_index_2043930_comb;
  wire [7:0] p1_array_index_2043931_comb;
  wire [7:0] p1_array_index_2043933_comb;
  wire [7:0] p1_array_index_2043934_comb;
  wire [7:0] p1_array_index_2043935_comb;
  wire [7:0] p1_array_index_2043936_comb;
  wire [7:0] p1_array_index_2043937_comb;
  wire [7:0] p1_array_index_2043938_comb;
  wire [7:0] p1_array_index_2043939_comb;
  wire [7:0] p1_array_index_2043941_comb;
  wire [7:0] p1_res7_comb;
  wire [7:0] p1_array_index_2043950_comb;
  wire [7:0] p1_array_index_2043951_comb;
  wire [7:0] p1_array_index_2043952_comb;
  wire [7:0] p1_array_index_2043953_comb;
  wire [7:0] p1_array_index_2043954_comb;
  wire [7:0] p1_array_index_2043955_comb;
  wire [7:0] p1_res7__2_comb;
  wire [7:0] p1_array_index_2043965_comb;
  wire [7:0] p1_array_index_2043966_comb;
  wire [7:0] p1_array_index_2043967_comb;
  wire [7:0] p1_array_index_2043968_comb;
  wire [7:0] p1_array_index_2043969_comb;
  wire [7:0] p1_res7__4_comb;
  wire [7:0] p1_array_index_2043979_comb;
  wire [7:0] p1_array_index_2043980_comb;
  wire [7:0] p1_array_index_2043981_comb;
  wire [7:0] p1_array_index_2043982_comb;
  wire [7:0] p1_array_index_2043983_comb;
  wire [7:0] p1_res7__6_comb;
  wire [7:0] p1_array_index_2043994_comb;
  wire [7:0] p1_array_index_2043995_comb;
  wire [7:0] p1_array_index_2043996_comb;
  wire [7:0] p1_array_index_2043997_comb;
  wire [7:0] p1_res7__8_comb;
  wire [7:0] p1_array_index_2044007_comb;
  wire [7:0] p1_array_index_2044008_comb;
  wire [7:0] p1_array_index_2044009_comb;
  wire [7:0] p1_array_index_2044010_comb;
  wire [7:0] p1_res7__10_comb;
  wire [7:0] p1_array_index_2044021_comb;
  wire [7:0] p1_array_index_2044022_comb;
  wire [7:0] p1_array_index_2044023_comb;
  wire [7:0] p1_res7__12_comb;
  wire [7:0] p1_array_index_2044033_comb;
  wire [7:0] p1_array_index_2044034_comb;
  wire [7:0] p1_array_index_2044035_comb;
  wire [7:0] p1_res7__14_comb;
  wire [7:0] p1_array_index_2044046_comb;
  wire [7:0] p1_array_index_2044047_comb;
  wire [7:0] p1_res7__16_comb;
  wire [7:0] p1_array_index_2044057_comb;
  wire [7:0] p1_array_index_2044058_comb;
  wire [7:0] p1_res7__18_comb;
  wire [7:0] p1_array_index_2044069_comb;
  wire [7:0] p1_res7__20_comb;
  wire [7:0] p1_array_index_2044079_comb;
  wire [7:0] p1_res7__22_comb;
  wire [7:0] p1_res7__24_comb;
  wire [7:0] p1_res7__26_comb;
  wire [7:0] p1_res7__28_comb;
  wire [7:0] p1_res7__30_comb;
  wire [127:0] p1_res_comb;
  wire [127:0] p1_bit_slice_2044119_comb;
  wire [127:0] p1_xor_2044120_comb;
  wire [127:0] p1_addedKey__33_comb;
  wire [7:0] p1_array_index_2044136_comb;
  wire [7:0] p1_array_index_2044137_comb;
  wire [7:0] p1_array_index_2044138_comb;
  wire [7:0] p1_array_index_2044139_comb;
  wire [7:0] p1_array_index_2044140_comb;
  wire [7:0] p1_array_index_2044141_comb;
  wire [7:0] p1_array_index_2044143_comb;
  wire [7:0] p1_array_index_2044145_comb;
  wire [7:0] p1_array_index_2044146_comb;
  wire [7:0] p1_array_index_2044147_comb;
  wire [7:0] p1_array_index_2044148_comb;
  wire [7:0] p1_array_index_2044149_comb;
  wire [7:0] p1_array_index_2044150_comb;
  wire [7:0] p1_array_index_2044152_comb;
  wire [7:0] p1_array_index_2044153_comb;
  wire [7:0] p1_array_index_2044154_comb;
  wire [7:0] p1_array_index_2044155_comb;
  wire [7:0] p1_array_index_2044156_comb;
  wire [7:0] p1_array_index_2044157_comb;
  wire [7:0] p1_array_index_2044158_comb;
  wire [7:0] p1_array_index_2044160_comb;
  wire [7:0] p1_res7__32_comb;
  wire [7:0] p1_array_index_2044169_comb;
  wire [7:0] p1_array_index_2044170_comb;
  wire [7:0] p1_array_index_2044171_comb;
  wire [7:0] p1_array_index_2044172_comb;
  wire [7:0] p1_array_index_2044173_comb;
  wire [7:0] p1_array_index_2044174_comb;
  wire [7:0] p1_res7__34_comb;
  wire [7:0] p1_array_index_2044184_comb;
  wire [7:0] p1_array_index_2044185_comb;
  wire [7:0] p1_array_index_2044186_comb;
  wire [7:0] p1_array_index_2044187_comb;
  wire [7:0] p1_array_index_2044188_comb;
  wire [7:0] p1_res7__36_comb;
  wire [7:0] p1_array_index_2044198_comb;
  wire [7:0] p1_array_index_2044199_comb;
  wire [7:0] p1_array_index_2044200_comb;
  wire [7:0] p1_array_index_2044201_comb;
  wire [7:0] p1_array_index_2044202_comb;
  wire [7:0] p1_res7__38_comb;
  wire [7:0] p1_array_index_2044213_comb;
  wire [7:0] p1_array_index_2044214_comb;
  wire [7:0] p1_array_index_2044215_comb;
  wire [7:0] p1_array_index_2044216_comb;
  wire [7:0] p1_res7__40_comb;
  wire [7:0] p1_array_index_2044226_comb;
  wire [7:0] p1_array_index_2044227_comb;
  wire [7:0] p1_array_index_2044228_comb;
  wire [7:0] p1_array_index_2044229_comb;
  wire [7:0] p1_res7__42_comb;
  wire [7:0] p1_array_index_2044240_comb;
  wire [7:0] p1_array_index_2044241_comb;
  wire [7:0] p1_array_index_2044242_comb;
  wire [7:0] p1_res7__44_comb;
  wire [7:0] p1_array_index_2044252_comb;
  wire [7:0] p1_array_index_2044253_comb;
  wire [7:0] p1_array_index_2044254_comb;
  wire [7:0] p1_res7__46_comb;
  wire [7:0] p1_array_index_2044265_comb;
  wire [7:0] p1_array_index_2044266_comb;
  wire [7:0] p1_res7__48_comb;
  wire [7:0] p1_array_index_2044276_comb;
  wire [7:0] p1_array_index_2044277_comb;
  wire [7:0] p1_res7__50_comb;
  wire [7:0] p1_array_index_2044288_comb;
  wire [7:0] p1_res7__52_comb;
  wire [7:0] p1_array_index_2044298_comb;
  wire [7:0] p1_res7__54_comb;
  wire [7:0] p1_res7__56_comb;
  wire [7:0] p1_res7__58_comb;
  wire [7:0] p1_res7__60_comb;
  wire [7:0] p1_res7__62_comb;
  wire [127:0] p1_res__1_comb;
  wire [127:0] p1_xor_2044338_comb;
  wire [127:0] p1_addedKey__34_comb;
  wire [7:0] p1_array_index_2044354_comb;
  wire [7:0] p1_array_index_2044355_comb;
  wire [7:0] p1_array_index_2044356_comb;
  wire [7:0] p1_array_index_2044357_comb;
  wire [7:0] p1_array_index_2044358_comb;
  wire [7:0] p1_array_index_2044359_comb;
  wire [7:0] p1_array_index_2044361_comb;
  wire [7:0] p1_array_index_2044363_comb;
  wire [7:0] p1_array_index_2044364_comb;
  wire [7:0] p1_array_index_2044365_comb;
  wire [7:0] p1_array_index_2044366_comb;
  wire [7:0] p1_array_index_2044367_comb;
  wire [7:0] p1_array_index_2044368_comb;
  wire [7:0] p1_array_index_2044370_comb;
  wire [7:0] p1_array_index_2044371_comb;
  wire [7:0] p1_array_index_2044372_comb;
  wire [7:0] p1_array_index_2044373_comb;
  wire [7:0] p1_array_index_2044374_comb;
  wire [7:0] p1_array_index_2044375_comb;
  wire [7:0] p1_array_index_2044376_comb;
  wire [7:0] p1_array_index_2044378_comb;
  wire [7:0] p1_res7__64_comb;
  wire [7:0] p1_array_index_2044387_comb;
  wire [7:0] p1_array_index_2044388_comb;
  wire [7:0] p1_array_index_2044389_comb;
  wire [7:0] p1_array_index_2044390_comb;
  wire [7:0] p1_array_index_2044391_comb;
  wire [7:0] p1_array_index_2044392_comb;
  wire [7:0] p1_res7__66_comb;
  wire [7:0] p1_array_index_2044402_comb;
  wire [7:0] p1_array_index_2044403_comb;
  wire [7:0] p1_array_index_2044404_comb;
  wire [7:0] p1_array_index_2044405_comb;
  wire [7:0] p1_array_index_2044406_comb;
  wire [7:0] p1_res7__68_comb;
  wire [7:0] p1_array_index_2044416_comb;
  wire [7:0] p1_array_index_2044417_comb;
  wire [7:0] p1_array_index_2044418_comb;
  wire [7:0] p1_array_index_2044419_comb;
  wire [7:0] p1_array_index_2044420_comb;
  wire [7:0] p1_res7__70_comb;
  wire [7:0] p1_array_index_2044431_comb;
  wire [7:0] p1_array_index_2044432_comb;
  wire [7:0] p1_array_index_2044433_comb;
  wire [7:0] p1_array_index_2044434_comb;
  wire [7:0] p1_res7__72_comb;
  wire [7:0] p1_array_index_2044444_comb;
  wire [7:0] p1_array_index_2044445_comb;
  wire [7:0] p1_array_index_2044446_comb;
  wire [7:0] p1_array_index_2044447_comb;
  wire [7:0] p1_res7__74_comb;
  wire [7:0] p1_array_index_2044458_comb;
  wire [7:0] p1_array_index_2044459_comb;
  wire [7:0] p1_array_index_2044460_comb;
  wire [7:0] p1_res7__76_comb;
  wire [7:0] p1_array_index_2044470_comb;
  wire [7:0] p1_array_index_2044471_comb;
  wire [7:0] p1_array_index_2044472_comb;
  wire [7:0] p1_res7__78_comb;
  wire [7:0] p1_array_index_2044483_comb;
  wire [7:0] p1_array_index_2044484_comb;
  wire [7:0] p1_res7__80_comb;
  wire [7:0] p1_array_index_2044494_comb;
  wire [7:0] p1_array_index_2044495_comb;
  wire [7:0] p1_res7__82_comb;
  wire [7:0] p1_array_index_2044506_comb;
  wire [7:0] p1_res7__84_comb;
  wire [7:0] p1_array_index_2044516_comb;
  wire [7:0] p1_res7__86_comb;
  wire [7:0] p1_res7__88_comb;
  wire [7:0] p1_res7__90_comb;
  wire [7:0] p1_res7__92_comb;
  wire [7:0] p1_res7__94_comb;
  wire [127:0] p1_res__2_comb;
  wire [127:0] p1_xor_2044556_comb;
  wire [127:0] p1_addedKey__35_comb;
  wire [7:0] p1_array_index_2044572_comb;
  wire [7:0] p1_array_index_2044573_comb;
  wire [7:0] p1_array_index_2044574_comb;
  wire [7:0] p1_array_index_2044575_comb;
  wire [7:0] p1_array_index_2044576_comb;
  wire [7:0] p1_array_index_2044577_comb;
  wire [7:0] p1_array_index_2044579_comb;
  wire [7:0] p1_array_index_2044581_comb;
  wire [7:0] p1_array_index_2044582_comb;
  wire [7:0] p1_array_index_2044583_comb;
  wire [7:0] p1_array_index_2044584_comb;
  wire [7:0] p1_array_index_2044585_comb;
  wire [7:0] p1_array_index_2044586_comb;
  wire [7:0] p1_array_index_2044588_comb;
  wire [7:0] p1_array_index_2044589_comb;
  wire [7:0] p1_array_index_2044590_comb;
  wire [7:0] p1_array_index_2044591_comb;
  wire [7:0] p1_array_index_2044592_comb;
  wire [7:0] p1_array_index_2044593_comb;
  wire [7:0] p1_array_index_2044594_comb;
  wire [7:0] p1_array_index_2044596_comb;
  wire [7:0] p1_res7__96_comb;
  wire [7:0] p1_array_index_2044605_comb;
  wire [7:0] p1_array_index_2044606_comb;
  wire [7:0] p1_array_index_2044607_comb;
  wire [7:0] p1_array_index_2044608_comb;
  wire [7:0] p1_array_index_2044609_comb;
  wire [7:0] p1_array_index_2044610_comb;
  wire [7:0] p1_res7__98_comb;
  wire [7:0] p1_array_index_2044620_comb;
  wire [7:0] p1_array_index_2044621_comb;
  wire [7:0] p1_array_index_2044622_comb;
  wire [7:0] p1_array_index_2044623_comb;
  wire [7:0] p1_array_index_2044624_comb;
  wire [7:0] p1_res7__100_comb;
  wire [7:0] p1_array_index_2044634_comb;
  wire [7:0] p1_array_index_2044635_comb;
  wire [7:0] p1_array_index_2044636_comb;
  wire [7:0] p1_array_index_2044637_comb;
  wire [7:0] p1_array_index_2044638_comb;
  wire [7:0] p1_res7__102_comb;
  wire [7:0] p1_array_index_2044649_comb;
  wire [7:0] p1_array_index_2044650_comb;
  wire [7:0] p1_array_index_2044651_comb;
  wire [7:0] p1_array_index_2044652_comb;
  wire [7:0] p1_res7__104_comb;
  wire [7:0] p1_array_index_2044662_comb;
  wire [7:0] p1_array_index_2044663_comb;
  wire [7:0] p1_array_index_2044664_comb;
  wire [7:0] p1_array_index_2044665_comb;
  wire [7:0] p1_res7__106_comb;
  wire [7:0] p1_array_index_2044676_comb;
  wire [7:0] p1_array_index_2044677_comb;
  wire [7:0] p1_array_index_2044678_comb;
  wire [7:0] p1_res7__108_comb;
  wire [7:0] p1_array_index_2044688_comb;
  wire [7:0] p1_array_index_2044689_comb;
  wire [7:0] p1_array_index_2044690_comb;
  wire [7:0] p1_res7__110_comb;
  wire [7:0] p1_array_index_2044701_comb;
  wire [7:0] p1_array_index_2044702_comb;
  wire [7:0] p1_res7__112_comb;
  wire [7:0] p1_array_index_2044712_comb;
  wire [7:0] p1_array_index_2044713_comb;
  wire [7:0] p1_res7__114_comb;
  wire [7:0] p1_array_index_2044724_comb;
  wire [7:0] p1_res7__116_comb;
  wire [7:0] p1_array_index_2044734_comb;
  wire [7:0] p1_res7__118_comb;
  wire [7:0] p1_res7__120_comb;
  wire [7:0] p1_res7__122_comb;
  wire [7:0] p1_res7__124_comb;
  wire [7:0] p1_res7__126_comb;
  wire [127:0] p1_res__3_comb;
  wire [127:0] p1_xor_2044774_comb;
  wire [127:0] p1_addedKey__36_comb;
  wire [7:0] p1_array_index_2044790_comb;
  wire [7:0] p1_array_index_2044791_comb;
  wire [7:0] p1_array_index_2044792_comb;
  wire [7:0] p1_array_index_2044793_comb;
  wire [7:0] p1_array_index_2044794_comb;
  wire [7:0] p1_array_index_2044795_comb;
  wire [7:0] p1_array_index_2044797_comb;
  wire [7:0] p1_array_index_2044799_comb;
  wire [7:0] p1_array_index_2044800_comb;
  wire [7:0] p1_array_index_2044801_comb;
  wire [7:0] p1_array_index_2044802_comb;
  wire [7:0] p1_array_index_2044803_comb;
  wire [7:0] p1_array_index_2044804_comb;
  wire [7:0] p1_array_index_2044806_comb;
  wire [7:0] p1_array_index_2044807_comb;
  wire [7:0] p1_array_index_2044808_comb;
  wire [7:0] p1_array_index_2044809_comb;
  wire [7:0] p1_array_index_2044810_comb;
  wire [7:0] p1_array_index_2044811_comb;
  wire [7:0] p1_array_index_2044812_comb;
  wire [7:0] p1_array_index_2044814_comb;
  wire [7:0] p1_res7__128_comb;
  wire [7:0] p1_array_index_2044823_comb;
  wire [7:0] p1_array_index_2044824_comb;
  wire [7:0] p1_array_index_2044825_comb;
  wire [7:0] p1_array_index_2044826_comb;
  wire [7:0] p1_array_index_2044827_comb;
  wire [7:0] p1_array_index_2044828_comb;
  wire [7:0] p1_res7__130_comb;
  wire [7:0] p1_array_index_2044838_comb;
  wire [7:0] p1_array_index_2044839_comb;
  wire [7:0] p1_array_index_2044840_comb;
  wire [7:0] p1_array_index_2044841_comb;
  wire [7:0] p1_array_index_2044842_comb;
  wire [7:0] p1_res7__132_comb;
  wire [7:0] p1_array_index_2044852_comb;
  wire [7:0] p1_array_index_2044853_comb;
  wire [7:0] p1_array_index_2044854_comb;
  wire [7:0] p1_array_index_2044855_comb;
  wire [7:0] p1_array_index_2044856_comb;
  wire [7:0] p1_res7__134_comb;
  wire [7:0] p1_array_index_2044867_comb;
  wire [7:0] p1_array_index_2044868_comb;
  wire [7:0] p1_array_index_2044869_comb;
  wire [7:0] p1_array_index_2044870_comb;
  wire [7:0] p1_res7__136_comb;
  wire [7:0] p1_array_index_2044880_comb;
  wire [7:0] p1_array_index_2044881_comb;
  wire [7:0] p1_array_index_2044882_comb;
  wire [7:0] p1_array_index_2044883_comb;
  wire [7:0] p1_res7__138_comb;
  wire [7:0] p1_array_index_2044894_comb;
  wire [7:0] p1_array_index_2044895_comb;
  wire [7:0] p1_array_index_2044896_comb;
  wire [7:0] p1_res7__140_comb;
  assign p1_bit_slice_2043893_comb = p0_key[255:128];
  assign p1_addedKey__32_comb = p1_bit_slice_2043893_comb ^ 128'h6ea2_7672_6c48_7ab8_5d27_bd10_dd84_9401;
  assign p1_array_index_2043911_comb = literal_2043896[p1_addedKey__32_comb[127:120]];
  assign p1_array_index_2043913_comb = literal_2043896[p1_addedKey__32_comb[119:112]];
  assign p1_array_index_2043915_comb = literal_2043896[p1_addedKey__32_comb[111:104]];
  assign p1_array_index_2043917_comb = literal_2043896[p1_addedKey__32_comb[103:96]];
  assign p1_array_index_2043919_comb = literal_2043896[p1_addedKey__32_comb[95:88]];
  assign p1_array_index_2043921_comb = literal_2043896[p1_addedKey__32_comb[87:80]];
  assign p1_array_index_2043924_comb = literal_2043896[p1_addedKey__32_comb[71:64]];
  assign p1_array_index_2043926_comb = literal_2043896[p1_addedKey__32_comb[55:48]];
  assign p1_array_index_2043927_comb = literal_2043896[p1_addedKey__32_comb[47:40]];
  assign p1_array_index_2043928_comb = literal_2043896[p1_addedKey__32_comb[39:32]];
  assign p1_array_index_2043929_comb = literal_2043896[p1_addedKey__32_comb[31:24]];
  assign p1_array_index_2043930_comb = literal_2043896[p1_addedKey__32_comb[23:16]];
  assign p1_array_index_2043931_comb = literal_2043896[p1_addedKey__32_comb[15:8]];
  assign p1_array_index_2043933_comb = literal_2043910[p1_array_index_2043911_comb];
  assign p1_array_index_2043934_comb = literal_2043912[p1_array_index_2043913_comb];
  assign p1_array_index_2043935_comb = literal_2043914[p1_array_index_2043915_comb];
  assign p1_array_index_2043936_comb = literal_2043916[p1_array_index_2043917_comb];
  assign p1_array_index_2043937_comb = literal_2043918[p1_array_index_2043919_comb];
  assign p1_array_index_2043938_comb = literal_2043920[p1_array_index_2043921_comb];
  assign p1_array_index_2043939_comb = literal_2043896[p1_addedKey__32_comb[79:72]];
  assign p1_array_index_2043941_comb = literal_2043896[p1_addedKey__32_comb[63:56]];
  assign p1_res7_comb = p1_array_index_2043933_comb ^ p1_array_index_2043934_comb ^ p1_array_index_2043935_comb ^ p1_array_index_2043936_comb ^ p1_array_index_2043937_comb ^ p1_array_index_2043938_comb ^ p1_array_index_2043939_comb ^ literal_2043923[p1_array_index_2043924_comb] ^ p1_array_index_2043941_comb ^ literal_2043920[p1_array_index_2043926_comb] ^ literal_2043918[p1_array_index_2043927_comb] ^ literal_2043916[p1_array_index_2043928_comb] ^ literal_2043914[p1_array_index_2043929_comb] ^ literal_2043912[p1_array_index_2043930_comb] ^ literal_2043910[p1_array_index_2043931_comb] ^ literal_2043896[p1_addedKey__32_comb[7:0]];
  assign p1_array_index_2043950_comb = literal_2043910[p1_res7_comb];
  assign p1_array_index_2043951_comb = literal_2043912[p1_array_index_2043911_comb];
  assign p1_array_index_2043952_comb = literal_2043914[p1_array_index_2043913_comb];
  assign p1_array_index_2043953_comb = literal_2043916[p1_array_index_2043915_comb];
  assign p1_array_index_2043954_comb = literal_2043918[p1_array_index_2043917_comb];
  assign p1_array_index_2043955_comb = literal_2043920[p1_array_index_2043919_comb];
  assign p1_res7__2_comb = p1_array_index_2043950_comb ^ p1_array_index_2043951_comb ^ p1_array_index_2043952_comb ^ p1_array_index_2043953_comb ^ p1_array_index_2043954_comb ^ p1_array_index_2043955_comb ^ p1_array_index_2043921_comb ^ literal_2043923[p1_array_index_2043939_comb] ^ p1_array_index_2043924_comb ^ literal_2043920[p1_array_index_2043941_comb] ^ literal_2043918[p1_array_index_2043926_comb] ^ literal_2043916[p1_array_index_2043927_comb] ^ literal_2043914[p1_array_index_2043928_comb] ^ literal_2043912[p1_array_index_2043929_comb] ^ literal_2043910[p1_array_index_2043930_comb] ^ p1_array_index_2043931_comb;
  assign p1_array_index_2043965_comb = literal_2043912[p1_res7_comb];
  assign p1_array_index_2043966_comb = literal_2043914[p1_array_index_2043911_comb];
  assign p1_array_index_2043967_comb = literal_2043916[p1_array_index_2043913_comb];
  assign p1_array_index_2043968_comb = literal_2043918[p1_array_index_2043915_comb];
  assign p1_array_index_2043969_comb = literal_2043920[p1_array_index_2043917_comb];
  assign p1_res7__4_comb = literal_2043910[p1_res7__2_comb] ^ p1_array_index_2043965_comb ^ p1_array_index_2043966_comb ^ p1_array_index_2043967_comb ^ p1_array_index_2043968_comb ^ p1_array_index_2043969_comb ^ p1_array_index_2043919_comb ^ literal_2043923[p1_array_index_2043921_comb] ^ p1_array_index_2043939_comb ^ literal_2043920[p1_array_index_2043924_comb] ^ literal_2043918[p1_array_index_2043941_comb] ^ literal_2043916[p1_array_index_2043926_comb] ^ literal_2043914[p1_array_index_2043927_comb] ^ literal_2043912[p1_array_index_2043928_comb] ^ literal_2043910[p1_array_index_2043929_comb] ^ p1_array_index_2043930_comb;
  assign p1_array_index_2043979_comb = literal_2043912[p1_res7__2_comb];
  assign p1_array_index_2043980_comb = literal_2043914[p1_res7_comb];
  assign p1_array_index_2043981_comb = literal_2043916[p1_array_index_2043911_comb];
  assign p1_array_index_2043982_comb = literal_2043918[p1_array_index_2043913_comb];
  assign p1_array_index_2043983_comb = literal_2043920[p1_array_index_2043915_comb];
  assign p1_res7__6_comb = literal_2043910[p1_res7__4_comb] ^ p1_array_index_2043979_comb ^ p1_array_index_2043980_comb ^ p1_array_index_2043981_comb ^ p1_array_index_2043982_comb ^ p1_array_index_2043983_comb ^ p1_array_index_2043917_comb ^ literal_2043923[p1_array_index_2043919_comb] ^ p1_array_index_2043921_comb ^ literal_2043920[p1_array_index_2043939_comb] ^ literal_2043918[p1_array_index_2043924_comb] ^ literal_2043916[p1_array_index_2043941_comb] ^ literal_2043914[p1_array_index_2043926_comb] ^ literal_2043912[p1_array_index_2043927_comb] ^ literal_2043910[p1_array_index_2043928_comb] ^ p1_array_index_2043929_comb;
  assign p1_array_index_2043994_comb = literal_2043914[p1_res7__2_comb];
  assign p1_array_index_2043995_comb = literal_2043916[p1_res7_comb];
  assign p1_array_index_2043996_comb = literal_2043918[p1_array_index_2043911_comb];
  assign p1_array_index_2043997_comb = literal_2043920[p1_array_index_2043913_comb];
  assign p1_res7__8_comb = literal_2043910[p1_res7__6_comb] ^ literal_2043912[p1_res7__4_comb] ^ p1_array_index_2043994_comb ^ p1_array_index_2043995_comb ^ p1_array_index_2043996_comb ^ p1_array_index_2043997_comb ^ p1_array_index_2043915_comb ^ literal_2043923[p1_array_index_2043917_comb] ^ p1_array_index_2043919_comb ^ p1_array_index_2043938_comb ^ literal_2043918[p1_array_index_2043939_comb] ^ literal_2043916[p1_array_index_2043924_comb] ^ literal_2043914[p1_array_index_2043941_comb] ^ literal_2043912[p1_array_index_2043926_comb] ^ literal_2043910[p1_array_index_2043927_comb] ^ p1_array_index_2043928_comb;
  assign p1_array_index_2044007_comb = literal_2043914[p1_res7__4_comb];
  assign p1_array_index_2044008_comb = literal_2043916[p1_res7__2_comb];
  assign p1_array_index_2044009_comb = literal_2043918[p1_res7_comb];
  assign p1_array_index_2044010_comb = literal_2043920[p1_array_index_2043911_comb];
  assign p1_res7__10_comb = literal_2043910[p1_res7__8_comb] ^ literal_2043912[p1_res7__6_comb] ^ p1_array_index_2044007_comb ^ p1_array_index_2044008_comb ^ p1_array_index_2044009_comb ^ p1_array_index_2044010_comb ^ p1_array_index_2043913_comb ^ literal_2043923[p1_array_index_2043915_comb] ^ p1_array_index_2043917_comb ^ p1_array_index_2043955_comb ^ literal_2043918[p1_array_index_2043921_comb] ^ literal_2043916[p1_array_index_2043939_comb] ^ literal_2043914[p1_array_index_2043924_comb] ^ literal_2043912[p1_array_index_2043941_comb] ^ literal_2043910[p1_array_index_2043926_comb] ^ p1_array_index_2043927_comb;
  assign p1_array_index_2044021_comb = literal_2043916[p1_res7__4_comb];
  assign p1_array_index_2044022_comb = literal_2043918[p1_res7__2_comb];
  assign p1_array_index_2044023_comb = literal_2043920[p1_res7_comb];
  assign p1_res7__12_comb = literal_2043910[p1_res7__10_comb] ^ literal_2043912[p1_res7__8_comb] ^ literal_2043914[p1_res7__6_comb] ^ p1_array_index_2044021_comb ^ p1_array_index_2044022_comb ^ p1_array_index_2044023_comb ^ p1_array_index_2043911_comb ^ literal_2043923[p1_array_index_2043913_comb] ^ p1_array_index_2043915_comb ^ p1_array_index_2043969_comb ^ p1_array_index_2043937_comb ^ literal_2043916[p1_array_index_2043921_comb] ^ literal_2043914[p1_array_index_2043939_comb] ^ literal_2043912[p1_array_index_2043924_comb] ^ literal_2043910[p1_array_index_2043941_comb] ^ p1_array_index_2043926_comb;
  assign p1_array_index_2044033_comb = literal_2043916[p1_res7__6_comb];
  assign p1_array_index_2044034_comb = literal_2043918[p1_res7__4_comb];
  assign p1_array_index_2044035_comb = literal_2043920[p1_res7__2_comb];
  assign p1_res7__14_comb = literal_2043910[p1_res7__12_comb] ^ literal_2043912[p1_res7__10_comb] ^ literal_2043914[p1_res7__8_comb] ^ p1_array_index_2044033_comb ^ p1_array_index_2044034_comb ^ p1_array_index_2044035_comb ^ p1_res7_comb ^ literal_2043923[p1_array_index_2043911_comb] ^ p1_array_index_2043913_comb ^ p1_array_index_2043983_comb ^ p1_array_index_2043954_comb ^ literal_2043916[p1_array_index_2043919_comb] ^ literal_2043914[p1_array_index_2043921_comb] ^ literal_2043912[p1_array_index_2043939_comb] ^ literal_2043910[p1_array_index_2043924_comb] ^ p1_array_index_2043941_comb;
  assign p1_array_index_2044046_comb = literal_2043918[p1_res7__6_comb];
  assign p1_array_index_2044047_comb = literal_2043920[p1_res7__4_comb];
  assign p1_res7__16_comb = literal_2043910[p1_res7__14_comb] ^ literal_2043912[p1_res7__12_comb] ^ literal_2043914[p1_res7__10_comb] ^ literal_2043916[p1_res7__8_comb] ^ p1_array_index_2044046_comb ^ p1_array_index_2044047_comb ^ p1_res7__2_comb ^ literal_2043923[p1_res7_comb] ^ p1_array_index_2043911_comb ^ p1_array_index_2043997_comb ^ p1_array_index_2043968_comb ^ p1_array_index_2043936_comb ^ literal_2043914[p1_array_index_2043919_comb] ^ literal_2043912[p1_array_index_2043921_comb] ^ literal_2043910[p1_array_index_2043939_comb] ^ p1_array_index_2043924_comb;
  assign p1_array_index_2044057_comb = literal_2043918[p1_res7__8_comb];
  assign p1_array_index_2044058_comb = literal_2043920[p1_res7__6_comb];
  assign p1_res7__18_comb = literal_2043910[p1_res7__16_comb] ^ literal_2043912[p1_res7__14_comb] ^ literal_2043914[p1_res7__12_comb] ^ literal_2043916[p1_res7__10_comb] ^ p1_array_index_2044057_comb ^ p1_array_index_2044058_comb ^ p1_res7__4_comb ^ literal_2043923[p1_res7__2_comb] ^ p1_res7_comb ^ p1_array_index_2044010_comb ^ p1_array_index_2043982_comb ^ p1_array_index_2043953_comb ^ literal_2043914[p1_array_index_2043917_comb] ^ literal_2043912[p1_array_index_2043919_comb] ^ literal_2043910[p1_array_index_2043921_comb] ^ p1_array_index_2043939_comb;
  assign p1_array_index_2044069_comb = literal_2043920[p1_res7__8_comb];
  assign p1_res7__20_comb = literal_2043910[p1_res7__18_comb] ^ literal_2043912[p1_res7__16_comb] ^ literal_2043914[p1_res7__14_comb] ^ literal_2043916[p1_res7__12_comb] ^ literal_2043918[p1_res7__10_comb] ^ p1_array_index_2044069_comb ^ p1_res7__6_comb ^ literal_2043923[p1_res7__4_comb] ^ p1_res7__2_comb ^ p1_array_index_2044023_comb ^ p1_array_index_2043996_comb ^ p1_array_index_2043967_comb ^ p1_array_index_2043935_comb ^ literal_2043912[p1_array_index_2043917_comb] ^ literal_2043910[p1_array_index_2043919_comb] ^ p1_array_index_2043921_comb;
  assign p1_array_index_2044079_comb = literal_2043920[p1_res7__10_comb];
  assign p1_res7__22_comb = literal_2043910[p1_res7__20_comb] ^ literal_2043912[p1_res7__18_comb] ^ literal_2043914[p1_res7__16_comb] ^ literal_2043916[p1_res7__14_comb] ^ literal_2043918[p1_res7__12_comb] ^ p1_array_index_2044079_comb ^ p1_res7__8_comb ^ literal_2043923[p1_res7__6_comb] ^ p1_res7__4_comb ^ p1_array_index_2044035_comb ^ p1_array_index_2044009_comb ^ p1_array_index_2043981_comb ^ p1_array_index_2043952_comb ^ literal_2043912[p1_array_index_2043915_comb] ^ literal_2043910[p1_array_index_2043917_comb] ^ p1_array_index_2043919_comb;
  assign p1_res7__24_comb = literal_2043910[p1_res7__22_comb] ^ literal_2043912[p1_res7__20_comb] ^ literal_2043914[p1_res7__18_comb] ^ literal_2043916[p1_res7__16_comb] ^ literal_2043918[p1_res7__14_comb] ^ literal_2043920[p1_res7__12_comb] ^ p1_res7__10_comb ^ literal_2043923[p1_res7__8_comb] ^ p1_res7__6_comb ^ p1_array_index_2044047_comb ^ p1_array_index_2044022_comb ^ p1_array_index_2043995_comb ^ p1_array_index_2043966_comb ^ p1_array_index_2043934_comb ^ literal_2043910[p1_array_index_2043915_comb] ^ p1_array_index_2043917_comb;
  assign p1_res7__26_comb = literal_2043910[p1_res7__24_comb] ^ literal_2043912[p1_res7__22_comb] ^ literal_2043914[p1_res7__20_comb] ^ literal_2043916[p1_res7__18_comb] ^ literal_2043918[p1_res7__16_comb] ^ literal_2043920[p1_res7__14_comb] ^ p1_res7__12_comb ^ literal_2043923[p1_res7__10_comb] ^ p1_res7__8_comb ^ p1_array_index_2044058_comb ^ p1_array_index_2044034_comb ^ p1_array_index_2044008_comb ^ p1_array_index_2043980_comb ^ p1_array_index_2043951_comb ^ literal_2043910[p1_array_index_2043913_comb] ^ p1_array_index_2043915_comb;
  assign p1_res7__28_comb = literal_2043910[p1_res7__26_comb] ^ literal_2043912[p1_res7__24_comb] ^ literal_2043914[p1_res7__22_comb] ^ literal_2043916[p1_res7__20_comb] ^ literal_2043918[p1_res7__18_comb] ^ literal_2043920[p1_res7__16_comb] ^ p1_res7__14_comb ^ literal_2043923[p1_res7__12_comb] ^ p1_res7__10_comb ^ p1_array_index_2044069_comb ^ p1_array_index_2044046_comb ^ p1_array_index_2044021_comb ^ p1_array_index_2043994_comb ^ p1_array_index_2043965_comb ^ p1_array_index_2043933_comb ^ p1_array_index_2043913_comb;
  assign p1_res7__30_comb = literal_2043910[p1_res7__28_comb] ^ literal_2043912[p1_res7__26_comb] ^ literal_2043914[p1_res7__24_comb] ^ literal_2043916[p1_res7__22_comb] ^ literal_2043918[p1_res7__20_comb] ^ literal_2043920[p1_res7__18_comb] ^ p1_res7__16_comb ^ literal_2043923[p1_res7__14_comb] ^ p1_res7__12_comb ^ p1_array_index_2044079_comb ^ p1_array_index_2044057_comb ^ p1_array_index_2044033_comb ^ p1_array_index_2044007_comb ^ p1_array_index_2043979_comb ^ p1_array_index_2043950_comb ^ p1_array_index_2043911_comb;
  assign p1_res_comb = {p1_res7__30_comb, p1_res7__28_comb, p1_res7__26_comb, p1_res7__24_comb, p1_res7__22_comb, p1_res7__20_comb, p1_res7__18_comb, p1_res7__16_comb, p1_res7__14_comb, p1_res7__12_comb, p1_res7__10_comb, p1_res7__8_comb, p1_res7__6_comb, p1_res7__4_comb, p1_res7__2_comb, p1_res7_comb};
  assign p1_bit_slice_2044119_comb = p0_key[127:0];
  assign p1_xor_2044120_comb = p1_res_comb ^ p1_bit_slice_2044119_comb;
  assign p1_addedKey__33_comb = p1_xor_2044120_comb ^ 128'hdc87_ece4_d890_f4b3_ba4e_b920_79cb_eb02;
  assign p1_array_index_2044136_comb = literal_2043896[p1_addedKey__33_comb[127:120]];
  assign p1_array_index_2044137_comb = literal_2043896[p1_addedKey__33_comb[119:112]];
  assign p1_array_index_2044138_comb = literal_2043896[p1_addedKey__33_comb[111:104]];
  assign p1_array_index_2044139_comb = literal_2043896[p1_addedKey__33_comb[103:96]];
  assign p1_array_index_2044140_comb = literal_2043896[p1_addedKey__33_comb[95:88]];
  assign p1_array_index_2044141_comb = literal_2043896[p1_addedKey__33_comb[87:80]];
  assign p1_array_index_2044143_comb = literal_2043896[p1_addedKey__33_comb[71:64]];
  assign p1_array_index_2044145_comb = literal_2043896[p1_addedKey__33_comb[55:48]];
  assign p1_array_index_2044146_comb = literal_2043896[p1_addedKey__33_comb[47:40]];
  assign p1_array_index_2044147_comb = literal_2043896[p1_addedKey__33_comb[39:32]];
  assign p1_array_index_2044148_comb = literal_2043896[p1_addedKey__33_comb[31:24]];
  assign p1_array_index_2044149_comb = literal_2043896[p1_addedKey__33_comb[23:16]];
  assign p1_array_index_2044150_comb = literal_2043896[p1_addedKey__33_comb[15:8]];
  assign p1_array_index_2044152_comb = literal_2043910[p1_array_index_2044136_comb];
  assign p1_array_index_2044153_comb = literal_2043912[p1_array_index_2044137_comb];
  assign p1_array_index_2044154_comb = literal_2043914[p1_array_index_2044138_comb];
  assign p1_array_index_2044155_comb = literal_2043916[p1_array_index_2044139_comb];
  assign p1_array_index_2044156_comb = literal_2043918[p1_array_index_2044140_comb];
  assign p1_array_index_2044157_comb = literal_2043920[p1_array_index_2044141_comb];
  assign p1_array_index_2044158_comb = literal_2043896[p1_addedKey__33_comb[79:72]];
  assign p1_array_index_2044160_comb = literal_2043896[p1_addedKey__33_comb[63:56]];
  assign p1_res7__32_comb = p1_array_index_2044152_comb ^ p1_array_index_2044153_comb ^ p1_array_index_2044154_comb ^ p1_array_index_2044155_comb ^ p1_array_index_2044156_comb ^ p1_array_index_2044157_comb ^ p1_array_index_2044158_comb ^ literal_2043923[p1_array_index_2044143_comb] ^ p1_array_index_2044160_comb ^ literal_2043920[p1_array_index_2044145_comb] ^ literal_2043918[p1_array_index_2044146_comb] ^ literal_2043916[p1_array_index_2044147_comb] ^ literal_2043914[p1_array_index_2044148_comb] ^ literal_2043912[p1_array_index_2044149_comb] ^ literal_2043910[p1_array_index_2044150_comb] ^ literal_2043896[p1_addedKey__33_comb[7:0]];
  assign p1_array_index_2044169_comb = literal_2043910[p1_res7__32_comb];
  assign p1_array_index_2044170_comb = literal_2043912[p1_array_index_2044136_comb];
  assign p1_array_index_2044171_comb = literal_2043914[p1_array_index_2044137_comb];
  assign p1_array_index_2044172_comb = literal_2043916[p1_array_index_2044138_comb];
  assign p1_array_index_2044173_comb = literal_2043918[p1_array_index_2044139_comb];
  assign p1_array_index_2044174_comb = literal_2043920[p1_array_index_2044140_comb];
  assign p1_res7__34_comb = p1_array_index_2044169_comb ^ p1_array_index_2044170_comb ^ p1_array_index_2044171_comb ^ p1_array_index_2044172_comb ^ p1_array_index_2044173_comb ^ p1_array_index_2044174_comb ^ p1_array_index_2044141_comb ^ literal_2043923[p1_array_index_2044158_comb] ^ p1_array_index_2044143_comb ^ literal_2043920[p1_array_index_2044160_comb] ^ literal_2043918[p1_array_index_2044145_comb] ^ literal_2043916[p1_array_index_2044146_comb] ^ literal_2043914[p1_array_index_2044147_comb] ^ literal_2043912[p1_array_index_2044148_comb] ^ literal_2043910[p1_array_index_2044149_comb] ^ p1_array_index_2044150_comb;
  assign p1_array_index_2044184_comb = literal_2043912[p1_res7__32_comb];
  assign p1_array_index_2044185_comb = literal_2043914[p1_array_index_2044136_comb];
  assign p1_array_index_2044186_comb = literal_2043916[p1_array_index_2044137_comb];
  assign p1_array_index_2044187_comb = literal_2043918[p1_array_index_2044138_comb];
  assign p1_array_index_2044188_comb = literal_2043920[p1_array_index_2044139_comb];
  assign p1_res7__36_comb = literal_2043910[p1_res7__34_comb] ^ p1_array_index_2044184_comb ^ p1_array_index_2044185_comb ^ p1_array_index_2044186_comb ^ p1_array_index_2044187_comb ^ p1_array_index_2044188_comb ^ p1_array_index_2044140_comb ^ literal_2043923[p1_array_index_2044141_comb] ^ p1_array_index_2044158_comb ^ literal_2043920[p1_array_index_2044143_comb] ^ literal_2043918[p1_array_index_2044160_comb] ^ literal_2043916[p1_array_index_2044145_comb] ^ literal_2043914[p1_array_index_2044146_comb] ^ literal_2043912[p1_array_index_2044147_comb] ^ literal_2043910[p1_array_index_2044148_comb] ^ p1_array_index_2044149_comb;
  assign p1_array_index_2044198_comb = literal_2043912[p1_res7__34_comb];
  assign p1_array_index_2044199_comb = literal_2043914[p1_res7__32_comb];
  assign p1_array_index_2044200_comb = literal_2043916[p1_array_index_2044136_comb];
  assign p1_array_index_2044201_comb = literal_2043918[p1_array_index_2044137_comb];
  assign p1_array_index_2044202_comb = literal_2043920[p1_array_index_2044138_comb];
  assign p1_res7__38_comb = literal_2043910[p1_res7__36_comb] ^ p1_array_index_2044198_comb ^ p1_array_index_2044199_comb ^ p1_array_index_2044200_comb ^ p1_array_index_2044201_comb ^ p1_array_index_2044202_comb ^ p1_array_index_2044139_comb ^ literal_2043923[p1_array_index_2044140_comb] ^ p1_array_index_2044141_comb ^ literal_2043920[p1_array_index_2044158_comb] ^ literal_2043918[p1_array_index_2044143_comb] ^ literal_2043916[p1_array_index_2044160_comb] ^ literal_2043914[p1_array_index_2044145_comb] ^ literal_2043912[p1_array_index_2044146_comb] ^ literal_2043910[p1_array_index_2044147_comb] ^ p1_array_index_2044148_comb;
  assign p1_array_index_2044213_comb = literal_2043914[p1_res7__34_comb];
  assign p1_array_index_2044214_comb = literal_2043916[p1_res7__32_comb];
  assign p1_array_index_2044215_comb = literal_2043918[p1_array_index_2044136_comb];
  assign p1_array_index_2044216_comb = literal_2043920[p1_array_index_2044137_comb];
  assign p1_res7__40_comb = literal_2043910[p1_res7__38_comb] ^ literal_2043912[p1_res7__36_comb] ^ p1_array_index_2044213_comb ^ p1_array_index_2044214_comb ^ p1_array_index_2044215_comb ^ p1_array_index_2044216_comb ^ p1_array_index_2044138_comb ^ literal_2043923[p1_array_index_2044139_comb] ^ p1_array_index_2044140_comb ^ p1_array_index_2044157_comb ^ literal_2043918[p1_array_index_2044158_comb] ^ literal_2043916[p1_array_index_2044143_comb] ^ literal_2043914[p1_array_index_2044160_comb] ^ literal_2043912[p1_array_index_2044145_comb] ^ literal_2043910[p1_array_index_2044146_comb] ^ p1_array_index_2044147_comb;
  assign p1_array_index_2044226_comb = literal_2043914[p1_res7__36_comb];
  assign p1_array_index_2044227_comb = literal_2043916[p1_res7__34_comb];
  assign p1_array_index_2044228_comb = literal_2043918[p1_res7__32_comb];
  assign p1_array_index_2044229_comb = literal_2043920[p1_array_index_2044136_comb];
  assign p1_res7__42_comb = literal_2043910[p1_res7__40_comb] ^ literal_2043912[p1_res7__38_comb] ^ p1_array_index_2044226_comb ^ p1_array_index_2044227_comb ^ p1_array_index_2044228_comb ^ p1_array_index_2044229_comb ^ p1_array_index_2044137_comb ^ literal_2043923[p1_array_index_2044138_comb] ^ p1_array_index_2044139_comb ^ p1_array_index_2044174_comb ^ literal_2043918[p1_array_index_2044141_comb] ^ literal_2043916[p1_array_index_2044158_comb] ^ literal_2043914[p1_array_index_2044143_comb] ^ literal_2043912[p1_array_index_2044160_comb] ^ literal_2043910[p1_array_index_2044145_comb] ^ p1_array_index_2044146_comb;
  assign p1_array_index_2044240_comb = literal_2043916[p1_res7__36_comb];
  assign p1_array_index_2044241_comb = literal_2043918[p1_res7__34_comb];
  assign p1_array_index_2044242_comb = literal_2043920[p1_res7__32_comb];
  assign p1_res7__44_comb = literal_2043910[p1_res7__42_comb] ^ literal_2043912[p1_res7__40_comb] ^ literal_2043914[p1_res7__38_comb] ^ p1_array_index_2044240_comb ^ p1_array_index_2044241_comb ^ p1_array_index_2044242_comb ^ p1_array_index_2044136_comb ^ literal_2043923[p1_array_index_2044137_comb] ^ p1_array_index_2044138_comb ^ p1_array_index_2044188_comb ^ p1_array_index_2044156_comb ^ literal_2043916[p1_array_index_2044141_comb] ^ literal_2043914[p1_array_index_2044158_comb] ^ literal_2043912[p1_array_index_2044143_comb] ^ literal_2043910[p1_array_index_2044160_comb] ^ p1_array_index_2044145_comb;
  assign p1_array_index_2044252_comb = literal_2043916[p1_res7__38_comb];
  assign p1_array_index_2044253_comb = literal_2043918[p1_res7__36_comb];
  assign p1_array_index_2044254_comb = literal_2043920[p1_res7__34_comb];
  assign p1_res7__46_comb = literal_2043910[p1_res7__44_comb] ^ literal_2043912[p1_res7__42_comb] ^ literal_2043914[p1_res7__40_comb] ^ p1_array_index_2044252_comb ^ p1_array_index_2044253_comb ^ p1_array_index_2044254_comb ^ p1_res7__32_comb ^ literal_2043923[p1_array_index_2044136_comb] ^ p1_array_index_2044137_comb ^ p1_array_index_2044202_comb ^ p1_array_index_2044173_comb ^ literal_2043916[p1_array_index_2044140_comb] ^ literal_2043914[p1_array_index_2044141_comb] ^ literal_2043912[p1_array_index_2044158_comb] ^ literal_2043910[p1_array_index_2044143_comb] ^ p1_array_index_2044160_comb;
  assign p1_array_index_2044265_comb = literal_2043918[p1_res7__38_comb];
  assign p1_array_index_2044266_comb = literal_2043920[p1_res7__36_comb];
  assign p1_res7__48_comb = literal_2043910[p1_res7__46_comb] ^ literal_2043912[p1_res7__44_comb] ^ literal_2043914[p1_res7__42_comb] ^ literal_2043916[p1_res7__40_comb] ^ p1_array_index_2044265_comb ^ p1_array_index_2044266_comb ^ p1_res7__34_comb ^ literal_2043923[p1_res7__32_comb] ^ p1_array_index_2044136_comb ^ p1_array_index_2044216_comb ^ p1_array_index_2044187_comb ^ p1_array_index_2044155_comb ^ literal_2043914[p1_array_index_2044140_comb] ^ literal_2043912[p1_array_index_2044141_comb] ^ literal_2043910[p1_array_index_2044158_comb] ^ p1_array_index_2044143_comb;
  assign p1_array_index_2044276_comb = literal_2043918[p1_res7__40_comb];
  assign p1_array_index_2044277_comb = literal_2043920[p1_res7__38_comb];
  assign p1_res7__50_comb = literal_2043910[p1_res7__48_comb] ^ literal_2043912[p1_res7__46_comb] ^ literal_2043914[p1_res7__44_comb] ^ literal_2043916[p1_res7__42_comb] ^ p1_array_index_2044276_comb ^ p1_array_index_2044277_comb ^ p1_res7__36_comb ^ literal_2043923[p1_res7__34_comb] ^ p1_res7__32_comb ^ p1_array_index_2044229_comb ^ p1_array_index_2044201_comb ^ p1_array_index_2044172_comb ^ literal_2043914[p1_array_index_2044139_comb] ^ literal_2043912[p1_array_index_2044140_comb] ^ literal_2043910[p1_array_index_2044141_comb] ^ p1_array_index_2044158_comb;
  assign p1_array_index_2044288_comb = literal_2043920[p1_res7__40_comb];
  assign p1_res7__52_comb = literal_2043910[p1_res7__50_comb] ^ literal_2043912[p1_res7__48_comb] ^ literal_2043914[p1_res7__46_comb] ^ literal_2043916[p1_res7__44_comb] ^ literal_2043918[p1_res7__42_comb] ^ p1_array_index_2044288_comb ^ p1_res7__38_comb ^ literal_2043923[p1_res7__36_comb] ^ p1_res7__34_comb ^ p1_array_index_2044242_comb ^ p1_array_index_2044215_comb ^ p1_array_index_2044186_comb ^ p1_array_index_2044154_comb ^ literal_2043912[p1_array_index_2044139_comb] ^ literal_2043910[p1_array_index_2044140_comb] ^ p1_array_index_2044141_comb;
  assign p1_array_index_2044298_comb = literal_2043920[p1_res7__42_comb];
  assign p1_res7__54_comb = literal_2043910[p1_res7__52_comb] ^ literal_2043912[p1_res7__50_comb] ^ literal_2043914[p1_res7__48_comb] ^ literal_2043916[p1_res7__46_comb] ^ literal_2043918[p1_res7__44_comb] ^ p1_array_index_2044298_comb ^ p1_res7__40_comb ^ literal_2043923[p1_res7__38_comb] ^ p1_res7__36_comb ^ p1_array_index_2044254_comb ^ p1_array_index_2044228_comb ^ p1_array_index_2044200_comb ^ p1_array_index_2044171_comb ^ literal_2043912[p1_array_index_2044138_comb] ^ literal_2043910[p1_array_index_2044139_comb] ^ p1_array_index_2044140_comb;
  assign p1_res7__56_comb = literal_2043910[p1_res7__54_comb] ^ literal_2043912[p1_res7__52_comb] ^ literal_2043914[p1_res7__50_comb] ^ literal_2043916[p1_res7__48_comb] ^ literal_2043918[p1_res7__46_comb] ^ literal_2043920[p1_res7__44_comb] ^ p1_res7__42_comb ^ literal_2043923[p1_res7__40_comb] ^ p1_res7__38_comb ^ p1_array_index_2044266_comb ^ p1_array_index_2044241_comb ^ p1_array_index_2044214_comb ^ p1_array_index_2044185_comb ^ p1_array_index_2044153_comb ^ literal_2043910[p1_array_index_2044138_comb] ^ p1_array_index_2044139_comb;
  assign p1_res7__58_comb = literal_2043910[p1_res7__56_comb] ^ literal_2043912[p1_res7__54_comb] ^ literal_2043914[p1_res7__52_comb] ^ literal_2043916[p1_res7__50_comb] ^ literal_2043918[p1_res7__48_comb] ^ literal_2043920[p1_res7__46_comb] ^ p1_res7__44_comb ^ literal_2043923[p1_res7__42_comb] ^ p1_res7__40_comb ^ p1_array_index_2044277_comb ^ p1_array_index_2044253_comb ^ p1_array_index_2044227_comb ^ p1_array_index_2044199_comb ^ p1_array_index_2044170_comb ^ literal_2043910[p1_array_index_2044137_comb] ^ p1_array_index_2044138_comb;
  assign p1_res7__60_comb = literal_2043910[p1_res7__58_comb] ^ literal_2043912[p1_res7__56_comb] ^ literal_2043914[p1_res7__54_comb] ^ literal_2043916[p1_res7__52_comb] ^ literal_2043918[p1_res7__50_comb] ^ literal_2043920[p1_res7__48_comb] ^ p1_res7__46_comb ^ literal_2043923[p1_res7__44_comb] ^ p1_res7__42_comb ^ p1_array_index_2044288_comb ^ p1_array_index_2044265_comb ^ p1_array_index_2044240_comb ^ p1_array_index_2044213_comb ^ p1_array_index_2044184_comb ^ p1_array_index_2044152_comb ^ p1_array_index_2044137_comb;
  assign p1_res7__62_comb = literal_2043910[p1_res7__60_comb] ^ literal_2043912[p1_res7__58_comb] ^ literal_2043914[p1_res7__56_comb] ^ literal_2043916[p1_res7__54_comb] ^ literal_2043918[p1_res7__52_comb] ^ literal_2043920[p1_res7__50_comb] ^ p1_res7__48_comb ^ literal_2043923[p1_res7__46_comb] ^ p1_res7__44_comb ^ p1_array_index_2044298_comb ^ p1_array_index_2044276_comb ^ p1_array_index_2044252_comb ^ p1_array_index_2044226_comb ^ p1_array_index_2044198_comb ^ p1_array_index_2044169_comb ^ p1_array_index_2044136_comb;
  assign p1_res__1_comb = {p1_res7__62_comb, p1_res7__60_comb, p1_res7__58_comb, p1_res7__56_comb, p1_res7__54_comb, p1_res7__52_comb, p1_res7__50_comb, p1_res7__48_comb, p1_res7__46_comb, p1_res7__44_comb, p1_res7__42_comb, p1_res7__40_comb, p1_res7__38_comb, p1_res7__36_comb, p1_res7__34_comb, p1_res7__32_comb};
  assign p1_xor_2044338_comb = p1_res__1_comb ^ p1_bit_slice_2043893_comb;
  assign p1_addedKey__34_comb = p1_xor_2044338_comb ^ 128'hb225_9a96_b4d8_8e0b_e769_0430_a44f_7f03;
  assign p1_array_index_2044354_comb = literal_2043896[p1_addedKey__34_comb[127:120]];
  assign p1_array_index_2044355_comb = literal_2043896[p1_addedKey__34_comb[119:112]];
  assign p1_array_index_2044356_comb = literal_2043896[p1_addedKey__34_comb[111:104]];
  assign p1_array_index_2044357_comb = literal_2043896[p1_addedKey__34_comb[103:96]];
  assign p1_array_index_2044358_comb = literal_2043896[p1_addedKey__34_comb[95:88]];
  assign p1_array_index_2044359_comb = literal_2043896[p1_addedKey__34_comb[87:80]];
  assign p1_array_index_2044361_comb = literal_2043896[p1_addedKey__34_comb[71:64]];
  assign p1_array_index_2044363_comb = literal_2043896[p1_addedKey__34_comb[55:48]];
  assign p1_array_index_2044364_comb = literal_2043896[p1_addedKey__34_comb[47:40]];
  assign p1_array_index_2044365_comb = literal_2043896[p1_addedKey__34_comb[39:32]];
  assign p1_array_index_2044366_comb = literal_2043896[p1_addedKey__34_comb[31:24]];
  assign p1_array_index_2044367_comb = literal_2043896[p1_addedKey__34_comb[23:16]];
  assign p1_array_index_2044368_comb = literal_2043896[p1_addedKey__34_comb[15:8]];
  assign p1_array_index_2044370_comb = literal_2043910[p1_array_index_2044354_comb];
  assign p1_array_index_2044371_comb = literal_2043912[p1_array_index_2044355_comb];
  assign p1_array_index_2044372_comb = literal_2043914[p1_array_index_2044356_comb];
  assign p1_array_index_2044373_comb = literal_2043916[p1_array_index_2044357_comb];
  assign p1_array_index_2044374_comb = literal_2043918[p1_array_index_2044358_comb];
  assign p1_array_index_2044375_comb = literal_2043920[p1_array_index_2044359_comb];
  assign p1_array_index_2044376_comb = literal_2043896[p1_addedKey__34_comb[79:72]];
  assign p1_array_index_2044378_comb = literal_2043896[p1_addedKey__34_comb[63:56]];
  assign p1_res7__64_comb = p1_array_index_2044370_comb ^ p1_array_index_2044371_comb ^ p1_array_index_2044372_comb ^ p1_array_index_2044373_comb ^ p1_array_index_2044374_comb ^ p1_array_index_2044375_comb ^ p1_array_index_2044376_comb ^ literal_2043923[p1_array_index_2044361_comb] ^ p1_array_index_2044378_comb ^ literal_2043920[p1_array_index_2044363_comb] ^ literal_2043918[p1_array_index_2044364_comb] ^ literal_2043916[p1_array_index_2044365_comb] ^ literal_2043914[p1_array_index_2044366_comb] ^ literal_2043912[p1_array_index_2044367_comb] ^ literal_2043910[p1_array_index_2044368_comb] ^ literal_2043896[p1_addedKey__34_comb[7:0]];
  assign p1_array_index_2044387_comb = literal_2043910[p1_res7__64_comb];
  assign p1_array_index_2044388_comb = literal_2043912[p1_array_index_2044354_comb];
  assign p1_array_index_2044389_comb = literal_2043914[p1_array_index_2044355_comb];
  assign p1_array_index_2044390_comb = literal_2043916[p1_array_index_2044356_comb];
  assign p1_array_index_2044391_comb = literal_2043918[p1_array_index_2044357_comb];
  assign p1_array_index_2044392_comb = literal_2043920[p1_array_index_2044358_comb];
  assign p1_res7__66_comb = p1_array_index_2044387_comb ^ p1_array_index_2044388_comb ^ p1_array_index_2044389_comb ^ p1_array_index_2044390_comb ^ p1_array_index_2044391_comb ^ p1_array_index_2044392_comb ^ p1_array_index_2044359_comb ^ literal_2043923[p1_array_index_2044376_comb] ^ p1_array_index_2044361_comb ^ literal_2043920[p1_array_index_2044378_comb] ^ literal_2043918[p1_array_index_2044363_comb] ^ literal_2043916[p1_array_index_2044364_comb] ^ literal_2043914[p1_array_index_2044365_comb] ^ literal_2043912[p1_array_index_2044366_comb] ^ literal_2043910[p1_array_index_2044367_comb] ^ p1_array_index_2044368_comb;
  assign p1_array_index_2044402_comb = literal_2043912[p1_res7__64_comb];
  assign p1_array_index_2044403_comb = literal_2043914[p1_array_index_2044354_comb];
  assign p1_array_index_2044404_comb = literal_2043916[p1_array_index_2044355_comb];
  assign p1_array_index_2044405_comb = literal_2043918[p1_array_index_2044356_comb];
  assign p1_array_index_2044406_comb = literal_2043920[p1_array_index_2044357_comb];
  assign p1_res7__68_comb = literal_2043910[p1_res7__66_comb] ^ p1_array_index_2044402_comb ^ p1_array_index_2044403_comb ^ p1_array_index_2044404_comb ^ p1_array_index_2044405_comb ^ p1_array_index_2044406_comb ^ p1_array_index_2044358_comb ^ literal_2043923[p1_array_index_2044359_comb] ^ p1_array_index_2044376_comb ^ literal_2043920[p1_array_index_2044361_comb] ^ literal_2043918[p1_array_index_2044378_comb] ^ literal_2043916[p1_array_index_2044363_comb] ^ literal_2043914[p1_array_index_2044364_comb] ^ literal_2043912[p1_array_index_2044365_comb] ^ literal_2043910[p1_array_index_2044366_comb] ^ p1_array_index_2044367_comb;
  assign p1_array_index_2044416_comb = literal_2043912[p1_res7__66_comb];
  assign p1_array_index_2044417_comb = literal_2043914[p1_res7__64_comb];
  assign p1_array_index_2044418_comb = literal_2043916[p1_array_index_2044354_comb];
  assign p1_array_index_2044419_comb = literal_2043918[p1_array_index_2044355_comb];
  assign p1_array_index_2044420_comb = literal_2043920[p1_array_index_2044356_comb];
  assign p1_res7__70_comb = literal_2043910[p1_res7__68_comb] ^ p1_array_index_2044416_comb ^ p1_array_index_2044417_comb ^ p1_array_index_2044418_comb ^ p1_array_index_2044419_comb ^ p1_array_index_2044420_comb ^ p1_array_index_2044357_comb ^ literal_2043923[p1_array_index_2044358_comb] ^ p1_array_index_2044359_comb ^ literal_2043920[p1_array_index_2044376_comb] ^ literal_2043918[p1_array_index_2044361_comb] ^ literal_2043916[p1_array_index_2044378_comb] ^ literal_2043914[p1_array_index_2044363_comb] ^ literal_2043912[p1_array_index_2044364_comb] ^ literal_2043910[p1_array_index_2044365_comb] ^ p1_array_index_2044366_comb;
  assign p1_array_index_2044431_comb = literal_2043914[p1_res7__66_comb];
  assign p1_array_index_2044432_comb = literal_2043916[p1_res7__64_comb];
  assign p1_array_index_2044433_comb = literal_2043918[p1_array_index_2044354_comb];
  assign p1_array_index_2044434_comb = literal_2043920[p1_array_index_2044355_comb];
  assign p1_res7__72_comb = literal_2043910[p1_res7__70_comb] ^ literal_2043912[p1_res7__68_comb] ^ p1_array_index_2044431_comb ^ p1_array_index_2044432_comb ^ p1_array_index_2044433_comb ^ p1_array_index_2044434_comb ^ p1_array_index_2044356_comb ^ literal_2043923[p1_array_index_2044357_comb] ^ p1_array_index_2044358_comb ^ p1_array_index_2044375_comb ^ literal_2043918[p1_array_index_2044376_comb] ^ literal_2043916[p1_array_index_2044361_comb] ^ literal_2043914[p1_array_index_2044378_comb] ^ literal_2043912[p1_array_index_2044363_comb] ^ literal_2043910[p1_array_index_2044364_comb] ^ p1_array_index_2044365_comb;
  assign p1_array_index_2044444_comb = literal_2043914[p1_res7__68_comb];
  assign p1_array_index_2044445_comb = literal_2043916[p1_res7__66_comb];
  assign p1_array_index_2044446_comb = literal_2043918[p1_res7__64_comb];
  assign p1_array_index_2044447_comb = literal_2043920[p1_array_index_2044354_comb];
  assign p1_res7__74_comb = literal_2043910[p1_res7__72_comb] ^ literal_2043912[p1_res7__70_comb] ^ p1_array_index_2044444_comb ^ p1_array_index_2044445_comb ^ p1_array_index_2044446_comb ^ p1_array_index_2044447_comb ^ p1_array_index_2044355_comb ^ literal_2043923[p1_array_index_2044356_comb] ^ p1_array_index_2044357_comb ^ p1_array_index_2044392_comb ^ literal_2043918[p1_array_index_2044359_comb] ^ literal_2043916[p1_array_index_2044376_comb] ^ literal_2043914[p1_array_index_2044361_comb] ^ literal_2043912[p1_array_index_2044378_comb] ^ literal_2043910[p1_array_index_2044363_comb] ^ p1_array_index_2044364_comb;
  assign p1_array_index_2044458_comb = literal_2043916[p1_res7__68_comb];
  assign p1_array_index_2044459_comb = literal_2043918[p1_res7__66_comb];
  assign p1_array_index_2044460_comb = literal_2043920[p1_res7__64_comb];
  assign p1_res7__76_comb = literal_2043910[p1_res7__74_comb] ^ literal_2043912[p1_res7__72_comb] ^ literal_2043914[p1_res7__70_comb] ^ p1_array_index_2044458_comb ^ p1_array_index_2044459_comb ^ p1_array_index_2044460_comb ^ p1_array_index_2044354_comb ^ literal_2043923[p1_array_index_2044355_comb] ^ p1_array_index_2044356_comb ^ p1_array_index_2044406_comb ^ p1_array_index_2044374_comb ^ literal_2043916[p1_array_index_2044359_comb] ^ literal_2043914[p1_array_index_2044376_comb] ^ literal_2043912[p1_array_index_2044361_comb] ^ literal_2043910[p1_array_index_2044378_comb] ^ p1_array_index_2044363_comb;
  assign p1_array_index_2044470_comb = literal_2043916[p1_res7__70_comb];
  assign p1_array_index_2044471_comb = literal_2043918[p1_res7__68_comb];
  assign p1_array_index_2044472_comb = literal_2043920[p1_res7__66_comb];
  assign p1_res7__78_comb = literal_2043910[p1_res7__76_comb] ^ literal_2043912[p1_res7__74_comb] ^ literal_2043914[p1_res7__72_comb] ^ p1_array_index_2044470_comb ^ p1_array_index_2044471_comb ^ p1_array_index_2044472_comb ^ p1_res7__64_comb ^ literal_2043923[p1_array_index_2044354_comb] ^ p1_array_index_2044355_comb ^ p1_array_index_2044420_comb ^ p1_array_index_2044391_comb ^ literal_2043916[p1_array_index_2044358_comb] ^ literal_2043914[p1_array_index_2044359_comb] ^ literal_2043912[p1_array_index_2044376_comb] ^ literal_2043910[p1_array_index_2044361_comb] ^ p1_array_index_2044378_comb;
  assign p1_array_index_2044483_comb = literal_2043918[p1_res7__70_comb];
  assign p1_array_index_2044484_comb = literal_2043920[p1_res7__68_comb];
  assign p1_res7__80_comb = literal_2043910[p1_res7__78_comb] ^ literal_2043912[p1_res7__76_comb] ^ literal_2043914[p1_res7__74_comb] ^ literal_2043916[p1_res7__72_comb] ^ p1_array_index_2044483_comb ^ p1_array_index_2044484_comb ^ p1_res7__66_comb ^ literal_2043923[p1_res7__64_comb] ^ p1_array_index_2044354_comb ^ p1_array_index_2044434_comb ^ p1_array_index_2044405_comb ^ p1_array_index_2044373_comb ^ literal_2043914[p1_array_index_2044358_comb] ^ literal_2043912[p1_array_index_2044359_comb] ^ literal_2043910[p1_array_index_2044376_comb] ^ p1_array_index_2044361_comb;
  assign p1_array_index_2044494_comb = literal_2043918[p1_res7__72_comb];
  assign p1_array_index_2044495_comb = literal_2043920[p1_res7__70_comb];
  assign p1_res7__82_comb = literal_2043910[p1_res7__80_comb] ^ literal_2043912[p1_res7__78_comb] ^ literal_2043914[p1_res7__76_comb] ^ literal_2043916[p1_res7__74_comb] ^ p1_array_index_2044494_comb ^ p1_array_index_2044495_comb ^ p1_res7__68_comb ^ literal_2043923[p1_res7__66_comb] ^ p1_res7__64_comb ^ p1_array_index_2044447_comb ^ p1_array_index_2044419_comb ^ p1_array_index_2044390_comb ^ literal_2043914[p1_array_index_2044357_comb] ^ literal_2043912[p1_array_index_2044358_comb] ^ literal_2043910[p1_array_index_2044359_comb] ^ p1_array_index_2044376_comb;
  assign p1_array_index_2044506_comb = literal_2043920[p1_res7__72_comb];
  assign p1_res7__84_comb = literal_2043910[p1_res7__82_comb] ^ literal_2043912[p1_res7__80_comb] ^ literal_2043914[p1_res7__78_comb] ^ literal_2043916[p1_res7__76_comb] ^ literal_2043918[p1_res7__74_comb] ^ p1_array_index_2044506_comb ^ p1_res7__70_comb ^ literal_2043923[p1_res7__68_comb] ^ p1_res7__66_comb ^ p1_array_index_2044460_comb ^ p1_array_index_2044433_comb ^ p1_array_index_2044404_comb ^ p1_array_index_2044372_comb ^ literal_2043912[p1_array_index_2044357_comb] ^ literal_2043910[p1_array_index_2044358_comb] ^ p1_array_index_2044359_comb;
  assign p1_array_index_2044516_comb = literal_2043920[p1_res7__74_comb];
  assign p1_res7__86_comb = literal_2043910[p1_res7__84_comb] ^ literal_2043912[p1_res7__82_comb] ^ literal_2043914[p1_res7__80_comb] ^ literal_2043916[p1_res7__78_comb] ^ literal_2043918[p1_res7__76_comb] ^ p1_array_index_2044516_comb ^ p1_res7__72_comb ^ literal_2043923[p1_res7__70_comb] ^ p1_res7__68_comb ^ p1_array_index_2044472_comb ^ p1_array_index_2044446_comb ^ p1_array_index_2044418_comb ^ p1_array_index_2044389_comb ^ literal_2043912[p1_array_index_2044356_comb] ^ literal_2043910[p1_array_index_2044357_comb] ^ p1_array_index_2044358_comb;
  assign p1_res7__88_comb = literal_2043910[p1_res7__86_comb] ^ literal_2043912[p1_res7__84_comb] ^ literal_2043914[p1_res7__82_comb] ^ literal_2043916[p1_res7__80_comb] ^ literal_2043918[p1_res7__78_comb] ^ literal_2043920[p1_res7__76_comb] ^ p1_res7__74_comb ^ literal_2043923[p1_res7__72_comb] ^ p1_res7__70_comb ^ p1_array_index_2044484_comb ^ p1_array_index_2044459_comb ^ p1_array_index_2044432_comb ^ p1_array_index_2044403_comb ^ p1_array_index_2044371_comb ^ literal_2043910[p1_array_index_2044356_comb] ^ p1_array_index_2044357_comb;
  assign p1_res7__90_comb = literal_2043910[p1_res7__88_comb] ^ literal_2043912[p1_res7__86_comb] ^ literal_2043914[p1_res7__84_comb] ^ literal_2043916[p1_res7__82_comb] ^ literal_2043918[p1_res7__80_comb] ^ literal_2043920[p1_res7__78_comb] ^ p1_res7__76_comb ^ literal_2043923[p1_res7__74_comb] ^ p1_res7__72_comb ^ p1_array_index_2044495_comb ^ p1_array_index_2044471_comb ^ p1_array_index_2044445_comb ^ p1_array_index_2044417_comb ^ p1_array_index_2044388_comb ^ literal_2043910[p1_array_index_2044355_comb] ^ p1_array_index_2044356_comb;
  assign p1_res7__92_comb = literal_2043910[p1_res7__90_comb] ^ literal_2043912[p1_res7__88_comb] ^ literal_2043914[p1_res7__86_comb] ^ literal_2043916[p1_res7__84_comb] ^ literal_2043918[p1_res7__82_comb] ^ literal_2043920[p1_res7__80_comb] ^ p1_res7__78_comb ^ literal_2043923[p1_res7__76_comb] ^ p1_res7__74_comb ^ p1_array_index_2044506_comb ^ p1_array_index_2044483_comb ^ p1_array_index_2044458_comb ^ p1_array_index_2044431_comb ^ p1_array_index_2044402_comb ^ p1_array_index_2044370_comb ^ p1_array_index_2044355_comb;
  assign p1_res7__94_comb = literal_2043910[p1_res7__92_comb] ^ literal_2043912[p1_res7__90_comb] ^ literal_2043914[p1_res7__88_comb] ^ literal_2043916[p1_res7__86_comb] ^ literal_2043918[p1_res7__84_comb] ^ literal_2043920[p1_res7__82_comb] ^ p1_res7__80_comb ^ literal_2043923[p1_res7__78_comb] ^ p1_res7__76_comb ^ p1_array_index_2044516_comb ^ p1_array_index_2044494_comb ^ p1_array_index_2044470_comb ^ p1_array_index_2044444_comb ^ p1_array_index_2044416_comb ^ p1_array_index_2044387_comb ^ p1_array_index_2044354_comb;
  assign p1_res__2_comb = {p1_res7__94_comb, p1_res7__92_comb, p1_res7__90_comb, p1_res7__88_comb, p1_res7__86_comb, p1_res7__84_comb, p1_res7__82_comb, p1_res7__80_comb, p1_res7__78_comb, p1_res7__76_comb, p1_res7__74_comb, p1_res7__72_comb, p1_res7__70_comb, p1_res7__68_comb, p1_res7__66_comb, p1_res7__64_comb};
  assign p1_xor_2044556_comb = p1_res__2_comb ^ p1_xor_2044120_comb;
  assign p1_addedKey__35_comb = p1_xor_2044556_comb ^ 128'h7bcd_1b0b_73e3_2ba5_b79c_b140_f255_1504;
  assign p1_array_index_2044572_comb = literal_2043896[p1_addedKey__35_comb[127:120]];
  assign p1_array_index_2044573_comb = literal_2043896[p1_addedKey__35_comb[119:112]];
  assign p1_array_index_2044574_comb = literal_2043896[p1_addedKey__35_comb[111:104]];
  assign p1_array_index_2044575_comb = literal_2043896[p1_addedKey__35_comb[103:96]];
  assign p1_array_index_2044576_comb = literal_2043896[p1_addedKey__35_comb[95:88]];
  assign p1_array_index_2044577_comb = literal_2043896[p1_addedKey__35_comb[87:80]];
  assign p1_array_index_2044579_comb = literal_2043896[p1_addedKey__35_comb[71:64]];
  assign p1_array_index_2044581_comb = literal_2043896[p1_addedKey__35_comb[55:48]];
  assign p1_array_index_2044582_comb = literal_2043896[p1_addedKey__35_comb[47:40]];
  assign p1_array_index_2044583_comb = literal_2043896[p1_addedKey__35_comb[39:32]];
  assign p1_array_index_2044584_comb = literal_2043896[p1_addedKey__35_comb[31:24]];
  assign p1_array_index_2044585_comb = literal_2043896[p1_addedKey__35_comb[23:16]];
  assign p1_array_index_2044586_comb = literal_2043896[p1_addedKey__35_comb[15:8]];
  assign p1_array_index_2044588_comb = literal_2043910[p1_array_index_2044572_comb];
  assign p1_array_index_2044589_comb = literal_2043912[p1_array_index_2044573_comb];
  assign p1_array_index_2044590_comb = literal_2043914[p1_array_index_2044574_comb];
  assign p1_array_index_2044591_comb = literal_2043916[p1_array_index_2044575_comb];
  assign p1_array_index_2044592_comb = literal_2043918[p1_array_index_2044576_comb];
  assign p1_array_index_2044593_comb = literal_2043920[p1_array_index_2044577_comb];
  assign p1_array_index_2044594_comb = literal_2043896[p1_addedKey__35_comb[79:72]];
  assign p1_array_index_2044596_comb = literal_2043896[p1_addedKey__35_comb[63:56]];
  assign p1_res7__96_comb = p1_array_index_2044588_comb ^ p1_array_index_2044589_comb ^ p1_array_index_2044590_comb ^ p1_array_index_2044591_comb ^ p1_array_index_2044592_comb ^ p1_array_index_2044593_comb ^ p1_array_index_2044594_comb ^ literal_2043923[p1_array_index_2044579_comb] ^ p1_array_index_2044596_comb ^ literal_2043920[p1_array_index_2044581_comb] ^ literal_2043918[p1_array_index_2044582_comb] ^ literal_2043916[p1_array_index_2044583_comb] ^ literal_2043914[p1_array_index_2044584_comb] ^ literal_2043912[p1_array_index_2044585_comb] ^ literal_2043910[p1_array_index_2044586_comb] ^ literal_2043896[p1_addedKey__35_comb[7:0]];
  assign p1_array_index_2044605_comb = literal_2043910[p1_res7__96_comb];
  assign p1_array_index_2044606_comb = literal_2043912[p1_array_index_2044572_comb];
  assign p1_array_index_2044607_comb = literal_2043914[p1_array_index_2044573_comb];
  assign p1_array_index_2044608_comb = literal_2043916[p1_array_index_2044574_comb];
  assign p1_array_index_2044609_comb = literal_2043918[p1_array_index_2044575_comb];
  assign p1_array_index_2044610_comb = literal_2043920[p1_array_index_2044576_comb];
  assign p1_res7__98_comb = p1_array_index_2044605_comb ^ p1_array_index_2044606_comb ^ p1_array_index_2044607_comb ^ p1_array_index_2044608_comb ^ p1_array_index_2044609_comb ^ p1_array_index_2044610_comb ^ p1_array_index_2044577_comb ^ literal_2043923[p1_array_index_2044594_comb] ^ p1_array_index_2044579_comb ^ literal_2043920[p1_array_index_2044596_comb] ^ literal_2043918[p1_array_index_2044581_comb] ^ literal_2043916[p1_array_index_2044582_comb] ^ literal_2043914[p1_array_index_2044583_comb] ^ literal_2043912[p1_array_index_2044584_comb] ^ literal_2043910[p1_array_index_2044585_comb] ^ p1_array_index_2044586_comb;
  assign p1_array_index_2044620_comb = literal_2043912[p1_res7__96_comb];
  assign p1_array_index_2044621_comb = literal_2043914[p1_array_index_2044572_comb];
  assign p1_array_index_2044622_comb = literal_2043916[p1_array_index_2044573_comb];
  assign p1_array_index_2044623_comb = literal_2043918[p1_array_index_2044574_comb];
  assign p1_array_index_2044624_comb = literal_2043920[p1_array_index_2044575_comb];
  assign p1_res7__100_comb = literal_2043910[p1_res7__98_comb] ^ p1_array_index_2044620_comb ^ p1_array_index_2044621_comb ^ p1_array_index_2044622_comb ^ p1_array_index_2044623_comb ^ p1_array_index_2044624_comb ^ p1_array_index_2044576_comb ^ literal_2043923[p1_array_index_2044577_comb] ^ p1_array_index_2044594_comb ^ literal_2043920[p1_array_index_2044579_comb] ^ literal_2043918[p1_array_index_2044596_comb] ^ literal_2043916[p1_array_index_2044581_comb] ^ literal_2043914[p1_array_index_2044582_comb] ^ literal_2043912[p1_array_index_2044583_comb] ^ literal_2043910[p1_array_index_2044584_comb] ^ p1_array_index_2044585_comb;
  assign p1_array_index_2044634_comb = literal_2043912[p1_res7__98_comb];
  assign p1_array_index_2044635_comb = literal_2043914[p1_res7__96_comb];
  assign p1_array_index_2044636_comb = literal_2043916[p1_array_index_2044572_comb];
  assign p1_array_index_2044637_comb = literal_2043918[p1_array_index_2044573_comb];
  assign p1_array_index_2044638_comb = literal_2043920[p1_array_index_2044574_comb];
  assign p1_res7__102_comb = literal_2043910[p1_res7__100_comb] ^ p1_array_index_2044634_comb ^ p1_array_index_2044635_comb ^ p1_array_index_2044636_comb ^ p1_array_index_2044637_comb ^ p1_array_index_2044638_comb ^ p1_array_index_2044575_comb ^ literal_2043923[p1_array_index_2044576_comb] ^ p1_array_index_2044577_comb ^ literal_2043920[p1_array_index_2044594_comb] ^ literal_2043918[p1_array_index_2044579_comb] ^ literal_2043916[p1_array_index_2044596_comb] ^ literal_2043914[p1_array_index_2044581_comb] ^ literal_2043912[p1_array_index_2044582_comb] ^ literal_2043910[p1_array_index_2044583_comb] ^ p1_array_index_2044584_comb;
  assign p1_array_index_2044649_comb = literal_2043914[p1_res7__98_comb];
  assign p1_array_index_2044650_comb = literal_2043916[p1_res7__96_comb];
  assign p1_array_index_2044651_comb = literal_2043918[p1_array_index_2044572_comb];
  assign p1_array_index_2044652_comb = literal_2043920[p1_array_index_2044573_comb];
  assign p1_res7__104_comb = literal_2043910[p1_res7__102_comb] ^ literal_2043912[p1_res7__100_comb] ^ p1_array_index_2044649_comb ^ p1_array_index_2044650_comb ^ p1_array_index_2044651_comb ^ p1_array_index_2044652_comb ^ p1_array_index_2044574_comb ^ literal_2043923[p1_array_index_2044575_comb] ^ p1_array_index_2044576_comb ^ p1_array_index_2044593_comb ^ literal_2043918[p1_array_index_2044594_comb] ^ literal_2043916[p1_array_index_2044579_comb] ^ literal_2043914[p1_array_index_2044596_comb] ^ literal_2043912[p1_array_index_2044581_comb] ^ literal_2043910[p1_array_index_2044582_comb] ^ p1_array_index_2044583_comb;
  assign p1_array_index_2044662_comb = literal_2043914[p1_res7__100_comb];
  assign p1_array_index_2044663_comb = literal_2043916[p1_res7__98_comb];
  assign p1_array_index_2044664_comb = literal_2043918[p1_res7__96_comb];
  assign p1_array_index_2044665_comb = literal_2043920[p1_array_index_2044572_comb];
  assign p1_res7__106_comb = literal_2043910[p1_res7__104_comb] ^ literal_2043912[p1_res7__102_comb] ^ p1_array_index_2044662_comb ^ p1_array_index_2044663_comb ^ p1_array_index_2044664_comb ^ p1_array_index_2044665_comb ^ p1_array_index_2044573_comb ^ literal_2043923[p1_array_index_2044574_comb] ^ p1_array_index_2044575_comb ^ p1_array_index_2044610_comb ^ literal_2043918[p1_array_index_2044577_comb] ^ literal_2043916[p1_array_index_2044594_comb] ^ literal_2043914[p1_array_index_2044579_comb] ^ literal_2043912[p1_array_index_2044596_comb] ^ literal_2043910[p1_array_index_2044581_comb] ^ p1_array_index_2044582_comb;
  assign p1_array_index_2044676_comb = literal_2043916[p1_res7__100_comb];
  assign p1_array_index_2044677_comb = literal_2043918[p1_res7__98_comb];
  assign p1_array_index_2044678_comb = literal_2043920[p1_res7__96_comb];
  assign p1_res7__108_comb = literal_2043910[p1_res7__106_comb] ^ literal_2043912[p1_res7__104_comb] ^ literal_2043914[p1_res7__102_comb] ^ p1_array_index_2044676_comb ^ p1_array_index_2044677_comb ^ p1_array_index_2044678_comb ^ p1_array_index_2044572_comb ^ literal_2043923[p1_array_index_2044573_comb] ^ p1_array_index_2044574_comb ^ p1_array_index_2044624_comb ^ p1_array_index_2044592_comb ^ literal_2043916[p1_array_index_2044577_comb] ^ literal_2043914[p1_array_index_2044594_comb] ^ literal_2043912[p1_array_index_2044579_comb] ^ literal_2043910[p1_array_index_2044596_comb] ^ p1_array_index_2044581_comb;
  assign p1_array_index_2044688_comb = literal_2043916[p1_res7__102_comb];
  assign p1_array_index_2044689_comb = literal_2043918[p1_res7__100_comb];
  assign p1_array_index_2044690_comb = literal_2043920[p1_res7__98_comb];
  assign p1_res7__110_comb = literal_2043910[p1_res7__108_comb] ^ literal_2043912[p1_res7__106_comb] ^ literal_2043914[p1_res7__104_comb] ^ p1_array_index_2044688_comb ^ p1_array_index_2044689_comb ^ p1_array_index_2044690_comb ^ p1_res7__96_comb ^ literal_2043923[p1_array_index_2044572_comb] ^ p1_array_index_2044573_comb ^ p1_array_index_2044638_comb ^ p1_array_index_2044609_comb ^ literal_2043916[p1_array_index_2044576_comb] ^ literal_2043914[p1_array_index_2044577_comb] ^ literal_2043912[p1_array_index_2044594_comb] ^ literal_2043910[p1_array_index_2044579_comb] ^ p1_array_index_2044596_comb;
  assign p1_array_index_2044701_comb = literal_2043918[p1_res7__102_comb];
  assign p1_array_index_2044702_comb = literal_2043920[p1_res7__100_comb];
  assign p1_res7__112_comb = literal_2043910[p1_res7__110_comb] ^ literal_2043912[p1_res7__108_comb] ^ literal_2043914[p1_res7__106_comb] ^ literal_2043916[p1_res7__104_comb] ^ p1_array_index_2044701_comb ^ p1_array_index_2044702_comb ^ p1_res7__98_comb ^ literal_2043923[p1_res7__96_comb] ^ p1_array_index_2044572_comb ^ p1_array_index_2044652_comb ^ p1_array_index_2044623_comb ^ p1_array_index_2044591_comb ^ literal_2043914[p1_array_index_2044576_comb] ^ literal_2043912[p1_array_index_2044577_comb] ^ literal_2043910[p1_array_index_2044594_comb] ^ p1_array_index_2044579_comb;
  assign p1_array_index_2044712_comb = literal_2043918[p1_res7__104_comb];
  assign p1_array_index_2044713_comb = literal_2043920[p1_res7__102_comb];
  assign p1_res7__114_comb = literal_2043910[p1_res7__112_comb] ^ literal_2043912[p1_res7__110_comb] ^ literal_2043914[p1_res7__108_comb] ^ literal_2043916[p1_res7__106_comb] ^ p1_array_index_2044712_comb ^ p1_array_index_2044713_comb ^ p1_res7__100_comb ^ literal_2043923[p1_res7__98_comb] ^ p1_res7__96_comb ^ p1_array_index_2044665_comb ^ p1_array_index_2044637_comb ^ p1_array_index_2044608_comb ^ literal_2043914[p1_array_index_2044575_comb] ^ literal_2043912[p1_array_index_2044576_comb] ^ literal_2043910[p1_array_index_2044577_comb] ^ p1_array_index_2044594_comb;
  assign p1_array_index_2044724_comb = literal_2043920[p1_res7__104_comb];
  assign p1_res7__116_comb = literal_2043910[p1_res7__114_comb] ^ literal_2043912[p1_res7__112_comb] ^ literal_2043914[p1_res7__110_comb] ^ literal_2043916[p1_res7__108_comb] ^ literal_2043918[p1_res7__106_comb] ^ p1_array_index_2044724_comb ^ p1_res7__102_comb ^ literal_2043923[p1_res7__100_comb] ^ p1_res7__98_comb ^ p1_array_index_2044678_comb ^ p1_array_index_2044651_comb ^ p1_array_index_2044622_comb ^ p1_array_index_2044590_comb ^ literal_2043912[p1_array_index_2044575_comb] ^ literal_2043910[p1_array_index_2044576_comb] ^ p1_array_index_2044577_comb;
  assign p1_array_index_2044734_comb = literal_2043920[p1_res7__106_comb];
  assign p1_res7__118_comb = literal_2043910[p1_res7__116_comb] ^ literal_2043912[p1_res7__114_comb] ^ literal_2043914[p1_res7__112_comb] ^ literal_2043916[p1_res7__110_comb] ^ literal_2043918[p1_res7__108_comb] ^ p1_array_index_2044734_comb ^ p1_res7__104_comb ^ literal_2043923[p1_res7__102_comb] ^ p1_res7__100_comb ^ p1_array_index_2044690_comb ^ p1_array_index_2044664_comb ^ p1_array_index_2044636_comb ^ p1_array_index_2044607_comb ^ literal_2043912[p1_array_index_2044574_comb] ^ literal_2043910[p1_array_index_2044575_comb] ^ p1_array_index_2044576_comb;
  assign p1_res7__120_comb = literal_2043910[p1_res7__118_comb] ^ literal_2043912[p1_res7__116_comb] ^ literal_2043914[p1_res7__114_comb] ^ literal_2043916[p1_res7__112_comb] ^ literal_2043918[p1_res7__110_comb] ^ literal_2043920[p1_res7__108_comb] ^ p1_res7__106_comb ^ literal_2043923[p1_res7__104_comb] ^ p1_res7__102_comb ^ p1_array_index_2044702_comb ^ p1_array_index_2044677_comb ^ p1_array_index_2044650_comb ^ p1_array_index_2044621_comb ^ p1_array_index_2044589_comb ^ literal_2043910[p1_array_index_2044574_comb] ^ p1_array_index_2044575_comb;
  assign p1_res7__122_comb = literal_2043910[p1_res7__120_comb] ^ literal_2043912[p1_res7__118_comb] ^ literal_2043914[p1_res7__116_comb] ^ literal_2043916[p1_res7__114_comb] ^ literal_2043918[p1_res7__112_comb] ^ literal_2043920[p1_res7__110_comb] ^ p1_res7__108_comb ^ literal_2043923[p1_res7__106_comb] ^ p1_res7__104_comb ^ p1_array_index_2044713_comb ^ p1_array_index_2044689_comb ^ p1_array_index_2044663_comb ^ p1_array_index_2044635_comb ^ p1_array_index_2044606_comb ^ literal_2043910[p1_array_index_2044573_comb] ^ p1_array_index_2044574_comb;
  assign p1_res7__124_comb = literal_2043910[p1_res7__122_comb] ^ literal_2043912[p1_res7__120_comb] ^ literal_2043914[p1_res7__118_comb] ^ literal_2043916[p1_res7__116_comb] ^ literal_2043918[p1_res7__114_comb] ^ literal_2043920[p1_res7__112_comb] ^ p1_res7__110_comb ^ literal_2043923[p1_res7__108_comb] ^ p1_res7__106_comb ^ p1_array_index_2044724_comb ^ p1_array_index_2044701_comb ^ p1_array_index_2044676_comb ^ p1_array_index_2044649_comb ^ p1_array_index_2044620_comb ^ p1_array_index_2044588_comb ^ p1_array_index_2044573_comb;
  assign p1_res7__126_comb = literal_2043910[p1_res7__124_comb] ^ literal_2043912[p1_res7__122_comb] ^ literal_2043914[p1_res7__120_comb] ^ literal_2043916[p1_res7__118_comb] ^ literal_2043918[p1_res7__116_comb] ^ literal_2043920[p1_res7__114_comb] ^ p1_res7__112_comb ^ literal_2043923[p1_res7__110_comb] ^ p1_res7__108_comb ^ p1_array_index_2044734_comb ^ p1_array_index_2044712_comb ^ p1_array_index_2044688_comb ^ p1_array_index_2044662_comb ^ p1_array_index_2044634_comb ^ p1_array_index_2044605_comb ^ p1_array_index_2044572_comb;
  assign p1_res__3_comb = {p1_res7__126_comb, p1_res7__124_comb, p1_res7__122_comb, p1_res7__120_comb, p1_res7__118_comb, p1_res7__116_comb, p1_res7__114_comb, p1_res7__112_comb, p1_res7__110_comb, p1_res7__108_comb, p1_res7__106_comb, p1_res7__104_comb, p1_res7__102_comb, p1_res7__100_comb, p1_res7__98_comb, p1_res7__96_comb};
  assign p1_xor_2044774_comb = p1_res__3_comb ^ p1_xor_2044338_comb;
  assign p1_addedKey__36_comb = p1_xor_2044774_comb ^ 128'h156f_6d79_1fab_511d_eabb_0c50_2fd1_8105;
  assign p1_array_index_2044790_comb = literal_2043896[p1_addedKey__36_comb[127:120]];
  assign p1_array_index_2044791_comb = literal_2043896[p1_addedKey__36_comb[119:112]];
  assign p1_array_index_2044792_comb = literal_2043896[p1_addedKey__36_comb[111:104]];
  assign p1_array_index_2044793_comb = literal_2043896[p1_addedKey__36_comb[103:96]];
  assign p1_array_index_2044794_comb = literal_2043896[p1_addedKey__36_comb[95:88]];
  assign p1_array_index_2044795_comb = literal_2043896[p1_addedKey__36_comb[87:80]];
  assign p1_array_index_2044797_comb = literal_2043896[p1_addedKey__36_comb[71:64]];
  assign p1_array_index_2044799_comb = literal_2043896[p1_addedKey__36_comb[55:48]];
  assign p1_array_index_2044800_comb = literal_2043896[p1_addedKey__36_comb[47:40]];
  assign p1_array_index_2044801_comb = literal_2043896[p1_addedKey__36_comb[39:32]];
  assign p1_array_index_2044802_comb = literal_2043896[p1_addedKey__36_comb[31:24]];
  assign p1_array_index_2044803_comb = literal_2043896[p1_addedKey__36_comb[23:16]];
  assign p1_array_index_2044804_comb = literal_2043896[p1_addedKey__36_comb[15:8]];
  assign p1_array_index_2044806_comb = literal_2043910[p1_array_index_2044790_comb];
  assign p1_array_index_2044807_comb = literal_2043912[p1_array_index_2044791_comb];
  assign p1_array_index_2044808_comb = literal_2043914[p1_array_index_2044792_comb];
  assign p1_array_index_2044809_comb = literal_2043916[p1_array_index_2044793_comb];
  assign p1_array_index_2044810_comb = literal_2043918[p1_array_index_2044794_comb];
  assign p1_array_index_2044811_comb = literal_2043920[p1_array_index_2044795_comb];
  assign p1_array_index_2044812_comb = literal_2043896[p1_addedKey__36_comb[79:72]];
  assign p1_array_index_2044814_comb = literal_2043896[p1_addedKey__36_comb[63:56]];
  assign p1_res7__128_comb = p1_array_index_2044806_comb ^ p1_array_index_2044807_comb ^ p1_array_index_2044808_comb ^ p1_array_index_2044809_comb ^ p1_array_index_2044810_comb ^ p1_array_index_2044811_comb ^ p1_array_index_2044812_comb ^ literal_2043923[p1_array_index_2044797_comb] ^ p1_array_index_2044814_comb ^ literal_2043920[p1_array_index_2044799_comb] ^ literal_2043918[p1_array_index_2044800_comb] ^ literal_2043916[p1_array_index_2044801_comb] ^ literal_2043914[p1_array_index_2044802_comb] ^ literal_2043912[p1_array_index_2044803_comb] ^ literal_2043910[p1_array_index_2044804_comb] ^ literal_2043896[p1_addedKey__36_comb[7:0]];
  assign p1_array_index_2044823_comb = literal_2043910[p1_res7__128_comb];
  assign p1_array_index_2044824_comb = literal_2043912[p1_array_index_2044790_comb];
  assign p1_array_index_2044825_comb = literal_2043914[p1_array_index_2044791_comb];
  assign p1_array_index_2044826_comb = literal_2043916[p1_array_index_2044792_comb];
  assign p1_array_index_2044827_comb = literal_2043918[p1_array_index_2044793_comb];
  assign p1_array_index_2044828_comb = literal_2043920[p1_array_index_2044794_comb];
  assign p1_res7__130_comb = p1_array_index_2044823_comb ^ p1_array_index_2044824_comb ^ p1_array_index_2044825_comb ^ p1_array_index_2044826_comb ^ p1_array_index_2044827_comb ^ p1_array_index_2044828_comb ^ p1_array_index_2044795_comb ^ literal_2043923[p1_array_index_2044812_comb] ^ p1_array_index_2044797_comb ^ literal_2043920[p1_array_index_2044814_comb] ^ literal_2043918[p1_array_index_2044799_comb] ^ literal_2043916[p1_array_index_2044800_comb] ^ literal_2043914[p1_array_index_2044801_comb] ^ literal_2043912[p1_array_index_2044802_comb] ^ literal_2043910[p1_array_index_2044803_comb] ^ p1_array_index_2044804_comb;
  assign p1_array_index_2044838_comb = literal_2043912[p1_res7__128_comb];
  assign p1_array_index_2044839_comb = literal_2043914[p1_array_index_2044790_comb];
  assign p1_array_index_2044840_comb = literal_2043916[p1_array_index_2044791_comb];
  assign p1_array_index_2044841_comb = literal_2043918[p1_array_index_2044792_comb];
  assign p1_array_index_2044842_comb = literal_2043920[p1_array_index_2044793_comb];
  assign p1_res7__132_comb = literal_2043910[p1_res7__130_comb] ^ p1_array_index_2044838_comb ^ p1_array_index_2044839_comb ^ p1_array_index_2044840_comb ^ p1_array_index_2044841_comb ^ p1_array_index_2044842_comb ^ p1_array_index_2044794_comb ^ literal_2043923[p1_array_index_2044795_comb] ^ p1_array_index_2044812_comb ^ literal_2043920[p1_array_index_2044797_comb] ^ literal_2043918[p1_array_index_2044814_comb] ^ literal_2043916[p1_array_index_2044799_comb] ^ literal_2043914[p1_array_index_2044800_comb] ^ literal_2043912[p1_array_index_2044801_comb] ^ literal_2043910[p1_array_index_2044802_comb] ^ p1_array_index_2044803_comb;
  assign p1_array_index_2044852_comb = literal_2043912[p1_res7__130_comb];
  assign p1_array_index_2044853_comb = literal_2043914[p1_res7__128_comb];
  assign p1_array_index_2044854_comb = literal_2043916[p1_array_index_2044790_comb];
  assign p1_array_index_2044855_comb = literal_2043918[p1_array_index_2044791_comb];
  assign p1_array_index_2044856_comb = literal_2043920[p1_array_index_2044792_comb];
  assign p1_res7__134_comb = literal_2043910[p1_res7__132_comb] ^ p1_array_index_2044852_comb ^ p1_array_index_2044853_comb ^ p1_array_index_2044854_comb ^ p1_array_index_2044855_comb ^ p1_array_index_2044856_comb ^ p1_array_index_2044793_comb ^ literal_2043923[p1_array_index_2044794_comb] ^ p1_array_index_2044795_comb ^ literal_2043920[p1_array_index_2044812_comb] ^ literal_2043918[p1_array_index_2044797_comb] ^ literal_2043916[p1_array_index_2044814_comb] ^ literal_2043914[p1_array_index_2044799_comb] ^ literal_2043912[p1_array_index_2044800_comb] ^ literal_2043910[p1_array_index_2044801_comb] ^ p1_array_index_2044802_comb;
  assign p1_array_index_2044867_comb = literal_2043914[p1_res7__130_comb];
  assign p1_array_index_2044868_comb = literal_2043916[p1_res7__128_comb];
  assign p1_array_index_2044869_comb = literal_2043918[p1_array_index_2044790_comb];
  assign p1_array_index_2044870_comb = literal_2043920[p1_array_index_2044791_comb];
  assign p1_res7__136_comb = literal_2043910[p1_res7__134_comb] ^ literal_2043912[p1_res7__132_comb] ^ p1_array_index_2044867_comb ^ p1_array_index_2044868_comb ^ p1_array_index_2044869_comb ^ p1_array_index_2044870_comb ^ p1_array_index_2044792_comb ^ literal_2043923[p1_array_index_2044793_comb] ^ p1_array_index_2044794_comb ^ p1_array_index_2044811_comb ^ literal_2043918[p1_array_index_2044812_comb] ^ literal_2043916[p1_array_index_2044797_comb] ^ literal_2043914[p1_array_index_2044814_comb] ^ literal_2043912[p1_array_index_2044799_comb] ^ literal_2043910[p1_array_index_2044800_comb] ^ p1_array_index_2044801_comb;
  assign p1_array_index_2044880_comb = literal_2043914[p1_res7__132_comb];
  assign p1_array_index_2044881_comb = literal_2043916[p1_res7__130_comb];
  assign p1_array_index_2044882_comb = literal_2043918[p1_res7__128_comb];
  assign p1_array_index_2044883_comb = literal_2043920[p1_array_index_2044790_comb];
  assign p1_res7__138_comb = literal_2043910[p1_res7__136_comb] ^ literal_2043912[p1_res7__134_comb] ^ p1_array_index_2044880_comb ^ p1_array_index_2044881_comb ^ p1_array_index_2044882_comb ^ p1_array_index_2044883_comb ^ p1_array_index_2044791_comb ^ literal_2043923[p1_array_index_2044792_comb] ^ p1_array_index_2044793_comb ^ p1_array_index_2044828_comb ^ literal_2043918[p1_array_index_2044795_comb] ^ literal_2043916[p1_array_index_2044812_comb] ^ literal_2043914[p1_array_index_2044797_comb] ^ literal_2043912[p1_array_index_2044814_comb] ^ literal_2043910[p1_array_index_2044799_comb] ^ p1_array_index_2044800_comb;
  assign p1_array_index_2044894_comb = literal_2043916[p1_res7__132_comb];
  assign p1_array_index_2044895_comb = literal_2043918[p1_res7__130_comb];
  assign p1_array_index_2044896_comb = literal_2043920[p1_res7__128_comb];
  assign p1_res7__140_comb = literal_2043910[p1_res7__138_comb] ^ literal_2043912[p1_res7__136_comb] ^ literal_2043914[p1_res7__134_comb] ^ p1_array_index_2044894_comb ^ p1_array_index_2044895_comb ^ p1_array_index_2044896_comb ^ p1_array_index_2044790_comb ^ literal_2043923[p1_array_index_2044791_comb] ^ p1_array_index_2044792_comb ^ p1_array_index_2044842_comb ^ p1_array_index_2044810_comb ^ literal_2043916[p1_array_index_2044795_comb] ^ literal_2043914[p1_array_index_2044812_comb] ^ literal_2043912[p1_array_index_2044797_comb] ^ literal_2043910[p1_array_index_2044814_comb] ^ p1_array_index_2044799_comb;

  // Registers for pipe stage 1:
  reg [127:0] p1_encoded;
  reg [127:0] p1_bit_slice_2043893;
  reg [127:0] p1_bit_slice_2044119;
  reg [127:0] p1_xor_2044556;
  reg [127:0] p1_xor_2044774;
  reg [7:0] p1_array_index_2044790;
  reg [7:0] p1_array_index_2044791;
  reg [7:0] p1_array_index_2044792;
  reg [7:0] p1_array_index_2044793;
  reg [7:0] p1_array_index_2044794;
  reg [7:0] p1_array_index_2044795;
  reg [7:0] p1_array_index_2044797;
  reg [7:0] p1_array_index_2044806;
  reg [7:0] p1_array_index_2044807;
  reg [7:0] p1_array_index_2044808;
  reg [7:0] p1_array_index_2044809;
  reg [7:0] p1_array_index_2044812;
  reg [7:0] p1_array_index_2044814;
  reg [7:0] p1_res7__128;
  reg [7:0] p1_array_index_2044823;
  reg [7:0] p1_array_index_2044824;
  reg [7:0] p1_array_index_2044825;
  reg [7:0] p1_array_index_2044826;
  reg [7:0] p1_array_index_2044827;
  reg [7:0] p1_res7__130;
  reg [7:0] p1_array_index_2044838;
  reg [7:0] p1_array_index_2044839;
  reg [7:0] p1_array_index_2044840;
  reg [7:0] p1_array_index_2044841;
  reg [7:0] p1_res7__132;
  reg [7:0] p1_array_index_2044852;
  reg [7:0] p1_array_index_2044853;
  reg [7:0] p1_array_index_2044854;
  reg [7:0] p1_array_index_2044855;
  reg [7:0] p1_array_index_2044856;
  reg [7:0] p1_res7__134;
  reg [7:0] p1_array_index_2044867;
  reg [7:0] p1_array_index_2044868;
  reg [7:0] p1_array_index_2044869;
  reg [7:0] p1_array_index_2044870;
  reg [7:0] p1_res7__136;
  reg [7:0] p1_array_index_2044880;
  reg [7:0] p1_array_index_2044881;
  reg [7:0] p1_array_index_2044882;
  reg [7:0] p1_array_index_2044883;
  reg [7:0] p1_res7__138;
  reg [7:0] p1_array_index_2044894;
  reg [7:0] p1_array_index_2044895;
  reg [7:0] p1_array_index_2044896;
  reg [7:0] p1_res7__140;
  reg [7:0] p2_literal_2043896[256];
  reg [7:0] p2_literal_2043910[256];
  reg [7:0] p2_literal_2043912[256];
  reg [7:0] p2_literal_2043914[256];
  reg [7:0] p2_literal_2043916[256];
  reg [7:0] p2_literal_2043918[256];
  reg [7:0] p2_literal_2043920[256];
  reg [7:0] p2_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p1_encoded <= p0_encoded;
    p1_bit_slice_2043893 <= p1_bit_slice_2043893_comb;
    p1_bit_slice_2044119 <= p1_bit_slice_2044119_comb;
    p1_xor_2044556 <= p1_xor_2044556_comb;
    p1_xor_2044774 <= p1_xor_2044774_comb;
    p1_array_index_2044790 <= p1_array_index_2044790_comb;
    p1_array_index_2044791 <= p1_array_index_2044791_comb;
    p1_array_index_2044792 <= p1_array_index_2044792_comb;
    p1_array_index_2044793 <= p1_array_index_2044793_comb;
    p1_array_index_2044794 <= p1_array_index_2044794_comb;
    p1_array_index_2044795 <= p1_array_index_2044795_comb;
    p1_array_index_2044797 <= p1_array_index_2044797_comb;
    p1_array_index_2044806 <= p1_array_index_2044806_comb;
    p1_array_index_2044807 <= p1_array_index_2044807_comb;
    p1_array_index_2044808 <= p1_array_index_2044808_comb;
    p1_array_index_2044809 <= p1_array_index_2044809_comb;
    p1_array_index_2044812 <= p1_array_index_2044812_comb;
    p1_array_index_2044814 <= p1_array_index_2044814_comb;
    p1_res7__128 <= p1_res7__128_comb;
    p1_array_index_2044823 <= p1_array_index_2044823_comb;
    p1_array_index_2044824 <= p1_array_index_2044824_comb;
    p1_array_index_2044825 <= p1_array_index_2044825_comb;
    p1_array_index_2044826 <= p1_array_index_2044826_comb;
    p1_array_index_2044827 <= p1_array_index_2044827_comb;
    p1_res7__130 <= p1_res7__130_comb;
    p1_array_index_2044838 <= p1_array_index_2044838_comb;
    p1_array_index_2044839 <= p1_array_index_2044839_comb;
    p1_array_index_2044840 <= p1_array_index_2044840_comb;
    p1_array_index_2044841 <= p1_array_index_2044841_comb;
    p1_res7__132 <= p1_res7__132_comb;
    p1_array_index_2044852 <= p1_array_index_2044852_comb;
    p1_array_index_2044853 <= p1_array_index_2044853_comb;
    p1_array_index_2044854 <= p1_array_index_2044854_comb;
    p1_array_index_2044855 <= p1_array_index_2044855_comb;
    p1_array_index_2044856 <= p1_array_index_2044856_comb;
    p1_res7__134 <= p1_res7__134_comb;
    p1_array_index_2044867 <= p1_array_index_2044867_comb;
    p1_array_index_2044868 <= p1_array_index_2044868_comb;
    p1_array_index_2044869 <= p1_array_index_2044869_comb;
    p1_array_index_2044870 <= p1_array_index_2044870_comb;
    p1_res7__136 <= p1_res7__136_comb;
    p1_array_index_2044880 <= p1_array_index_2044880_comb;
    p1_array_index_2044881 <= p1_array_index_2044881_comb;
    p1_array_index_2044882 <= p1_array_index_2044882_comb;
    p1_array_index_2044883 <= p1_array_index_2044883_comb;
    p1_res7__138 <= p1_res7__138_comb;
    p1_array_index_2044894 <= p1_array_index_2044894_comb;
    p1_array_index_2044895 <= p1_array_index_2044895_comb;
    p1_array_index_2044896 <= p1_array_index_2044896_comb;
    p1_res7__140 <= p1_res7__140_comb;
    p2_literal_2043896 <= p1_literal_2043896;
    p2_literal_2043910 <= p1_literal_2043910;
    p2_literal_2043912 <= p1_literal_2043912;
    p2_literal_2043914 <= p1_literal_2043914;
    p2_literal_2043916 <= p1_literal_2043916;
    p2_literal_2043918 <= p1_literal_2043918;
    p2_literal_2043920 <= p1_literal_2043920;
    p2_literal_2043923 <= p1_literal_2043923;
  end

  // ===== Pipe stage 2:
  wire [7:0] p2_array_index_2045022_comb;
  wire [7:0] p2_array_index_2045023_comb;
  wire [7:0] p2_array_index_2045024_comb;
  wire [7:0] p2_res7__142_comb;
  wire [7:0] p2_array_index_2045035_comb;
  wire [7:0] p2_array_index_2045036_comb;
  wire [7:0] p2_res7__144_comb;
  wire [7:0] p2_array_index_2045046_comb;
  wire [7:0] p2_array_index_2045047_comb;
  wire [7:0] p2_res7__146_comb;
  wire [7:0] p2_array_index_2045058_comb;
  wire [7:0] p2_res7__148_comb;
  wire [7:0] p2_array_index_2045068_comb;
  wire [7:0] p2_res7__150_comb;
  wire [7:0] p2_res7__152_comb;
  wire [7:0] p2_res7__154_comb;
  wire [7:0] p2_res7__156_comb;
  wire [7:0] p2_res7__158_comb;
  wire [127:0] p2_res__4_comb;
  wire [127:0] p2_xor_2045108_comb;
  wire [127:0] p2_addedKey__37_comb;
  wire [7:0] p2_array_index_2045124_comb;
  wire [7:0] p2_array_index_2045125_comb;
  wire [7:0] p2_array_index_2045126_comb;
  wire [7:0] p2_array_index_2045127_comb;
  wire [7:0] p2_array_index_2045128_comb;
  wire [7:0] p2_array_index_2045129_comb;
  wire [7:0] p2_array_index_2045131_comb;
  wire [7:0] p2_array_index_2045133_comb;
  wire [7:0] p2_array_index_2045134_comb;
  wire [7:0] p2_array_index_2045135_comb;
  wire [7:0] p2_array_index_2045136_comb;
  wire [7:0] p2_array_index_2045137_comb;
  wire [7:0] p2_array_index_2045138_comb;
  wire [7:0] p2_array_index_2045140_comb;
  wire [7:0] p2_array_index_2045141_comb;
  wire [7:0] p2_array_index_2045142_comb;
  wire [7:0] p2_array_index_2045143_comb;
  wire [7:0] p2_array_index_2045144_comb;
  wire [7:0] p2_array_index_2045145_comb;
  wire [7:0] p2_array_index_2045146_comb;
  wire [7:0] p2_array_index_2045148_comb;
  wire [7:0] p2_res7__160_comb;
  wire [7:0] p2_array_index_2045157_comb;
  wire [7:0] p2_array_index_2045158_comb;
  wire [7:0] p2_array_index_2045159_comb;
  wire [7:0] p2_array_index_2045160_comb;
  wire [7:0] p2_array_index_2045161_comb;
  wire [7:0] p2_array_index_2045162_comb;
  wire [7:0] p2_res7__162_comb;
  wire [7:0] p2_array_index_2045172_comb;
  wire [7:0] p2_array_index_2045173_comb;
  wire [7:0] p2_array_index_2045174_comb;
  wire [7:0] p2_array_index_2045175_comb;
  wire [7:0] p2_array_index_2045176_comb;
  wire [7:0] p2_res7__164_comb;
  wire [7:0] p2_array_index_2045186_comb;
  wire [7:0] p2_array_index_2045187_comb;
  wire [7:0] p2_array_index_2045188_comb;
  wire [7:0] p2_array_index_2045189_comb;
  wire [7:0] p2_array_index_2045190_comb;
  wire [7:0] p2_res7__166_comb;
  wire [7:0] p2_array_index_2045201_comb;
  wire [7:0] p2_array_index_2045202_comb;
  wire [7:0] p2_array_index_2045203_comb;
  wire [7:0] p2_array_index_2045204_comb;
  wire [7:0] p2_res7__168_comb;
  wire [7:0] p2_array_index_2045214_comb;
  wire [7:0] p2_array_index_2045215_comb;
  wire [7:0] p2_array_index_2045216_comb;
  wire [7:0] p2_array_index_2045217_comb;
  wire [7:0] p2_res7__170_comb;
  wire [7:0] p2_array_index_2045228_comb;
  wire [7:0] p2_array_index_2045229_comb;
  wire [7:0] p2_array_index_2045230_comb;
  wire [7:0] p2_res7__172_comb;
  wire [7:0] p2_array_index_2045240_comb;
  wire [7:0] p2_array_index_2045241_comb;
  wire [7:0] p2_array_index_2045242_comb;
  wire [7:0] p2_res7__174_comb;
  wire [7:0] p2_array_index_2045253_comb;
  wire [7:0] p2_array_index_2045254_comb;
  wire [7:0] p2_res7__176_comb;
  wire [7:0] p2_array_index_2045264_comb;
  wire [7:0] p2_array_index_2045265_comb;
  wire [7:0] p2_res7__178_comb;
  wire [7:0] p2_array_index_2045276_comb;
  wire [7:0] p2_res7__180_comb;
  wire [7:0] p2_array_index_2045286_comb;
  wire [7:0] p2_res7__182_comb;
  wire [7:0] p2_res7__184_comb;
  wire [7:0] p2_res7__186_comb;
  wire [7:0] p2_res7__188_comb;
  wire [7:0] p2_res7__190_comb;
  wire [127:0] p2_res__5_comb;
  wire [127:0] p2_xor_2045326_comb;
  wire [127:0] p2_addedKey__38_comb;
  wire [7:0] p2_array_index_2045342_comb;
  wire [7:0] p2_array_index_2045343_comb;
  wire [7:0] p2_array_index_2045344_comb;
  wire [7:0] p2_array_index_2045345_comb;
  wire [7:0] p2_array_index_2045346_comb;
  wire [7:0] p2_array_index_2045347_comb;
  wire [7:0] p2_array_index_2045349_comb;
  wire [7:0] p2_array_index_2045351_comb;
  wire [7:0] p2_array_index_2045352_comb;
  wire [7:0] p2_array_index_2045353_comb;
  wire [7:0] p2_array_index_2045354_comb;
  wire [7:0] p2_array_index_2045355_comb;
  wire [7:0] p2_array_index_2045356_comb;
  wire [7:0] p2_array_index_2045358_comb;
  wire [7:0] p2_array_index_2045359_comb;
  wire [7:0] p2_array_index_2045360_comb;
  wire [7:0] p2_array_index_2045361_comb;
  wire [7:0] p2_array_index_2045362_comb;
  wire [7:0] p2_array_index_2045363_comb;
  wire [7:0] p2_array_index_2045364_comb;
  wire [7:0] p2_array_index_2045366_comb;
  wire [7:0] p2_res7__192_comb;
  wire [7:0] p2_array_index_2045375_comb;
  wire [7:0] p2_array_index_2045376_comb;
  wire [7:0] p2_array_index_2045377_comb;
  wire [7:0] p2_array_index_2045378_comb;
  wire [7:0] p2_array_index_2045379_comb;
  wire [7:0] p2_array_index_2045380_comb;
  wire [7:0] p2_res7__194_comb;
  wire [7:0] p2_array_index_2045390_comb;
  wire [7:0] p2_array_index_2045391_comb;
  wire [7:0] p2_array_index_2045392_comb;
  wire [7:0] p2_array_index_2045393_comb;
  wire [7:0] p2_array_index_2045394_comb;
  wire [7:0] p2_res7__196_comb;
  wire [7:0] p2_array_index_2045404_comb;
  wire [7:0] p2_array_index_2045405_comb;
  wire [7:0] p2_array_index_2045406_comb;
  wire [7:0] p2_array_index_2045407_comb;
  wire [7:0] p2_array_index_2045408_comb;
  wire [7:0] p2_res7__198_comb;
  wire [7:0] p2_array_index_2045419_comb;
  wire [7:0] p2_array_index_2045420_comb;
  wire [7:0] p2_array_index_2045421_comb;
  wire [7:0] p2_array_index_2045422_comb;
  wire [7:0] p2_res7__200_comb;
  wire [7:0] p2_array_index_2045432_comb;
  wire [7:0] p2_array_index_2045433_comb;
  wire [7:0] p2_array_index_2045434_comb;
  wire [7:0] p2_array_index_2045435_comb;
  wire [7:0] p2_res7__202_comb;
  wire [7:0] p2_array_index_2045446_comb;
  wire [7:0] p2_array_index_2045447_comb;
  wire [7:0] p2_array_index_2045448_comb;
  wire [7:0] p2_res7__204_comb;
  wire [7:0] p2_array_index_2045458_comb;
  wire [7:0] p2_array_index_2045459_comb;
  wire [7:0] p2_array_index_2045460_comb;
  wire [7:0] p2_res7__206_comb;
  wire [7:0] p2_array_index_2045471_comb;
  wire [7:0] p2_array_index_2045472_comb;
  wire [7:0] p2_res7__208_comb;
  wire [7:0] p2_array_index_2045482_comb;
  wire [7:0] p2_array_index_2045483_comb;
  wire [7:0] p2_res7__210_comb;
  wire [7:0] p2_array_index_2045494_comb;
  wire [7:0] p2_res7__212_comb;
  wire [7:0] p2_array_index_2045504_comb;
  wire [7:0] p2_res7__214_comb;
  wire [7:0] p2_res7__216_comb;
  wire [7:0] p2_res7__218_comb;
  wire [7:0] p2_res7__220_comb;
  wire [7:0] p2_res7__222_comb;
  wire [127:0] p2_res__6_comb;
  wire [127:0] p2_k3_comb;
  wire [127:0] p2_addedKey__39_comb;
  wire [7:0] p2_array_index_2045560_comb;
  wire [7:0] p2_array_index_2045561_comb;
  wire [7:0] p2_array_index_2045562_comb;
  wire [7:0] p2_array_index_2045563_comb;
  wire [7:0] p2_array_index_2045564_comb;
  wire [7:0] p2_array_index_2045565_comb;
  wire [7:0] p2_array_index_2045567_comb;
  wire [7:0] p2_array_index_2045569_comb;
  wire [7:0] p2_array_index_2045570_comb;
  wire [7:0] p2_array_index_2045571_comb;
  wire [7:0] p2_array_index_2045572_comb;
  wire [7:0] p2_array_index_2045573_comb;
  wire [7:0] p2_array_index_2045574_comb;
  wire [7:0] p2_array_index_2045576_comb;
  wire [7:0] p2_array_index_2045577_comb;
  wire [7:0] p2_array_index_2045578_comb;
  wire [7:0] p2_array_index_2045579_comb;
  wire [7:0] p2_array_index_2045580_comb;
  wire [7:0] p2_array_index_2045581_comb;
  wire [7:0] p2_array_index_2045582_comb;
  wire [7:0] p2_array_index_2045584_comb;
  wire [7:0] p2_res7__224_comb;
  wire [7:0] p2_array_index_2045593_comb;
  wire [7:0] p2_array_index_2045594_comb;
  wire [7:0] p2_array_index_2045595_comb;
  wire [7:0] p2_array_index_2045596_comb;
  wire [7:0] p2_array_index_2045597_comb;
  wire [7:0] p2_array_index_2045598_comb;
  wire [7:0] p2_res7__226_comb;
  wire [7:0] p2_array_index_2045608_comb;
  wire [7:0] p2_array_index_2045609_comb;
  wire [7:0] p2_array_index_2045610_comb;
  wire [7:0] p2_array_index_2045611_comb;
  wire [7:0] p2_array_index_2045612_comb;
  wire [7:0] p2_res7__228_comb;
  wire [7:0] p2_array_index_2045622_comb;
  wire [7:0] p2_array_index_2045623_comb;
  wire [7:0] p2_array_index_2045624_comb;
  wire [7:0] p2_array_index_2045625_comb;
  wire [7:0] p2_array_index_2045626_comb;
  wire [7:0] p2_res7__230_comb;
  wire [7:0] p2_array_index_2045637_comb;
  wire [7:0] p2_array_index_2045638_comb;
  wire [7:0] p2_array_index_2045639_comb;
  wire [7:0] p2_array_index_2045640_comb;
  wire [7:0] p2_res7__232_comb;
  wire [7:0] p2_array_index_2045650_comb;
  wire [7:0] p2_array_index_2045651_comb;
  wire [7:0] p2_array_index_2045652_comb;
  wire [7:0] p2_array_index_2045653_comb;
  wire [7:0] p2_res7__234_comb;
  wire [7:0] p2_array_index_2045664_comb;
  wire [7:0] p2_array_index_2045665_comb;
  wire [7:0] p2_array_index_2045666_comb;
  wire [7:0] p2_res7__236_comb;
  wire [7:0] p2_array_index_2045676_comb;
  wire [7:0] p2_array_index_2045677_comb;
  wire [7:0] p2_array_index_2045678_comb;
  wire [7:0] p2_res7__238_comb;
  wire [7:0] p2_array_index_2045689_comb;
  wire [7:0] p2_array_index_2045690_comb;
  wire [7:0] p2_res7__240_comb;
  wire [7:0] p2_array_index_2045700_comb;
  wire [7:0] p2_array_index_2045701_comb;
  wire [7:0] p2_res7__242_comb;
  wire [7:0] p2_array_index_2045712_comb;
  wire [7:0] p2_res7__244_comb;
  wire [7:0] p2_array_index_2045722_comb;
  wire [7:0] p2_res7__246_comb;
  wire [7:0] p2_res7__248_comb;
  wire [7:0] p2_res7__250_comb;
  wire [7:0] p2_res7__252_comb;
  wire [7:0] p2_res7__254_comb;
  wire [127:0] p2_res__7_comb;
  wire [127:0] p2_k2_comb;
  wire [127:0] p2_addedKey__40_comb;
  wire [7:0] p2_array_index_2045778_comb;
  wire [7:0] p2_array_index_2045779_comb;
  wire [7:0] p2_array_index_2045780_comb;
  wire [7:0] p2_array_index_2045781_comb;
  wire [7:0] p2_array_index_2045782_comb;
  wire [7:0] p2_array_index_2045783_comb;
  wire [7:0] p2_array_index_2045785_comb;
  wire [7:0] p2_array_index_2045787_comb;
  wire [7:0] p2_array_index_2045788_comb;
  wire [7:0] p2_array_index_2045789_comb;
  wire [7:0] p2_array_index_2045790_comb;
  wire [7:0] p2_array_index_2045791_comb;
  wire [7:0] p2_array_index_2045792_comb;
  wire [7:0] p2_array_index_2045794_comb;
  wire [7:0] p2_array_index_2045795_comb;
  wire [7:0] p2_array_index_2045796_comb;
  wire [7:0] p2_array_index_2045797_comb;
  wire [7:0] p2_array_index_2045798_comb;
  wire [7:0] p2_array_index_2045799_comb;
  wire [7:0] p2_array_index_2045800_comb;
  wire [7:0] p2_array_index_2045802_comb;
  wire [7:0] p2_res7__256_comb;
  wire [7:0] p2_array_index_2045811_comb;
  wire [7:0] p2_array_index_2045812_comb;
  wire [7:0] p2_array_index_2045813_comb;
  wire [7:0] p2_array_index_2045814_comb;
  wire [7:0] p2_array_index_2045815_comb;
  wire [7:0] p2_array_index_2045816_comb;
  wire [7:0] p2_res7__258_comb;
  wire [7:0] p2_array_index_2045826_comb;
  wire [7:0] p2_array_index_2045827_comb;
  wire [7:0] p2_array_index_2045828_comb;
  wire [7:0] p2_array_index_2045829_comb;
  wire [7:0] p2_array_index_2045830_comb;
  wire [7:0] p2_res7__260_comb;
  wire [7:0] p2_array_index_2045840_comb;
  wire [7:0] p2_array_index_2045841_comb;
  wire [7:0] p2_array_index_2045842_comb;
  wire [7:0] p2_array_index_2045843_comb;
  wire [7:0] p2_array_index_2045844_comb;
  wire [7:0] p2_res7__262_comb;
  wire [7:0] p2_array_index_2045855_comb;
  wire [7:0] p2_array_index_2045856_comb;
  wire [7:0] p2_array_index_2045857_comb;
  wire [7:0] p2_array_index_2045858_comb;
  wire [7:0] p2_res7__264_comb;
  wire [7:0] p2_array_index_2045868_comb;
  wire [7:0] p2_array_index_2045869_comb;
  wire [7:0] p2_array_index_2045870_comb;
  wire [7:0] p2_array_index_2045871_comb;
  wire [7:0] p2_res7__266_comb;
  wire [7:0] p2_array_index_2045882_comb;
  wire [7:0] p2_array_index_2045883_comb;
  wire [7:0] p2_array_index_2045884_comb;
  wire [7:0] p2_res7__268_comb;
  wire [7:0] p2_array_index_2045894_comb;
  wire [7:0] p2_array_index_2045895_comb;
  wire [7:0] p2_array_index_2045896_comb;
  wire [7:0] p2_res7__270_comb;
  wire [7:0] p2_array_index_2045907_comb;
  wire [7:0] p2_array_index_2045908_comb;
  wire [7:0] p2_res7__272_comb;
  wire [7:0] p2_array_index_2045918_comb;
  wire [7:0] p2_array_index_2045919_comb;
  wire [7:0] p2_res7__274_comb;
  wire [7:0] p2_array_index_2045930_comb;
  wire [7:0] p2_res7__276_comb;
  wire [7:0] p2_array_index_2045940_comb;
  wire [7:0] p2_res7__278_comb;
  wire [7:0] p2_res7__280_comb;
  wire [7:0] p2_res7__282_comb;
  wire [7:0] p2_array_index_2045963_comb;
  wire [7:0] p2_array_index_2045964_comb;
  wire [7:0] p2_array_index_2045965_comb;
  wire [7:0] p2_array_index_2045966_comb;
  wire [7:0] p2_array_index_2045967_comb;
  wire [7:0] p2_array_index_2045968_comb;
  wire [7:0] p2_array_index_2045969_comb;
  assign p2_array_index_2045022_comb = p1_literal_2043916[p1_res7__134];
  assign p2_array_index_2045023_comb = p1_literal_2043918[p1_res7__132];
  assign p2_array_index_2045024_comb = p1_literal_2043920[p1_res7__130];
  assign p2_res7__142_comb = p1_literal_2043910[p1_res7__140] ^ p1_literal_2043912[p1_res7__138] ^ p1_literal_2043914[p1_res7__136] ^ p2_array_index_2045022_comb ^ p2_array_index_2045023_comb ^ p2_array_index_2045024_comb ^ p1_res7__128 ^ p1_literal_2043923[p1_array_index_2044790] ^ p1_array_index_2044791 ^ p1_array_index_2044856 ^ p1_array_index_2044827 ^ p1_literal_2043916[p1_array_index_2044794] ^ p1_literal_2043914[p1_array_index_2044795] ^ p1_literal_2043912[p1_array_index_2044812] ^ p1_literal_2043910[p1_array_index_2044797] ^ p1_array_index_2044814;
  assign p2_array_index_2045035_comb = p1_literal_2043918[p1_res7__134];
  assign p2_array_index_2045036_comb = p1_literal_2043920[p1_res7__132];
  assign p2_res7__144_comb = p1_literal_2043910[p2_res7__142_comb] ^ p1_literal_2043912[p1_res7__140] ^ p1_literal_2043914[p1_res7__138] ^ p1_literal_2043916[p1_res7__136] ^ p2_array_index_2045035_comb ^ p2_array_index_2045036_comb ^ p1_res7__130 ^ p1_literal_2043923[p1_res7__128] ^ p1_array_index_2044790 ^ p1_array_index_2044870 ^ p1_array_index_2044841 ^ p1_array_index_2044809 ^ p1_literal_2043914[p1_array_index_2044794] ^ p1_literal_2043912[p1_array_index_2044795] ^ p1_literal_2043910[p1_array_index_2044812] ^ p1_array_index_2044797;
  assign p2_array_index_2045046_comb = p1_literal_2043918[p1_res7__136];
  assign p2_array_index_2045047_comb = p1_literal_2043920[p1_res7__134];
  assign p2_res7__146_comb = p1_literal_2043910[p2_res7__144_comb] ^ p1_literal_2043912[p2_res7__142_comb] ^ p1_literal_2043914[p1_res7__140] ^ p1_literal_2043916[p1_res7__138] ^ p2_array_index_2045046_comb ^ p2_array_index_2045047_comb ^ p1_res7__132 ^ p1_literal_2043923[p1_res7__130] ^ p1_res7__128 ^ p1_array_index_2044883 ^ p1_array_index_2044855 ^ p1_array_index_2044826 ^ p1_literal_2043914[p1_array_index_2044793] ^ p1_literal_2043912[p1_array_index_2044794] ^ p1_literal_2043910[p1_array_index_2044795] ^ p1_array_index_2044812;
  assign p2_array_index_2045058_comb = p1_literal_2043920[p1_res7__136];
  assign p2_res7__148_comb = p1_literal_2043910[p2_res7__146_comb] ^ p1_literal_2043912[p2_res7__144_comb] ^ p1_literal_2043914[p2_res7__142_comb] ^ p1_literal_2043916[p1_res7__140] ^ p1_literal_2043918[p1_res7__138] ^ p2_array_index_2045058_comb ^ p1_res7__134 ^ p1_literal_2043923[p1_res7__132] ^ p1_res7__130 ^ p1_array_index_2044896 ^ p1_array_index_2044869 ^ p1_array_index_2044840 ^ p1_array_index_2044808 ^ p1_literal_2043912[p1_array_index_2044793] ^ p1_literal_2043910[p1_array_index_2044794] ^ p1_array_index_2044795;
  assign p2_array_index_2045068_comb = p1_literal_2043920[p1_res7__138];
  assign p2_res7__150_comb = p1_literal_2043910[p2_res7__148_comb] ^ p1_literal_2043912[p2_res7__146_comb] ^ p1_literal_2043914[p2_res7__144_comb] ^ p1_literal_2043916[p2_res7__142_comb] ^ p1_literal_2043918[p1_res7__140] ^ p2_array_index_2045068_comb ^ p1_res7__136 ^ p1_literal_2043923[p1_res7__134] ^ p1_res7__132 ^ p2_array_index_2045024_comb ^ p1_array_index_2044882 ^ p1_array_index_2044854 ^ p1_array_index_2044825 ^ p1_literal_2043912[p1_array_index_2044792] ^ p1_literal_2043910[p1_array_index_2044793] ^ p1_array_index_2044794;
  assign p2_res7__152_comb = p1_literal_2043910[p2_res7__150_comb] ^ p1_literal_2043912[p2_res7__148_comb] ^ p1_literal_2043914[p2_res7__146_comb] ^ p1_literal_2043916[p2_res7__144_comb] ^ p1_literal_2043918[p2_res7__142_comb] ^ p1_literal_2043920[p1_res7__140] ^ p1_res7__138 ^ p1_literal_2043923[p1_res7__136] ^ p1_res7__134 ^ p2_array_index_2045036_comb ^ p1_array_index_2044895 ^ p1_array_index_2044868 ^ p1_array_index_2044839 ^ p1_array_index_2044807 ^ p1_literal_2043910[p1_array_index_2044792] ^ p1_array_index_2044793;
  assign p2_res7__154_comb = p1_literal_2043910[p2_res7__152_comb] ^ p1_literal_2043912[p2_res7__150_comb] ^ p1_literal_2043914[p2_res7__148_comb] ^ p1_literal_2043916[p2_res7__146_comb] ^ p1_literal_2043918[p2_res7__144_comb] ^ p1_literal_2043920[p2_res7__142_comb] ^ p1_res7__140 ^ p1_literal_2043923[p1_res7__138] ^ p1_res7__136 ^ p2_array_index_2045047_comb ^ p2_array_index_2045023_comb ^ p1_array_index_2044881 ^ p1_array_index_2044853 ^ p1_array_index_2044824 ^ p1_literal_2043910[p1_array_index_2044791] ^ p1_array_index_2044792;
  assign p2_res7__156_comb = p1_literal_2043910[p2_res7__154_comb] ^ p1_literal_2043912[p2_res7__152_comb] ^ p1_literal_2043914[p2_res7__150_comb] ^ p1_literal_2043916[p2_res7__148_comb] ^ p1_literal_2043918[p2_res7__146_comb] ^ p1_literal_2043920[p2_res7__144_comb] ^ p2_res7__142_comb ^ p1_literal_2043923[p1_res7__140] ^ p1_res7__138 ^ p2_array_index_2045058_comb ^ p2_array_index_2045035_comb ^ p1_array_index_2044894 ^ p1_array_index_2044867 ^ p1_array_index_2044838 ^ p1_array_index_2044806 ^ p1_array_index_2044791;
  assign p2_res7__158_comb = p1_literal_2043910[p2_res7__156_comb] ^ p1_literal_2043912[p2_res7__154_comb] ^ p1_literal_2043914[p2_res7__152_comb] ^ p1_literal_2043916[p2_res7__150_comb] ^ p1_literal_2043918[p2_res7__148_comb] ^ p1_literal_2043920[p2_res7__146_comb] ^ p2_res7__144_comb ^ p1_literal_2043923[p2_res7__142_comb] ^ p1_res7__140 ^ p2_array_index_2045068_comb ^ p2_array_index_2045046_comb ^ p2_array_index_2045022_comb ^ p1_array_index_2044880 ^ p1_array_index_2044852 ^ p1_array_index_2044823 ^ p1_array_index_2044790;
  assign p2_res__4_comb = {p2_res7__158_comb, p2_res7__156_comb, p2_res7__154_comb, p2_res7__152_comb, p2_res7__150_comb, p2_res7__148_comb, p2_res7__146_comb, p2_res7__144_comb, p2_res7__142_comb, p1_res7__140, p1_res7__138, p1_res7__136, p1_res7__134, p1_res7__132, p1_res7__130, p1_res7__128};
  assign p2_xor_2045108_comb = p2_res__4_comb ^ p1_xor_2044556;
  assign p2_addedKey__37_comb = p2_xor_2045108_comb ^ 128'ha74a_f7ef_ab73_df16_0dd2_0860_8b9e_fe06;
  assign p2_array_index_2045124_comb = p1_literal_2043896[p2_addedKey__37_comb[127:120]];
  assign p2_array_index_2045125_comb = p1_literal_2043896[p2_addedKey__37_comb[119:112]];
  assign p2_array_index_2045126_comb = p1_literal_2043896[p2_addedKey__37_comb[111:104]];
  assign p2_array_index_2045127_comb = p1_literal_2043896[p2_addedKey__37_comb[103:96]];
  assign p2_array_index_2045128_comb = p1_literal_2043896[p2_addedKey__37_comb[95:88]];
  assign p2_array_index_2045129_comb = p1_literal_2043896[p2_addedKey__37_comb[87:80]];
  assign p2_array_index_2045131_comb = p1_literal_2043896[p2_addedKey__37_comb[71:64]];
  assign p2_array_index_2045133_comb = p1_literal_2043896[p2_addedKey__37_comb[55:48]];
  assign p2_array_index_2045134_comb = p1_literal_2043896[p2_addedKey__37_comb[47:40]];
  assign p2_array_index_2045135_comb = p1_literal_2043896[p2_addedKey__37_comb[39:32]];
  assign p2_array_index_2045136_comb = p1_literal_2043896[p2_addedKey__37_comb[31:24]];
  assign p2_array_index_2045137_comb = p1_literal_2043896[p2_addedKey__37_comb[23:16]];
  assign p2_array_index_2045138_comb = p1_literal_2043896[p2_addedKey__37_comb[15:8]];
  assign p2_array_index_2045140_comb = p1_literal_2043910[p2_array_index_2045124_comb];
  assign p2_array_index_2045141_comb = p1_literal_2043912[p2_array_index_2045125_comb];
  assign p2_array_index_2045142_comb = p1_literal_2043914[p2_array_index_2045126_comb];
  assign p2_array_index_2045143_comb = p1_literal_2043916[p2_array_index_2045127_comb];
  assign p2_array_index_2045144_comb = p1_literal_2043918[p2_array_index_2045128_comb];
  assign p2_array_index_2045145_comb = p1_literal_2043920[p2_array_index_2045129_comb];
  assign p2_array_index_2045146_comb = p1_literal_2043896[p2_addedKey__37_comb[79:72]];
  assign p2_array_index_2045148_comb = p1_literal_2043896[p2_addedKey__37_comb[63:56]];
  assign p2_res7__160_comb = p2_array_index_2045140_comb ^ p2_array_index_2045141_comb ^ p2_array_index_2045142_comb ^ p2_array_index_2045143_comb ^ p2_array_index_2045144_comb ^ p2_array_index_2045145_comb ^ p2_array_index_2045146_comb ^ p1_literal_2043923[p2_array_index_2045131_comb] ^ p2_array_index_2045148_comb ^ p1_literal_2043920[p2_array_index_2045133_comb] ^ p1_literal_2043918[p2_array_index_2045134_comb] ^ p1_literal_2043916[p2_array_index_2045135_comb] ^ p1_literal_2043914[p2_array_index_2045136_comb] ^ p1_literal_2043912[p2_array_index_2045137_comb] ^ p1_literal_2043910[p2_array_index_2045138_comb] ^ p1_literal_2043896[p2_addedKey__37_comb[7:0]];
  assign p2_array_index_2045157_comb = p1_literal_2043910[p2_res7__160_comb];
  assign p2_array_index_2045158_comb = p1_literal_2043912[p2_array_index_2045124_comb];
  assign p2_array_index_2045159_comb = p1_literal_2043914[p2_array_index_2045125_comb];
  assign p2_array_index_2045160_comb = p1_literal_2043916[p2_array_index_2045126_comb];
  assign p2_array_index_2045161_comb = p1_literal_2043918[p2_array_index_2045127_comb];
  assign p2_array_index_2045162_comb = p1_literal_2043920[p2_array_index_2045128_comb];
  assign p2_res7__162_comb = p2_array_index_2045157_comb ^ p2_array_index_2045158_comb ^ p2_array_index_2045159_comb ^ p2_array_index_2045160_comb ^ p2_array_index_2045161_comb ^ p2_array_index_2045162_comb ^ p2_array_index_2045129_comb ^ p1_literal_2043923[p2_array_index_2045146_comb] ^ p2_array_index_2045131_comb ^ p1_literal_2043920[p2_array_index_2045148_comb] ^ p1_literal_2043918[p2_array_index_2045133_comb] ^ p1_literal_2043916[p2_array_index_2045134_comb] ^ p1_literal_2043914[p2_array_index_2045135_comb] ^ p1_literal_2043912[p2_array_index_2045136_comb] ^ p1_literal_2043910[p2_array_index_2045137_comb] ^ p2_array_index_2045138_comb;
  assign p2_array_index_2045172_comb = p1_literal_2043912[p2_res7__160_comb];
  assign p2_array_index_2045173_comb = p1_literal_2043914[p2_array_index_2045124_comb];
  assign p2_array_index_2045174_comb = p1_literal_2043916[p2_array_index_2045125_comb];
  assign p2_array_index_2045175_comb = p1_literal_2043918[p2_array_index_2045126_comb];
  assign p2_array_index_2045176_comb = p1_literal_2043920[p2_array_index_2045127_comb];
  assign p2_res7__164_comb = p1_literal_2043910[p2_res7__162_comb] ^ p2_array_index_2045172_comb ^ p2_array_index_2045173_comb ^ p2_array_index_2045174_comb ^ p2_array_index_2045175_comb ^ p2_array_index_2045176_comb ^ p2_array_index_2045128_comb ^ p1_literal_2043923[p2_array_index_2045129_comb] ^ p2_array_index_2045146_comb ^ p1_literal_2043920[p2_array_index_2045131_comb] ^ p1_literal_2043918[p2_array_index_2045148_comb] ^ p1_literal_2043916[p2_array_index_2045133_comb] ^ p1_literal_2043914[p2_array_index_2045134_comb] ^ p1_literal_2043912[p2_array_index_2045135_comb] ^ p1_literal_2043910[p2_array_index_2045136_comb] ^ p2_array_index_2045137_comb;
  assign p2_array_index_2045186_comb = p1_literal_2043912[p2_res7__162_comb];
  assign p2_array_index_2045187_comb = p1_literal_2043914[p2_res7__160_comb];
  assign p2_array_index_2045188_comb = p1_literal_2043916[p2_array_index_2045124_comb];
  assign p2_array_index_2045189_comb = p1_literal_2043918[p2_array_index_2045125_comb];
  assign p2_array_index_2045190_comb = p1_literal_2043920[p2_array_index_2045126_comb];
  assign p2_res7__166_comb = p1_literal_2043910[p2_res7__164_comb] ^ p2_array_index_2045186_comb ^ p2_array_index_2045187_comb ^ p2_array_index_2045188_comb ^ p2_array_index_2045189_comb ^ p2_array_index_2045190_comb ^ p2_array_index_2045127_comb ^ p1_literal_2043923[p2_array_index_2045128_comb] ^ p2_array_index_2045129_comb ^ p1_literal_2043920[p2_array_index_2045146_comb] ^ p1_literal_2043918[p2_array_index_2045131_comb] ^ p1_literal_2043916[p2_array_index_2045148_comb] ^ p1_literal_2043914[p2_array_index_2045133_comb] ^ p1_literal_2043912[p2_array_index_2045134_comb] ^ p1_literal_2043910[p2_array_index_2045135_comb] ^ p2_array_index_2045136_comb;
  assign p2_array_index_2045201_comb = p1_literal_2043914[p2_res7__162_comb];
  assign p2_array_index_2045202_comb = p1_literal_2043916[p2_res7__160_comb];
  assign p2_array_index_2045203_comb = p1_literal_2043918[p2_array_index_2045124_comb];
  assign p2_array_index_2045204_comb = p1_literal_2043920[p2_array_index_2045125_comb];
  assign p2_res7__168_comb = p1_literal_2043910[p2_res7__166_comb] ^ p1_literal_2043912[p2_res7__164_comb] ^ p2_array_index_2045201_comb ^ p2_array_index_2045202_comb ^ p2_array_index_2045203_comb ^ p2_array_index_2045204_comb ^ p2_array_index_2045126_comb ^ p1_literal_2043923[p2_array_index_2045127_comb] ^ p2_array_index_2045128_comb ^ p2_array_index_2045145_comb ^ p1_literal_2043918[p2_array_index_2045146_comb] ^ p1_literal_2043916[p2_array_index_2045131_comb] ^ p1_literal_2043914[p2_array_index_2045148_comb] ^ p1_literal_2043912[p2_array_index_2045133_comb] ^ p1_literal_2043910[p2_array_index_2045134_comb] ^ p2_array_index_2045135_comb;
  assign p2_array_index_2045214_comb = p1_literal_2043914[p2_res7__164_comb];
  assign p2_array_index_2045215_comb = p1_literal_2043916[p2_res7__162_comb];
  assign p2_array_index_2045216_comb = p1_literal_2043918[p2_res7__160_comb];
  assign p2_array_index_2045217_comb = p1_literal_2043920[p2_array_index_2045124_comb];
  assign p2_res7__170_comb = p1_literal_2043910[p2_res7__168_comb] ^ p1_literal_2043912[p2_res7__166_comb] ^ p2_array_index_2045214_comb ^ p2_array_index_2045215_comb ^ p2_array_index_2045216_comb ^ p2_array_index_2045217_comb ^ p2_array_index_2045125_comb ^ p1_literal_2043923[p2_array_index_2045126_comb] ^ p2_array_index_2045127_comb ^ p2_array_index_2045162_comb ^ p1_literal_2043918[p2_array_index_2045129_comb] ^ p1_literal_2043916[p2_array_index_2045146_comb] ^ p1_literal_2043914[p2_array_index_2045131_comb] ^ p1_literal_2043912[p2_array_index_2045148_comb] ^ p1_literal_2043910[p2_array_index_2045133_comb] ^ p2_array_index_2045134_comb;
  assign p2_array_index_2045228_comb = p1_literal_2043916[p2_res7__164_comb];
  assign p2_array_index_2045229_comb = p1_literal_2043918[p2_res7__162_comb];
  assign p2_array_index_2045230_comb = p1_literal_2043920[p2_res7__160_comb];
  assign p2_res7__172_comb = p1_literal_2043910[p2_res7__170_comb] ^ p1_literal_2043912[p2_res7__168_comb] ^ p1_literal_2043914[p2_res7__166_comb] ^ p2_array_index_2045228_comb ^ p2_array_index_2045229_comb ^ p2_array_index_2045230_comb ^ p2_array_index_2045124_comb ^ p1_literal_2043923[p2_array_index_2045125_comb] ^ p2_array_index_2045126_comb ^ p2_array_index_2045176_comb ^ p2_array_index_2045144_comb ^ p1_literal_2043916[p2_array_index_2045129_comb] ^ p1_literal_2043914[p2_array_index_2045146_comb] ^ p1_literal_2043912[p2_array_index_2045131_comb] ^ p1_literal_2043910[p2_array_index_2045148_comb] ^ p2_array_index_2045133_comb;
  assign p2_array_index_2045240_comb = p1_literal_2043916[p2_res7__166_comb];
  assign p2_array_index_2045241_comb = p1_literal_2043918[p2_res7__164_comb];
  assign p2_array_index_2045242_comb = p1_literal_2043920[p2_res7__162_comb];
  assign p2_res7__174_comb = p1_literal_2043910[p2_res7__172_comb] ^ p1_literal_2043912[p2_res7__170_comb] ^ p1_literal_2043914[p2_res7__168_comb] ^ p2_array_index_2045240_comb ^ p2_array_index_2045241_comb ^ p2_array_index_2045242_comb ^ p2_res7__160_comb ^ p1_literal_2043923[p2_array_index_2045124_comb] ^ p2_array_index_2045125_comb ^ p2_array_index_2045190_comb ^ p2_array_index_2045161_comb ^ p1_literal_2043916[p2_array_index_2045128_comb] ^ p1_literal_2043914[p2_array_index_2045129_comb] ^ p1_literal_2043912[p2_array_index_2045146_comb] ^ p1_literal_2043910[p2_array_index_2045131_comb] ^ p2_array_index_2045148_comb;
  assign p2_array_index_2045253_comb = p1_literal_2043918[p2_res7__166_comb];
  assign p2_array_index_2045254_comb = p1_literal_2043920[p2_res7__164_comb];
  assign p2_res7__176_comb = p1_literal_2043910[p2_res7__174_comb] ^ p1_literal_2043912[p2_res7__172_comb] ^ p1_literal_2043914[p2_res7__170_comb] ^ p1_literal_2043916[p2_res7__168_comb] ^ p2_array_index_2045253_comb ^ p2_array_index_2045254_comb ^ p2_res7__162_comb ^ p1_literal_2043923[p2_res7__160_comb] ^ p2_array_index_2045124_comb ^ p2_array_index_2045204_comb ^ p2_array_index_2045175_comb ^ p2_array_index_2045143_comb ^ p1_literal_2043914[p2_array_index_2045128_comb] ^ p1_literal_2043912[p2_array_index_2045129_comb] ^ p1_literal_2043910[p2_array_index_2045146_comb] ^ p2_array_index_2045131_comb;
  assign p2_array_index_2045264_comb = p1_literal_2043918[p2_res7__168_comb];
  assign p2_array_index_2045265_comb = p1_literal_2043920[p2_res7__166_comb];
  assign p2_res7__178_comb = p1_literal_2043910[p2_res7__176_comb] ^ p1_literal_2043912[p2_res7__174_comb] ^ p1_literal_2043914[p2_res7__172_comb] ^ p1_literal_2043916[p2_res7__170_comb] ^ p2_array_index_2045264_comb ^ p2_array_index_2045265_comb ^ p2_res7__164_comb ^ p1_literal_2043923[p2_res7__162_comb] ^ p2_res7__160_comb ^ p2_array_index_2045217_comb ^ p2_array_index_2045189_comb ^ p2_array_index_2045160_comb ^ p1_literal_2043914[p2_array_index_2045127_comb] ^ p1_literal_2043912[p2_array_index_2045128_comb] ^ p1_literal_2043910[p2_array_index_2045129_comb] ^ p2_array_index_2045146_comb;
  assign p2_array_index_2045276_comb = p1_literal_2043920[p2_res7__168_comb];
  assign p2_res7__180_comb = p1_literal_2043910[p2_res7__178_comb] ^ p1_literal_2043912[p2_res7__176_comb] ^ p1_literal_2043914[p2_res7__174_comb] ^ p1_literal_2043916[p2_res7__172_comb] ^ p1_literal_2043918[p2_res7__170_comb] ^ p2_array_index_2045276_comb ^ p2_res7__166_comb ^ p1_literal_2043923[p2_res7__164_comb] ^ p2_res7__162_comb ^ p2_array_index_2045230_comb ^ p2_array_index_2045203_comb ^ p2_array_index_2045174_comb ^ p2_array_index_2045142_comb ^ p1_literal_2043912[p2_array_index_2045127_comb] ^ p1_literal_2043910[p2_array_index_2045128_comb] ^ p2_array_index_2045129_comb;
  assign p2_array_index_2045286_comb = p1_literal_2043920[p2_res7__170_comb];
  assign p2_res7__182_comb = p1_literal_2043910[p2_res7__180_comb] ^ p1_literal_2043912[p2_res7__178_comb] ^ p1_literal_2043914[p2_res7__176_comb] ^ p1_literal_2043916[p2_res7__174_comb] ^ p1_literal_2043918[p2_res7__172_comb] ^ p2_array_index_2045286_comb ^ p2_res7__168_comb ^ p1_literal_2043923[p2_res7__166_comb] ^ p2_res7__164_comb ^ p2_array_index_2045242_comb ^ p2_array_index_2045216_comb ^ p2_array_index_2045188_comb ^ p2_array_index_2045159_comb ^ p1_literal_2043912[p2_array_index_2045126_comb] ^ p1_literal_2043910[p2_array_index_2045127_comb] ^ p2_array_index_2045128_comb;
  assign p2_res7__184_comb = p1_literal_2043910[p2_res7__182_comb] ^ p1_literal_2043912[p2_res7__180_comb] ^ p1_literal_2043914[p2_res7__178_comb] ^ p1_literal_2043916[p2_res7__176_comb] ^ p1_literal_2043918[p2_res7__174_comb] ^ p1_literal_2043920[p2_res7__172_comb] ^ p2_res7__170_comb ^ p1_literal_2043923[p2_res7__168_comb] ^ p2_res7__166_comb ^ p2_array_index_2045254_comb ^ p2_array_index_2045229_comb ^ p2_array_index_2045202_comb ^ p2_array_index_2045173_comb ^ p2_array_index_2045141_comb ^ p1_literal_2043910[p2_array_index_2045126_comb] ^ p2_array_index_2045127_comb;
  assign p2_res7__186_comb = p1_literal_2043910[p2_res7__184_comb] ^ p1_literal_2043912[p2_res7__182_comb] ^ p1_literal_2043914[p2_res7__180_comb] ^ p1_literal_2043916[p2_res7__178_comb] ^ p1_literal_2043918[p2_res7__176_comb] ^ p1_literal_2043920[p2_res7__174_comb] ^ p2_res7__172_comb ^ p1_literal_2043923[p2_res7__170_comb] ^ p2_res7__168_comb ^ p2_array_index_2045265_comb ^ p2_array_index_2045241_comb ^ p2_array_index_2045215_comb ^ p2_array_index_2045187_comb ^ p2_array_index_2045158_comb ^ p1_literal_2043910[p2_array_index_2045125_comb] ^ p2_array_index_2045126_comb;
  assign p2_res7__188_comb = p1_literal_2043910[p2_res7__186_comb] ^ p1_literal_2043912[p2_res7__184_comb] ^ p1_literal_2043914[p2_res7__182_comb] ^ p1_literal_2043916[p2_res7__180_comb] ^ p1_literal_2043918[p2_res7__178_comb] ^ p1_literal_2043920[p2_res7__176_comb] ^ p2_res7__174_comb ^ p1_literal_2043923[p2_res7__172_comb] ^ p2_res7__170_comb ^ p2_array_index_2045276_comb ^ p2_array_index_2045253_comb ^ p2_array_index_2045228_comb ^ p2_array_index_2045201_comb ^ p2_array_index_2045172_comb ^ p2_array_index_2045140_comb ^ p2_array_index_2045125_comb;
  assign p2_res7__190_comb = p1_literal_2043910[p2_res7__188_comb] ^ p1_literal_2043912[p2_res7__186_comb] ^ p1_literal_2043914[p2_res7__184_comb] ^ p1_literal_2043916[p2_res7__182_comb] ^ p1_literal_2043918[p2_res7__180_comb] ^ p1_literal_2043920[p2_res7__178_comb] ^ p2_res7__176_comb ^ p1_literal_2043923[p2_res7__174_comb] ^ p2_res7__172_comb ^ p2_array_index_2045286_comb ^ p2_array_index_2045264_comb ^ p2_array_index_2045240_comb ^ p2_array_index_2045214_comb ^ p2_array_index_2045186_comb ^ p2_array_index_2045157_comb ^ p2_array_index_2045124_comb;
  assign p2_res__5_comb = {p2_res7__190_comb, p2_res7__188_comb, p2_res7__186_comb, p2_res7__184_comb, p2_res7__182_comb, p2_res7__180_comb, p2_res7__178_comb, p2_res7__176_comb, p2_res7__174_comb, p2_res7__172_comb, p2_res7__170_comb, p2_res7__168_comb, p2_res7__166_comb, p2_res7__164_comb, p2_res7__162_comb, p2_res7__160_comb};
  assign p2_xor_2045326_comb = p2_res__5_comb ^ p1_xor_2044774;
  assign p2_addedKey__38_comb = p2_xor_2045326_comb ^ 128'hc9e8_819d_c73b_a5ae_50f5_b570_561a_6a07;
  assign p2_array_index_2045342_comb = p1_literal_2043896[p2_addedKey__38_comb[127:120]];
  assign p2_array_index_2045343_comb = p1_literal_2043896[p2_addedKey__38_comb[119:112]];
  assign p2_array_index_2045344_comb = p1_literal_2043896[p2_addedKey__38_comb[111:104]];
  assign p2_array_index_2045345_comb = p1_literal_2043896[p2_addedKey__38_comb[103:96]];
  assign p2_array_index_2045346_comb = p1_literal_2043896[p2_addedKey__38_comb[95:88]];
  assign p2_array_index_2045347_comb = p1_literal_2043896[p2_addedKey__38_comb[87:80]];
  assign p2_array_index_2045349_comb = p1_literal_2043896[p2_addedKey__38_comb[71:64]];
  assign p2_array_index_2045351_comb = p1_literal_2043896[p2_addedKey__38_comb[55:48]];
  assign p2_array_index_2045352_comb = p1_literal_2043896[p2_addedKey__38_comb[47:40]];
  assign p2_array_index_2045353_comb = p1_literal_2043896[p2_addedKey__38_comb[39:32]];
  assign p2_array_index_2045354_comb = p1_literal_2043896[p2_addedKey__38_comb[31:24]];
  assign p2_array_index_2045355_comb = p1_literal_2043896[p2_addedKey__38_comb[23:16]];
  assign p2_array_index_2045356_comb = p1_literal_2043896[p2_addedKey__38_comb[15:8]];
  assign p2_array_index_2045358_comb = p1_literal_2043910[p2_array_index_2045342_comb];
  assign p2_array_index_2045359_comb = p1_literal_2043912[p2_array_index_2045343_comb];
  assign p2_array_index_2045360_comb = p1_literal_2043914[p2_array_index_2045344_comb];
  assign p2_array_index_2045361_comb = p1_literal_2043916[p2_array_index_2045345_comb];
  assign p2_array_index_2045362_comb = p1_literal_2043918[p2_array_index_2045346_comb];
  assign p2_array_index_2045363_comb = p1_literal_2043920[p2_array_index_2045347_comb];
  assign p2_array_index_2045364_comb = p1_literal_2043896[p2_addedKey__38_comb[79:72]];
  assign p2_array_index_2045366_comb = p1_literal_2043896[p2_addedKey__38_comb[63:56]];
  assign p2_res7__192_comb = p2_array_index_2045358_comb ^ p2_array_index_2045359_comb ^ p2_array_index_2045360_comb ^ p2_array_index_2045361_comb ^ p2_array_index_2045362_comb ^ p2_array_index_2045363_comb ^ p2_array_index_2045364_comb ^ p1_literal_2043923[p2_array_index_2045349_comb] ^ p2_array_index_2045366_comb ^ p1_literal_2043920[p2_array_index_2045351_comb] ^ p1_literal_2043918[p2_array_index_2045352_comb] ^ p1_literal_2043916[p2_array_index_2045353_comb] ^ p1_literal_2043914[p2_array_index_2045354_comb] ^ p1_literal_2043912[p2_array_index_2045355_comb] ^ p1_literal_2043910[p2_array_index_2045356_comb] ^ p1_literal_2043896[p2_addedKey__38_comb[7:0]];
  assign p2_array_index_2045375_comb = p1_literal_2043910[p2_res7__192_comb];
  assign p2_array_index_2045376_comb = p1_literal_2043912[p2_array_index_2045342_comb];
  assign p2_array_index_2045377_comb = p1_literal_2043914[p2_array_index_2045343_comb];
  assign p2_array_index_2045378_comb = p1_literal_2043916[p2_array_index_2045344_comb];
  assign p2_array_index_2045379_comb = p1_literal_2043918[p2_array_index_2045345_comb];
  assign p2_array_index_2045380_comb = p1_literal_2043920[p2_array_index_2045346_comb];
  assign p2_res7__194_comb = p2_array_index_2045375_comb ^ p2_array_index_2045376_comb ^ p2_array_index_2045377_comb ^ p2_array_index_2045378_comb ^ p2_array_index_2045379_comb ^ p2_array_index_2045380_comb ^ p2_array_index_2045347_comb ^ p1_literal_2043923[p2_array_index_2045364_comb] ^ p2_array_index_2045349_comb ^ p1_literal_2043920[p2_array_index_2045366_comb] ^ p1_literal_2043918[p2_array_index_2045351_comb] ^ p1_literal_2043916[p2_array_index_2045352_comb] ^ p1_literal_2043914[p2_array_index_2045353_comb] ^ p1_literal_2043912[p2_array_index_2045354_comb] ^ p1_literal_2043910[p2_array_index_2045355_comb] ^ p2_array_index_2045356_comb;
  assign p2_array_index_2045390_comb = p1_literal_2043912[p2_res7__192_comb];
  assign p2_array_index_2045391_comb = p1_literal_2043914[p2_array_index_2045342_comb];
  assign p2_array_index_2045392_comb = p1_literal_2043916[p2_array_index_2045343_comb];
  assign p2_array_index_2045393_comb = p1_literal_2043918[p2_array_index_2045344_comb];
  assign p2_array_index_2045394_comb = p1_literal_2043920[p2_array_index_2045345_comb];
  assign p2_res7__196_comb = p1_literal_2043910[p2_res7__194_comb] ^ p2_array_index_2045390_comb ^ p2_array_index_2045391_comb ^ p2_array_index_2045392_comb ^ p2_array_index_2045393_comb ^ p2_array_index_2045394_comb ^ p2_array_index_2045346_comb ^ p1_literal_2043923[p2_array_index_2045347_comb] ^ p2_array_index_2045364_comb ^ p1_literal_2043920[p2_array_index_2045349_comb] ^ p1_literal_2043918[p2_array_index_2045366_comb] ^ p1_literal_2043916[p2_array_index_2045351_comb] ^ p1_literal_2043914[p2_array_index_2045352_comb] ^ p1_literal_2043912[p2_array_index_2045353_comb] ^ p1_literal_2043910[p2_array_index_2045354_comb] ^ p2_array_index_2045355_comb;
  assign p2_array_index_2045404_comb = p1_literal_2043912[p2_res7__194_comb];
  assign p2_array_index_2045405_comb = p1_literal_2043914[p2_res7__192_comb];
  assign p2_array_index_2045406_comb = p1_literal_2043916[p2_array_index_2045342_comb];
  assign p2_array_index_2045407_comb = p1_literal_2043918[p2_array_index_2045343_comb];
  assign p2_array_index_2045408_comb = p1_literal_2043920[p2_array_index_2045344_comb];
  assign p2_res7__198_comb = p1_literal_2043910[p2_res7__196_comb] ^ p2_array_index_2045404_comb ^ p2_array_index_2045405_comb ^ p2_array_index_2045406_comb ^ p2_array_index_2045407_comb ^ p2_array_index_2045408_comb ^ p2_array_index_2045345_comb ^ p1_literal_2043923[p2_array_index_2045346_comb] ^ p2_array_index_2045347_comb ^ p1_literal_2043920[p2_array_index_2045364_comb] ^ p1_literal_2043918[p2_array_index_2045349_comb] ^ p1_literal_2043916[p2_array_index_2045366_comb] ^ p1_literal_2043914[p2_array_index_2045351_comb] ^ p1_literal_2043912[p2_array_index_2045352_comb] ^ p1_literal_2043910[p2_array_index_2045353_comb] ^ p2_array_index_2045354_comb;
  assign p2_array_index_2045419_comb = p1_literal_2043914[p2_res7__194_comb];
  assign p2_array_index_2045420_comb = p1_literal_2043916[p2_res7__192_comb];
  assign p2_array_index_2045421_comb = p1_literal_2043918[p2_array_index_2045342_comb];
  assign p2_array_index_2045422_comb = p1_literal_2043920[p2_array_index_2045343_comb];
  assign p2_res7__200_comb = p1_literal_2043910[p2_res7__198_comb] ^ p1_literal_2043912[p2_res7__196_comb] ^ p2_array_index_2045419_comb ^ p2_array_index_2045420_comb ^ p2_array_index_2045421_comb ^ p2_array_index_2045422_comb ^ p2_array_index_2045344_comb ^ p1_literal_2043923[p2_array_index_2045345_comb] ^ p2_array_index_2045346_comb ^ p2_array_index_2045363_comb ^ p1_literal_2043918[p2_array_index_2045364_comb] ^ p1_literal_2043916[p2_array_index_2045349_comb] ^ p1_literal_2043914[p2_array_index_2045366_comb] ^ p1_literal_2043912[p2_array_index_2045351_comb] ^ p1_literal_2043910[p2_array_index_2045352_comb] ^ p2_array_index_2045353_comb;
  assign p2_array_index_2045432_comb = p1_literal_2043914[p2_res7__196_comb];
  assign p2_array_index_2045433_comb = p1_literal_2043916[p2_res7__194_comb];
  assign p2_array_index_2045434_comb = p1_literal_2043918[p2_res7__192_comb];
  assign p2_array_index_2045435_comb = p1_literal_2043920[p2_array_index_2045342_comb];
  assign p2_res7__202_comb = p1_literal_2043910[p2_res7__200_comb] ^ p1_literal_2043912[p2_res7__198_comb] ^ p2_array_index_2045432_comb ^ p2_array_index_2045433_comb ^ p2_array_index_2045434_comb ^ p2_array_index_2045435_comb ^ p2_array_index_2045343_comb ^ p1_literal_2043923[p2_array_index_2045344_comb] ^ p2_array_index_2045345_comb ^ p2_array_index_2045380_comb ^ p1_literal_2043918[p2_array_index_2045347_comb] ^ p1_literal_2043916[p2_array_index_2045364_comb] ^ p1_literal_2043914[p2_array_index_2045349_comb] ^ p1_literal_2043912[p2_array_index_2045366_comb] ^ p1_literal_2043910[p2_array_index_2045351_comb] ^ p2_array_index_2045352_comb;
  assign p2_array_index_2045446_comb = p1_literal_2043916[p2_res7__196_comb];
  assign p2_array_index_2045447_comb = p1_literal_2043918[p2_res7__194_comb];
  assign p2_array_index_2045448_comb = p1_literal_2043920[p2_res7__192_comb];
  assign p2_res7__204_comb = p1_literal_2043910[p2_res7__202_comb] ^ p1_literal_2043912[p2_res7__200_comb] ^ p1_literal_2043914[p2_res7__198_comb] ^ p2_array_index_2045446_comb ^ p2_array_index_2045447_comb ^ p2_array_index_2045448_comb ^ p2_array_index_2045342_comb ^ p1_literal_2043923[p2_array_index_2045343_comb] ^ p2_array_index_2045344_comb ^ p2_array_index_2045394_comb ^ p2_array_index_2045362_comb ^ p1_literal_2043916[p2_array_index_2045347_comb] ^ p1_literal_2043914[p2_array_index_2045364_comb] ^ p1_literal_2043912[p2_array_index_2045349_comb] ^ p1_literal_2043910[p2_array_index_2045366_comb] ^ p2_array_index_2045351_comb;
  assign p2_array_index_2045458_comb = p1_literal_2043916[p2_res7__198_comb];
  assign p2_array_index_2045459_comb = p1_literal_2043918[p2_res7__196_comb];
  assign p2_array_index_2045460_comb = p1_literal_2043920[p2_res7__194_comb];
  assign p2_res7__206_comb = p1_literal_2043910[p2_res7__204_comb] ^ p1_literal_2043912[p2_res7__202_comb] ^ p1_literal_2043914[p2_res7__200_comb] ^ p2_array_index_2045458_comb ^ p2_array_index_2045459_comb ^ p2_array_index_2045460_comb ^ p2_res7__192_comb ^ p1_literal_2043923[p2_array_index_2045342_comb] ^ p2_array_index_2045343_comb ^ p2_array_index_2045408_comb ^ p2_array_index_2045379_comb ^ p1_literal_2043916[p2_array_index_2045346_comb] ^ p1_literal_2043914[p2_array_index_2045347_comb] ^ p1_literal_2043912[p2_array_index_2045364_comb] ^ p1_literal_2043910[p2_array_index_2045349_comb] ^ p2_array_index_2045366_comb;
  assign p2_array_index_2045471_comb = p1_literal_2043918[p2_res7__198_comb];
  assign p2_array_index_2045472_comb = p1_literal_2043920[p2_res7__196_comb];
  assign p2_res7__208_comb = p1_literal_2043910[p2_res7__206_comb] ^ p1_literal_2043912[p2_res7__204_comb] ^ p1_literal_2043914[p2_res7__202_comb] ^ p1_literal_2043916[p2_res7__200_comb] ^ p2_array_index_2045471_comb ^ p2_array_index_2045472_comb ^ p2_res7__194_comb ^ p1_literal_2043923[p2_res7__192_comb] ^ p2_array_index_2045342_comb ^ p2_array_index_2045422_comb ^ p2_array_index_2045393_comb ^ p2_array_index_2045361_comb ^ p1_literal_2043914[p2_array_index_2045346_comb] ^ p1_literal_2043912[p2_array_index_2045347_comb] ^ p1_literal_2043910[p2_array_index_2045364_comb] ^ p2_array_index_2045349_comb;
  assign p2_array_index_2045482_comb = p1_literal_2043918[p2_res7__200_comb];
  assign p2_array_index_2045483_comb = p1_literal_2043920[p2_res7__198_comb];
  assign p2_res7__210_comb = p1_literal_2043910[p2_res7__208_comb] ^ p1_literal_2043912[p2_res7__206_comb] ^ p1_literal_2043914[p2_res7__204_comb] ^ p1_literal_2043916[p2_res7__202_comb] ^ p2_array_index_2045482_comb ^ p2_array_index_2045483_comb ^ p2_res7__196_comb ^ p1_literal_2043923[p2_res7__194_comb] ^ p2_res7__192_comb ^ p2_array_index_2045435_comb ^ p2_array_index_2045407_comb ^ p2_array_index_2045378_comb ^ p1_literal_2043914[p2_array_index_2045345_comb] ^ p1_literal_2043912[p2_array_index_2045346_comb] ^ p1_literal_2043910[p2_array_index_2045347_comb] ^ p2_array_index_2045364_comb;
  assign p2_array_index_2045494_comb = p1_literal_2043920[p2_res7__200_comb];
  assign p2_res7__212_comb = p1_literal_2043910[p2_res7__210_comb] ^ p1_literal_2043912[p2_res7__208_comb] ^ p1_literal_2043914[p2_res7__206_comb] ^ p1_literal_2043916[p2_res7__204_comb] ^ p1_literal_2043918[p2_res7__202_comb] ^ p2_array_index_2045494_comb ^ p2_res7__198_comb ^ p1_literal_2043923[p2_res7__196_comb] ^ p2_res7__194_comb ^ p2_array_index_2045448_comb ^ p2_array_index_2045421_comb ^ p2_array_index_2045392_comb ^ p2_array_index_2045360_comb ^ p1_literal_2043912[p2_array_index_2045345_comb] ^ p1_literal_2043910[p2_array_index_2045346_comb] ^ p2_array_index_2045347_comb;
  assign p2_array_index_2045504_comb = p1_literal_2043920[p2_res7__202_comb];
  assign p2_res7__214_comb = p1_literal_2043910[p2_res7__212_comb] ^ p1_literal_2043912[p2_res7__210_comb] ^ p1_literal_2043914[p2_res7__208_comb] ^ p1_literal_2043916[p2_res7__206_comb] ^ p1_literal_2043918[p2_res7__204_comb] ^ p2_array_index_2045504_comb ^ p2_res7__200_comb ^ p1_literal_2043923[p2_res7__198_comb] ^ p2_res7__196_comb ^ p2_array_index_2045460_comb ^ p2_array_index_2045434_comb ^ p2_array_index_2045406_comb ^ p2_array_index_2045377_comb ^ p1_literal_2043912[p2_array_index_2045344_comb] ^ p1_literal_2043910[p2_array_index_2045345_comb] ^ p2_array_index_2045346_comb;
  assign p2_res7__216_comb = p1_literal_2043910[p2_res7__214_comb] ^ p1_literal_2043912[p2_res7__212_comb] ^ p1_literal_2043914[p2_res7__210_comb] ^ p1_literal_2043916[p2_res7__208_comb] ^ p1_literal_2043918[p2_res7__206_comb] ^ p1_literal_2043920[p2_res7__204_comb] ^ p2_res7__202_comb ^ p1_literal_2043923[p2_res7__200_comb] ^ p2_res7__198_comb ^ p2_array_index_2045472_comb ^ p2_array_index_2045447_comb ^ p2_array_index_2045420_comb ^ p2_array_index_2045391_comb ^ p2_array_index_2045359_comb ^ p1_literal_2043910[p2_array_index_2045344_comb] ^ p2_array_index_2045345_comb;
  assign p2_res7__218_comb = p1_literal_2043910[p2_res7__216_comb] ^ p1_literal_2043912[p2_res7__214_comb] ^ p1_literal_2043914[p2_res7__212_comb] ^ p1_literal_2043916[p2_res7__210_comb] ^ p1_literal_2043918[p2_res7__208_comb] ^ p1_literal_2043920[p2_res7__206_comb] ^ p2_res7__204_comb ^ p1_literal_2043923[p2_res7__202_comb] ^ p2_res7__200_comb ^ p2_array_index_2045483_comb ^ p2_array_index_2045459_comb ^ p2_array_index_2045433_comb ^ p2_array_index_2045405_comb ^ p2_array_index_2045376_comb ^ p1_literal_2043910[p2_array_index_2045343_comb] ^ p2_array_index_2045344_comb;
  assign p2_res7__220_comb = p1_literal_2043910[p2_res7__218_comb] ^ p1_literal_2043912[p2_res7__216_comb] ^ p1_literal_2043914[p2_res7__214_comb] ^ p1_literal_2043916[p2_res7__212_comb] ^ p1_literal_2043918[p2_res7__210_comb] ^ p1_literal_2043920[p2_res7__208_comb] ^ p2_res7__206_comb ^ p1_literal_2043923[p2_res7__204_comb] ^ p2_res7__202_comb ^ p2_array_index_2045494_comb ^ p2_array_index_2045471_comb ^ p2_array_index_2045446_comb ^ p2_array_index_2045419_comb ^ p2_array_index_2045390_comb ^ p2_array_index_2045358_comb ^ p2_array_index_2045343_comb;
  assign p2_res7__222_comb = p1_literal_2043910[p2_res7__220_comb] ^ p1_literal_2043912[p2_res7__218_comb] ^ p1_literal_2043914[p2_res7__216_comb] ^ p1_literal_2043916[p2_res7__214_comb] ^ p1_literal_2043918[p2_res7__212_comb] ^ p1_literal_2043920[p2_res7__210_comb] ^ p2_res7__208_comb ^ p1_literal_2043923[p2_res7__206_comb] ^ p2_res7__204_comb ^ p2_array_index_2045504_comb ^ p2_array_index_2045482_comb ^ p2_array_index_2045458_comb ^ p2_array_index_2045432_comb ^ p2_array_index_2045404_comb ^ p2_array_index_2045375_comb ^ p2_array_index_2045342_comb;
  assign p2_res__6_comb = {p2_res7__222_comb, p2_res7__220_comb, p2_res7__218_comb, p2_res7__216_comb, p2_res7__214_comb, p2_res7__212_comb, p2_res7__210_comb, p2_res7__208_comb, p2_res7__206_comb, p2_res7__204_comb, p2_res7__202_comb, p2_res7__200_comb, p2_res7__198_comb, p2_res7__196_comb, p2_res7__194_comb, p2_res7__192_comb};
  assign p2_k3_comb = p2_res__6_comb ^ p2_xor_2045108_comb;
  assign p2_addedKey__39_comb = p2_k3_comb ^ 128'hf659_3616_e605_5689_adfb_a180_27aa_2a08;
  assign p2_array_index_2045560_comb = p1_literal_2043896[p2_addedKey__39_comb[127:120]];
  assign p2_array_index_2045561_comb = p1_literal_2043896[p2_addedKey__39_comb[119:112]];
  assign p2_array_index_2045562_comb = p1_literal_2043896[p2_addedKey__39_comb[111:104]];
  assign p2_array_index_2045563_comb = p1_literal_2043896[p2_addedKey__39_comb[103:96]];
  assign p2_array_index_2045564_comb = p1_literal_2043896[p2_addedKey__39_comb[95:88]];
  assign p2_array_index_2045565_comb = p1_literal_2043896[p2_addedKey__39_comb[87:80]];
  assign p2_array_index_2045567_comb = p1_literal_2043896[p2_addedKey__39_comb[71:64]];
  assign p2_array_index_2045569_comb = p1_literal_2043896[p2_addedKey__39_comb[55:48]];
  assign p2_array_index_2045570_comb = p1_literal_2043896[p2_addedKey__39_comb[47:40]];
  assign p2_array_index_2045571_comb = p1_literal_2043896[p2_addedKey__39_comb[39:32]];
  assign p2_array_index_2045572_comb = p1_literal_2043896[p2_addedKey__39_comb[31:24]];
  assign p2_array_index_2045573_comb = p1_literal_2043896[p2_addedKey__39_comb[23:16]];
  assign p2_array_index_2045574_comb = p1_literal_2043896[p2_addedKey__39_comb[15:8]];
  assign p2_array_index_2045576_comb = p1_literal_2043910[p2_array_index_2045560_comb];
  assign p2_array_index_2045577_comb = p1_literal_2043912[p2_array_index_2045561_comb];
  assign p2_array_index_2045578_comb = p1_literal_2043914[p2_array_index_2045562_comb];
  assign p2_array_index_2045579_comb = p1_literal_2043916[p2_array_index_2045563_comb];
  assign p2_array_index_2045580_comb = p1_literal_2043918[p2_array_index_2045564_comb];
  assign p2_array_index_2045581_comb = p1_literal_2043920[p2_array_index_2045565_comb];
  assign p2_array_index_2045582_comb = p1_literal_2043896[p2_addedKey__39_comb[79:72]];
  assign p2_array_index_2045584_comb = p1_literal_2043896[p2_addedKey__39_comb[63:56]];
  assign p2_res7__224_comb = p2_array_index_2045576_comb ^ p2_array_index_2045577_comb ^ p2_array_index_2045578_comb ^ p2_array_index_2045579_comb ^ p2_array_index_2045580_comb ^ p2_array_index_2045581_comb ^ p2_array_index_2045582_comb ^ p1_literal_2043923[p2_array_index_2045567_comb] ^ p2_array_index_2045584_comb ^ p1_literal_2043920[p2_array_index_2045569_comb] ^ p1_literal_2043918[p2_array_index_2045570_comb] ^ p1_literal_2043916[p2_array_index_2045571_comb] ^ p1_literal_2043914[p2_array_index_2045572_comb] ^ p1_literal_2043912[p2_array_index_2045573_comb] ^ p1_literal_2043910[p2_array_index_2045574_comb] ^ p1_literal_2043896[p2_addedKey__39_comb[7:0]];
  assign p2_array_index_2045593_comb = p1_literal_2043910[p2_res7__224_comb];
  assign p2_array_index_2045594_comb = p1_literal_2043912[p2_array_index_2045560_comb];
  assign p2_array_index_2045595_comb = p1_literal_2043914[p2_array_index_2045561_comb];
  assign p2_array_index_2045596_comb = p1_literal_2043916[p2_array_index_2045562_comb];
  assign p2_array_index_2045597_comb = p1_literal_2043918[p2_array_index_2045563_comb];
  assign p2_array_index_2045598_comb = p1_literal_2043920[p2_array_index_2045564_comb];
  assign p2_res7__226_comb = p2_array_index_2045593_comb ^ p2_array_index_2045594_comb ^ p2_array_index_2045595_comb ^ p2_array_index_2045596_comb ^ p2_array_index_2045597_comb ^ p2_array_index_2045598_comb ^ p2_array_index_2045565_comb ^ p1_literal_2043923[p2_array_index_2045582_comb] ^ p2_array_index_2045567_comb ^ p1_literal_2043920[p2_array_index_2045584_comb] ^ p1_literal_2043918[p2_array_index_2045569_comb] ^ p1_literal_2043916[p2_array_index_2045570_comb] ^ p1_literal_2043914[p2_array_index_2045571_comb] ^ p1_literal_2043912[p2_array_index_2045572_comb] ^ p1_literal_2043910[p2_array_index_2045573_comb] ^ p2_array_index_2045574_comb;
  assign p2_array_index_2045608_comb = p1_literal_2043912[p2_res7__224_comb];
  assign p2_array_index_2045609_comb = p1_literal_2043914[p2_array_index_2045560_comb];
  assign p2_array_index_2045610_comb = p1_literal_2043916[p2_array_index_2045561_comb];
  assign p2_array_index_2045611_comb = p1_literal_2043918[p2_array_index_2045562_comb];
  assign p2_array_index_2045612_comb = p1_literal_2043920[p2_array_index_2045563_comb];
  assign p2_res7__228_comb = p1_literal_2043910[p2_res7__226_comb] ^ p2_array_index_2045608_comb ^ p2_array_index_2045609_comb ^ p2_array_index_2045610_comb ^ p2_array_index_2045611_comb ^ p2_array_index_2045612_comb ^ p2_array_index_2045564_comb ^ p1_literal_2043923[p2_array_index_2045565_comb] ^ p2_array_index_2045582_comb ^ p1_literal_2043920[p2_array_index_2045567_comb] ^ p1_literal_2043918[p2_array_index_2045584_comb] ^ p1_literal_2043916[p2_array_index_2045569_comb] ^ p1_literal_2043914[p2_array_index_2045570_comb] ^ p1_literal_2043912[p2_array_index_2045571_comb] ^ p1_literal_2043910[p2_array_index_2045572_comb] ^ p2_array_index_2045573_comb;
  assign p2_array_index_2045622_comb = p1_literal_2043912[p2_res7__226_comb];
  assign p2_array_index_2045623_comb = p1_literal_2043914[p2_res7__224_comb];
  assign p2_array_index_2045624_comb = p1_literal_2043916[p2_array_index_2045560_comb];
  assign p2_array_index_2045625_comb = p1_literal_2043918[p2_array_index_2045561_comb];
  assign p2_array_index_2045626_comb = p1_literal_2043920[p2_array_index_2045562_comb];
  assign p2_res7__230_comb = p1_literal_2043910[p2_res7__228_comb] ^ p2_array_index_2045622_comb ^ p2_array_index_2045623_comb ^ p2_array_index_2045624_comb ^ p2_array_index_2045625_comb ^ p2_array_index_2045626_comb ^ p2_array_index_2045563_comb ^ p1_literal_2043923[p2_array_index_2045564_comb] ^ p2_array_index_2045565_comb ^ p1_literal_2043920[p2_array_index_2045582_comb] ^ p1_literal_2043918[p2_array_index_2045567_comb] ^ p1_literal_2043916[p2_array_index_2045584_comb] ^ p1_literal_2043914[p2_array_index_2045569_comb] ^ p1_literal_2043912[p2_array_index_2045570_comb] ^ p1_literal_2043910[p2_array_index_2045571_comb] ^ p2_array_index_2045572_comb;
  assign p2_array_index_2045637_comb = p1_literal_2043914[p2_res7__226_comb];
  assign p2_array_index_2045638_comb = p1_literal_2043916[p2_res7__224_comb];
  assign p2_array_index_2045639_comb = p1_literal_2043918[p2_array_index_2045560_comb];
  assign p2_array_index_2045640_comb = p1_literal_2043920[p2_array_index_2045561_comb];
  assign p2_res7__232_comb = p1_literal_2043910[p2_res7__230_comb] ^ p1_literal_2043912[p2_res7__228_comb] ^ p2_array_index_2045637_comb ^ p2_array_index_2045638_comb ^ p2_array_index_2045639_comb ^ p2_array_index_2045640_comb ^ p2_array_index_2045562_comb ^ p1_literal_2043923[p2_array_index_2045563_comb] ^ p2_array_index_2045564_comb ^ p2_array_index_2045581_comb ^ p1_literal_2043918[p2_array_index_2045582_comb] ^ p1_literal_2043916[p2_array_index_2045567_comb] ^ p1_literal_2043914[p2_array_index_2045584_comb] ^ p1_literal_2043912[p2_array_index_2045569_comb] ^ p1_literal_2043910[p2_array_index_2045570_comb] ^ p2_array_index_2045571_comb;
  assign p2_array_index_2045650_comb = p1_literal_2043914[p2_res7__228_comb];
  assign p2_array_index_2045651_comb = p1_literal_2043916[p2_res7__226_comb];
  assign p2_array_index_2045652_comb = p1_literal_2043918[p2_res7__224_comb];
  assign p2_array_index_2045653_comb = p1_literal_2043920[p2_array_index_2045560_comb];
  assign p2_res7__234_comb = p1_literal_2043910[p2_res7__232_comb] ^ p1_literal_2043912[p2_res7__230_comb] ^ p2_array_index_2045650_comb ^ p2_array_index_2045651_comb ^ p2_array_index_2045652_comb ^ p2_array_index_2045653_comb ^ p2_array_index_2045561_comb ^ p1_literal_2043923[p2_array_index_2045562_comb] ^ p2_array_index_2045563_comb ^ p2_array_index_2045598_comb ^ p1_literal_2043918[p2_array_index_2045565_comb] ^ p1_literal_2043916[p2_array_index_2045582_comb] ^ p1_literal_2043914[p2_array_index_2045567_comb] ^ p1_literal_2043912[p2_array_index_2045584_comb] ^ p1_literal_2043910[p2_array_index_2045569_comb] ^ p2_array_index_2045570_comb;
  assign p2_array_index_2045664_comb = p1_literal_2043916[p2_res7__228_comb];
  assign p2_array_index_2045665_comb = p1_literal_2043918[p2_res7__226_comb];
  assign p2_array_index_2045666_comb = p1_literal_2043920[p2_res7__224_comb];
  assign p2_res7__236_comb = p1_literal_2043910[p2_res7__234_comb] ^ p1_literal_2043912[p2_res7__232_comb] ^ p1_literal_2043914[p2_res7__230_comb] ^ p2_array_index_2045664_comb ^ p2_array_index_2045665_comb ^ p2_array_index_2045666_comb ^ p2_array_index_2045560_comb ^ p1_literal_2043923[p2_array_index_2045561_comb] ^ p2_array_index_2045562_comb ^ p2_array_index_2045612_comb ^ p2_array_index_2045580_comb ^ p1_literal_2043916[p2_array_index_2045565_comb] ^ p1_literal_2043914[p2_array_index_2045582_comb] ^ p1_literal_2043912[p2_array_index_2045567_comb] ^ p1_literal_2043910[p2_array_index_2045584_comb] ^ p2_array_index_2045569_comb;
  assign p2_array_index_2045676_comb = p1_literal_2043916[p2_res7__230_comb];
  assign p2_array_index_2045677_comb = p1_literal_2043918[p2_res7__228_comb];
  assign p2_array_index_2045678_comb = p1_literal_2043920[p2_res7__226_comb];
  assign p2_res7__238_comb = p1_literal_2043910[p2_res7__236_comb] ^ p1_literal_2043912[p2_res7__234_comb] ^ p1_literal_2043914[p2_res7__232_comb] ^ p2_array_index_2045676_comb ^ p2_array_index_2045677_comb ^ p2_array_index_2045678_comb ^ p2_res7__224_comb ^ p1_literal_2043923[p2_array_index_2045560_comb] ^ p2_array_index_2045561_comb ^ p2_array_index_2045626_comb ^ p2_array_index_2045597_comb ^ p1_literal_2043916[p2_array_index_2045564_comb] ^ p1_literal_2043914[p2_array_index_2045565_comb] ^ p1_literal_2043912[p2_array_index_2045582_comb] ^ p1_literal_2043910[p2_array_index_2045567_comb] ^ p2_array_index_2045584_comb;
  assign p2_array_index_2045689_comb = p1_literal_2043918[p2_res7__230_comb];
  assign p2_array_index_2045690_comb = p1_literal_2043920[p2_res7__228_comb];
  assign p2_res7__240_comb = p1_literal_2043910[p2_res7__238_comb] ^ p1_literal_2043912[p2_res7__236_comb] ^ p1_literal_2043914[p2_res7__234_comb] ^ p1_literal_2043916[p2_res7__232_comb] ^ p2_array_index_2045689_comb ^ p2_array_index_2045690_comb ^ p2_res7__226_comb ^ p1_literal_2043923[p2_res7__224_comb] ^ p2_array_index_2045560_comb ^ p2_array_index_2045640_comb ^ p2_array_index_2045611_comb ^ p2_array_index_2045579_comb ^ p1_literal_2043914[p2_array_index_2045564_comb] ^ p1_literal_2043912[p2_array_index_2045565_comb] ^ p1_literal_2043910[p2_array_index_2045582_comb] ^ p2_array_index_2045567_comb;
  assign p2_array_index_2045700_comb = p1_literal_2043918[p2_res7__232_comb];
  assign p2_array_index_2045701_comb = p1_literal_2043920[p2_res7__230_comb];
  assign p2_res7__242_comb = p1_literal_2043910[p2_res7__240_comb] ^ p1_literal_2043912[p2_res7__238_comb] ^ p1_literal_2043914[p2_res7__236_comb] ^ p1_literal_2043916[p2_res7__234_comb] ^ p2_array_index_2045700_comb ^ p2_array_index_2045701_comb ^ p2_res7__228_comb ^ p1_literal_2043923[p2_res7__226_comb] ^ p2_res7__224_comb ^ p2_array_index_2045653_comb ^ p2_array_index_2045625_comb ^ p2_array_index_2045596_comb ^ p1_literal_2043914[p2_array_index_2045563_comb] ^ p1_literal_2043912[p2_array_index_2045564_comb] ^ p1_literal_2043910[p2_array_index_2045565_comb] ^ p2_array_index_2045582_comb;
  assign p2_array_index_2045712_comb = p1_literal_2043920[p2_res7__232_comb];
  assign p2_res7__244_comb = p1_literal_2043910[p2_res7__242_comb] ^ p1_literal_2043912[p2_res7__240_comb] ^ p1_literal_2043914[p2_res7__238_comb] ^ p1_literal_2043916[p2_res7__236_comb] ^ p1_literal_2043918[p2_res7__234_comb] ^ p2_array_index_2045712_comb ^ p2_res7__230_comb ^ p1_literal_2043923[p2_res7__228_comb] ^ p2_res7__226_comb ^ p2_array_index_2045666_comb ^ p2_array_index_2045639_comb ^ p2_array_index_2045610_comb ^ p2_array_index_2045578_comb ^ p1_literal_2043912[p2_array_index_2045563_comb] ^ p1_literal_2043910[p2_array_index_2045564_comb] ^ p2_array_index_2045565_comb;
  assign p2_array_index_2045722_comb = p1_literal_2043920[p2_res7__234_comb];
  assign p2_res7__246_comb = p1_literal_2043910[p2_res7__244_comb] ^ p1_literal_2043912[p2_res7__242_comb] ^ p1_literal_2043914[p2_res7__240_comb] ^ p1_literal_2043916[p2_res7__238_comb] ^ p1_literal_2043918[p2_res7__236_comb] ^ p2_array_index_2045722_comb ^ p2_res7__232_comb ^ p1_literal_2043923[p2_res7__230_comb] ^ p2_res7__228_comb ^ p2_array_index_2045678_comb ^ p2_array_index_2045652_comb ^ p2_array_index_2045624_comb ^ p2_array_index_2045595_comb ^ p1_literal_2043912[p2_array_index_2045562_comb] ^ p1_literal_2043910[p2_array_index_2045563_comb] ^ p2_array_index_2045564_comb;
  assign p2_res7__248_comb = p1_literal_2043910[p2_res7__246_comb] ^ p1_literal_2043912[p2_res7__244_comb] ^ p1_literal_2043914[p2_res7__242_comb] ^ p1_literal_2043916[p2_res7__240_comb] ^ p1_literal_2043918[p2_res7__238_comb] ^ p1_literal_2043920[p2_res7__236_comb] ^ p2_res7__234_comb ^ p1_literal_2043923[p2_res7__232_comb] ^ p2_res7__230_comb ^ p2_array_index_2045690_comb ^ p2_array_index_2045665_comb ^ p2_array_index_2045638_comb ^ p2_array_index_2045609_comb ^ p2_array_index_2045577_comb ^ p1_literal_2043910[p2_array_index_2045562_comb] ^ p2_array_index_2045563_comb;
  assign p2_res7__250_comb = p1_literal_2043910[p2_res7__248_comb] ^ p1_literal_2043912[p2_res7__246_comb] ^ p1_literal_2043914[p2_res7__244_comb] ^ p1_literal_2043916[p2_res7__242_comb] ^ p1_literal_2043918[p2_res7__240_comb] ^ p1_literal_2043920[p2_res7__238_comb] ^ p2_res7__236_comb ^ p1_literal_2043923[p2_res7__234_comb] ^ p2_res7__232_comb ^ p2_array_index_2045701_comb ^ p2_array_index_2045677_comb ^ p2_array_index_2045651_comb ^ p2_array_index_2045623_comb ^ p2_array_index_2045594_comb ^ p1_literal_2043910[p2_array_index_2045561_comb] ^ p2_array_index_2045562_comb;
  assign p2_res7__252_comb = p1_literal_2043910[p2_res7__250_comb] ^ p1_literal_2043912[p2_res7__248_comb] ^ p1_literal_2043914[p2_res7__246_comb] ^ p1_literal_2043916[p2_res7__244_comb] ^ p1_literal_2043918[p2_res7__242_comb] ^ p1_literal_2043920[p2_res7__240_comb] ^ p2_res7__238_comb ^ p1_literal_2043923[p2_res7__236_comb] ^ p2_res7__234_comb ^ p2_array_index_2045712_comb ^ p2_array_index_2045689_comb ^ p2_array_index_2045664_comb ^ p2_array_index_2045637_comb ^ p2_array_index_2045608_comb ^ p2_array_index_2045576_comb ^ p2_array_index_2045561_comb;
  assign p2_res7__254_comb = p1_literal_2043910[p2_res7__252_comb] ^ p1_literal_2043912[p2_res7__250_comb] ^ p1_literal_2043914[p2_res7__248_comb] ^ p1_literal_2043916[p2_res7__246_comb] ^ p1_literal_2043918[p2_res7__244_comb] ^ p1_literal_2043920[p2_res7__242_comb] ^ p2_res7__240_comb ^ p1_literal_2043923[p2_res7__238_comb] ^ p2_res7__236_comb ^ p2_array_index_2045722_comb ^ p2_array_index_2045700_comb ^ p2_array_index_2045676_comb ^ p2_array_index_2045650_comb ^ p2_array_index_2045622_comb ^ p2_array_index_2045593_comb ^ p2_array_index_2045560_comb;
  assign p2_res__7_comb = {p2_res7__254_comb, p2_res7__252_comb, p2_res7__250_comb, p2_res7__248_comb, p2_res7__246_comb, p2_res7__244_comb, p2_res7__242_comb, p2_res7__240_comb, p2_res7__238_comb, p2_res7__236_comb, p2_res7__234_comb, p2_res7__232_comb, p2_res7__230_comb, p2_res7__228_comb, p2_res7__226_comb, p2_res7__224_comb};
  assign p2_k2_comb = p2_res__7_comb ^ p2_xor_2045326_comb;
  assign p2_addedKey__40_comb = p2_k2_comb ^ 128'h98fb_4064_8a4d_2c31_f0dc_1c90_fa2e_be09;
  assign p2_array_index_2045778_comb = p1_literal_2043896[p2_addedKey__40_comb[127:120]];
  assign p2_array_index_2045779_comb = p1_literal_2043896[p2_addedKey__40_comb[119:112]];
  assign p2_array_index_2045780_comb = p1_literal_2043896[p2_addedKey__40_comb[111:104]];
  assign p2_array_index_2045781_comb = p1_literal_2043896[p2_addedKey__40_comb[103:96]];
  assign p2_array_index_2045782_comb = p1_literal_2043896[p2_addedKey__40_comb[95:88]];
  assign p2_array_index_2045783_comb = p1_literal_2043896[p2_addedKey__40_comb[87:80]];
  assign p2_array_index_2045785_comb = p1_literal_2043896[p2_addedKey__40_comb[71:64]];
  assign p2_array_index_2045787_comb = p1_literal_2043896[p2_addedKey__40_comb[55:48]];
  assign p2_array_index_2045788_comb = p1_literal_2043896[p2_addedKey__40_comb[47:40]];
  assign p2_array_index_2045789_comb = p1_literal_2043896[p2_addedKey__40_comb[39:32]];
  assign p2_array_index_2045790_comb = p1_literal_2043896[p2_addedKey__40_comb[31:24]];
  assign p2_array_index_2045791_comb = p1_literal_2043896[p2_addedKey__40_comb[23:16]];
  assign p2_array_index_2045792_comb = p1_literal_2043896[p2_addedKey__40_comb[15:8]];
  assign p2_array_index_2045794_comb = p1_literal_2043910[p2_array_index_2045778_comb];
  assign p2_array_index_2045795_comb = p1_literal_2043912[p2_array_index_2045779_comb];
  assign p2_array_index_2045796_comb = p1_literal_2043914[p2_array_index_2045780_comb];
  assign p2_array_index_2045797_comb = p1_literal_2043916[p2_array_index_2045781_comb];
  assign p2_array_index_2045798_comb = p1_literal_2043918[p2_array_index_2045782_comb];
  assign p2_array_index_2045799_comb = p1_literal_2043920[p2_array_index_2045783_comb];
  assign p2_array_index_2045800_comb = p1_literal_2043896[p2_addedKey__40_comb[79:72]];
  assign p2_array_index_2045802_comb = p1_literal_2043896[p2_addedKey__40_comb[63:56]];
  assign p2_res7__256_comb = p2_array_index_2045794_comb ^ p2_array_index_2045795_comb ^ p2_array_index_2045796_comb ^ p2_array_index_2045797_comb ^ p2_array_index_2045798_comb ^ p2_array_index_2045799_comb ^ p2_array_index_2045800_comb ^ p1_literal_2043923[p2_array_index_2045785_comb] ^ p2_array_index_2045802_comb ^ p1_literal_2043920[p2_array_index_2045787_comb] ^ p1_literal_2043918[p2_array_index_2045788_comb] ^ p1_literal_2043916[p2_array_index_2045789_comb] ^ p1_literal_2043914[p2_array_index_2045790_comb] ^ p1_literal_2043912[p2_array_index_2045791_comb] ^ p1_literal_2043910[p2_array_index_2045792_comb] ^ p1_literal_2043896[p2_addedKey__40_comb[7:0]];
  assign p2_array_index_2045811_comb = p1_literal_2043910[p2_res7__256_comb];
  assign p2_array_index_2045812_comb = p1_literal_2043912[p2_array_index_2045778_comb];
  assign p2_array_index_2045813_comb = p1_literal_2043914[p2_array_index_2045779_comb];
  assign p2_array_index_2045814_comb = p1_literal_2043916[p2_array_index_2045780_comb];
  assign p2_array_index_2045815_comb = p1_literal_2043918[p2_array_index_2045781_comb];
  assign p2_array_index_2045816_comb = p1_literal_2043920[p2_array_index_2045782_comb];
  assign p2_res7__258_comb = p2_array_index_2045811_comb ^ p2_array_index_2045812_comb ^ p2_array_index_2045813_comb ^ p2_array_index_2045814_comb ^ p2_array_index_2045815_comb ^ p2_array_index_2045816_comb ^ p2_array_index_2045783_comb ^ p1_literal_2043923[p2_array_index_2045800_comb] ^ p2_array_index_2045785_comb ^ p1_literal_2043920[p2_array_index_2045802_comb] ^ p1_literal_2043918[p2_array_index_2045787_comb] ^ p1_literal_2043916[p2_array_index_2045788_comb] ^ p1_literal_2043914[p2_array_index_2045789_comb] ^ p1_literal_2043912[p2_array_index_2045790_comb] ^ p1_literal_2043910[p2_array_index_2045791_comb] ^ p2_array_index_2045792_comb;
  assign p2_array_index_2045826_comb = p1_literal_2043912[p2_res7__256_comb];
  assign p2_array_index_2045827_comb = p1_literal_2043914[p2_array_index_2045778_comb];
  assign p2_array_index_2045828_comb = p1_literal_2043916[p2_array_index_2045779_comb];
  assign p2_array_index_2045829_comb = p1_literal_2043918[p2_array_index_2045780_comb];
  assign p2_array_index_2045830_comb = p1_literal_2043920[p2_array_index_2045781_comb];
  assign p2_res7__260_comb = p1_literal_2043910[p2_res7__258_comb] ^ p2_array_index_2045826_comb ^ p2_array_index_2045827_comb ^ p2_array_index_2045828_comb ^ p2_array_index_2045829_comb ^ p2_array_index_2045830_comb ^ p2_array_index_2045782_comb ^ p1_literal_2043923[p2_array_index_2045783_comb] ^ p2_array_index_2045800_comb ^ p1_literal_2043920[p2_array_index_2045785_comb] ^ p1_literal_2043918[p2_array_index_2045802_comb] ^ p1_literal_2043916[p2_array_index_2045787_comb] ^ p1_literal_2043914[p2_array_index_2045788_comb] ^ p1_literal_2043912[p2_array_index_2045789_comb] ^ p1_literal_2043910[p2_array_index_2045790_comb] ^ p2_array_index_2045791_comb;
  assign p2_array_index_2045840_comb = p1_literal_2043912[p2_res7__258_comb];
  assign p2_array_index_2045841_comb = p1_literal_2043914[p2_res7__256_comb];
  assign p2_array_index_2045842_comb = p1_literal_2043916[p2_array_index_2045778_comb];
  assign p2_array_index_2045843_comb = p1_literal_2043918[p2_array_index_2045779_comb];
  assign p2_array_index_2045844_comb = p1_literal_2043920[p2_array_index_2045780_comb];
  assign p2_res7__262_comb = p1_literal_2043910[p2_res7__260_comb] ^ p2_array_index_2045840_comb ^ p2_array_index_2045841_comb ^ p2_array_index_2045842_comb ^ p2_array_index_2045843_comb ^ p2_array_index_2045844_comb ^ p2_array_index_2045781_comb ^ p1_literal_2043923[p2_array_index_2045782_comb] ^ p2_array_index_2045783_comb ^ p1_literal_2043920[p2_array_index_2045800_comb] ^ p1_literal_2043918[p2_array_index_2045785_comb] ^ p1_literal_2043916[p2_array_index_2045802_comb] ^ p1_literal_2043914[p2_array_index_2045787_comb] ^ p1_literal_2043912[p2_array_index_2045788_comb] ^ p1_literal_2043910[p2_array_index_2045789_comb] ^ p2_array_index_2045790_comb;
  assign p2_array_index_2045855_comb = p1_literal_2043914[p2_res7__258_comb];
  assign p2_array_index_2045856_comb = p1_literal_2043916[p2_res7__256_comb];
  assign p2_array_index_2045857_comb = p1_literal_2043918[p2_array_index_2045778_comb];
  assign p2_array_index_2045858_comb = p1_literal_2043920[p2_array_index_2045779_comb];
  assign p2_res7__264_comb = p1_literal_2043910[p2_res7__262_comb] ^ p1_literal_2043912[p2_res7__260_comb] ^ p2_array_index_2045855_comb ^ p2_array_index_2045856_comb ^ p2_array_index_2045857_comb ^ p2_array_index_2045858_comb ^ p2_array_index_2045780_comb ^ p1_literal_2043923[p2_array_index_2045781_comb] ^ p2_array_index_2045782_comb ^ p2_array_index_2045799_comb ^ p1_literal_2043918[p2_array_index_2045800_comb] ^ p1_literal_2043916[p2_array_index_2045785_comb] ^ p1_literal_2043914[p2_array_index_2045802_comb] ^ p1_literal_2043912[p2_array_index_2045787_comb] ^ p1_literal_2043910[p2_array_index_2045788_comb] ^ p2_array_index_2045789_comb;
  assign p2_array_index_2045868_comb = p1_literal_2043914[p2_res7__260_comb];
  assign p2_array_index_2045869_comb = p1_literal_2043916[p2_res7__258_comb];
  assign p2_array_index_2045870_comb = p1_literal_2043918[p2_res7__256_comb];
  assign p2_array_index_2045871_comb = p1_literal_2043920[p2_array_index_2045778_comb];
  assign p2_res7__266_comb = p1_literal_2043910[p2_res7__264_comb] ^ p1_literal_2043912[p2_res7__262_comb] ^ p2_array_index_2045868_comb ^ p2_array_index_2045869_comb ^ p2_array_index_2045870_comb ^ p2_array_index_2045871_comb ^ p2_array_index_2045779_comb ^ p1_literal_2043923[p2_array_index_2045780_comb] ^ p2_array_index_2045781_comb ^ p2_array_index_2045816_comb ^ p1_literal_2043918[p2_array_index_2045783_comb] ^ p1_literal_2043916[p2_array_index_2045800_comb] ^ p1_literal_2043914[p2_array_index_2045785_comb] ^ p1_literal_2043912[p2_array_index_2045802_comb] ^ p1_literal_2043910[p2_array_index_2045787_comb] ^ p2_array_index_2045788_comb;
  assign p2_array_index_2045882_comb = p1_literal_2043916[p2_res7__260_comb];
  assign p2_array_index_2045883_comb = p1_literal_2043918[p2_res7__258_comb];
  assign p2_array_index_2045884_comb = p1_literal_2043920[p2_res7__256_comb];
  assign p2_res7__268_comb = p1_literal_2043910[p2_res7__266_comb] ^ p1_literal_2043912[p2_res7__264_comb] ^ p1_literal_2043914[p2_res7__262_comb] ^ p2_array_index_2045882_comb ^ p2_array_index_2045883_comb ^ p2_array_index_2045884_comb ^ p2_array_index_2045778_comb ^ p1_literal_2043923[p2_array_index_2045779_comb] ^ p2_array_index_2045780_comb ^ p2_array_index_2045830_comb ^ p2_array_index_2045798_comb ^ p1_literal_2043916[p2_array_index_2045783_comb] ^ p1_literal_2043914[p2_array_index_2045800_comb] ^ p1_literal_2043912[p2_array_index_2045785_comb] ^ p1_literal_2043910[p2_array_index_2045802_comb] ^ p2_array_index_2045787_comb;
  assign p2_array_index_2045894_comb = p1_literal_2043916[p2_res7__262_comb];
  assign p2_array_index_2045895_comb = p1_literal_2043918[p2_res7__260_comb];
  assign p2_array_index_2045896_comb = p1_literal_2043920[p2_res7__258_comb];
  assign p2_res7__270_comb = p1_literal_2043910[p2_res7__268_comb] ^ p1_literal_2043912[p2_res7__266_comb] ^ p1_literal_2043914[p2_res7__264_comb] ^ p2_array_index_2045894_comb ^ p2_array_index_2045895_comb ^ p2_array_index_2045896_comb ^ p2_res7__256_comb ^ p1_literal_2043923[p2_array_index_2045778_comb] ^ p2_array_index_2045779_comb ^ p2_array_index_2045844_comb ^ p2_array_index_2045815_comb ^ p1_literal_2043916[p2_array_index_2045782_comb] ^ p1_literal_2043914[p2_array_index_2045783_comb] ^ p1_literal_2043912[p2_array_index_2045800_comb] ^ p1_literal_2043910[p2_array_index_2045785_comb] ^ p2_array_index_2045802_comb;
  assign p2_array_index_2045907_comb = p1_literal_2043918[p2_res7__262_comb];
  assign p2_array_index_2045908_comb = p1_literal_2043920[p2_res7__260_comb];
  assign p2_res7__272_comb = p1_literal_2043910[p2_res7__270_comb] ^ p1_literal_2043912[p2_res7__268_comb] ^ p1_literal_2043914[p2_res7__266_comb] ^ p1_literal_2043916[p2_res7__264_comb] ^ p2_array_index_2045907_comb ^ p2_array_index_2045908_comb ^ p2_res7__258_comb ^ p1_literal_2043923[p2_res7__256_comb] ^ p2_array_index_2045778_comb ^ p2_array_index_2045858_comb ^ p2_array_index_2045829_comb ^ p2_array_index_2045797_comb ^ p1_literal_2043914[p2_array_index_2045782_comb] ^ p1_literal_2043912[p2_array_index_2045783_comb] ^ p1_literal_2043910[p2_array_index_2045800_comb] ^ p2_array_index_2045785_comb;
  assign p2_array_index_2045918_comb = p1_literal_2043918[p2_res7__264_comb];
  assign p2_array_index_2045919_comb = p1_literal_2043920[p2_res7__262_comb];
  assign p2_res7__274_comb = p1_literal_2043910[p2_res7__272_comb] ^ p1_literal_2043912[p2_res7__270_comb] ^ p1_literal_2043914[p2_res7__268_comb] ^ p1_literal_2043916[p2_res7__266_comb] ^ p2_array_index_2045918_comb ^ p2_array_index_2045919_comb ^ p2_res7__260_comb ^ p1_literal_2043923[p2_res7__258_comb] ^ p2_res7__256_comb ^ p2_array_index_2045871_comb ^ p2_array_index_2045843_comb ^ p2_array_index_2045814_comb ^ p1_literal_2043914[p2_array_index_2045781_comb] ^ p1_literal_2043912[p2_array_index_2045782_comb] ^ p1_literal_2043910[p2_array_index_2045783_comb] ^ p2_array_index_2045800_comb;
  assign p2_array_index_2045930_comb = p1_literal_2043920[p2_res7__264_comb];
  assign p2_res7__276_comb = p1_literal_2043910[p2_res7__274_comb] ^ p1_literal_2043912[p2_res7__272_comb] ^ p1_literal_2043914[p2_res7__270_comb] ^ p1_literal_2043916[p2_res7__268_comb] ^ p1_literal_2043918[p2_res7__266_comb] ^ p2_array_index_2045930_comb ^ p2_res7__262_comb ^ p1_literal_2043923[p2_res7__260_comb] ^ p2_res7__258_comb ^ p2_array_index_2045884_comb ^ p2_array_index_2045857_comb ^ p2_array_index_2045828_comb ^ p2_array_index_2045796_comb ^ p1_literal_2043912[p2_array_index_2045781_comb] ^ p1_literal_2043910[p2_array_index_2045782_comb] ^ p2_array_index_2045783_comb;
  assign p2_array_index_2045940_comb = p1_literal_2043920[p2_res7__266_comb];
  assign p2_res7__278_comb = p1_literal_2043910[p2_res7__276_comb] ^ p1_literal_2043912[p2_res7__274_comb] ^ p1_literal_2043914[p2_res7__272_comb] ^ p1_literal_2043916[p2_res7__270_comb] ^ p1_literal_2043918[p2_res7__268_comb] ^ p2_array_index_2045940_comb ^ p2_res7__264_comb ^ p1_literal_2043923[p2_res7__262_comb] ^ p2_res7__260_comb ^ p2_array_index_2045896_comb ^ p2_array_index_2045870_comb ^ p2_array_index_2045842_comb ^ p2_array_index_2045813_comb ^ p1_literal_2043912[p2_array_index_2045780_comb] ^ p1_literal_2043910[p2_array_index_2045781_comb] ^ p2_array_index_2045782_comb;
  assign p2_res7__280_comb = p1_literal_2043910[p2_res7__278_comb] ^ p1_literal_2043912[p2_res7__276_comb] ^ p1_literal_2043914[p2_res7__274_comb] ^ p1_literal_2043916[p2_res7__272_comb] ^ p1_literal_2043918[p2_res7__270_comb] ^ p1_literal_2043920[p2_res7__268_comb] ^ p2_res7__266_comb ^ p1_literal_2043923[p2_res7__264_comb] ^ p2_res7__262_comb ^ p2_array_index_2045908_comb ^ p2_array_index_2045883_comb ^ p2_array_index_2045856_comb ^ p2_array_index_2045827_comb ^ p2_array_index_2045795_comb ^ p1_literal_2043910[p2_array_index_2045780_comb] ^ p2_array_index_2045781_comb;
  assign p2_res7__282_comb = p1_literal_2043910[p2_res7__280_comb] ^ p1_literal_2043912[p2_res7__278_comb] ^ p1_literal_2043914[p2_res7__276_comb] ^ p1_literal_2043916[p2_res7__274_comb] ^ p1_literal_2043918[p2_res7__272_comb] ^ p1_literal_2043920[p2_res7__270_comb] ^ p2_res7__268_comb ^ p1_literal_2043923[p2_res7__266_comb] ^ p2_res7__264_comb ^ p2_array_index_2045919_comb ^ p2_array_index_2045895_comb ^ p2_array_index_2045869_comb ^ p2_array_index_2045841_comb ^ p2_array_index_2045812_comb ^ p1_literal_2043910[p2_array_index_2045779_comb] ^ p2_array_index_2045780_comb;
  assign p2_array_index_2045963_comb = p1_literal_2043910[p2_res7__282_comb];
  assign p2_array_index_2045964_comb = p1_literal_2043912[p2_res7__280_comb];
  assign p2_array_index_2045965_comb = p1_literal_2043914[p2_res7__278_comb];
  assign p2_array_index_2045966_comb = p1_literal_2043916[p2_res7__276_comb];
  assign p2_array_index_2045967_comb = p1_literal_2043918[p2_res7__274_comb];
  assign p2_array_index_2045968_comb = p1_literal_2043920[p2_res7__272_comb];
  assign p2_array_index_2045969_comb = p1_literal_2043923[p2_res7__268_comb];

  // Registers for pipe stage 2:
  reg [127:0] p2_encoded;
  reg [127:0] p2_bit_slice_2043893;
  reg [127:0] p2_bit_slice_2044119;
  reg [127:0] p2_k3;
  reg [127:0] p2_k2;
  reg [7:0] p2_array_index_2045778;
  reg [7:0] p2_array_index_2045779;
  reg [7:0] p2_array_index_2045794;
  reg [7:0] p2_res7__256;
  reg [7:0] p2_array_index_2045811;
  reg [7:0] p2_res7__258;
  reg [7:0] p2_array_index_2045826;
  reg [7:0] p2_res7__260;
  reg [7:0] p2_array_index_2045840;
  reg [7:0] p2_res7__262;
  reg [7:0] p2_array_index_2045855;
  reg [7:0] p2_res7__264;
  reg [7:0] p2_array_index_2045868;
  reg [7:0] p2_res7__266;
  reg [7:0] p2_array_index_2045882;
  reg [7:0] p2_res7__268;
  reg [7:0] p2_array_index_2045894;
  reg [7:0] p2_res7__270;
  reg [7:0] p2_array_index_2045907;
  reg [7:0] p2_res7__272;
  reg [7:0] p2_array_index_2045918;
  reg [7:0] p2_res7__274;
  reg [7:0] p2_array_index_2045930;
  reg [7:0] p2_res7__276;
  reg [7:0] p2_array_index_2045940;
  reg [7:0] p2_res7__278;
  reg [7:0] p2_res7__280;
  reg [7:0] p2_res7__282;
  reg [7:0] p2_array_index_2045963;
  reg [7:0] p2_array_index_2045964;
  reg [7:0] p2_array_index_2045965;
  reg [7:0] p2_array_index_2045966;
  reg [7:0] p2_array_index_2045967;
  reg [7:0] p2_array_index_2045968;
  reg [7:0] p2_array_index_2045969;
  reg [7:0] p3_literal_2043896[256];
  reg [7:0] p3_literal_2043910[256];
  reg [7:0] p3_literal_2043912[256];
  reg [7:0] p3_literal_2043914[256];
  reg [7:0] p3_literal_2043916[256];
  reg [7:0] p3_literal_2043918[256];
  reg [7:0] p3_literal_2043920[256];
  reg [7:0] p3_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p2_encoded <= p1_encoded;
    p2_bit_slice_2043893 <= p1_bit_slice_2043893;
    p2_bit_slice_2044119 <= p1_bit_slice_2044119;
    p2_k3 <= p2_k3_comb;
    p2_k2 <= p2_k2_comb;
    p2_array_index_2045778 <= p2_array_index_2045778_comb;
    p2_array_index_2045779 <= p2_array_index_2045779_comb;
    p2_array_index_2045794 <= p2_array_index_2045794_comb;
    p2_res7__256 <= p2_res7__256_comb;
    p2_array_index_2045811 <= p2_array_index_2045811_comb;
    p2_res7__258 <= p2_res7__258_comb;
    p2_array_index_2045826 <= p2_array_index_2045826_comb;
    p2_res7__260 <= p2_res7__260_comb;
    p2_array_index_2045840 <= p2_array_index_2045840_comb;
    p2_res7__262 <= p2_res7__262_comb;
    p2_array_index_2045855 <= p2_array_index_2045855_comb;
    p2_res7__264 <= p2_res7__264_comb;
    p2_array_index_2045868 <= p2_array_index_2045868_comb;
    p2_res7__266 <= p2_res7__266_comb;
    p2_array_index_2045882 <= p2_array_index_2045882_comb;
    p2_res7__268 <= p2_res7__268_comb;
    p2_array_index_2045894 <= p2_array_index_2045894_comb;
    p2_res7__270 <= p2_res7__270_comb;
    p2_array_index_2045907 <= p2_array_index_2045907_comb;
    p2_res7__272 <= p2_res7__272_comb;
    p2_array_index_2045918 <= p2_array_index_2045918_comb;
    p2_res7__274 <= p2_res7__274_comb;
    p2_array_index_2045930 <= p2_array_index_2045930_comb;
    p2_res7__276 <= p2_res7__276_comb;
    p2_array_index_2045940 <= p2_array_index_2045940_comb;
    p2_res7__278 <= p2_res7__278_comb;
    p2_res7__280 <= p2_res7__280_comb;
    p2_res7__282 <= p2_res7__282_comb;
    p2_array_index_2045963 <= p2_array_index_2045963_comb;
    p2_array_index_2045964 <= p2_array_index_2045964_comb;
    p2_array_index_2045965 <= p2_array_index_2045965_comb;
    p2_array_index_2045966 <= p2_array_index_2045966_comb;
    p2_array_index_2045967 <= p2_array_index_2045967_comb;
    p2_array_index_2045968 <= p2_array_index_2045968_comb;
    p2_array_index_2045969 <= p2_array_index_2045969_comb;
    p3_literal_2043896 <= p2_literal_2043896;
    p3_literal_2043910 <= p2_literal_2043910;
    p3_literal_2043912 <= p2_literal_2043912;
    p3_literal_2043914 <= p2_literal_2043914;
    p3_literal_2043916 <= p2_literal_2043916;
    p3_literal_2043918 <= p2_literal_2043918;
    p3_literal_2043920 <= p2_literal_2043920;
    p3_literal_2043923 <= p2_literal_2043923;
  end

  // ===== Pipe stage 3:
  wire [7:0] p3_res7__284_comb;
  wire [7:0] p3_res7__286_comb;
  wire [127:0] p3_res__8_comb;
  wire [127:0] p3_xor_2046076_comb;
  wire [127:0] p3_addedKey__41_comb;
  wire [7:0] p3_array_index_2046092_comb;
  wire [7:0] p3_array_index_2046093_comb;
  wire [7:0] p3_array_index_2046094_comb;
  wire [7:0] p3_array_index_2046095_comb;
  wire [7:0] p3_array_index_2046096_comb;
  wire [7:0] p3_array_index_2046097_comb;
  wire [7:0] p3_array_index_2046099_comb;
  wire [7:0] p3_array_index_2046101_comb;
  wire [7:0] p3_array_index_2046102_comb;
  wire [7:0] p3_array_index_2046103_comb;
  wire [7:0] p3_array_index_2046104_comb;
  wire [7:0] p3_array_index_2046105_comb;
  wire [7:0] p3_array_index_2046106_comb;
  wire [7:0] p3_array_index_2046108_comb;
  wire [7:0] p3_array_index_2046109_comb;
  wire [7:0] p3_array_index_2046110_comb;
  wire [7:0] p3_array_index_2046111_comb;
  wire [7:0] p3_array_index_2046112_comb;
  wire [7:0] p3_array_index_2046113_comb;
  wire [7:0] p3_array_index_2046114_comb;
  wire [7:0] p3_array_index_2046116_comb;
  wire [7:0] p3_res7__288_comb;
  wire [7:0] p3_array_index_2046125_comb;
  wire [7:0] p3_array_index_2046126_comb;
  wire [7:0] p3_array_index_2046127_comb;
  wire [7:0] p3_array_index_2046128_comb;
  wire [7:0] p3_array_index_2046129_comb;
  wire [7:0] p3_array_index_2046130_comb;
  wire [7:0] p3_res7__290_comb;
  wire [7:0] p3_array_index_2046140_comb;
  wire [7:0] p3_array_index_2046141_comb;
  wire [7:0] p3_array_index_2046142_comb;
  wire [7:0] p3_array_index_2046143_comb;
  wire [7:0] p3_array_index_2046144_comb;
  wire [7:0] p3_res7__292_comb;
  wire [7:0] p3_array_index_2046154_comb;
  wire [7:0] p3_array_index_2046155_comb;
  wire [7:0] p3_array_index_2046156_comb;
  wire [7:0] p3_array_index_2046157_comb;
  wire [7:0] p3_array_index_2046158_comb;
  wire [7:0] p3_res7__294_comb;
  wire [7:0] p3_array_index_2046169_comb;
  wire [7:0] p3_array_index_2046170_comb;
  wire [7:0] p3_array_index_2046171_comb;
  wire [7:0] p3_array_index_2046172_comb;
  wire [7:0] p3_res7__296_comb;
  wire [7:0] p3_array_index_2046182_comb;
  wire [7:0] p3_array_index_2046183_comb;
  wire [7:0] p3_array_index_2046184_comb;
  wire [7:0] p3_array_index_2046185_comb;
  wire [7:0] p3_res7__298_comb;
  wire [7:0] p3_array_index_2046196_comb;
  wire [7:0] p3_array_index_2046197_comb;
  wire [7:0] p3_array_index_2046198_comb;
  wire [7:0] p3_res7__300_comb;
  wire [7:0] p3_array_index_2046208_comb;
  wire [7:0] p3_array_index_2046209_comb;
  wire [7:0] p3_array_index_2046210_comb;
  wire [7:0] p3_res7__302_comb;
  wire [7:0] p3_array_index_2046221_comb;
  wire [7:0] p3_array_index_2046222_comb;
  wire [7:0] p3_res7__304_comb;
  wire [7:0] p3_array_index_2046232_comb;
  wire [7:0] p3_array_index_2046233_comb;
  wire [7:0] p3_res7__306_comb;
  wire [7:0] p3_array_index_2046244_comb;
  wire [7:0] p3_res7__308_comb;
  wire [7:0] p3_array_index_2046254_comb;
  wire [7:0] p3_res7__310_comb;
  wire [7:0] p3_res7__312_comb;
  wire [7:0] p3_res7__314_comb;
  wire [7:0] p3_res7__316_comb;
  wire [7:0] p3_res7__318_comb;
  wire [127:0] p3_res__9_comb;
  wire [127:0] p3_xor_2046294_comb;
  wire [127:0] p3_addedKey__42_comb;
  wire [7:0] p3_array_index_2046310_comb;
  wire [7:0] p3_array_index_2046311_comb;
  wire [7:0] p3_array_index_2046312_comb;
  wire [7:0] p3_array_index_2046313_comb;
  wire [7:0] p3_array_index_2046314_comb;
  wire [7:0] p3_array_index_2046315_comb;
  wire [7:0] p3_array_index_2046317_comb;
  wire [7:0] p3_array_index_2046319_comb;
  wire [7:0] p3_array_index_2046320_comb;
  wire [7:0] p3_array_index_2046321_comb;
  wire [7:0] p3_array_index_2046322_comb;
  wire [7:0] p3_array_index_2046323_comb;
  wire [7:0] p3_array_index_2046324_comb;
  wire [7:0] p3_array_index_2046326_comb;
  wire [7:0] p3_array_index_2046327_comb;
  wire [7:0] p3_array_index_2046328_comb;
  wire [7:0] p3_array_index_2046329_comb;
  wire [7:0] p3_array_index_2046330_comb;
  wire [7:0] p3_array_index_2046331_comb;
  wire [7:0] p3_array_index_2046332_comb;
  wire [7:0] p3_array_index_2046334_comb;
  wire [7:0] p3_res7__320_comb;
  wire [7:0] p3_array_index_2046343_comb;
  wire [7:0] p3_array_index_2046344_comb;
  wire [7:0] p3_array_index_2046345_comb;
  wire [7:0] p3_array_index_2046346_comb;
  wire [7:0] p3_array_index_2046347_comb;
  wire [7:0] p3_array_index_2046348_comb;
  wire [7:0] p3_res7__322_comb;
  wire [7:0] p3_array_index_2046358_comb;
  wire [7:0] p3_array_index_2046359_comb;
  wire [7:0] p3_array_index_2046360_comb;
  wire [7:0] p3_array_index_2046361_comb;
  wire [7:0] p3_array_index_2046362_comb;
  wire [7:0] p3_res7__324_comb;
  wire [7:0] p3_array_index_2046372_comb;
  wire [7:0] p3_array_index_2046373_comb;
  wire [7:0] p3_array_index_2046374_comb;
  wire [7:0] p3_array_index_2046375_comb;
  wire [7:0] p3_array_index_2046376_comb;
  wire [7:0] p3_res7__326_comb;
  wire [7:0] p3_array_index_2046387_comb;
  wire [7:0] p3_array_index_2046388_comb;
  wire [7:0] p3_array_index_2046389_comb;
  wire [7:0] p3_array_index_2046390_comb;
  wire [7:0] p3_res7__328_comb;
  wire [7:0] p3_array_index_2046400_comb;
  wire [7:0] p3_array_index_2046401_comb;
  wire [7:0] p3_array_index_2046402_comb;
  wire [7:0] p3_array_index_2046403_comb;
  wire [7:0] p3_res7__330_comb;
  wire [7:0] p3_array_index_2046414_comb;
  wire [7:0] p3_array_index_2046415_comb;
  wire [7:0] p3_array_index_2046416_comb;
  wire [7:0] p3_res7__332_comb;
  wire [7:0] p3_array_index_2046426_comb;
  wire [7:0] p3_array_index_2046427_comb;
  wire [7:0] p3_array_index_2046428_comb;
  wire [7:0] p3_res7__334_comb;
  wire [7:0] p3_array_index_2046439_comb;
  wire [7:0] p3_array_index_2046440_comb;
  wire [7:0] p3_res7__336_comb;
  wire [7:0] p3_array_index_2046450_comb;
  wire [7:0] p3_array_index_2046451_comb;
  wire [7:0] p3_res7__338_comb;
  wire [7:0] p3_array_index_2046462_comb;
  wire [7:0] p3_res7__340_comb;
  wire [7:0] p3_array_index_2046472_comb;
  wire [7:0] p3_res7__342_comb;
  wire [7:0] p3_res7__344_comb;
  wire [7:0] p3_res7__346_comb;
  wire [7:0] p3_res7__348_comb;
  wire [7:0] p3_res7__350_comb;
  wire [127:0] p3_res__10_comb;
  wire [127:0] p3_xor_2046512_comb;
  wire [127:0] p3_addedKey__43_comb;
  wire [7:0] p3_array_index_2046528_comb;
  wire [7:0] p3_array_index_2046529_comb;
  wire [7:0] p3_array_index_2046530_comb;
  wire [7:0] p3_array_index_2046531_comb;
  wire [7:0] p3_array_index_2046532_comb;
  wire [7:0] p3_array_index_2046533_comb;
  wire [7:0] p3_array_index_2046535_comb;
  wire [7:0] p3_array_index_2046537_comb;
  wire [7:0] p3_array_index_2046538_comb;
  wire [7:0] p3_array_index_2046539_comb;
  wire [7:0] p3_array_index_2046540_comb;
  wire [7:0] p3_array_index_2046541_comb;
  wire [7:0] p3_array_index_2046542_comb;
  wire [7:0] p3_array_index_2046544_comb;
  wire [7:0] p3_array_index_2046545_comb;
  wire [7:0] p3_array_index_2046546_comb;
  wire [7:0] p3_array_index_2046547_comb;
  wire [7:0] p3_array_index_2046548_comb;
  wire [7:0] p3_array_index_2046549_comb;
  wire [7:0] p3_array_index_2046550_comb;
  wire [7:0] p3_array_index_2046552_comb;
  wire [7:0] p3_res7__352_comb;
  wire [7:0] p3_array_index_2046561_comb;
  wire [7:0] p3_array_index_2046562_comb;
  wire [7:0] p3_array_index_2046563_comb;
  wire [7:0] p3_array_index_2046564_comb;
  wire [7:0] p3_array_index_2046565_comb;
  wire [7:0] p3_array_index_2046566_comb;
  wire [7:0] p3_res7__354_comb;
  wire [7:0] p3_array_index_2046576_comb;
  wire [7:0] p3_array_index_2046577_comb;
  wire [7:0] p3_array_index_2046578_comb;
  wire [7:0] p3_array_index_2046579_comb;
  wire [7:0] p3_array_index_2046580_comb;
  wire [7:0] p3_res7__356_comb;
  wire [7:0] p3_array_index_2046590_comb;
  wire [7:0] p3_array_index_2046591_comb;
  wire [7:0] p3_array_index_2046592_comb;
  wire [7:0] p3_array_index_2046593_comb;
  wire [7:0] p3_array_index_2046594_comb;
  wire [7:0] p3_res7__358_comb;
  wire [7:0] p3_array_index_2046605_comb;
  wire [7:0] p3_array_index_2046606_comb;
  wire [7:0] p3_array_index_2046607_comb;
  wire [7:0] p3_array_index_2046608_comb;
  wire [7:0] p3_res7__360_comb;
  wire [7:0] p3_array_index_2046618_comb;
  wire [7:0] p3_array_index_2046619_comb;
  wire [7:0] p3_array_index_2046620_comb;
  wire [7:0] p3_array_index_2046621_comb;
  wire [7:0] p3_res7__362_comb;
  wire [7:0] p3_array_index_2046632_comb;
  wire [7:0] p3_array_index_2046633_comb;
  wire [7:0] p3_array_index_2046634_comb;
  wire [7:0] p3_res7__364_comb;
  wire [7:0] p3_array_index_2046644_comb;
  wire [7:0] p3_array_index_2046645_comb;
  wire [7:0] p3_array_index_2046646_comb;
  wire [7:0] p3_res7__366_comb;
  wire [7:0] p3_array_index_2046657_comb;
  wire [7:0] p3_array_index_2046658_comb;
  wire [7:0] p3_res7__368_comb;
  wire [7:0] p3_array_index_2046668_comb;
  wire [7:0] p3_array_index_2046669_comb;
  wire [7:0] p3_res7__370_comb;
  wire [7:0] p3_array_index_2046680_comb;
  wire [7:0] p3_res7__372_comb;
  wire [7:0] p3_array_index_2046690_comb;
  wire [7:0] p3_res7__374_comb;
  wire [7:0] p3_res7__376_comb;
  wire [7:0] p3_res7__378_comb;
  wire [7:0] p3_res7__380_comb;
  wire [7:0] p3_res7__382_comb;
  wire [127:0] p3_res__11_comb;
  wire [127:0] p3_xor_2046730_comb;
  wire [127:0] p3_addedKey__44_comb;
  wire [7:0] p3_array_index_2046746_comb;
  wire [7:0] p3_array_index_2046747_comb;
  wire [7:0] p3_array_index_2046748_comb;
  wire [7:0] p3_array_index_2046749_comb;
  wire [7:0] p3_array_index_2046750_comb;
  wire [7:0] p3_array_index_2046751_comb;
  wire [7:0] p3_array_index_2046753_comb;
  wire [7:0] p3_array_index_2046755_comb;
  wire [7:0] p3_array_index_2046756_comb;
  wire [7:0] p3_array_index_2046757_comb;
  wire [7:0] p3_array_index_2046758_comb;
  wire [7:0] p3_array_index_2046759_comb;
  wire [7:0] p3_array_index_2046760_comb;
  wire [7:0] p3_array_index_2046762_comb;
  wire [7:0] p3_array_index_2046763_comb;
  wire [7:0] p3_array_index_2046764_comb;
  wire [7:0] p3_array_index_2046765_comb;
  wire [7:0] p3_array_index_2046766_comb;
  wire [7:0] p3_array_index_2046767_comb;
  wire [7:0] p3_array_index_2046768_comb;
  wire [7:0] p3_array_index_2046770_comb;
  wire [7:0] p3_res7__384_comb;
  wire [7:0] p3_array_index_2046779_comb;
  wire [7:0] p3_array_index_2046780_comb;
  wire [7:0] p3_array_index_2046781_comb;
  wire [7:0] p3_array_index_2046782_comb;
  wire [7:0] p3_array_index_2046783_comb;
  wire [7:0] p3_array_index_2046784_comb;
  wire [7:0] p3_res7__386_comb;
  wire [7:0] p3_array_index_2046794_comb;
  wire [7:0] p3_array_index_2046795_comb;
  wire [7:0] p3_array_index_2046796_comb;
  wire [7:0] p3_array_index_2046797_comb;
  wire [7:0] p3_array_index_2046798_comb;
  wire [7:0] p3_res7__388_comb;
  wire [7:0] p3_array_index_2046808_comb;
  wire [7:0] p3_array_index_2046809_comb;
  wire [7:0] p3_array_index_2046810_comb;
  wire [7:0] p3_array_index_2046811_comb;
  wire [7:0] p3_array_index_2046812_comb;
  wire [7:0] p3_res7__390_comb;
  wire [7:0] p3_array_index_2046823_comb;
  wire [7:0] p3_array_index_2046824_comb;
  wire [7:0] p3_array_index_2046825_comb;
  wire [7:0] p3_array_index_2046826_comb;
  wire [7:0] p3_res7__392_comb;
  wire [7:0] p3_array_index_2046836_comb;
  wire [7:0] p3_array_index_2046837_comb;
  wire [7:0] p3_array_index_2046838_comb;
  wire [7:0] p3_array_index_2046839_comb;
  wire [7:0] p3_res7__394_comb;
  wire [7:0] p3_array_index_2046850_comb;
  wire [7:0] p3_array_index_2046851_comb;
  wire [7:0] p3_array_index_2046852_comb;
  wire [7:0] p3_res7__396_comb;
  wire [7:0] p3_array_index_2046862_comb;
  wire [7:0] p3_array_index_2046863_comb;
  wire [7:0] p3_array_index_2046864_comb;
  wire [7:0] p3_res7__398_comb;
  wire [7:0] p3_array_index_2046875_comb;
  wire [7:0] p3_array_index_2046876_comb;
  wire [7:0] p3_res7__400_comb;
  wire [7:0] p3_array_index_2046886_comb;
  wire [7:0] p3_array_index_2046887_comb;
  wire [7:0] p3_res7__402_comb;
  wire [7:0] p3_array_index_2046898_comb;
  wire [7:0] p3_res7__404_comb;
  wire [7:0] p3_array_index_2046908_comb;
  wire [7:0] p3_res7__406_comb;
  wire [7:0] p3_res7__408_comb;
  wire [7:0] p3_res7__410_comb;
  wire [7:0] p3_res7__412_comb;
  wire [7:0] p3_res7__414_comb;
  wire [127:0] p3_res__12_comb;
  wire [127:0] p3_xor_2046948_comb;
  wire [127:0] p3_addedKey__45_comb;
  wire [7:0] p3_array_index_2046964_comb;
  wire [7:0] p3_array_index_2046965_comb;
  wire [7:0] p3_array_index_2046966_comb;
  wire [7:0] p3_array_index_2046967_comb;
  wire [7:0] p3_array_index_2046968_comb;
  wire [7:0] p3_array_index_2046969_comb;
  wire [7:0] p3_array_index_2046971_comb;
  wire [7:0] p3_array_index_2046973_comb;
  wire [7:0] p3_array_index_2046974_comb;
  wire [7:0] p3_array_index_2046975_comb;
  wire [7:0] p3_array_index_2046976_comb;
  wire [7:0] p3_array_index_2046977_comb;
  wire [7:0] p3_array_index_2046978_comb;
  wire [7:0] p3_array_index_2046980_comb;
  wire [7:0] p3_array_index_2046981_comb;
  wire [7:0] p3_array_index_2046982_comb;
  wire [7:0] p3_array_index_2046983_comb;
  wire [7:0] p3_array_index_2046984_comb;
  wire [7:0] p3_array_index_2046985_comb;
  wire [7:0] p3_array_index_2046986_comb;
  wire [7:0] p3_array_index_2046988_comb;
  wire [7:0] p3_res7__416_comb;
  wire [7:0] p3_array_index_2046997_comb;
  wire [7:0] p3_array_index_2046998_comb;
  wire [7:0] p3_array_index_2046999_comb;
  wire [7:0] p3_array_index_2047000_comb;
  wire [7:0] p3_array_index_2047001_comb;
  wire [7:0] p3_array_index_2047002_comb;
  wire [7:0] p3_res7__418_comb;
  wire [7:0] p3_array_index_2047012_comb;
  wire [7:0] p3_array_index_2047013_comb;
  wire [7:0] p3_array_index_2047014_comb;
  wire [7:0] p3_array_index_2047015_comb;
  wire [7:0] p3_array_index_2047016_comb;
  wire [7:0] p3_res7__420_comb;
  wire [7:0] p3_array_index_2047026_comb;
  wire [7:0] p3_array_index_2047027_comb;
  wire [7:0] p3_array_index_2047028_comb;
  wire [7:0] p3_array_index_2047029_comb;
  wire [7:0] p3_array_index_2047030_comb;
  wire [7:0] p3_res7__422_comb;
  wire [7:0] p3_array_index_2047041_comb;
  wire [7:0] p3_array_index_2047042_comb;
  wire [7:0] p3_array_index_2047043_comb;
  wire [7:0] p3_array_index_2047044_comb;
  wire [7:0] p3_res7__424_comb;
  assign p3_res7__284_comb = p2_array_index_2045963 ^ p2_array_index_2045964 ^ p2_array_index_2045965 ^ p2_array_index_2045966 ^ p2_array_index_2045967 ^ p2_array_index_2045968 ^ p2_res7__270 ^ p2_array_index_2045969 ^ p2_res7__266 ^ p2_array_index_2045930 ^ p2_array_index_2045907 ^ p2_array_index_2045882 ^ p2_array_index_2045855 ^ p2_array_index_2045826 ^ p2_array_index_2045794 ^ p2_array_index_2045779;
  assign p3_res7__286_comb = p2_literal_2043910[p3_res7__284_comb] ^ p2_literal_2043912[p2_res7__282] ^ p2_literal_2043914[p2_res7__280] ^ p2_literal_2043916[p2_res7__278] ^ p2_literal_2043918[p2_res7__276] ^ p2_literal_2043920[p2_res7__274] ^ p2_res7__272 ^ p2_literal_2043923[p2_res7__270] ^ p2_res7__268 ^ p2_array_index_2045940 ^ p2_array_index_2045918 ^ p2_array_index_2045894 ^ p2_array_index_2045868 ^ p2_array_index_2045840 ^ p2_array_index_2045811 ^ p2_array_index_2045778;
  assign p3_res__8_comb = {p3_res7__286_comb, p3_res7__284_comb, p2_res7__282, p2_res7__280, p2_res7__278, p2_res7__276, p2_res7__274, p2_res7__272, p2_res7__270, p2_res7__268, p2_res7__266, p2_res7__264, p2_res7__262, p2_res7__260, p2_res7__258, p2_res7__256};
  assign p3_xor_2046076_comb = p3_res__8_comb ^ p2_k3;
  assign p3_addedKey__41_comb = p3_xor_2046076_comb ^ 128'h2ade_daf2_3e95_a23a_17b5_18a0_5e61_c10a;
  assign p3_array_index_2046092_comb = p2_literal_2043896[p3_addedKey__41_comb[127:120]];
  assign p3_array_index_2046093_comb = p2_literal_2043896[p3_addedKey__41_comb[119:112]];
  assign p3_array_index_2046094_comb = p2_literal_2043896[p3_addedKey__41_comb[111:104]];
  assign p3_array_index_2046095_comb = p2_literal_2043896[p3_addedKey__41_comb[103:96]];
  assign p3_array_index_2046096_comb = p2_literal_2043896[p3_addedKey__41_comb[95:88]];
  assign p3_array_index_2046097_comb = p2_literal_2043896[p3_addedKey__41_comb[87:80]];
  assign p3_array_index_2046099_comb = p2_literal_2043896[p3_addedKey__41_comb[71:64]];
  assign p3_array_index_2046101_comb = p2_literal_2043896[p3_addedKey__41_comb[55:48]];
  assign p3_array_index_2046102_comb = p2_literal_2043896[p3_addedKey__41_comb[47:40]];
  assign p3_array_index_2046103_comb = p2_literal_2043896[p3_addedKey__41_comb[39:32]];
  assign p3_array_index_2046104_comb = p2_literal_2043896[p3_addedKey__41_comb[31:24]];
  assign p3_array_index_2046105_comb = p2_literal_2043896[p3_addedKey__41_comb[23:16]];
  assign p3_array_index_2046106_comb = p2_literal_2043896[p3_addedKey__41_comb[15:8]];
  assign p3_array_index_2046108_comb = p2_literal_2043910[p3_array_index_2046092_comb];
  assign p3_array_index_2046109_comb = p2_literal_2043912[p3_array_index_2046093_comb];
  assign p3_array_index_2046110_comb = p2_literal_2043914[p3_array_index_2046094_comb];
  assign p3_array_index_2046111_comb = p2_literal_2043916[p3_array_index_2046095_comb];
  assign p3_array_index_2046112_comb = p2_literal_2043918[p3_array_index_2046096_comb];
  assign p3_array_index_2046113_comb = p2_literal_2043920[p3_array_index_2046097_comb];
  assign p3_array_index_2046114_comb = p2_literal_2043896[p3_addedKey__41_comb[79:72]];
  assign p3_array_index_2046116_comb = p2_literal_2043896[p3_addedKey__41_comb[63:56]];
  assign p3_res7__288_comb = p3_array_index_2046108_comb ^ p3_array_index_2046109_comb ^ p3_array_index_2046110_comb ^ p3_array_index_2046111_comb ^ p3_array_index_2046112_comb ^ p3_array_index_2046113_comb ^ p3_array_index_2046114_comb ^ p2_literal_2043923[p3_array_index_2046099_comb] ^ p3_array_index_2046116_comb ^ p2_literal_2043920[p3_array_index_2046101_comb] ^ p2_literal_2043918[p3_array_index_2046102_comb] ^ p2_literal_2043916[p3_array_index_2046103_comb] ^ p2_literal_2043914[p3_array_index_2046104_comb] ^ p2_literal_2043912[p3_array_index_2046105_comb] ^ p2_literal_2043910[p3_array_index_2046106_comb] ^ p2_literal_2043896[p3_addedKey__41_comb[7:0]];
  assign p3_array_index_2046125_comb = p2_literal_2043910[p3_res7__288_comb];
  assign p3_array_index_2046126_comb = p2_literal_2043912[p3_array_index_2046092_comb];
  assign p3_array_index_2046127_comb = p2_literal_2043914[p3_array_index_2046093_comb];
  assign p3_array_index_2046128_comb = p2_literal_2043916[p3_array_index_2046094_comb];
  assign p3_array_index_2046129_comb = p2_literal_2043918[p3_array_index_2046095_comb];
  assign p3_array_index_2046130_comb = p2_literal_2043920[p3_array_index_2046096_comb];
  assign p3_res7__290_comb = p3_array_index_2046125_comb ^ p3_array_index_2046126_comb ^ p3_array_index_2046127_comb ^ p3_array_index_2046128_comb ^ p3_array_index_2046129_comb ^ p3_array_index_2046130_comb ^ p3_array_index_2046097_comb ^ p2_literal_2043923[p3_array_index_2046114_comb] ^ p3_array_index_2046099_comb ^ p2_literal_2043920[p3_array_index_2046116_comb] ^ p2_literal_2043918[p3_array_index_2046101_comb] ^ p2_literal_2043916[p3_array_index_2046102_comb] ^ p2_literal_2043914[p3_array_index_2046103_comb] ^ p2_literal_2043912[p3_array_index_2046104_comb] ^ p2_literal_2043910[p3_array_index_2046105_comb] ^ p3_array_index_2046106_comb;
  assign p3_array_index_2046140_comb = p2_literal_2043912[p3_res7__288_comb];
  assign p3_array_index_2046141_comb = p2_literal_2043914[p3_array_index_2046092_comb];
  assign p3_array_index_2046142_comb = p2_literal_2043916[p3_array_index_2046093_comb];
  assign p3_array_index_2046143_comb = p2_literal_2043918[p3_array_index_2046094_comb];
  assign p3_array_index_2046144_comb = p2_literal_2043920[p3_array_index_2046095_comb];
  assign p3_res7__292_comb = p2_literal_2043910[p3_res7__290_comb] ^ p3_array_index_2046140_comb ^ p3_array_index_2046141_comb ^ p3_array_index_2046142_comb ^ p3_array_index_2046143_comb ^ p3_array_index_2046144_comb ^ p3_array_index_2046096_comb ^ p2_literal_2043923[p3_array_index_2046097_comb] ^ p3_array_index_2046114_comb ^ p2_literal_2043920[p3_array_index_2046099_comb] ^ p2_literal_2043918[p3_array_index_2046116_comb] ^ p2_literal_2043916[p3_array_index_2046101_comb] ^ p2_literal_2043914[p3_array_index_2046102_comb] ^ p2_literal_2043912[p3_array_index_2046103_comb] ^ p2_literal_2043910[p3_array_index_2046104_comb] ^ p3_array_index_2046105_comb;
  assign p3_array_index_2046154_comb = p2_literal_2043912[p3_res7__290_comb];
  assign p3_array_index_2046155_comb = p2_literal_2043914[p3_res7__288_comb];
  assign p3_array_index_2046156_comb = p2_literal_2043916[p3_array_index_2046092_comb];
  assign p3_array_index_2046157_comb = p2_literal_2043918[p3_array_index_2046093_comb];
  assign p3_array_index_2046158_comb = p2_literal_2043920[p3_array_index_2046094_comb];
  assign p3_res7__294_comb = p2_literal_2043910[p3_res7__292_comb] ^ p3_array_index_2046154_comb ^ p3_array_index_2046155_comb ^ p3_array_index_2046156_comb ^ p3_array_index_2046157_comb ^ p3_array_index_2046158_comb ^ p3_array_index_2046095_comb ^ p2_literal_2043923[p3_array_index_2046096_comb] ^ p3_array_index_2046097_comb ^ p2_literal_2043920[p3_array_index_2046114_comb] ^ p2_literal_2043918[p3_array_index_2046099_comb] ^ p2_literal_2043916[p3_array_index_2046116_comb] ^ p2_literal_2043914[p3_array_index_2046101_comb] ^ p2_literal_2043912[p3_array_index_2046102_comb] ^ p2_literal_2043910[p3_array_index_2046103_comb] ^ p3_array_index_2046104_comb;
  assign p3_array_index_2046169_comb = p2_literal_2043914[p3_res7__290_comb];
  assign p3_array_index_2046170_comb = p2_literal_2043916[p3_res7__288_comb];
  assign p3_array_index_2046171_comb = p2_literal_2043918[p3_array_index_2046092_comb];
  assign p3_array_index_2046172_comb = p2_literal_2043920[p3_array_index_2046093_comb];
  assign p3_res7__296_comb = p2_literal_2043910[p3_res7__294_comb] ^ p2_literal_2043912[p3_res7__292_comb] ^ p3_array_index_2046169_comb ^ p3_array_index_2046170_comb ^ p3_array_index_2046171_comb ^ p3_array_index_2046172_comb ^ p3_array_index_2046094_comb ^ p2_literal_2043923[p3_array_index_2046095_comb] ^ p3_array_index_2046096_comb ^ p3_array_index_2046113_comb ^ p2_literal_2043918[p3_array_index_2046114_comb] ^ p2_literal_2043916[p3_array_index_2046099_comb] ^ p2_literal_2043914[p3_array_index_2046116_comb] ^ p2_literal_2043912[p3_array_index_2046101_comb] ^ p2_literal_2043910[p3_array_index_2046102_comb] ^ p3_array_index_2046103_comb;
  assign p3_array_index_2046182_comb = p2_literal_2043914[p3_res7__292_comb];
  assign p3_array_index_2046183_comb = p2_literal_2043916[p3_res7__290_comb];
  assign p3_array_index_2046184_comb = p2_literal_2043918[p3_res7__288_comb];
  assign p3_array_index_2046185_comb = p2_literal_2043920[p3_array_index_2046092_comb];
  assign p3_res7__298_comb = p2_literal_2043910[p3_res7__296_comb] ^ p2_literal_2043912[p3_res7__294_comb] ^ p3_array_index_2046182_comb ^ p3_array_index_2046183_comb ^ p3_array_index_2046184_comb ^ p3_array_index_2046185_comb ^ p3_array_index_2046093_comb ^ p2_literal_2043923[p3_array_index_2046094_comb] ^ p3_array_index_2046095_comb ^ p3_array_index_2046130_comb ^ p2_literal_2043918[p3_array_index_2046097_comb] ^ p2_literal_2043916[p3_array_index_2046114_comb] ^ p2_literal_2043914[p3_array_index_2046099_comb] ^ p2_literal_2043912[p3_array_index_2046116_comb] ^ p2_literal_2043910[p3_array_index_2046101_comb] ^ p3_array_index_2046102_comb;
  assign p3_array_index_2046196_comb = p2_literal_2043916[p3_res7__292_comb];
  assign p3_array_index_2046197_comb = p2_literal_2043918[p3_res7__290_comb];
  assign p3_array_index_2046198_comb = p2_literal_2043920[p3_res7__288_comb];
  assign p3_res7__300_comb = p2_literal_2043910[p3_res7__298_comb] ^ p2_literal_2043912[p3_res7__296_comb] ^ p2_literal_2043914[p3_res7__294_comb] ^ p3_array_index_2046196_comb ^ p3_array_index_2046197_comb ^ p3_array_index_2046198_comb ^ p3_array_index_2046092_comb ^ p2_literal_2043923[p3_array_index_2046093_comb] ^ p3_array_index_2046094_comb ^ p3_array_index_2046144_comb ^ p3_array_index_2046112_comb ^ p2_literal_2043916[p3_array_index_2046097_comb] ^ p2_literal_2043914[p3_array_index_2046114_comb] ^ p2_literal_2043912[p3_array_index_2046099_comb] ^ p2_literal_2043910[p3_array_index_2046116_comb] ^ p3_array_index_2046101_comb;
  assign p3_array_index_2046208_comb = p2_literal_2043916[p3_res7__294_comb];
  assign p3_array_index_2046209_comb = p2_literal_2043918[p3_res7__292_comb];
  assign p3_array_index_2046210_comb = p2_literal_2043920[p3_res7__290_comb];
  assign p3_res7__302_comb = p2_literal_2043910[p3_res7__300_comb] ^ p2_literal_2043912[p3_res7__298_comb] ^ p2_literal_2043914[p3_res7__296_comb] ^ p3_array_index_2046208_comb ^ p3_array_index_2046209_comb ^ p3_array_index_2046210_comb ^ p3_res7__288_comb ^ p2_literal_2043923[p3_array_index_2046092_comb] ^ p3_array_index_2046093_comb ^ p3_array_index_2046158_comb ^ p3_array_index_2046129_comb ^ p2_literal_2043916[p3_array_index_2046096_comb] ^ p2_literal_2043914[p3_array_index_2046097_comb] ^ p2_literal_2043912[p3_array_index_2046114_comb] ^ p2_literal_2043910[p3_array_index_2046099_comb] ^ p3_array_index_2046116_comb;
  assign p3_array_index_2046221_comb = p2_literal_2043918[p3_res7__294_comb];
  assign p3_array_index_2046222_comb = p2_literal_2043920[p3_res7__292_comb];
  assign p3_res7__304_comb = p2_literal_2043910[p3_res7__302_comb] ^ p2_literal_2043912[p3_res7__300_comb] ^ p2_literal_2043914[p3_res7__298_comb] ^ p2_literal_2043916[p3_res7__296_comb] ^ p3_array_index_2046221_comb ^ p3_array_index_2046222_comb ^ p3_res7__290_comb ^ p2_literal_2043923[p3_res7__288_comb] ^ p3_array_index_2046092_comb ^ p3_array_index_2046172_comb ^ p3_array_index_2046143_comb ^ p3_array_index_2046111_comb ^ p2_literal_2043914[p3_array_index_2046096_comb] ^ p2_literal_2043912[p3_array_index_2046097_comb] ^ p2_literal_2043910[p3_array_index_2046114_comb] ^ p3_array_index_2046099_comb;
  assign p3_array_index_2046232_comb = p2_literal_2043918[p3_res7__296_comb];
  assign p3_array_index_2046233_comb = p2_literal_2043920[p3_res7__294_comb];
  assign p3_res7__306_comb = p2_literal_2043910[p3_res7__304_comb] ^ p2_literal_2043912[p3_res7__302_comb] ^ p2_literal_2043914[p3_res7__300_comb] ^ p2_literal_2043916[p3_res7__298_comb] ^ p3_array_index_2046232_comb ^ p3_array_index_2046233_comb ^ p3_res7__292_comb ^ p2_literal_2043923[p3_res7__290_comb] ^ p3_res7__288_comb ^ p3_array_index_2046185_comb ^ p3_array_index_2046157_comb ^ p3_array_index_2046128_comb ^ p2_literal_2043914[p3_array_index_2046095_comb] ^ p2_literal_2043912[p3_array_index_2046096_comb] ^ p2_literal_2043910[p3_array_index_2046097_comb] ^ p3_array_index_2046114_comb;
  assign p3_array_index_2046244_comb = p2_literal_2043920[p3_res7__296_comb];
  assign p3_res7__308_comb = p2_literal_2043910[p3_res7__306_comb] ^ p2_literal_2043912[p3_res7__304_comb] ^ p2_literal_2043914[p3_res7__302_comb] ^ p2_literal_2043916[p3_res7__300_comb] ^ p2_literal_2043918[p3_res7__298_comb] ^ p3_array_index_2046244_comb ^ p3_res7__294_comb ^ p2_literal_2043923[p3_res7__292_comb] ^ p3_res7__290_comb ^ p3_array_index_2046198_comb ^ p3_array_index_2046171_comb ^ p3_array_index_2046142_comb ^ p3_array_index_2046110_comb ^ p2_literal_2043912[p3_array_index_2046095_comb] ^ p2_literal_2043910[p3_array_index_2046096_comb] ^ p3_array_index_2046097_comb;
  assign p3_array_index_2046254_comb = p2_literal_2043920[p3_res7__298_comb];
  assign p3_res7__310_comb = p2_literal_2043910[p3_res7__308_comb] ^ p2_literal_2043912[p3_res7__306_comb] ^ p2_literal_2043914[p3_res7__304_comb] ^ p2_literal_2043916[p3_res7__302_comb] ^ p2_literal_2043918[p3_res7__300_comb] ^ p3_array_index_2046254_comb ^ p3_res7__296_comb ^ p2_literal_2043923[p3_res7__294_comb] ^ p3_res7__292_comb ^ p3_array_index_2046210_comb ^ p3_array_index_2046184_comb ^ p3_array_index_2046156_comb ^ p3_array_index_2046127_comb ^ p2_literal_2043912[p3_array_index_2046094_comb] ^ p2_literal_2043910[p3_array_index_2046095_comb] ^ p3_array_index_2046096_comb;
  assign p3_res7__312_comb = p2_literal_2043910[p3_res7__310_comb] ^ p2_literal_2043912[p3_res7__308_comb] ^ p2_literal_2043914[p3_res7__306_comb] ^ p2_literal_2043916[p3_res7__304_comb] ^ p2_literal_2043918[p3_res7__302_comb] ^ p2_literal_2043920[p3_res7__300_comb] ^ p3_res7__298_comb ^ p2_literal_2043923[p3_res7__296_comb] ^ p3_res7__294_comb ^ p3_array_index_2046222_comb ^ p3_array_index_2046197_comb ^ p3_array_index_2046170_comb ^ p3_array_index_2046141_comb ^ p3_array_index_2046109_comb ^ p2_literal_2043910[p3_array_index_2046094_comb] ^ p3_array_index_2046095_comb;
  assign p3_res7__314_comb = p2_literal_2043910[p3_res7__312_comb] ^ p2_literal_2043912[p3_res7__310_comb] ^ p2_literal_2043914[p3_res7__308_comb] ^ p2_literal_2043916[p3_res7__306_comb] ^ p2_literal_2043918[p3_res7__304_comb] ^ p2_literal_2043920[p3_res7__302_comb] ^ p3_res7__300_comb ^ p2_literal_2043923[p3_res7__298_comb] ^ p3_res7__296_comb ^ p3_array_index_2046233_comb ^ p3_array_index_2046209_comb ^ p3_array_index_2046183_comb ^ p3_array_index_2046155_comb ^ p3_array_index_2046126_comb ^ p2_literal_2043910[p3_array_index_2046093_comb] ^ p3_array_index_2046094_comb;
  assign p3_res7__316_comb = p2_literal_2043910[p3_res7__314_comb] ^ p2_literal_2043912[p3_res7__312_comb] ^ p2_literal_2043914[p3_res7__310_comb] ^ p2_literal_2043916[p3_res7__308_comb] ^ p2_literal_2043918[p3_res7__306_comb] ^ p2_literal_2043920[p3_res7__304_comb] ^ p3_res7__302_comb ^ p2_literal_2043923[p3_res7__300_comb] ^ p3_res7__298_comb ^ p3_array_index_2046244_comb ^ p3_array_index_2046221_comb ^ p3_array_index_2046196_comb ^ p3_array_index_2046169_comb ^ p3_array_index_2046140_comb ^ p3_array_index_2046108_comb ^ p3_array_index_2046093_comb;
  assign p3_res7__318_comb = p2_literal_2043910[p3_res7__316_comb] ^ p2_literal_2043912[p3_res7__314_comb] ^ p2_literal_2043914[p3_res7__312_comb] ^ p2_literal_2043916[p3_res7__310_comb] ^ p2_literal_2043918[p3_res7__308_comb] ^ p2_literal_2043920[p3_res7__306_comb] ^ p3_res7__304_comb ^ p2_literal_2043923[p3_res7__302_comb] ^ p3_res7__300_comb ^ p3_array_index_2046254_comb ^ p3_array_index_2046232_comb ^ p3_array_index_2046208_comb ^ p3_array_index_2046182_comb ^ p3_array_index_2046154_comb ^ p3_array_index_2046125_comb ^ p3_array_index_2046092_comb;
  assign p3_res__9_comb = {p3_res7__318_comb, p3_res7__316_comb, p3_res7__314_comb, p3_res7__312_comb, p3_res7__310_comb, p3_res7__308_comb, p3_res7__306_comb, p3_res7__304_comb, p3_res7__302_comb, p3_res7__300_comb, p3_res7__298_comb, p3_res7__296_comb, p3_res7__294_comb, p3_res7__292_comb, p3_res7__290_comb, p3_res7__288_comb};
  assign p3_xor_2046294_comb = p3_res__9_comb ^ p2_k2;
  assign p3_addedKey__42_comb = p3_xor_2046294_comb ^ 128'h447c_ac80_52dd_d882_4a92_a5b0_83e5_550b;
  assign p3_array_index_2046310_comb = p2_literal_2043896[p3_addedKey__42_comb[127:120]];
  assign p3_array_index_2046311_comb = p2_literal_2043896[p3_addedKey__42_comb[119:112]];
  assign p3_array_index_2046312_comb = p2_literal_2043896[p3_addedKey__42_comb[111:104]];
  assign p3_array_index_2046313_comb = p2_literal_2043896[p3_addedKey__42_comb[103:96]];
  assign p3_array_index_2046314_comb = p2_literal_2043896[p3_addedKey__42_comb[95:88]];
  assign p3_array_index_2046315_comb = p2_literal_2043896[p3_addedKey__42_comb[87:80]];
  assign p3_array_index_2046317_comb = p2_literal_2043896[p3_addedKey__42_comb[71:64]];
  assign p3_array_index_2046319_comb = p2_literal_2043896[p3_addedKey__42_comb[55:48]];
  assign p3_array_index_2046320_comb = p2_literal_2043896[p3_addedKey__42_comb[47:40]];
  assign p3_array_index_2046321_comb = p2_literal_2043896[p3_addedKey__42_comb[39:32]];
  assign p3_array_index_2046322_comb = p2_literal_2043896[p3_addedKey__42_comb[31:24]];
  assign p3_array_index_2046323_comb = p2_literal_2043896[p3_addedKey__42_comb[23:16]];
  assign p3_array_index_2046324_comb = p2_literal_2043896[p3_addedKey__42_comb[15:8]];
  assign p3_array_index_2046326_comb = p2_literal_2043910[p3_array_index_2046310_comb];
  assign p3_array_index_2046327_comb = p2_literal_2043912[p3_array_index_2046311_comb];
  assign p3_array_index_2046328_comb = p2_literal_2043914[p3_array_index_2046312_comb];
  assign p3_array_index_2046329_comb = p2_literal_2043916[p3_array_index_2046313_comb];
  assign p3_array_index_2046330_comb = p2_literal_2043918[p3_array_index_2046314_comb];
  assign p3_array_index_2046331_comb = p2_literal_2043920[p3_array_index_2046315_comb];
  assign p3_array_index_2046332_comb = p2_literal_2043896[p3_addedKey__42_comb[79:72]];
  assign p3_array_index_2046334_comb = p2_literal_2043896[p3_addedKey__42_comb[63:56]];
  assign p3_res7__320_comb = p3_array_index_2046326_comb ^ p3_array_index_2046327_comb ^ p3_array_index_2046328_comb ^ p3_array_index_2046329_comb ^ p3_array_index_2046330_comb ^ p3_array_index_2046331_comb ^ p3_array_index_2046332_comb ^ p2_literal_2043923[p3_array_index_2046317_comb] ^ p3_array_index_2046334_comb ^ p2_literal_2043920[p3_array_index_2046319_comb] ^ p2_literal_2043918[p3_array_index_2046320_comb] ^ p2_literal_2043916[p3_array_index_2046321_comb] ^ p2_literal_2043914[p3_array_index_2046322_comb] ^ p2_literal_2043912[p3_array_index_2046323_comb] ^ p2_literal_2043910[p3_array_index_2046324_comb] ^ p2_literal_2043896[p3_addedKey__42_comb[7:0]];
  assign p3_array_index_2046343_comb = p2_literal_2043910[p3_res7__320_comb];
  assign p3_array_index_2046344_comb = p2_literal_2043912[p3_array_index_2046310_comb];
  assign p3_array_index_2046345_comb = p2_literal_2043914[p3_array_index_2046311_comb];
  assign p3_array_index_2046346_comb = p2_literal_2043916[p3_array_index_2046312_comb];
  assign p3_array_index_2046347_comb = p2_literal_2043918[p3_array_index_2046313_comb];
  assign p3_array_index_2046348_comb = p2_literal_2043920[p3_array_index_2046314_comb];
  assign p3_res7__322_comb = p3_array_index_2046343_comb ^ p3_array_index_2046344_comb ^ p3_array_index_2046345_comb ^ p3_array_index_2046346_comb ^ p3_array_index_2046347_comb ^ p3_array_index_2046348_comb ^ p3_array_index_2046315_comb ^ p2_literal_2043923[p3_array_index_2046332_comb] ^ p3_array_index_2046317_comb ^ p2_literal_2043920[p3_array_index_2046334_comb] ^ p2_literal_2043918[p3_array_index_2046319_comb] ^ p2_literal_2043916[p3_array_index_2046320_comb] ^ p2_literal_2043914[p3_array_index_2046321_comb] ^ p2_literal_2043912[p3_array_index_2046322_comb] ^ p2_literal_2043910[p3_array_index_2046323_comb] ^ p3_array_index_2046324_comb;
  assign p3_array_index_2046358_comb = p2_literal_2043912[p3_res7__320_comb];
  assign p3_array_index_2046359_comb = p2_literal_2043914[p3_array_index_2046310_comb];
  assign p3_array_index_2046360_comb = p2_literal_2043916[p3_array_index_2046311_comb];
  assign p3_array_index_2046361_comb = p2_literal_2043918[p3_array_index_2046312_comb];
  assign p3_array_index_2046362_comb = p2_literal_2043920[p3_array_index_2046313_comb];
  assign p3_res7__324_comb = p2_literal_2043910[p3_res7__322_comb] ^ p3_array_index_2046358_comb ^ p3_array_index_2046359_comb ^ p3_array_index_2046360_comb ^ p3_array_index_2046361_comb ^ p3_array_index_2046362_comb ^ p3_array_index_2046314_comb ^ p2_literal_2043923[p3_array_index_2046315_comb] ^ p3_array_index_2046332_comb ^ p2_literal_2043920[p3_array_index_2046317_comb] ^ p2_literal_2043918[p3_array_index_2046334_comb] ^ p2_literal_2043916[p3_array_index_2046319_comb] ^ p2_literal_2043914[p3_array_index_2046320_comb] ^ p2_literal_2043912[p3_array_index_2046321_comb] ^ p2_literal_2043910[p3_array_index_2046322_comb] ^ p3_array_index_2046323_comb;
  assign p3_array_index_2046372_comb = p2_literal_2043912[p3_res7__322_comb];
  assign p3_array_index_2046373_comb = p2_literal_2043914[p3_res7__320_comb];
  assign p3_array_index_2046374_comb = p2_literal_2043916[p3_array_index_2046310_comb];
  assign p3_array_index_2046375_comb = p2_literal_2043918[p3_array_index_2046311_comb];
  assign p3_array_index_2046376_comb = p2_literal_2043920[p3_array_index_2046312_comb];
  assign p3_res7__326_comb = p2_literal_2043910[p3_res7__324_comb] ^ p3_array_index_2046372_comb ^ p3_array_index_2046373_comb ^ p3_array_index_2046374_comb ^ p3_array_index_2046375_comb ^ p3_array_index_2046376_comb ^ p3_array_index_2046313_comb ^ p2_literal_2043923[p3_array_index_2046314_comb] ^ p3_array_index_2046315_comb ^ p2_literal_2043920[p3_array_index_2046332_comb] ^ p2_literal_2043918[p3_array_index_2046317_comb] ^ p2_literal_2043916[p3_array_index_2046334_comb] ^ p2_literal_2043914[p3_array_index_2046319_comb] ^ p2_literal_2043912[p3_array_index_2046320_comb] ^ p2_literal_2043910[p3_array_index_2046321_comb] ^ p3_array_index_2046322_comb;
  assign p3_array_index_2046387_comb = p2_literal_2043914[p3_res7__322_comb];
  assign p3_array_index_2046388_comb = p2_literal_2043916[p3_res7__320_comb];
  assign p3_array_index_2046389_comb = p2_literal_2043918[p3_array_index_2046310_comb];
  assign p3_array_index_2046390_comb = p2_literal_2043920[p3_array_index_2046311_comb];
  assign p3_res7__328_comb = p2_literal_2043910[p3_res7__326_comb] ^ p2_literal_2043912[p3_res7__324_comb] ^ p3_array_index_2046387_comb ^ p3_array_index_2046388_comb ^ p3_array_index_2046389_comb ^ p3_array_index_2046390_comb ^ p3_array_index_2046312_comb ^ p2_literal_2043923[p3_array_index_2046313_comb] ^ p3_array_index_2046314_comb ^ p3_array_index_2046331_comb ^ p2_literal_2043918[p3_array_index_2046332_comb] ^ p2_literal_2043916[p3_array_index_2046317_comb] ^ p2_literal_2043914[p3_array_index_2046334_comb] ^ p2_literal_2043912[p3_array_index_2046319_comb] ^ p2_literal_2043910[p3_array_index_2046320_comb] ^ p3_array_index_2046321_comb;
  assign p3_array_index_2046400_comb = p2_literal_2043914[p3_res7__324_comb];
  assign p3_array_index_2046401_comb = p2_literal_2043916[p3_res7__322_comb];
  assign p3_array_index_2046402_comb = p2_literal_2043918[p3_res7__320_comb];
  assign p3_array_index_2046403_comb = p2_literal_2043920[p3_array_index_2046310_comb];
  assign p3_res7__330_comb = p2_literal_2043910[p3_res7__328_comb] ^ p2_literal_2043912[p3_res7__326_comb] ^ p3_array_index_2046400_comb ^ p3_array_index_2046401_comb ^ p3_array_index_2046402_comb ^ p3_array_index_2046403_comb ^ p3_array_index_2046311_comb ^ p2_literal_2043923[p3_array_index_2046312_comb] ^ p3_array_index_2046313_comb ^ p3_array_index_2046348_comb ^ p2_literal_2043918[p3_array_index_2046315_comb] ^ p2_literal_2043916[p3_array_index_2046332_comb] ^ p2_literal_2043914[p3_array_index_2046317_comb] ^ p2_literal_2043912[p3_array_index_2046334_comb] ^ p2_literal_2043910[p3_array_index_2046319_comb] ^ p3_array_index_2046320_comb;
  assign p3_array_index_2046414_comb = p2_literal_2043916[p3_res7__324_comb];
  assign p3_array_index_2046415_comb = p2_literal_2043918[p3_res7__322_comb];
  assign p3_array_index_2046416_comb = p2_literal_2043920[p3_res7__320_comb];
  assign p3_res7__332_comb = p2_literal_2043910[p3_res7__330_comb] ^ p2_literal_2043912[p3_res7__328_comb] ^ p2_literal_2043914[p3_res7__326_comb] ^ p3_array_index_2046414_comb ^ p3_array_index_2046415_comb ^ p3_array_index_2046416_comb ^ p3_array_index_2046310_comb ^ p2_literal_2043923[p3_array_index_2046311_comb] ^ p3_array_index_2046312_comb ^ p3_array_index_2046362_comb ^ p3_array_index_2046330_comb ^ p2_literal_2043916[p3_array_index_2046315_comb] ^ p2_literal_2043914[p3_array_index_2046332_comb] ^ p2_literal_2043912[p3_array_index_2046317_comb] ^ p2_literal_2043910[p3_array_index_2046334_comb] ^ p3_array_index_2046319_comb;
  assign p3_array_index_2046426_comb = p2_literal_2043916[p3_res7__326_comb];
  assign p3_array_index_2046427_comb = p2_literal_2043918[p3_res7__324_comb];
  assign p3_array_index_2046428_comb = p2_literal_2043920[p3_res7__322_comb];
  assign p3_res7__334_comb = p2_literal_2043910[p3_res7__332_comb] ^ p2_literal_2043912[p3_res7__330_comb] ^ p2_literal_2043914[p3_res7__328_comb] ^ p3_array_index_2046426_comb ^ p3_array_index_2046427_comb ^ p3_array_index_2046428_comb ^ p3_res7__320_comb ^ p2_literal_2043923[p3_array_index_2046310_comb] ^ p3_array_index_2046311_comb ^ p3_array_index_2046376_comb ^ p3_array_index_2046347_comb ^ p2_literal_2043916[p3_array_index_2046314_comb] ^ p2_literal_2043914[p3_array_index_2046315_comb] ^ p2_literal_2043912[p3_array_index_2046332_comb] ^ p2_literal_2043910[p3_array_index_2046317_comb] ^ p3_array_index_2046334_comb;
  assign p3_array_index_2046439_comb = p2_literal_2043918[p3_res7__326_comb];
  assign p3_array_index_2046440_comb = p2_literal_2043920[p3_res7__324_comb];
  assign p3_res7__336_comb = p2_literal_2043910[p3_res7__334_comb] ^ p2_literal_2043912[p3_res7__332_comb] ^ p2_literal_2043914[p3_res7__330_comb] ^ p2_literal_2043916[p3_res7__328_comb] ^ p3_array_index_2046439_comb ^ p3_array_index_2046440_comb ^ p3_res7__322_comb ^ p2_literal_2043923[p3_res7__320_comb] ^ p3_array_index_2046310_comb ^ p3_array_index_2046390_comb ^ p3_array_index_2046361_comb ^ p3_array_index_2046329_comb ^ p2_literal_2043914[p3_array_index_2046314_comb] ^ p2_literal_2043912[p3_array_index_2046315_comb] ^ p2_literal_2043910[p3_array_index_2046332_comb] ^ p3_array_index_2046317_comb;
  assign p3_array_index_2046450_comb = p2_literal_2043918[p3_res7__328_comb];
  assign p3_array_index_2046451_comb = p2_literal_2043920[p3_res7__326_comb];
  assign p3_res7__338_comb = p2_literal_2043910[p3_res7__336_comb] ^ p2_literal_2043912[p3_res7__334_comb] ^ p2_literal_2043914[p3_res7__332_comb] ^ p2_literal_2043916[p3_res7__330_comb] ^ p3_array_index_2046450_comb ^ p3_array_index_2046451_comb ^ p3_res7__324_comb ^ p2_literal_2043923[p3_res7__322_comb] ^ p3_res7__320_comb ^ p3_array_index_2046403_comb ^ p3_array_index_2046375_comb ^ p3_array_index_2046346_comb ^ p2_literal_2043914[p3_array_index_2046313_comb] ^ p2_literal_2043912[p3_array_index_2046314_comb] ^ p2_literal_2043910[p3_array_index_2046315_comb] ^ p3_array_index_2046332_comb;
  assign p3_array_index_2046462_comb = p2_literal_2043920[p3_res7__328_comb];
  assign p3_res7__340_comb = p2_literal_2043910[p3_res7__338_comb] ^ p2_literal_2043912[p3_res7__336_comb] ^ p2_literal_2043914[p3_res7__334_comb] ^ p2_literal_2043916[p3_res7__332_comb] ^ p2_literal_2043918[p3_res7__330_comb] ^ p3_array_index_2046462_comb ^ p3_res7__326_comb ^ p2_literal_2043923[p3_res7__324_comb] ^ p3_res7__322_comb ^ p3_array_index_2046416_comb ^ p3_array_index_2046389_comb ^ p3_array_index_2046360_comb ^ p3_array_index_2046328_comb ^ p2_literal_2043912[p3_array_index_2046313_comb] ^ p2_literal_2043910[p3_array_index_2046314_comb] ^ p3_array_index_2046315_comb;
  assign p3_array_index_2046472_comb = p2_literal_2043920[p3_res7__330_comb];
  assign p3_res7__342_comb = p2_literal_2043910[p3_res7__340_comb] ^ p2_literal_2043912[p3_res7__338_comb] ^ p2_literal_2043914[p3_res7__336_comb] ^ p2_literal_2043916[p3_res7__334_comb] ^ p2_literal_2043918[p3_res7__332_comb] ^ p3_array_index_2046472_comb ^ p3_res7__328_comb ^ p2_literal_2043923[p3_res7__326_comb] ^ p3_res7__324_comb ^ p3_array_index_2046428_comb ^ p3_array_index_2046402_comb ^ p3_array_index_2046374_comb ^ p3_array_index_2046345_comb ^ p2_literal_2043912[p3_array_index_2046312_comb] ^ p2_literal_2043910[p3_array_index_2046313_comb] ^ p3_array_index_2046314_comb;
  assign p3_res7__344_comb = p2_literal_2043910[p3_res7__342_comb] ^ p2_literal_2043912[p3_res7__340_comb] ^ p2_literal_2043914[p3_res7__338_comb] ^ p2_literal_2043916[p3_res7__336_comb] ^ p2_literal_2043918[p3_res7__334_comb] ^ p2_literal_2043920[p3_res7__332_comb] ^ p3_res7__330_comb ^ p2_literal_2043923[p3_res7__328_comb] ^ p3_res7__326_comb ^ p3_array_index_2046440_comb ^ p3_array_index_2046415_comb ^ p3_array_index_2046388_comb ^ p3_array_index_2046359_comb ^ p3_array_index_2046327_comb ^ p2_literal_2043910[p3_array_index_2046312_comb] ^ p3_array_index_2046313_comb;
  assign p3_res7__346_comb = p2_literal_2043910[p3_res7__344_comb] ^ p2_literal_2043912[p3_res7__342_comb] ^ p2_literal_2043914[p3_res7__340_comb] ^ p2_literal_2043916[p3_res7__338_comb] ^ p2_literal_2043918[p3_res7__336_comb] ^ p2_literal_2043920[p3_res7__334_comb] ^ p3_res7__332_comb ^ p2_literal_2043923[p3_res7__330_comb] ^ p3_res7__328_comb ^ p3_array_index_2046451_comb ^ p3_array_index_2046427_comb ^ p3_array_index_2046401_comb ^ p3_array_index_2046373_comb ^ p3_array_index_2046344_comb ^ p2_literal_2043910[p3_array_index_2046311_comb] ^ p3_array_index_2046312_comb;
  assign p3_res7__348_comb = p2_literal_2043910[p3_res7__346_comb] ^ p2_literal_2043912[p3_res7__344_comb] ^ p2_literal_2043914[p3_res7__342_comb] ^ p2_literal_2043916[p3_res7__340_comb] ^ p2_literal_2043918[p3_res7__338_comb] ^ p2_literal_2043920[p3_res7__336_comb] ^ p3_res7__334_comb ^ p2_literal_2043923[p3_res7__332_comb] ^ p3_res7__330_comb ^ p3_array_index_2046462_comb ^ p3_array_index_2046439_comb ^ p3_array_index_2046414_comb ^ p3_array_index_2046387_comb ^ p3_array_index_2046358_comb ^ p3_array_index_2046326_comb ^ p3_array_index_2046311_comb;
  assign p3_res7__350_comb = p2_literal_2043910[p3_res7__348_comb] ^ p2_literal_2043912[p3_res7__346_comb] ^ p2_literal_2043914[p3_res7__344_comb] ^ p2_literal_2043916[p3_res7__342_comb] ^ p2_literal_2043918[p3_res7__340_comb] ^ p2_literal_2043920[p3_res7__338_comb] ^ p3_res7__336_comb ^ p2_literal_2043923[p3_res7__334_comb] ^ p3_res7__332_comb ^ p3_array_index_2046472_comb ^ p3_array_index_2046450_comb ^ p3_array_index_2046426_comb ^ p3_array_index_2046400_comb ^ p3_array_index_2046372_comb ^ p3_array_index_2046343_comb ^ p3_array_index_2046310_comb;
  assign p3_res__10_comb = {p3_res7__350_comb, p3_res7__348_comb, p3_res7__346_comb, p3_res7__344_comb, p3_res7__342_comb, p3_res7__340_comb, p3_res7__338_comb, p3_res7__336_comb, p3_res7__334_comb, p3_res7__332_comb, p3_res7__330_comb, p3_res7__328_comb, p3_res7__326_comb, p3_res7__324_comb, p3_res7__322_comb, p3_res7__320_comb};
  assign p3_xor_2046512_comb = p3_res__10_comb ^ p3_xor_2046076_comb;
  assign p3_addedKey__43_comb = p3_xor_2046512_comb ^ 128'h8d94_2d1d_95e6_7d2c_1a67_10c0_d5ff_3f0c;
  assign p3_array_index_2046528_comb = p2_literal_2043896[p3_addedKey__43_comb[127:120]];
  assign p3_array_index_2046529_comb = p2_literal_2043896[p3_addedKey__43_comb[119:112]];
  assign p3_array_index_2046530_comb = p2_literal_2043896[p3_addedKey__43_comb[111:104]];
  assign p3_array_index_2046531_comb = p2_literal_2043896[p3_addedKey__43_comb[103:96]];
  assign p3_array_index_2046532_comb = p2_literal_2043896[p3_addedKey__43_comb[95:88]];
  assign p3_array_index_2046533_comb = p2_literal_2043896[p3_addedKey__43_comb[87:80]];
  assign p3_array_index_2046535_comb = p2_literal_2043896[p3_addedKey__43_comb[71:64]];
  assign p3_array_index_2046537_comb = p2_literal_2043896[p3_addedKey__43_comb[55:48]];
  assign p3_array_index_2046538_comb = p2_literal_2043896[p3_addedKey__43_comb[47:40]];
  assign p3_array_index_2046539_comb = p2_literal_2043896[p3_addedKey__43_comb[39:32]];
  assign p3_array_index_2046540_comb = p2_literal_2043896[p3_addedKey__43_comb[31:24]];
  assign p3_array_index_2046541_comb = p2_literal_2043896[p3_addedKey__43_comb[23:16]];
  assign p3_array_index_2046542_comb = p2_literal_2043896[p3_addedKey__43_comb[15:8]];
  assign p3_array_index_2046544_comb = p2_literal_2043910[p3_array_index_2046528_comb];
  assign p3_array_index_2046545_comb = p2_literal_2043912[p3_array_index_2046529_comb];
  assign p3_array_index_2046546_comb = p2_literal_2043914[p3_array_index_2046530_comb];
  assign p3_array_index_2046547_comb = p2_literal_2043916[p3_array_index_2046531_comb];
  assign p3_array_index_2046548_comb = p2_literal_2043918[p3_array_index_2046532_comb];
  assign p3_array_index_2046549_comb = p2_literal_2043920[p3_array_index_2046533_comb];
  assign p3_array_index_2046550_comb = p2_literal_2043896[p3_addedKey__43_comb[79:72]];
  assign p3_array_index_2046552_comb = p2_literal_2043896[p3_addedKey__43_comb[63:56]];
  assign p3_res7__352_comb = p3_array_index_2046544_comb ^ p3_array_index_2046545_comb ^ p3_array_index_2046546_comb ^ p3_array_index_2046547_comb ^ p3_array_index_2046548_comb ^ p3_array_index_2046549_comb ^ p3_array_index_2046550_comb ^ p2_literal_2043923[p3_array_index_2046535_comb] ^ p3_array_index_2046552_comb ^ p2_literal_2043920[p3_array_index_2046537_comb] ^ p2_literal_2043918[p3_array_index_2046538_comb] ^ p2_literal_2043916[p3_array_index_2046539_comb] ^ p2_literal_2043914[p3_array_index_2046540_comb] ^ p2_literal_2043912[p3_array_index_2046541_comb] ^ p2_literal_2043910[p3_array_index_2046542_comb] ^ p2_literal_2043896[p3_addedKey__43_comb[7:0]];
  assign p3_array_index_2046561_comb = p2_literal_2043910[p3_res7__352_comb];
  assign p3_array_index_2046562_comb = p2_literal_2043912[p3_array_index_2046528_comb];
  assign p3_array_index_2046563_comb = p2_literal_2043914[p3_array_index_2046529_comb];
  assign p3_array_index_2046564_comb = p2_literal_2043916[p3_array_index_2046530_comb];
  assign p3_array_index_2046565_comb = p2_literal_2043918[p3_array_index_2046531_comb];
  assign p3_array_index_2046566_comb = p2_literal_2043920[p3_array_index_2046532_comb];
  assign p3_res7__354_comb = p3_array_index_2046561_comb ^ p3_array_index_2046562_comb ^ p3_array_index_2046563_comb ^ p3_array_index_2046564_comb ^ p3_array_index_2046565_comb ^ p3_array_index_2046566_comb ^ p3_array_index_2046533_comb ^ p2_literal_2043923[p3_array_index_2046550_comb] ^ p3_array_index_2046535_comb ^ p2_literal_2043920[p3_array_index_2046552_comb] ^ p2_literal_2043918[p3_array_index_2046537_comb] ^ p2_literal_2043916[p3_array_index_2046538_comb] ^ p2_literal_2043914[p3_array_index_2046539_comb] ^ p2_literal_2043912[p3_array_index_2046540_comb] ^ p2_literal_2043910[p3_array_index_2046541_comb] ^ p3_array_index_2046542_comb;
  assign p3_array_index_2046576_comb = p2_literal_2043912[p3_res7__352_comb];
  assign p3_array_index_2046577_comb = p2_literal_2043914[p3_array_index_2046528_comb];
  assign p3_array_index_2046578_comb = p2_literal_2043916[p3_array_index_2046529_comb];
  assign p3_array_index_2046579_comb = p2_literal_2043918[p3_array_index_2046530_comb];
  assign p3_array_index_2046580_comb = p2_literal_2043920[p3_array_index_2046531_comb];
  assign p3_res7__356_comb = p2_literal_2043910[p3_res7__354_comb] ^ p3_array_index_2046576_comb ^ p3_array_index_2046577_comb ^ p3_array_index_2046578_comb ^ p3_array_index_2046579_comb ^ p3_array_index_2046580_comb ^ p3_array_index_2046532_comb ^ p2_literal_2043923[p3_array_index_2046533_comb] ^ p3_array_index_2046550_comb ^ p2_literal_2043920[p3_array_index_2046535_comb] ^ p2_literal_2043918[p3_array_index_2046552_comb] ^ p2_literal_2043916[p3_array_index_2046537_comb] ^ p2_literal_2043914[p3_array_index_2046538_comb] ^ p2_literal_2043912[p3_array_index_2046539_comb] ^ p2_literal_2043910[p3_array_index_2046540_comb] ^ p3_array_index_2046541_comb;
  assign p3_array_index_2046590_comb = p2_literal_2043912[p3_res7__354_comb];
  assign p3_array_index_2046591_comb = p2_literal_2043914[p3_res7__352_comb];
  assign p3_array_index_2046592_comb = p2_literal_2043916[p3_array_index_2046528_comb];
  assign p3_array_index_2046593_comb = p2_literal_2043918[p3_array_index_2046529_comb];
  assign p3_array_index_2046594_comb = p2_literal_2043920[p3_array_index_2046530_comb];
  assign p3_res7__358_comb = p2_literal_2043910[p3_res7__356_comb] ^ p3_array_index_2046590_comb ^ p3_array_index_2046591_comb ^ p3_array_index_2046592_comb ^ p3_array_index_2046593_comb ^ p3_array_index_2046594_comb ^ p3_array_index_2046531_comb ^ p2_literal_2043923[p3_array_index_2046532_comb] ^ p3_array_index_2046533_comb ^ p2_literal_2043920[p3_array_index_2046550_comb] ^ p2_literal_2043918[p3_array_index_2046535_comb] ^ p2_literal_2043916[p3_array_index_2046552_comb] ^ p2_literal_2043914[p3_array_index_2046537_comb] ^ p2_literal_2043912[p3_array_index_2046538_comb] ^ p2_literal_2043910[p3_array_index_2046539_comb] ^ p3_array_index_2046540_comb;
  assign p3_array_index_2046605_comb = p2_literal_2043914[p3_res7__354_comb];
  assign p3_array_index_2046606_comb = p2_literal_2043916[p3_res7__352_comb];
  assign p3_array_index_2046607_comb = p2_literal_2043918[p3_array_index_2046528_comb];
  assign p3_array_index_2046608_comb = p2_literal_2043920[p3_array_index_2046529_comb];
  assign p3_res7__360_comb = p2_literal_2043910[p3_res7__358_comb] ^ p2_literal_2043912[p3_res7__356_comb] ^ p3_array_index_2046605_comb ^ p3_array_index_2046606_comb ^ p3_array_index_2046607_comb ^ p3_array_index_2046608_comb ^ p3_array_index_2046530_comb ^ p2_literal_2043923[p3_array_index_2046531_comb] ^ p3_array_index_2046532_comb ^ p3_array_index_2046549_comb ^ p2_literal_2043918[p3_array_index_2046550_comb] ^ p2_literal_2043916[p3_array_index_2046535_comb] ^ p2_literal_2043914[p3_array_index_2046552_comb] ^ p2_literal_2043912[p3_array_index_2046537_comb] ^ p2_literal_2043910[p3_array_index_2046538_comb] ^ p3_array_index_2046539_comb;
  assign p3_array_index_2046618_comb = p2_literal_2043914[p3_res7__356_comb];
  assign p3_array_index_2046619_comb = p2_literal_2043916[p3_res7__354_comb];
  assign p3_array_index_2046620_comb = p2_literal_2043918[p3_res7__352_comb];
  assign p3_array_index_2046621_comb = p2_literal_2043920[p3_array_index_2046528_comb];
  assign p3_res7__362_comb = p2_literal_2043910[p3_res7__360_comb] ^ p2_literal_2043912[p3_res7__358_comb] ^ p3_array_index_2046618_comb ^ p3_array_index_2046619_comb ^ p3_array_index_2046620_comb ^ p3_array_index_2046621_comb ^ p3_array_index_2046529_comb ^ p2_literal_2043923[p3_array_index_2046530_comb] ^ p3_array_index_2046531_comb ^ p3_array_index_2046566_comb ^ p2_literal_2043918[p3_array_index_2046533_comb] ^ p2_literal_2043916[p3_array_index_2046550_comb] ^ p2_literal_2043914[p3_array_index_2046535_comb] ^ p2_literal_2043912[p3_array_index_2046552_comb] ^ p2_literal_2043910[p3_array_index_2046537_comb] ^ p3_array_index_2046538_comb;
  assign p3_array_index_2046632_comb = p2_literal_2043916[p3_res7__356_comb];
  assign p3_array_index_2046633_comb = p2_literal_2043918[p3_res7__354_comb];
  assign p3_array_index_2046634_comb = p2_literal_2043920[p3_res7__352_comb];
  assign p3_res7__364_comb = p2_literal_2043910[p3_res7__362_comb] ^ p2_literal_2043912[p3_res7__360_comb] ^ p2_literal_2043914[p3_res7__358_comb] ^ p3_array_index_2046632_comb ^ p3_array_index_2046633_comb ^ p3_array_index_2046634_comb ^ p3_array_index_2046528_comb ^ p2_literal_2043923[p3_array_index_2046529_comb] ^ p3_array_index_2046530_comb ^ p3_array_index_2046580_comb ^ p3_array_index_2046548_comb ^ p2_literal_2043916[p3_array_index_2046533_comb] ^ p2_literal_2043914[p3_array_index_2046550_comb] ^ p2_literal_2043912[p3_array_index_2046535_comb] ^ p2_literal_2043910[p3_array_index_2046552_comb] ^ p3_array_index_2046537_comb;
  assign p3_array_index_2046644_comb = p2_literal_2043916[p3_res7__358_comb];
  assign p3_array_index_2046645_comb = p2_literal_2043918[p3_res7__356_comb];
  assign p3_array_index_2046646_comb = p2_literal_2043920[p3_res7__354_comb];
  assign p3_res7__366_comb = p2_literal_2043910[p3_res7__364_comb] ^ p2_literal_2043912[p3_res7__362_comb] ^ p2_literal_2043914[p3_res7__360_comb] ^ p3_array_index_2046644_comb ^ p3_array_index_2046645_comb ^ p3_array_index_2046646_comb ^ p3_res7__352_comb ^ p2_literal_2043923[p3_array_index_2046528_comb] ^ p3_array_index_2046529_comb ^ p3_array_index_2046594_comb ^ p3_array_index_2046565_comb ^ p2_literal_2043916[p3_array_index_2046532_comb] ^ p2_literal_2043914[p3_array_index_2046533_comb] ^ p2_literal_2043912[p3_array_index_2046550_comb] ^ p2_literal_2043910[p3_array_index_2046535_comb] ^ p3_array_index_2046552_comb;
  assign p3_array_index_2046657_comb = p2_literal_2043918[p3_res7__358_comb];
  assign p3_array_index_2046658_comb = p2_literal_2043920[p3_res7__356_comb];
  assign p3_res7__368_comb = p2_literal_2043910[p3_res7__366_comb] ^ p2_literal_2043912[p3_res7__364_comb] ^ p2_literal_2043914[p3_res7__362_comb] ^ p2_literal_2043916[p3_res7__360_comb] ^ p3_array_index_2046657_comb ^ p3_array_index_2046658_comb ^ p3_res7__354_comb ^ p2_literal_2043923[p3_res7__352_comb] ^ p3_array_index_2046528_comb ^ p3_array_index_2046608_comb ^ p3_array_index_2046579_comb ^ p3_array_index_2046547_comb ^ p2_literal_2043914[p3_array_index_2046532_comb] ^ p2_literal_2043912[p3_array_index_2046533_comb] ^ p2_literal_2043910[p3_array_index_2046550_comb] ^ p3_array_index_2046535_comb;
  assign p3_array_index_2046668_comb = p2_literal_2043918[p3_res7__360_comb];
  assign p3_array_index_2046669_comb = p2_literal_2043920[p3_res7__358_comb];
  assign p3_res7__370_comb = p2_literal_2043910[p3_res7__368_comb] ^ p2_literal_2043912[p3_res7__366_comb] ^ p2_literal_2043914[p3_res7__364_comb] ^ p2_literal_2043916[p3_res7__362_comb] ^ p3_array_index_2046668_comb ^ p3_array_index_2046669_comb ^ p3_res7__356_comb ^ p2_literal_2043923[p3_res7__354_comb] ^ p3_res7__352_comb ^ p3_array_index_2046621_comb ^ p3_array_index_2046593_comb ^ p3_array_index_2046564_comb ^ p2_literal_2043914[p3_array_index_2046531_comb] ^ p2_literal_2043912[p3_array_index_2046532_comb] ^ p2_literal_2043910[p3_array_index_2046533_comb] ^ p3_array_index_2046550_comb;
  assign p3_array_index_2046680_comb = p2_literal_2043920[p3_res7__360_comb];
  assign p3_res7__372_comb = p2_literal_2043910[p3_res7__370_comb] ^ p2_literal_2043912[p3_res7__368_comb] ^ p2_literal_2043914[p3_res7__366_comb] ^ p2_literal_2043916[p3_res7__364_comb] ^ p2_literal_2043918[p3_res7__362_comb] ^ p3_array_index_2046680_comb ^ p3_res7__358_comb ^ p2_literal_2043923[p3_res7__356_comb] ^ p3_res7__354_comb ^ p3_array_index_2046634_comb ^ p3_array_index_2046607_comb ^ p3_array_index_2046578_comb ^ p3_array_index_2046546_comb ^ p2_literal_2043912[p3_array_index_2046531_comb] ^ p2_literal_2043910[p3_array_index_2046532_comb] ^ p3_array_index_2046533_comb;
  assign p3_array_index_2046690_comb = p2_literal_2043920[p3_res7__362_comb];
  assign p3_res7__374_comb = p2_literal_2043910[p3_res7__372_comb] ^ p2_literal_2043912[p3_res7__370_comb] ^ p2_literal_2043914[p3_res7__368_comb] ^ p2_literal_2043916[p3_res7__366_comb] ^ p2_literal_2043918[p3_res7__364_comb] ^ p3_array_index_2046690_comb ^ p3_res7__360_comb ^ p2_literal_2043923[p3_res7__358_comb] ^ p3_res7__356_comb ^ p3_array_index_2046646_comb ^ p3_array_index_2046620_comb ^ p3_array_index_2046592_comb ^ p3_array_index_2046563_comb ^ p2_literal_2043912[p3_array_index_2046530_comb] ^ p2_literal_2043910[p3_array_index_2046531_comb] ^ p3_array_index_2046532_comb;
  assign p3_res7__376_comb = p2_literal_2043910[p3_res7__374_comb] ^ p2_literal_2043912[p3_res7__372_comb] ^ p2_literal_2043914[p3_res7__370_comb] ^ p2_literal_2043916[p3_res7__368_comb] ^ p2_literal_2043918[p3_res7__366_comb] ^ p2_literal_2043920[p3_res7__364_comb] ^ p3_res7__362_comb ^ p2_literal_2043923[p3_res7__360_comb] ^ p3_res7__358_comb ^ p3_array_index_2046658_comb ^ p3_array_index_2046633_comb ^ p3_array_index_2046606_comb ^ p3_array_index_2046577_comb ^ p3_array_index_2046545_comb ^ p2_literal_2043910[p3_array_index_2046530_comb] ^ p3_array_index_2046531_comb;
  assign p3_res7__378_comb = p2_literal_2043910[p3_res7__376_comb] ^ p2_literal_2043912[p3_res7__374_comb] ^ p2_literal_2043914[p3_res7__372_comb] ^ p2_literal_2043916[p3_res7__370_comb] ^ p2_literal_2043918[p3_res7__368_comb] ^ p2_literal_2043920[p3_res7__366_comb] ^ p3_res7__364_comb ^ p2_literal_2043923[p3_res7__362_comb] ^ p3_res7__360_comb ^ p3_array_index_2046669_comb ^ p3_array_index_2046645_comb ^ p3_array_index_2046619_comb ^ p3_array_index_2046591_comb ^ p3_array_index_2046562_comb ^ p2_literal_2043910[p3_array_index_2046529_comb] ^ p3_array_index_2046530_comb;
  assign p3_res7__380_comb = p2_literal_2043910[p3_res7__378_comb] ^ p2_literal_2043912[p3_res7__376_comb] ^ p2_literal_2043914[p3_res7__374_comb] ^ p2_literal_2043916[p3_res7__372_comb] ^ p2_literal_2043918[p3_res7__370_comb] ^ p2_literal_2043920[p3_res7__368_comb] ^ p3_res7__366_comb ^ p2_literal_2043923[p3_res7__364_comb] ^ p3_res7__362_comb ^ p3_array_index_2046680_comb ^ p3_array_index_2046657_comb ^ p3_array_index_2046632_comb ^ p3_array_index_2046605_comb ^ p3_array_index_2046576_comb ^ p3_array_index_2046544_comb ^ p3_array_index_2046529_comb;
  assign p3_res7__382_comb = p2_literal_2043910[p3_res7__380_comb] ^ p2_literal_2043912[p3_res7__378_comb] ^ p2_literal_2043914[p3_res7__376_comb] ^ p2_literal_2043916[p3_res7__374_comb] ^ p2_literal_2043918[p3_res7__372_comb] ^ p2_literal_2043920[p3_res7__370_comb] ^ p3_res7__368_comb ^ p2_literal_2043923[p3_res7__366_comb] ^ p3_res7__364_comb ^ p3_array_index_2046690_comb ^ p3_array_index_2046668_comb ^ p3_array_index_2046644_comb ^ p3_array_index_2046618_comb ^ p3_array_index_2046590_comb ^ p3_array_index_2046561_comb ^ p3_array_index_2046528_comb;
  assign p3_res__11_comb = {p3_res7__382_comb, p3_res7__380_comb, p3_res7__378_comb, p3_res7__376_comb, p3_res7__374_comb, p3_res7__372_comb, p3_res7__370_comb, p3_res7__368_comb, p3_res7__366_comb, p3_res7__364_comb, p3_res7__362_comb, p3_res7__360_comb, p3_res7__358_comb, p3_res7__356_comb, p3_res7__354_comb, p3_res7__352_comb};
  assign p3_xor_2046730_comb = p3_res__11_comb ^ p3_xor_2046294_comb;
  assign p3_addedKey__44_comb = p3_xor_2046730_comb ^ 128'he336_5b6f_f9ae_0794_4740_add0_087b_ab0d;
  assign p3_array_index_2046746_comb = p2_literal_2043896[p3_addedKey__44_comb[127:120]];
  assign p3_array_index_2046747_comb = p2_literal_2043896[p3_addedKey__44_comb[119:112]];
  assign p3_array_index_2046748_comb = p2_literal_2043896[p3_addedKey__44_comb[111:104]];
  assign p3_array_index_2046749_comb = p2_literal_2043896[p3_addedKey__44_comb[103:96]];
  assign p3_array_index_2046750_comb = p2_literal_2043896[p3_addedKey__44_comb[95:88]];
  assign p3_array_index_2046751_comb = p2_literal_2043896[p3_addedKey__44_comb[87:80]];
  assign p3_array_index_2046753_comb = p2_literal_2043896[p3_addedKey__44_comb[71:64]];
  assign p3_array_index_2046755_comb = p2_literal_2043896[p3_addedKey__44_comb[55:48]];
  assign p3_array_index_2046756_comb = p2_literal_2043896[p3_addedKey__44_comb[47:40]];
  assign p3_array_index_2046757_comb = p2_literal_2043896[p3_addedKey__44_comb[39:32]];
  assign p3_array_index_2046758_comb = p2_literal_2043896[p3_addedKey__44_comb[31:24]];
  assign p3_array_index_2046759_comb = p2_literal_2043896[p3_addedKey__44_comb[23:16]];
  assign p3_array_index_2046760_comb = p2_literal_2043896[p3_addedKey__44_comb[15:8]];
  assign p3_array_index_2046762_comb = p2_literal_2043910[p3_array_index_2046746_comb];
  assign p3_array_index_2046763_comb = p2_literal_2043912[p3_array_index_2046747_comb];
  assign p3_array_index_2046764_comb = p2_literal_2043914[p3_array_index_2046748_comb];
  assign p3_array_index_2046765_comb = p2_literal_2043916[p3_array_index_2046749_comb];
  assign p3_array_index_2046766_comb = p2_literal_2043918[p3_array_index_2046750_comb];
  assign p3_array_index_2046767_comb = p2_literal_2043920[p3_array_index_2046751_comb];
  assign p3_array_index_2046768_comb = p2_literal_2043896[p3_addedKey__44_comb[79:72]];
  assign p3_array_index_2046770_comb = p2_literal_2043896[p3_addedKey__44_comb[63:56]];
  assign p3_res7__384_comb = p3_array_index_2046762_comb ^ p3_array_index_2046763_comb ^ p3_array_index_2046764_comb ^ p3_array_index_2046765_comb ^ p3_array_index_2046766_comb ^ p3_array_index_2046767_comb ^ p3_array_index_2046768_comb ^ p2_literal_2043923[p3_array_index_2046753_comb] ^ p3_array_index_2046770_comb ^ p2_literal_2043920[p3_array_index_2046755_comb] ^ p2_literal_2043918[p3_array_index_2046756_comb] ^ p2_literal_2043916[p3_array_index_2046757_comb] ^ p2_literal_2043914[p3_array_index_2046758_comb] ^ p2_literal_2043912[p3_array_index_2046759_comb] ^ p2_literal_2043910[p3_array_index_2046760_comb] ^ p2_literal_2043896[p3_addedKey__44_comb[7:0]];
  assign p3_array_index_2046779_comb = p2_literal_2043910[p3_res7__384_comb];
  assign p3_array_index_2046780_comb = p2_literal_2043912[p3_array_index_2046746_comb];
  assign p3_array_index_2046781_comb = p2_literal_2043914[p3_array_index_2046747_comb];
  assign p3_array_index_2046782_comb = p2_literal_2043916[p3_array_index_2046748_comb];
  assign p3_array_index_2046783_comb = p2_literal_2043918[p3_array_index_2046749_comb];
  assign p3_array_index_2046784_comb = p2_literal_2043920[p3_array_index_2046750_comb];
  assign p3_res7__386_comb = p3_array_index_2046779_comb ^ p3_array_index_2046780_comb ^ p3_array_index_2046781_comb ^ p3_array_index_2046782_comb ^ p3_array_index_2046783_comb ^ p3_array_index_2046784_comb ^ p3_array_index_2046751_comb ^ p2_literal_2043923[p3_array_index_2046768_comb] ^ p3_array_index_2046753_comb ^ p2_literal_2043920[p3_array_index_2046770_comb] ^ p2_literal_2043918[p3_array_index_2046755_comb] ^ p2_literal_2043916[p3_array_index_2046756_comb] ^ p2_literal_2043914[p3_array_index_2046757_comb] ^ p2_literal_2043912[p3_array_index_2046758_comb] ^ p2_literal_2043910[p3_array_index_2046759_comb] ^ p3_array_index_2046760_comb;
  assign p3_array_index_2046794_comb = p2_literal_2043912[p3_res7__384_comb];
  assign p3_array_index_2046795_comb = p2_literal_2043914[p3_array_index_2046746_comb];
  assign p3_array_index_2046796_comb = p2_literal_2043916[p3_array_index_2046747_comb];
  assign p3_array_index_2046797_comb = p2_literal_2043918[p3_array_index_2046748_comb];
  assign p3_array_index_2046798_comb = p2_literal_2043920[p3_array_index_2046749_comb];
  assign p3_res7__388_comb = p2_literal_2043910[p3_res7__386_comb] ^ p3_array_index_2046794_comb ^ p3_array_index_2046795_comb ^ p3_array_index_2046796_comb ^ p3_array_index_2046797_comb ^ p3_array_index_2046798_comb ^ p3_array_index_2046750_comb ^ p2_literal_2043923[p3_array_index_2046751_comb] ^ p3_array_index_2046768_comb ^ p2_literal_2043920[p3_array_index_2046753_comb] ^ p2_literal_2043918[p3_array_index_2046770_comb] ^ p2_literal_2043916[p3_array_index_2046755_comb] ^ p2_literal_2043914[p3_array_index_2046756_comb] ^ p2_literal_2043912[p3_array_index_2046757_comb] ^ p2_literal_2043910[p3_array_index_2046758_comb] ^ p3_array_index_2046759_comb;
  assign p3_array_index_2046808_comb = p2_literal_2043912[p3_res7__386_comb];
  assign p3_array_index_2046809_comb = p2_literal_2043914[p3_res7__384_comb];
  assign p3_array_index_2046810_comb = p2_literal_2043916[p3_array_index_2046746_comb];
  assign p3_array_index_2046811_comb = p2_literal_2043918[p3_array_index_2046747_comb];
  assign p3_array_index_2046812_comb = p2_literal_2043920[p3_array_index_2046748_comb];
  assign p3_res7__390_comb = p2_literal_2043910[p3_res7__388_comb] ^ p3_array_index_2046808_comb ^ p3_array_index_2046809_comb ^ p3_array_index_2046810_comb ^ p3_array_index_2046811_comb ^ p3_array_index_2046812_comb ^ p3_array_index_2046749_comb ^ p2_literal_2043923[p3_array_index_2046750_comb] ^ p3_array_index_2046751_comb ^ p2_literal_2043920[p3_array_index_2046768_comb] ^ p2_literal_2043918[p3_array_index_2046753_comb] ^ p2_literal_2043916[p3_array_index_2046770_comb] ^ p2_literal_2043914[p3_array_index_2046755_comb] ^ p2_literal_2043912[p3_array_index_2046756_comb] ^ p2_literal_2043910[p3_array_index_2046757_comb] ^ p3_array_index_2046758_comb;
  assign p3_array_index_2046823_comb = p2_literal_2043914[p3_res7__386_comb];
  assign p3_array_index_2046824_comb = p2_literal_2043916[p3_res7__384_comb];
  assign p3_array_index_2046825_comb = p2_literal_2043918[p3_array_index_2046746_comb];
  assign p3_array_index_2046826_comb = p2_literal_2043920[p3_array_index_2046747_comb];
  assign p3_res7__392_comb = p2_literal_2043910[p3_res7__390_comb] ^ p2_literal_2043912[p3_res7__388_comb] ^ p3_array_index_2046823_comb ^ p3_array_index_2046824_comb ^ p3_array_index_2046825_comb ^ p3_array_index_2046826_comb ^ p3_array_index_2046748_comb ^ p2_literal_2043923[p3_array_index_2046749_comb] ^ p3_array_index_2046750_comb ^ p3_array_index_2046767_comb ^ p2_literal_2043918[p3_array_index_2046768_comb] ^ p2_literal_2043916[p3_array_index_2046753_comb] ^ p2_literal_2043914[p3_array_index_2046770_comb] ^ p2_literal_2043912[p3_array_index_2046755_comb] ^ p2_literal_2043910[p3_array_index_2046756_comb] ^ p3_array_index_2046757_comb;
  assign p3_array_index_2046836_comb = p2_literal_2043914[p3_res7__388_comb];
  assign p3_array_index_2046837_comb = p2_literal_2043916[p3_res7__386_comb];
  assign p3_array_index_2046838_comb = p2_literal_2043918[p3_res7__384_comb];
  assign p3_array_index_2046839_comb = p2_literal_2043920[p3_array_index_2046746_comb];
  assign p3_res7__394_comb = p2_literal_2043910[p3_res7__392_comb] ^ p2_literal_2043912[p3_res7__390_comb] ^ p3_array_index_2046836_comb ^ p3_array_index_2046837_comb ^ p3_array_index_2046838_comb ^ p3_array_index_2046839_comb ^ p3_array_index_2046747_comb ^ p2_literal_2043923[p3_array_index_2046748_comb] ^ p3_array_index_2046749_comb ^ p3_array_index_2046784_comb ^ p2_literal_2043918[p3_array_index_2046751_comb] ^ p2_literal_2043916[p3_array_index_2046768_comb] ^ p2_literal_2043914[p3_array_index_2046753_comb] ^ p2_literal_2043912[p3_array_index_2046770_comb] ^ p2_literal_2043910[p3_array_index_2046755_comb] ^ p3_array_index_2046756_comb;
  assign p3_array_index_2046850_comb = p2_literal_2043916[p3_res7__388_comb];
  assign p3_array_index_2046851_comb = p2_literal_2043918[p3_res7__386_comb];
  assign p3_array_index_2046852_comb = p2_literal_2043920[p3_res7__384_comb];
  assign p3_res7__396_comb = p2_literal_2043910[p3_res7__394_comb] ^ p2_literal_2043912[p3_res7__392_comb] ^ p2_literal_2043914[p3_res7__390_comb] ^ p3_array_index_2046850_comb ^ p3_array_index_2046851_comb ^ p3_array_index_2046852_comb ^ p3_array_index_2046746_comb ^ p2_literal_2043923[p3_array_index_2046747_comb] ^ p3_array_index_2046748_comb ^ p3_array_index_2046798_comb ^ p3_array_index_2046766_comb ^ p2_literal_2043916[p3_array_index_2046751_comb] ^ p2_literal_2043914[p3_array_index_2046768_comb] ^ p2_literal_2043912[p3_array_index_2046753_comb] ^ p2_literal_2043910[p3_array_index_2046770_comb] ^ p3_array_index_2046755_comb;
  assign p3_array_index_2046862_comb = p2_literal_2043916[p3_res7__390_comb];
  assign p3_array_index_2046863_comb = p2_literal_2043918[p3_res7__388_comb];
  assign p3_array_index_2046864_comb = p2_literal_2043920[p3_res7__386_comb];
  assign p3_res7__398_comb = p2_literal_2043910[p3_res7__396_comb] ^ p2_literal_2043912[p3_res7__394_comb] ^ p2_literal_2043914[p3_res7__392_comb] ^ p3_array_index_2046862_comb ^ p3_array_index_2046863_comb ^ p3_array_index_2046864_comb ^ p3_res7__384_comb ^ p2_literal_2043923[p3_array_index_2046746_comb] ^ p3_array_index_2046747_comb ^ p3_array_index_2046812_comb ^ p3_array_index_2046783_comb ^ p2_literal_2043916[p3_array_index_2046750_comb] ^ p2_literal_2043914[p3_array_index_2046751_comb] ^ p2_literal_2043912[p3_array_index_2046768_comb] ^ p2_literal_2043910[p3_array_index_2046753_comb] ^ p3_array_index_2046770_comb;
  assign p3_array_index_2046875_comb = p2_literal_2043918[p3_res7__390_comb];
  assign p3_array_index_2046876_comb = p2_literal_2043920[p3_res7__388_comb];
  assign p3_res7__400_comb = p2_literal_2043910[p3_res7__398_comb] ^ p2_literal_2043912[p3_res7__396_comb] ^ p2_literal_2043914[p3_res7__394_comb] ^ p2_literal_2043916[p3_res7__392_comb] ^ p3_array_index_2046875_comb ^ p3_array_index_2046876_comb ^ p3_res7__386_comb ^ p2_literal_2043923[p3_res7__384_comb] ^ p3_array_index_2046746_comb ^ p3_array_index_2046826_comb ^ p3_array_index_2046797_comb ^ p3_array_index_2046765_comb ^ p2_literal_2043914[p3_array_index_2046750_comb] ^ p2_literal_2043912[p3_array_index_2046751_comb] ^ p2_literal_2043910[p3_array_index_2046768_comb] ^ p3_array_index_2046753_comb;
  assign p3_array_index_2046886_comb = p2_literal_2043918[p3_res7__392_comb];
  assign p3_array_index_2046887_comb = p2_literal_2043920[p3_res7__390_comb];
  assign p3_res7__402_comb = p2_literal_2043910[p3_res7__400_comb] ^ p2_literal_2043912[p3_res7__398_comb] ^ p2_literal_2043914[p3_res7__396_comb] ^ p2_literal_2043916[p3_res7__394_comb] ^ p3_array_index_2046886_comb ^ p3_array_index_2046887_comb ^ p3_res7__388_comb ^ p2_literal_2043923[p3_res7__386_comb] ^ p3_res7__384_comb ^ p3_array_index_2046839_comb ^ p3_array_index_2046811_comb ^ p3_array_index_2046782_comb ^ p2_literal_2043914[p3_array_index_2046749_comb] ^ p2_literal_2043912[p3_array_index_2046750_comb] ^ p2_literal_2043910[p3_array_index_2046751_comb] ^ p3_array_index_2046768_comb;
  assign p3_array_index_2046898_comb = p2_literal_2043920[p3_res7__392_comb];
  assign p3_res7__404_comb = p2_literal_2043910[p3_res7__402_comb] ^ p2_literal_2043912[p3_res7__400_comb] ^ p2_literal_2043914[p3_res7__398_comb] ^ p2_literal_2043916[p3_res7__396_comb] ^ p2_literal_2043918[p3_res7__394_comb] ^ p3_array_index_2046898_comb ^ p3_res7__390_comb ^ p2_literal_2043923[p3_res7__388_comb] ^ p3_res7__386_comb ^ p3_array_index_2046852_comb ^ p3_array_index_2046825_comb ^ p3_array_index_2046796_comb ^ p3_array_index_2046764_comb ^ p2_literal_2043912[p3_array_index_2046749_comb] ^ p2_literal_2043910[p3_array_index_2046750_comb] ^ p3_array_index_2046751_comb;
  assign p3_array_index_2046908_comb = p2_literal_2043920[p3_res7__394_comb];
  assign p3_res7__406_comb = p2_literal_2043910[p3_res7__404_comb] ^ p2_literal_2043912[p3_res7__402_comb] ^ p2_literal_2043914[p3_res7__400_comb] ^ p2_literal_2043916[p3_res7__398_comb] ^ p2_literal_2043918[p3_res7__396_comb] ^ p3_array_index_2046908_comb ^ p3_res7__392_comb ^ p2_literal_2043923[p3_res7__390_comb] ^ p3_res7__388_comb ^ p3_array_index_2046864_comb ^ p3_array_index_2046838_comb ^ p3_array_index_2046810_comb ^ p3_array_index_2046781_comb ^ p2_literal_2043912[p3_array_index_2046748_comb] ^ p2_literal_2043910[p3_array_index_2046749_comb] ^ p3_array_index_2046750_comb;
  assign p3_res7__408_comb = p2_literal_2043910[p3_res7__406_comb] ^ p2_literal_2043912[p3_res7__404_comb] ^ p2_literal_2043914[p3_res7__402_comb] ^ p2_literal_2043916[p3_res7__400_comb] ^ p2_literal_2043918[p3_res7__398_comb] ^ p2_literal_2043920[p3_res7__396_comb] ^ p3_res7__394_comb ^ p2_literal_2043923[p3_res7__392_comb] ^ p3_res7__390_comb ^ p3_array_index_2046876_comb ^ p3_array_index_2046851_comb ^ p3_array_index_2046824_comb ^ p3_array_index_2046795_comb ^ p3_array_index_2046763_comb ^ p2_literal_2043910[p3_array_index_2046748_comb] ^ p3_array_index_2046749_comb;
  assign p3_res7__410_comb = p2_literal_2043910[p3_res7__408_comb] ^ p2_literal_2043912[p3_res7__406_comb] ^ p2_literal_2043914[p3_res7__404_comb] ^ p2_literal_2043916[p3_res7__402_comb] ^ p2_literal_2043918[p3_res7__400_comb] ^ p2_literal_2043920[p3_res7__398_comb] ^ p3_res7__396_comb ^ p2_literal_2043923[p3_res7__394_comb] ^ p3_res7__392_comb ^ p3_array_index_2046887_comb ^ p3_array_index_2046863_comb ^ p3_array_index_2046837_comb ^ p3_array_index_2046809_comb ^ p3_array_index_2046780_comb ^ p2_literal_2043910[p3_array_index_2046747_comb] ^ p3_array_index_2046748_comb;
  assign p3_res7__412_comb = p2_literal_2043910[p3_res7__410_comb] ^ p2_literal_2043912[p3_res7__408_comb] ^ p2_literal_2043914[p3_res7__406_comb] ^ p2_literal_2043916[p3_res7__404_comb] ^ p2_literal_2043918[p3_res7__402_comb] ^ p2_literal_2043920[p3_res7__400_comb] ^ p3_res7__398_comb ^ p2_literal_2043923[p3_res7__396_comb] ^ p3_res7__394_comb ^ p3_array_index_2046898_comb ^ p3_array_index_2046875_comb ^ p3_array_index_2046850_comb ^ p3_array_index_2046823_comb ^ p3_array_index_2046794_comb ^ p3_array_index_2046762_comb ^ p3_array_index_2046747_comb;
  assign p3_res7__414_comb = p2_literal_2043910[p3_res7__412_comb] ^ p2_literal_2043912[p3_res7__410_comb] ^ p2_literal_2043914[p3_res7__408_comb] ^ p2_literal_2043916[p3_res7__406_comb] ^ p2_literal_2043918[p3_res7__404_comb] ^ p2_literal_2043920[p3_res7__402_comb] ^ p3_res7__400_comb ^ p2_literal_2043923[p3_res7__398_comb] ^ p3_res7__396_comb ^ p3_array_index_2046908_comb ^ p3_array_index_2046886_comb ^ p3_array_index_2046862_comb ^ p3_array_index_2046836_comb ^ p3_array_index_2046808_comb ^ p3_array_index_2046779_comb ^ p3_array_index_2046746_comb;
  assign p3_res__12_comb = {p3_res7__414_comb, p3_res7__412_comb, p3_res7__410_comb, p3_res7__408_comb, p3_res7__406_comb, p3_res7__404_comb, p3_res7__402_comb, p3_res7__400_comb, p3_res7__398_comb, p3_res7__396_comb, p3_res7__394_comb, p3_res7__392_comb, p3_res7__390_comb, p3_res7__388_comb, p3_res7__386_comb, p3_res7__384_comb};
  assign p3_xor_2046948_comb = p3_res__12_comb ^ p3_xor_2046512_comb;
  assign p3_addedKey__45_comb = p3_xor_2046948_comb ^ 128'h5113_c1f9_4d76_899f_a029_a9e0_ac34_d40e;
  assign p3_array_index_2046964_comb = p2_literal_2043896[p3_addedKey__45_comb[127:120]];
  assign p3_array_index_2046965_comb = p2_literal_2043896[p3_addedKey__45_comb[119:112]];
  assign p3_array_index_2046966_comb = p2_literal_2043896[p3_addedKey__45_comb[111:104]];
  assign p3_array_index_2046967_comb = p2_literal_2043896[p3_addedKey__45_comb[103:96]];
  assign p3_array_index_2046968_comb = p2_literal_2043896[p3_addedKey__45_comb[95:88]];
  assign p3_array_index_2046969_comb = p2_literal_2043896[p3_addedKey__45_comb[87:80]];
  assign p3_array_index_2046971_comb = p2_literal_2043896[p3_addedKey__45_comb[71:64]];
  assign p3_array_index_2046973_comb = p2_literal_2043896[p3_addedKey__45_comb[55:48]];
  assign p3_array_index_2046974_comb = p2_literal_2043896[p3_addedKey__45_comb[47:40]];
  assign p3_array_index_2046975_comb = p2_literal_2043896[p3_addedKey__45_comb[39:32]];
  assign p3_array_index_2046976_comb = p2_literal_2043896[p3_addedKey__45_comb[31:24]];
  assign p3_array_index_2046977_comb = p2_literal_2043896[p3_addedKey__45_comb[23:16]];
  assign p3_array_index_2046978_comb = p2_literal_2043896[p3_addedKey__45_comb[15:8]];
  assign p3_array_index_2046980_comb = p2_literal_2043910[p3_array_index_2046964_comb];
  assign p3_array_index_2046981_comb = p2_literal_2043912[p3_array_index_2046965_comb];
  assign p3_array_index_2046982_comb = p2_literal_2043914[p3_array_index_2046966_comb];
  assign p3_array_index_2046983_comb = p2_literal_2043916[p3_array_index_2046967_comb];
  assign p3_array_index_2046984_comb = p2_literal_2043918[p3_array_index_2046968_comb];
  assign p3_array_index_2046985_comb = p2_literal_2043920[p3_array_index_2046969_comb];
  assign p3_array_index_2046986_comb = p2_literal_2043896[p3_addedKey__45_comb[79:72]];
  assign p3_array_index_2046988_comb = p2_literal_2043896[p3_addedKey__45_comb[63:56]];
  assign p3_res7__416_comb = p3_array_index_2046980_comb ^ p3_array_index_2046981_comb ^ p3_array_index_2046982_comb ^ p3_array_index_2046983_comb ^ p3_array_index_2046984_comb ^ p3_array_index_2046985_comb ^ p3_array_index_2046986_comb ^ p2_literal_2043923[p3_array_index_2046971_comb] ^ p3_array_index_2046988_comb ^ p2_literal_2043920[p3_array_index_2046973_comb] ^ p2_literal_2043918[p3_array_index_2046974_comb] ^ p2_literal_2043916[p3_array_index_2046975_comb] ^ p2_literal_2043914[p3_array_index_2046976_comb] ^ p2_literal_2043912[p3_array_index_2046977_comb] ^ p2_literal_2043910[p3_array_index_2046978_comb] ^ p2_literal_2043896[p3_addedKey__45_comb[7:0]];
  assign p3_array_index_2046997_comb = p2_literal_2043910[p3_res7__416_comb];
  assign p3_array_index_2046998_comb = p2_literal_2043912[p3_array_index_2046964_comb];
  assign p3_array_index_2046999_comb = p2_literal_2043914[p3_array_index_2046965_comb];
  assign p3_array_index_2047000_comb = p2_literal_2043916[p3_array_index_2046966_comb];
  assign p3_array_index_2047001_comb = p2_literal_2043918[p3_array_index_2046967_comb];
  assign p3_array_index_2047002_comb = p2_literal_2043920[p3_array_index_2046968_comb];
  assign p3_res7__418_comb = p3_array_index_2046997_comb ^ p3_array_index_2046998_comb ^ p3_array_index_2046999_comb ^ p3_array_index_2047000_comb ^ p3_array_index_2047001_comb ^ p3_array_index_2047002_comb ^ p3_array_index_2046969_comb ^ p2_literal_2043923[p3_array_index_2046986_comb] ^ p3_array_index_2046971_comb ^ p2_literal_2043920[p3_array_index_2046988_comb] ^ p2_literal_2043918[p3_array_index_2046973_comb] ^ p2_literal_2043916[p3_array_index_2046974_comb] ^ p2_literal_2043914[p3_array_index_2046975_comb] ^ p2_literal_2043912[p3_array_index_2046976_comb] ^ p2_literal_2043910[p3_array_index_2046977_comb] ^ p3_array_index_2046978_comb;
  assign p3_array_index_2047012_comb = p2_literal_2043912[p3_res7__416_comb];
  assign p3_array_index_2047013_comb = p2_literal_2043914[p3_array_index_2046964_comb];
  assign p3_array_index_2047014_comb = p2_literal_2043916[p3_array_index_2046965_comb];
  assign p3_array_index_2047015_comb = p2_literal_2043918[p3_array_index_2046966_comb];
  assign p3_array_index_2047016_comb = p2_literal_2043920[p3_array_index_2046967_comb];
  assign p3_res7__420_comb = p2_literal_2043910[p3_res7__418_comb] ^ p3_array_index_2047012_comb ^ p3_array_index_2047013_comb ^ p3_array_index_2047014_comb ^ p3_array_index_2047015_comb ^ p3_array_index_2047016_comb ^ p3_array_index_2046968_comb ^ p2_literal_2043923[p3_array_index_2046969_comb] ^ p3_array_index_2046986_comb ^ p2_literal_2043920[p3_array_index_2046971_comb] ^ p2_literal_2043918[p3_array_index_2046988_comb] ^ p2_literal_2043916[p3_array_index_2046973_comb] ^ p2_literal_2043914[p3_array_index_2046974_comb] ^ p2_literal_2043912[p3_array_index_2046975_comb] ^ p2_literal_2043910[p3_array_index_2046976_comb] ^ p3_array_index_2046977_comb;
  assign p3_array_index_2047026_comb = p2_literal_2043912[p3_res7__418_comb];
  assign p3_array_index_2047027_comb = p2_literal_2043914[p3_res7__416_comb];
  assign p3_array_index_2047028_comb = p2_literal_2043916[p3_array_index_2046964_comb];
  assign p3_array_index_2047029_comb = p2_literal_2043918[p3_array_index_2046965_comb];
  assign p3_array_index_2047030_comb = p2_literal_2043920[p3_array_index_2046966_comb];
  assign p3_res7__422_comb = p2_literal_2043910[p3_res7__420_comb] ^ p3_array_index_2047026_comb ^ p3_array_index_2047027_comb ^ p3_array_index_2047028_comb ^ p3_array_index_2047029_comb ^ p3_array_index_2047030_comb ^ p3_array_index_2046967_comb ^ p2_literal_2043923[p3_array_index_2046968_comb] ^ p3_array_index_2046969_comb ^ p2_literal_2043920[p3_array_index_2046986_comb] ^ p2_literal_2043918[p3_array_index_2046971_comb] ^ p2_literal_2043916[p3_array_index_2046988_comb] ^ p2_literal_2043914[p3_array_index_2046973_comb] ^ p2_literal_2043912[p3_array_index_2046974_comb] ^ p2_literal_2043910[p3_array_index_2046975_comb] ^ p3_array_index_2046976_comb;
  assign p3_array_index_2047041_comb = p2_literal_2043914[p3_res7__418_comb];
  assign p3_array_index_2047042_comb = p2_literal_2043916[p3_res7__416_comb];
  assign p3_array_index_2047043_comb = p2_literal_2043918[p3_array_index_2046964_comb];
  assign p3_array_index_2047044_comb = p2_literal_2043920[p3_array_index_2046965_comb];
  assign p3_res7__424_comb = p2_literal_2043910[p3_res7__422_comb] ^ p2_literal_2043912[p3_res7__420_comb] ^ p3_array_index_2047041_comb ^ p3_array_index_2047042_comb ^ p3_array_index_2047043_comb ^ p3_array_index_2047044_comb ^ p3_array_index_2046966_comb ^ p2_literal_2043923[p3_array_index_2046967_comb] ^ p3_array_index_2046968_comb ^ p3_array_index_2046985_comb ^ p2_literal_2043918[p3_array_index_2046986_comb] ^ p2_literal_2043916[p3_array_index_2046971_comb] ^ p2_literal_2043914[p3_array_index_2046988_comb] ^ p2_literal_2043912[p3_array_index_2046973_comb] ^ p2_literal_2043910[p3_array_index_2046974_comb] ^ p3_array_index_2046975_comb;

  // Registers for pipe stage 3:
  reg [127:0] p3_encoded;
  reg [127:0] p3_bit_slice_2043893;
  reg [127:0] p3_bit_slice_2044119;
  reg [127:0] p3_k3;
  reg [127:0] p3_k2;
  reg [127:0] p3_xor_2046730;
  reg [127:0] p3_xor_2046948;
  reg [7:0] p3_array_index_2046964;
  reg [7:0] p3_array_index_2046965;
  reg [7:0] p3_array_index_2046966;
  reg [7:0] p3_array_index_2046967;
  reg [7:0] p3_array_index_2046968;
  reg [7:0] p3_array_index_2046969;
  reg [7:0] p3_array_index_2046971;
  reg [7:0] p3_array_index_2046973;
  reg [7:0] p3_array_index_2046974;
  reg [7:0] p3_array_index_2046980;
  reg [7:0] p3_array_index_2046981;
  reg [7:0] p3_array_index_2046982;
  reg [7:0] p3_array_index_2046983;
  reg [7:0] p3_array_index_2046984;
  reg [7:0] p3_array_index_2046986;
  reg [7:0] p3_array_index_2046988;
  reg [7:0] p3_res7__416;
  reg [7:0] p3_array_index_2046997;
  reg [7:0] p3_array_index_2046998;
  reg [7:0] p3_array_index_2046999;
  reg [7:0] p3_array_index_2047000;
  reg [7:0] p3_array_index_2047001;
  reg [7:0] p3_array_index_2047002;
  reg [7:0] p3_res7__418;
  reg [7:0] p3_array_index_2047012;
  reg [7:0] p3_array_index_2047013;
  reg [7:0] p3_array_index_2047014;
  reg [7:0] p3_array_index_2047015;
  reg [7:0] p3_array_index_2047016;
  reg [7:0] p3_res7__420;
  reg [7:0] p3_array_index_2047026;
  reg [7:0] p3_array_index_2047027;
  reg [7:0] p3_array_index_2047028;
  reg [7:0] p3_array_index_2047029;
  reg [7:0] p3_array_index_2047030;
  reg [7:0] p3_res7__422;
  reg [7:0] p3_array_index_2047041;
  reg [7:0] p3_array_index_2047042;
  reg [7:0] p3_array_index_2047043;
  reg [7:0] p3_array_index_2047044;
  reg [7:0] p3_res7__424;
  reg [7:0] p4_literal_2043896[256];
  reg [7:0] p4_literal_2043910[256];
  reg [7:0] p4_literal_2043912[256];
  reg [7:0] p4_literal_2043914[256];
  reg [7:0] p4_literal_2043916[256];
  reg [7:0] p4_literal_2043918[256];
  reg [7:0] p4_literal_2043920[256];
  reg [7:0] p4_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p3_encoded <= p2_encoded;
    p3_bit_slice_2043893 <= p2_bit_slice_2043893;
    p3_bit_slice_2044119 <= p2_bit_slice_2044119;
    p3_k3 <= p2_k3;
    p3_k2 <= p2_k2;
    p3_xor_2046730 <= p3_xor_2046730_comb;
    p3_xor_2046948 <= p3_xor_2046948_comb;
    p3_array_index_2046964 <= p3_array_index_2046964_comb;
    p3_array_index_2046965 <= p3_array_index_2046965_comb;
    p3_array_index_2046966 <= p3_array_index_2046966_comb;
    p3_array_index_2046967 <= p3_array_index_2046967_comb;
    p3_array_index_2046968 <= p3_array_index_2046968_comb;
    p3_array_index_2046969 <= p3_array_index_2046969_comb;
    p3_array_index_2046971 <= p3_array_index_2046971_comb;
    p3_array_index_2046973 <= p3_array_index_2046973_comb;
    p3_array_index_2046974 <= p3_array_index_2046974_comb;
    p3_array_index_2046980 <= p3_array_index_2046980_comb;
    p3_array_index_2046981 <= p3_array_index_2046981_comb;
    p3_array_index_2046982 <= p3_array_index_2046982_comb;
    p3_array_index_2046983 <= p3_array_index_2046983_comb;
    p3_array_index_2046984 <= p3_array_index_2046984_comb;
    p3_array_index_2046986 <= p3_array_index_2046986_comb;
    p3_array_index_2046988 <= p3_array_index_2046988_comb;
    p3_res7__416 <= p3_res7__416_comb;
    p3_array_index_2046997 <= p3_array_index_2046997_comb;
    p3_array_index_2046998 <= p3_array_index_2046998_comb;
    p3_array_index_2046999 <= p3_array_index_2046999_comb;
    p3_array_index_2047000 <= p3_array_index_2047000_comb;
    p3_array_index_2047001 <= p3_array_index_2047001_comb;
    p3_array_index_2047002 <= p3_array_index_2047002_comb;
    p3_res7__418 <= p3_res7__418_comb;
    p3_array_index_2047012 <= p3_array_index_2047012_comb;
    p3_array_index_2047013 <= p3_array_index_2047013_comb;
    p3_array_index_2047014 <= p3_array_index_2047014_comb;
    p3_array_index_2047015 <= p3_array_index_2047015_comb;
    p3_array_index_2047016 <= p3_array_index_2047016_comb;
    p3_res7__420 <= p3_res7__420_comb;
    p3_array_index_2047026 <= p3_array_index_2047026_comb;
    p3_array_index_2047027 <= p3_array_index_2047027_comb;
    p3_array_index_2047028 <= p3_array_index_2047028_comb;
    p3_array_index_2047029 <= p3_array_index_2047029_comb;
    p3_array_index_2047030 <= p3_array_index_2047030_comb;
    p3_res7__422 <= p3_res7__422_comb;
    p3_array_index_2047041 <= p3_array_index_2047041_comb;
    p3_array_index_2047042 <= p3_array_index_2047042_comb;
    p3_array_index_2047043 <= p3_array_index_2047043_comb;
    p3_array_index_2047044 <= p3_array_index_2047044_comb;
    p3_res7__424 <= p3_res7__424_comb;
    p4_literal_2043896 <= p3_literal_2043896;
    p4_literal_2043910 <= p3_literal_2043910;
    p4_literal_2043912 <= p3_literal_2043912;
    p4_literal_2043914 <= p3_literal_2043914;
    p4_literal_2043916 <= p3_literal_2043916;
    p4_literal_2043918 <= p3_literal_2043918;
    p4_literal_2043920 <= p3_literal_2043920;
    p4_literal_2043923 <= p3_literal_2043923;
  end

  // ===== Pipe stage 4:
  wire [7:0] p4_array_index_2047166_comb;
  wire [7:0] p4_array_index_2047167_comb;
  wire [7:0] p4_array_index_2047168_comb;
  wire [7:0] p4_array_index_2047169_comb;
  wire [7:0] p4_res7__426_comb;
  wire [7:0] p4_array_index_2047180_comb;
  wire [7:0] p4_array_index_2047181_comb;
  wire [7:0] p4_array_index_2047182_comb;
  wire [7:0] p4_res7__428_comb;
  wire [7:0] p4_array_index_2047192_comb;
  wire [7:0] p4_array_index_2047193_comb;
  wire [7:0] p4_array_index_2047194_comb;
  wire [7:0] p4_res7__430_comb;
  wire [7:0] p4_array_index_2047205_comb;
  wire [7:0] p4_array_index_2047206_comb;
  wire [7:0] p4_res7__432_comb;
  wire [7:0] p4_array_index_2047216_comb;
  wire [7:0] p4_array_index_2047217_comb;
  wire [7:0] p4_res7__434_comb;
  wire [7:0] p4_array_index_2047228_comb;
  wire [7:0] p4_res7__436_comb;
  wire [7:0] p4_array_index_2047238_comb;
  wire [7:0] p4_res7__438_comb;
  wire [7:0] p4_res7__440_comb;
  wire [7:0] p4_res7__442_comb;
  wire [7:0] p4_res7__444_comb;
  wire [7:0] p4_res7__446_comb;
  wire [127:0] p4_res__13_comb;
  wire [127:0] p4_xor_2047278_comb;
  wire [127:0] p4_addedKey__46_comb;
  wire [7:0] p4_array_index_2047294_comb;
  wire [7:0] p4_array_index_2047295_comb;
  wire [7:0] p4_array_index_2047296_comb;
  wire [7:0] p4_array_index_2047297_comb;
  wire [7:0] p4_array_index_2047298_comb;
  wire [7:0] p4_array_index_2047299_comb;
  wire [7:0] p4_array_index_2047301_comb;
  wire [7:0] p4_array_index_2047303_comb;
  wire [7:0] p4_array_index_2047304_comb;
  wire [7:0] p4_array_index_2047305_comb;
  wire [7:0] p4_array_index_2047306_comb;
  wire [7:0] p4_array_index_2047307_comb;
  wire [7:0] p4_array_index_2047308_comb;
  wire [7:0] p4_array_index_2047310_comb;
  wire [7:0] p4_array_index_2047311_comb;
  wire [7:0] p4_array_index_2047312_comb;
  wire [7:0] p4_array_index_2047313_comb;
  wire [7:0] p4_array_index_2047314_comb;
  wire [7:0] p4_array_index_2047315_comb;
  wire [7:0] p4_array_index_2047316_comb;
  wire [7:0] p4_array_index_2047318_comb;
  wire [7:0] p4_res7__448_comb;
  wire [7:0] p4_array_index_2047327_comb;
  wire [7:0] p4_array_index_2047328_comb;
  wire [7:0] p4_array_index_2047329_comb;
  wire [7:0] p4_array_index_2047330_comb;
  wire [7:0] p4_array_index_2047331_comb;
  wire [7:0] p4_array_index_2047332_comb;
  wire [7:0] p4_res7__450_comb;
  wire [7:0] p4_array_index_2047342_comb;
  wire [7:0] p4_array_index_2047343_comb;
  wire [7:0] p4_array_index_2047344_comb;
  wire [7:0] p4_array_index_2047345_comb;
  wire [7:0] p4_array_index_2047346_comb;
  wire [7:0] p4_res7__452_comb;
  wire [7:0] p4_array_index_2047356_comb;
  wire [7:0] p4_array_index_2047357_comb;
  wire [7:0] p4_array_index_2047358_comb;
  wire [7:0] p4_array_index_2047359_comb;
  wire [7:0] p4_array_index_2047360_comb;
  wire [7:0] p4_res7__454_comb;
  wire [7:0] p4_array_index_2047371_comb;
  wire [7:0] p4_array_index_2047372_comb;
  wire [7:0] p4_array_index_2047373_comb;
  wire [7:0] p4_array_index_2047374_comb;
  wire [7:0] p4_res7__456_comb;
  wire [7:0] p4_array_index_2047384_comb;
  wire [7:0] p4_array_index_2047385_comb;
  wire [7:0] p4_array_index_2047386_comb;
  wire [7:0] p4_array_index_2047387_comb;
  wire [7:0] p4_res7__458_comb;
  wire [7:0] p4_array_index_2047398_comb;
  wire [7:0] p4_array_index_2047399_comb;
  wire [7:0] p4_array_index_2047400_comb;
  wire [7:0] p4_res7__460_comb;
  wire [7:0] p4_array_index_2047410_comb;
  wire [7:0] p4_array_index_2047411_comb;
  wire [7:0] p4_array_index_2047412_comb;
  wire [7:0] p4_res7__462_comb;
  wire [7:0] p4_array_index_2047423_comb;
  wire [7:0] p4_array_index_2047424_comb;
  wire [7:0] p4_res7__464_comb;
  wire [7:0] p4_array_index_2047434_comb;
  wire [7:0] p4_array_index_2047435_comb;
  wire [7:0] p4_res7__466_comb;
  wire [7:0] p4_array_index_2047446_comb;
  wire [7:0] p4_res7__468_comb;
  wire [7:0] p4_array_index_2047456_comb;
  wire [7:0] p4_res7__470_comb;
  wire [7:0] p4_res7__472_comb;
  wire [7:0] p4_res7__474_comb;
  wire [7:0] p4_res7__476_comb;
  wire [7:0] p4_res7__478_comb;
  wire [127:0] p4_res__14_comb;
  wire [127:0] p4_k5_comb;
  wire [127:0] p4_addedKey__47_comb;
  wire [7:0] p4_array_index_2047512_comb;
  wire [7:0] p4_array_index_2047513_comb;
  wire [7:0] p4_array_index_2047514_comb;
  wire [7:0] p4_array_index_2047515_comb;
  wire [7:0] p4_array_index_2047516_comb;
  wire [7:0] p4_array_index_2047517_comb;
  wire [7:0] p4_array_index_2047519_comb;
  wire [7:0] p4_array_index_2047521_comb;
  wire [7:0] p4_array_index_2047522_comb;
  wire [7:0] p4_array_index_2047523_comb;
  wire [7:0] p4_array_index_2047524_comb;
  wire [7:0] p4_array_index_2047525_comb;
  wire [7:0] p4_array_index_2047526_comb;
  wire [7:0] p4_array_index_2047528_comb;
  wire [7:0] p4_array_index_2047529_comb;
  wire [7:0] p4_array_index_2047530_comb;
  wire [7:0] p4_array_index_2047531_comb;
  wire [7:0] p4_array_index_2047532_comb;
  wire [7:0] p4_array_index_2047533_comb;
  wire [7:0] p4_array_index_2047534_comb;
  wire [7:0] p4_array_index_2047536_comb;
  wire [7:0] p4_res7__480_comb;
  wire [7:0] p4_array_index_2047545_comb;
  wire [7:0] p4_array_index_2047546_comb;
  wire [7:0] p4_array_index_2047547_comb;
  wire [7:0] p4_array_index_2047548_comb;
  wire [7:0] p4_array_index_2047549_comb;
  wire [7:0] p4_array_index_2047550_comb;
  wire [7:0] p4_res7__482_comb;
  wire [7:0] p4_array_index_2047560_comb;
  wire [7:0] p4_array_index_2047561_comb;
  wire [7:0] p4_array_index_2047562_comb;
  wire [7:0] p4_array_index_2047563_comb;
  wire [7:0] p4_array_index_2047564_comb;
  wire [7:0] p4_res7__484_comb;
  wire [7:0] p4_array_index_2047574_comb;
  wire [7:0] p4_array_index_2047575_comb;
  wire [7:0] p4_array_index_2047576_comb;
  wire [7:0] p4_array_index_2047577_comb;
  wire [7:0] p4_array_index_2047578_comb;
  wire [7:0] p4_res7__486_comb;
  wire [7:0] p4_array_index_2047589_comb;
  wire [7:0] p4_array_index_2047590_comb;
  wire [7:0] p4_array_index_2047591_comb;
  wire [7:0] p4_array_index_2047592_comb;
  wire [7:0] p4_res7__488_comb;
  wire [7:0] p4_array_index_2047602_comb;
  wire [7:0] p4_array_index_2047603_comb;
  wire [7:0] p4_array_index_2047604_comb;
  wire [7:0] p4_array_index_2047605_comb;
  wire [7:0] p4_res7__490_comb;
  wire [7:0] p4_array_index_2047616_comb;
  wire [7:0] p4_array_index_2047617_comb;
  wire [7:0] p4_array_index_2047618_comb;
  wire [7:0] p4_res7__492_comb;
  wire [7:0] p4_array_index_2047628_comb;
  wire [7:0] p4_array_index_2047629_comb;
  wire [7:0] p4_array_index_2047630_comb;
  wire [7:0] p4_res7__494_comb;
  wire [7:0] p4_array_index_2047641_comb;
  wire [7:0] p4_array_index_2047642_comb;
  wire [7:0] p4_res7__496_comb;
  wire [7:0] p4_array_index_2047652_comb;
  wire [7:0] p4_array_index_2047653_comb;
  wire [7:0] p4_res7__498_comb;
  wire [7:0] p4_array_index_2047664_comb;
  wire [7:0] p4_res7__500_comb;
  wire [7:0] p4_array_index_2047674_comb;
  wire [7:0] p4_res7__502_comb;
  wire [7:0] p4_res7__504_comb;
  wire [7:0] p4_res7__506_comb;
  wire [7:0] p4_res7__508_comb;
  wire [7:0] p4_res7__510_comb;
  wire [127:0] p4_res__15_comb;
  wire [127:0] p4_k4_comb;
  wire [127:0] p4_addedKey__48_comb;
  wire [7:0] p4_array_index_2047730_comb;
  wire [7:0] p4_array_index_2047731_comb;
  wire [7:0] p4_array_index_2047732_comb;
  wire [7:0] p4_array_index_2047733_comb;
  wire [7:0] p4_array_index_2047734_comb;
  wire [7:0] p4_array_index_2047735_comb;
  wire [7:0] p4_array_index_2047737_comb;
  wire [7:0] p4_array_index_2047739_comb;
  wire [7:0] p4_array_index_2047740_comb;
  wire [7:0] p4_array_index_2047741_comb;
  wire [7:0] p4_array_index_2047742_comb;
  wire [7:0] p4_array_index_2047743_comb;
  wire [7:0] p4_array_index_2047744_comb;
  wire [7:0] p4_array_index_2047746_comb;
  wire [7:0] p4_array_index_2047747_comb;
  wire [7:0] p4_array_index_2047748_comb;
  wire [7:0] p4_array_index_2047749_comb;
  wire [7:0] p4_array_index_2047750_comb;
  wire [7:0] p4_array_index_2047751_comb;
  wire [7:0] p4_array_index_2047752_comb;
  wire [7:0] p4_array_index_2047754_comb;
  wire [7:0] p4_res7__512_comb;
  wire [7:0] p4_array_index_2047763_comb;
  wire [7:0] p4_array_index_2047764_comb;
  wire [7:0] p4_array_index_2047765_comb;
  wire [7:0] p4_array_index_2047766_comb;
  wire [7:0] p4_array_index_2047767_comb;
  wire [7:0] p4_array_index_2047768_comb;
  wire [7:0] p4_res7__514_comb;
  wire [7:0] p4_array_index_2047778_comb;
  wire [7:0] p4_array_index_2047779_comb;
  wire [7:0] p4_array_index_2047780_comb;
  wire [7:0] p4_array_index_2047781_comb;
  wire [7:0] p4_array_index_2047782_comb;
  wire [7:0] p4_res7__516_comb;
  wire [7:0] p4_array_index_2047792_comb;
  wire [7:0] p4_array_index_2047793_comb;
  wire [7:0] p4_array_index_2047794_comb;
  wire [7:0] p4_array_index_2047795_comb;
  wire [7:0] p4_array_index_2047796_comb;
  wire [7:0] p4_res7__518_comb;
  wire [7:0] p4_array_index_2047807_comb;
  wire [7:0] p4_array_index_2047808_comb;
  wire [7:0] p4_array_index_2047809_comb;
  wire [7:0] p4_array_index_2047810_comb;
  wire [7:0] p4_res7__520_comb;
  wire [7:0] p4_array_index_2047820_comb;
  wire [7:0] p4_array_index_2047821_comb;
  wire [7:0] p4_array_index_2047822_comb;
  wire [7:0] p4_array_index_2047823_comb;
  wire [7:0] p4_res7__522_comb;
  wire [7:0] p4_array_index_2047834_comb;
  wire [7:0] p4_array_index_2047835_comb;
  wire [7:0] p4_array_index_2047836_comb;
  wire [7:0] p4_res7__524_comb;
  wire [7:0] p4_array_index_2047846_comb;
  wire [7:0] p4_array_index_2047847_comb;
  wire [7:0] p4_array_index_2047848_comb;
  wire [7:0] p4_res7__526_comb;
  wire [7:0] p4_array_index_2047859_comb;
  wire [7:0] p4_array_index_2047860_comb;
  wire [7:0] p4_res7__528_comb;
  wire [7:0] p4_array_index_2047870_comb;
  wire [7:0] p4_array_index_2047871_comb;
  wire [7:0] p4_res7__530_comb;
  wire [7:0] p4_array_index_2047882_comb;
  wire [7:0] p4_res7__532_comb;
  wire [7:0] p4_array_index_2047892_comb;
  wire [7:0] p4_res7__534_comb;
  wire [7:0] p4_res7__536_comb;
  wire [7:0] p4_res7__538_comb;
  wire [7:0] p4_res7__540_comb;
  wire [7:0] p4_res7__542_comb;
  wire [127:0] p4_res__16_comb;
  wire [127:0] p4_xor_2047932_comb;
  wire [127:0] p4_addedKey__49_comb;
  wire [7:0] p4_array_index_2047948_comb;
  wire [7:0] p4_array_index_2047949_comb;
  wire [7:0] p4_array_index_2047950_comb;
  wire [7:0] p4_array_index_2047951_comb;
  wire [7:0] p4_array_index_2047952_comb;
  wire [7:0] p4_array_index_2047953_comb;
  wire [7:0] p4_array_index_2047955_comb;
  wire [7:0] p4_array_index_2047957_comb;
  wire [7:0] p4_array_index_2047958_comb;
  wire [7:0] p4_array_index_2047959_comb;
  wire [7:0] p4_array_index_2047960_comb;
  wire [7:0] p4_array_index_2047961_comb;
  wire [7:0] p4_array_index_2047962_comb;
  wire [7:0] p4_array_index_2047964_comb;
  wire [7:0] p4_array_index_2047965_comb;
  wire [7:0] p4_array_index_2047966_comb;
  wire [7:0] p4_array_index_2047967_comb;
  wire [7:0] p4_array_index_2047968_comb;
  wire [7:0] p4_array_index_2047969_comb;
  wire [7:0] p4_array_index_2047970_comb;
  wire [7:0] p4_array_index_2047972_comb;
  wire [7:0] p4_res7__544_comb;
  wire [7:0] p4_array_index_2047981_comb;
  wire [7:0] p4_array_index_2047982_comb;
  wire [7:0] p4_array_index_2047983_comb;
  wire [7:0] p4_array_index_2047984_comb;
  wire [7:0] p4_array_index_2047985_comb;
  wire [7:0] p4_array_index_2047986_comb;
  wire [7:0] p4_res7__546_comb;
  wire [7:0] p4_array_index_2047996_comb;
  wire [7:0] p4_array_index_2047997_comb;
  wire [7:0] p4_array_index_2047998_comb;
  wire [7:0] p4_array_index_2047999_comb;
  wire [7:0] p4_array_index_2048000_comb;
  wire [7:0] p4_res7__548_comb;
  wire [7:0] p4_array_index_2048010_comb;
  wire [7:0] p4_array_index_2048011_comb;
  wire [7:0] p4_array_index_2048012_comb;
  wire [7:0] p4_array_index_2048013_comb;
  wire [7:0] p4_array_index_2048014_comb;
  wire [7:0] p4_res7__550_comb;
  wire [7:0] p4_array_index_2048025_comb;
  wire [7:0] p4_array_index_2048026_comb;
  wire [7:0] p4_array_index_2048027_comb;
  wire [7:0] p4_array_index_2048028_comb;
  wire [7:0] p4_res7__552_comb;
  wire [7:0] p4_array_index_2048038_comb;
  wire [7:0] p4_array_index_2048039_comb;
  wire [7:0] p4_array_index_2048040_comb;
  wire [7:0] p4_array_index_2048041_comb;
  wire [7:0] p4_res7__554_comb;
  wire [7:0] p4_array_index_2048052_comb;
  wire [7:0] p4_array_index_2048053_comb;
  wire [7:0] p4_array_index_2048054_comb;
  wire [7:0] p4_res7__556_comb;
  wire [7:0] p4_array_index_2048064_comb;
  wire [7:0] p4_array_index_2048065_comb;
  wire [7:0] p4_array_index_2048066_comb;
  wire [7:0] p4_res7__558_comb;
  wire [7:0] p4_array_index_2048077_comb;
  wire [7:0] p4_array_index_2048078_comb;
  wire [7:0] p4_res7__560_comb;
  wire [7:0] p4_array_index_2048088_comb;
  wire [7:0] p4_array_index_2048089_comb;
  wire [7:0] p4_res7__562_comb;
  wire [7:0] p4_array_index_2048100_comb;
  wire [7:0] p4_res7__564_comb;
  wire [7:0] p4_array_index_2048110_comb;
  wire [7:0] p4_res7__566_comb;
  wire [7:0] p4_array_index_2048115_comb;
  wire [7:0] p4_array_index_2048116_comb;
  wire [7:0] p4_array_index_2048117_comb;
  wire [7:0] p4_array_index_2048118_comb;
  wire [7:0] p4_array_index_2048119_comb;
  wire [7:0] p4_array_index_2048120_comb;
  wire [7:0] p4_array_index_2048121_comb;
  wire [7:0] p4_array_index_2048122_comb;
  assign p4_array_index_2047166_comb = p3_literal_2043914[p3_res7__420];
  assign p4_array_index_2047167_comb = p3_literal_2043916[p3_res7__418];
  assign p4_array_index_2047168_comb = p3_literal_2043918[p3_res7__416];
  assign p4_array_index_2047169_comb = p3_literal_2043920[p3_array_index_2046964];
  assign p4_res7__426_comb = p3_literal_2043910[p3_res7__424] ^ p3_literal_2043912[p3_res7__422] ^ p4_array_index_2047166_comb ^ p4_array_index_2047167_comb ^ p4_array_index_2047168_comb ^ p4_array_index_2047169_comb ^ p3_array_index_2046965 ^ p3_literal_2043923[p3_array_index_2046966] ^ p3_array_index_2046967 ^ p3_array_index_2047002 ^ p3_literal_2043918[p3_array_index_2046969] ^ p3_literal_2043916[p3_array_index_2046986] ^ p3_literal_2043914[p3_array_index_2046971] ^ p3_literal_2043912[p3_array_index_2046988] ^ p3_literal_2043910[p3_array_index_2046973] ^ p3_array_index_2046974;
  assign p4_array_index_2047180_comb = p3_literal_2043916[p3_res7__420];
  assign p4_array_index_2047181_comb = p3_literal_2043918[p3_res7__418];
  assign p4_array_index_2047182_comb = p3_literal_2043920[p3_res7__416];
  assign p4_res7__428_comb = p3_literal_2043910[p4_res7__426_comb] ^ p3_literal_2043912[p3_res7__424] ^ p3_literal_2043914[p3_res7__422] ^ p4_array_index_2047180_comb ^ p4_array_index_2047181_comb ^ p4_array_index_2047182_comb ^ p3_array_index_2046964 ^ p3_literal_2043923[p3_array_index_2046965] ^ p3_array_index_2046966 ^ p3_array_index_2047016 ^ p3_array_index_2046984 ^ p3_literal_2043916[p3_array_index_2046969] ^ p3_literal_2043914[p3_array_index_2046986] ^ p3_literal_2043912[p3_array_index_2046971] ^ p3_literal_2043910[p3_array_index_2046988] ^ p3_array_index_2046973;
  assign p4_array_index_2047192_comb = p3_literal_2043916[p3_res7__422];
  assign p4_array_index_2047193_comb = p3_literal_2043918[p3_res7__420];
  assign p4_array_index_2047194_comb = p3_literal_2043920[p3_res7__418];
  assign p4_res7__430_comb = p3_literal_2043910[p4_res7__428_comb] ^ p3_literal_2043912[p4_res7__426_comb] ^ p3_literal_2043914[p3_res7__424] ^ p4_array_index_2047192_comb ^ p4_array_index_2047193_comb ^ p4_array_index_2047194_comb ^ p3_res7__416 ^ p3_literal_2043923[p3_array_index_2046964] ^ p3_array_index_2046965 ^ p3_array_index_2047030 ^ p3_array_index_2047001 ^ p3_literal_2043916[p3_array_index_2046968] ^ p3_literal_2043914[p3_array_index_2046969] ^ p3_literal_2043912[p3_array_index_2046986] ^ p3_literal_2043910[p3_array_index_2046971] ^ p3_array_index_2046988;
  assign p4_array_index_2047205_comb = p3_literal_2043918[p3_res7__422];
  assign p4_array_index_2047206_comb = p3_literal_2043920[p3_res7__420];
  assign p4_res7__432_comb = p3_literal_2043910[p4_res7__430_comb] ^ p3_literal_2043912[p4_res7__428_comb] ^ p3_literal_2043914[p4_res7__426_comb] ^ p3_literal_2043916[p3_res7__424] ^ p4_array_index_2047205_comb ^ p4_array_index_2047206_comb ^ p3_res7__418 ^ p3_literal_2043923[p3_res7__416] ^ p3_array_index_2046964 ^ p3_array_index_2047044 ^ p3_array_index_2047015 ^ p3_array_index_2046983 ^ p3_literal_2043914[p3_array_index_2046968] ^ p3_literal_2043912[p3_array_index_2046969] ^ p3_literal_2043910[p3_array_index_2046986] ^ p3_array_index_2046971;
  assign p4_array_index_2047216_comb = p3_literal_2043918[p3_res7__424];
  assign p4_array_index_2047217_comb = p3_literal_2043920[p3_res7__422];
  assign p4_res7__434_comb = p3_literal_2043910[p4_res7__432_comb] ^ p3_literal_2043912[p4_res7__430_comb] ^ p3_literal_2043914[p4_res7__428_comb] ^ p3_literal_2043916[p4_res7__426_comb] ^ p4_array_index_2047216_comb ^ p4_array_index_2047217_comb ^ p3_res7__420 ^ p3_literal_2043923[p3_res7__418] ^ p3_res7__416 ^ p4_array_index_2047169_comb ^ p3_array_index_2047029 ^ p3_array_index_2047000 ^ p3_literal_2043914[p3_array_index_2046967] ^ p3_literal_2043912[p3_array_index_2046968] ^ p3_literal_2043910[p3_array_index_2046969] ^ p3_array_index_2046986;
  assign p4_array_index_2047228_comb = p3_literal_2043920[p3_res7__424];
  assign p4_res7__436_comb = p3_literal_2043910[p4_res7__434_comb] ^ p3_literal_2043912[p4_res7__432_comb] ^ p3_literal_2043914[p4_res7__430_comb] ^ p3_literal_2043916[p4_res7__428_comb] ^ p3_literal_2043918[p4_res7__426_comb] ^ p4_array_index_2047228_comb ^ p3_res7__422 ^ p3_literal_2043923[p3_res7__420] ^ p3_res7__418 ^ p4_array_index_2047182_comb ^ p3_array_index_2047043 ^ p3_array_index_2047014 ^ p3_array_index_2046982 ^ p3_literal_2043912[p3_array_index_2046967] ^ p3_literal_2043910[p3_array_index_2046968] ^ p3_array_index_2046969;
  assign p4_array_index_2047238_comb = p3_literal_2043920[p4_res7__426_comb];
  assign p4_res7__438_comb = p3_literal_2043910[p4_res7__436_comb] ^ p3_literal_2043912[p4_res7__434_comb] ^ p3_literal_2043914[p4_res7__432_comb] ^ p3_literal_2043916[p4_res7__430_comb] ^ p3_literal_2043918[p4_res7__428_comb] ^ p4_array_index_2047238_comb ^ p3_res7__424 ^ p3_literal_2043923[p3_res7__422] ^ p3_res7__420 ^ p4_array_index_2047194_comb ^ p4_array_index_2047168_comb ^ p3_array_index_2047028 ^ p3_array_index_2046999 ^ p3_literal_2043912[p3_array_index_2046966] ^ p3_literal_2043910[p3_array_index_2046967] ^ p3_array_index_2046968;
  assign p4_res7__440_comb = p3_literal_2043910[p4_res7__438_comb] ^ p3_literal_2043912[p4_res7__436_comb] ^ p3_literal_2043914[p4_res7__434_comb] ^ p3_literal_2043916[p4_res7__432_comb] ^ p3_literal_2043918[p4_res7__430_comb] ^ p3_literal_2043920[p4_res7__428_comb] ^ p4_res7__426_comb ^ p3_literal_2043923[p3_res7__424] ^ p3_res7__422 ^ p4_array_index_2047206_comb ^ p4_array_index_2047181_comb ^ p3_array_index_2047042 ^ p3_array_index_2047013 ^ p3_array_index_2046981 ^ p3_literal_2043910[p3_array_index_2046966] ^ p3_array_index_2046967;
  assign p4_res7__442_comb = p3_literal_2043910[p4_res7__440_comb] ^ p3_literal_2043912[p4_res7__438_comb] ^ p3_literal_2043914[p4_res7__436_comb] ^ p3_literal_2043916[p4_res7__434_comb] ^ p3_literal_2043918[p4_res7__432_comb] ^ p3_literal_2043920[p4_res7__430_comb] ^ p4_res7__428_comb ^ p3_literal_2043923[p4_res7__426_comb] ^ p3_res7__424 ^ p4_array_index_2047217_comb ^ p4_array_index_2047193_comb ^ p4_array_index_2047167_comb ^ p3_array_index_2047027 ^ p3_array_index_2046998 ^ p3_literal_2043910[p3_array_index_2046965] ^ p3_array_index_2046966;
  assign p4_res7__444_comb = p3_literal_2043910[p4_res7__442_comb] ^ p3_literal_2043912[p4_res7__440_comb] ^ p3_literal_2043914[p4_res7__438_comb] ^ p3_literal_2043916[p4_res7__436_comb] ^ p3_literal_2043918[p4_res7__434_comb] ^ p3_literal_2043920[p4_res7__432_comb] ^ p4_res7__430_comb ^ p3_literal_2043923[p4_res7__428_comb] ^ p4_res7__426_comb ^ p4_array_index_2047228_comb ^ p4_array_index_2047205_comb ^ p4_array_index_2047180_comb ^ p3_array_index_2047041 ^ p3_array_index_2047012 ^ p3_array_index_2046980 ^ p3_array_index_2046965;
  assign p4_res7__446_comb = p3_literal_2043910[p4_res7__444_comb] ^ p3_literal_2043912[p4_res7__442_comb] ^ p3_literal_2043914[p4_res7__440_comb] ^ p3_literal_2043916[p4_res7__438_comb] ^ p3_literal_2043918[p4_res7__436_comb] ^ p3_literal_2043920[p4_res7__434_comb] ^ p4_res7__432_comb ^ p3_literal_2043923[p4_res7__430_comb] ^ p4_res7__428_comb ^ p4_array_index_2047238_comb ^ p4_array_index_2047216_comb ^ p4_array_index_2047192_comb ^ p4_array_index_2047166_comb ^ p3_array_index_2047026 ^ p3_array_index_2046997 ^ p3_array_index_2046964;
  assign p4_res__13_comb = {p4_res7__446_comb, p4_res7__444_comb, p4_res7__442_comb, p4_res7__440_comb, p4_res7__438_comb, p4_res7__436_comb, p4_res7__434_comb, p4_res7__432_comb, p4_res7__430_comb, p4_res7__428_comb, p4_res7__426_comb, p3_res7__424, p3_res7__422, p3_res7__420, p3_res7__418, p3_res7__416};
  assign p4_xor_2047278_comb = p4_res__13_comb ^ p3_xor_2046730;
  assign p4_addedKey__46_comb = p4_xor_2047278_comb ^ 128'h3fb1_b78b_213e_f327_fd0e_14f0_71b0_400f;
  assign p4_array_index_2047294_comb = p3_literal_2043896[p4_addedKey__46_comb[127:120]];
  assign p4_array_index_2047295_comb = p3_literal_2043896[p4_addedKey__46_comb[119:112]];
  assign p4_array_index_2047296_comb = p3_literal_2043896[p4_addedKey__46_comb[111:104]];
  assign p4_array_index_2047297_comb = p3_literal_2043896[p4_addedKey__46_comb[103:96]];
  assign p4_array_index_2047298_comb = p3_literal_2043896[p4_addedKey__46_comb[95:88]];
  assign p4_array_index_2047299_comb = p3_literal_2043896[p4_addedKey__46_comb[87:80]];
  assign p4_array_index_2047301_comb = p3_literal_2043896[p4_addedKey__46_comb[71:64]];
  assign p4_array_index_2047303_comb = p3_literal_2043896[p4_addedKey__46_comb[55:48]];
  assign p4_array_index_2047304_comb = p3_literal_2043896[p4_addedKey__46_comb[47:40]];
  assign p4_array_index_2047305_comb = p3_literal_2043896[p4_addedKey__46_comb[39:32]];
  assign p4_array_index_2047306_comb = p3_literal_2043896[p4_addedKey__46_comb[31:24]];
  assign p4_array_index_2047307_comb = p3_literal_2043896[p4_addedKey__46_comb[23:16]];
  assign p4_array_index_2047308_comb = p3_literal_2043896[p4_addedKey__46_comb[15:8]];
  assign p4_array_index_2047310_comb = p3_literal_2043910[p4_array_index_2047294_comb];
  assign p4_array_index_2047311_comb = p3_literal_2043912[p4_array_index_2047295_comb];
  assign p4_array_index_2047312_comb = p3_literal_2043914[p4_array_index_2047296_comb];
  assign p4_array_index_2047313_comb = p3_literal_2043916[p4_array_index_2047297_comb];
  assign p4_array_index_2047314_comb = p3_literal_2043918[p4_array_index_2047298_comb];
  assign p4_array_index_2047315_comb = p3_literal_2043920[p4_array_index_2047299_comb];
  assign p4_array_index_2047316_comb = p3_literal_2043896[p4_addedKey__46_comb[79:72]];
  assign p4_array_index_2047318_comb = p3_literal_2043896[p4_addedKey__46_comb[63:56]];
  assign p4_res7__448_comb = p4_array_index_2047310_comb ^ p4_array_index_2047311_comb ^ p4_array_index_2047312_comb ^ p4_array_index_2047313_comb ^ p4_array_index_2047314_comb ^ p4_array_index_2047315_comb ^ p4_array_index_2047316_comb ^ p3_literal_2043923[p4_array_index_2047301_comb] ^ p4_array_index_2047318_comb ^ p3_literal_2043920[p4_array_index_2047303_comb] ^ p3_literal_2043918[p4_array_index_2047304_comb] ^ p3_literal_2043916[p4_array_index_2047305_comb] ^ p3_literal_2043914[p4_array_index_2047306_comb] ^ p3_literal_2043912[p4_array_index_2047307_comb] ^ p3_literal_2043910[p4_array_index_2047308_comb] ^ p3_literal_2043896[p4_addedKey__46_comb[7:0]];
  assign p4_array_index_2047327_comb = p3_literal_2043910[p4_res7__448_comb];
  assign p4_array_index_2047328_comb = p3_literal_2043912[p4_array_index_2047294_comb];
  assign p4_array_index_2047329_comb = p3_literal_2043914[p4_array_index_2047295_comb];
  assign p4_array_index_2047330_comb = p3_literal_2043916[p4_array_index_2047296_comb];
  assign p4_array_index_2047331_comb = p3_literal_2043918[p4_array_index_2047297_comb];
  assign p4_array_index_2047332_comb = p3_literal_2043920[p4_array_index_2047298_comb];
  assign p4_res7__450_comb = p4_array_index_2047327_comb ^ p4_array_index_2047328_comb ^ p4_array_index_2047329_comb ^ p4_array_index_2047330_comb ^ p4_array_index_2047331_comb ^ p4_array_index_2047332_comb ^ p4_array_index_2047299_comb ^ p3_literal_2043923[p4_array_index_2047316_comb] ^ p4_array_index_2047301_comb ^ p3_literal_2043920[p4_array_index_2047318_comb] ^ p3_literal_2043918[p4_array_index_2047303_comb] ^ p3_literal_2043916[p4_array_index_2047304_comb] ^ p3_literal_2043914[p4_array_index_2047305_comb] ^ p3_literal_2043912[p4_array_index_2047306_comb] ^ p3_literal_2043910[p4_array_index_2047307_comb] ^ p4_array_index_2047308_comb;
  assign p4_array_index_2047342_comb = p3_literal_2043912[p4_res7__448_comb];
  assign p4_array_index_2047343_comb = p3_literal_2043914[p4_array_index_2047294_comb];
  assign p4_array_index_2047344_comb = p3_literal_2043916[p4_array_index_2047295_comb];
  assign p4_array_index_2047345_comb = p3_literal_2043918[p4_array_index_2047296_comb];
  assign p4_array_index_2047346_comb = p3_literal_2043920[p4_array_index_2047297_comb];
  assign p4_res7__452_comb = p3_literal_2043910[p4_res7__450_comb] ^ p4_array_index_2047342_comb ^ p4_array_index_2047343_comb ^ p4_array_index_2047344_comb ^ p4_array_index_2047345_comb ^ p4_array_index_2047346_comb ^ p4_array_index_2047298_comb ^ p3_literal_2043923[p4_array_index_2047299_comb] ^ p4_array_index_2047316_comb ^ p3_literal_2043920[p4_array_index_2047301_comb] ^ p3_literal_2043918[p4_array_index_2047318_comb] ^ p3_literal_2043916[p4_array_index_2047303_comb] ^ p3_literal_2043914[p4_array_index_2047304_comb] ^ p3_literal_2043912[p4_array_index_2047305_comb] ^ p3_literal_2043910[p4_array_index_2047306_comb] ^ p4_array_index_2047307_comb;
  assign p4_array_index_2047356_comb = p3_literal_2043912[p4_res7__450_comb];
  assign p4_array_index_2047357_comb = p3_literal_2043914[p4_res7__448_comb];
  assign p4_array_index_2047358_comb = p3_literal_2043916[p4_array_index_2047294_comb];
  assign p4_array_index_2047359_comb = p3_literal_2043918[p4_array_index_2047295_comb];
  assign p4_array_index_2047360_comb = p3_literal_2043920[p4_array_index_2047296_comb];
  assign p4_res7__454_comb = p3_literal_2043910[p4_res7__452_comb] ^ p4_array_index_2047356_comb ^ p4_array_index_2047357_comb ^ p4_array_index_2047358_comb ^ p4_array_index_2047359_comb ^ p4_array_index_2047360_comb ^ p4_array_index_2047297_comb ^ p3_literal_2043923[p4_array_index_2047298_comb] ^ p4_array_index_2047299_comb ^ p3_literal_2043920[p4_array_index_2047316_comb] ^ p3_literal_2043918[p4_array_index_2047301_comb] ^ p3_literal_2043916[p4_array_index_2047318_comb] ^ p3_literal_2043914[p4_array_index_2047303_comb] ^ p3_literal_2043912[p4_array_index_2047304_comb] ^ p3_literal_2043910[p4_array_index_2047305_comb] ^ p4_array_index_2047306_comb;
  assign p4_array_index_2047371_comb = p3_literal_2043914[p4_res7__450_comb];
  assign p4_array_index_2047372_comb = p3_literal_2043916[p4_res7__448_comb];
  assign p4_array_index_2047373_comb = p3_literal_2043918[p4_array_index_2047294_comb];
  assign p4_array_index_2047374_comb = p3_literal_2043920[p4_array_index_2047295_comb];
  assign p4_res7__456_comb = p3_literal_2043910[p4_res7__454_comb] ^ p3_literal_2043912[p4_res7__452_comb] ^ p4_array_index_2047371_comb ^ p4_array_index_2047372_comb ^ p4_array_index_2047373_comb ^ p4_array_index_2047374_comb ^ p4_array_index_2047296_comb ^ p3_literal_2043923[p4_array_index_2047297_comb] ^ p4_array_index_2047298_comb ^ p4_array_index_2047315_comb ^ p3_literal_2043918[p4_array_index_2047316_comb] ^ p3_literal_2043916[p4_array_index_2047301_comb] ^ p3_literal_2043914[p4_array_index_2047318_comb] ^ p3_literal_2043912[p4_array_index_2047303_comb] ^ p3_literal_2043910[p4_array_index_2047304_comb] ^ p4_array_index_2047305_comb;
  assign p4_array_index_2047384_comb = p3_literal_2043914[p4_res7__452_comb];
  assign p4_array_index_2047385_comb = p3_literal_2043916[p4_res7__450_comb];
  assign p4_array_index_2047386_comb = p3_literal_2043918[p4_res7__448_comb];
  assign p4_array_index_2047387_comb = p3_literal_2043920[p4_array_index_2047294_comb];
  assign p4_res7__458_comb = p3_literal_2043910[p4_res7__456_comb] ^ p3_literal_2043912[p4_res7__454_comb] ^ p4_array_index_2047384_comb ^ p4_array_index_2047385_comb ^ p4_array_index_2047386_comb ^ p4_array_index_2047387_comb ^ p4_array_index_2047295_comb ^ p3_literal_2043923[p4_array_index_2047296_comb] ^ p4_array_index_2047297_comb ^ p4_array_index_2047332_comb ^ p3_literal_2043918[p4_array_index_2047299_comb] ^ p3_literal_2043916[p4_array_index_2047316_comb] ^ p3_literal_2043914[p4_array_index_2047301_comb] ^ p3_literal_2043912[p4_array_index_2047318_comb] ^ p3_literal_2043910[p4_array_index_2047303_comb] ^ p4_array_index_2047304_comb;
  assign p4_array_index_2047398_comb = p3_literal_2043916[p4_res7__452_comb];
  assign p4_array_index_2047399_comb = p3_literal_2043918[p4_res7__450_comb];
  assign p4_array_index_2047400_comb = p3_literal_2043920[p4_res7__448_comb];
  assign p4_res7__460_comb = p3_literal_2043910[p4_res7__458_comb] ^ p3_literal_2043912[p4_res7__456_comb] ^ p3_literal_2043914[p4_res7__454_comb] ^ p4_array_index_2047398_comb ^ p4_array_index_2047399_comb ^ p4_array_index_2047400_comb ^ p4_array_index_2047294_comb ^ p3_literal_2043923[p4_array_index_2047295_comb] ^ p4_array_index_2047296_comb ^ p4_array_index_2047346_comb ^ p4_array_index_2047314_comb ^ p3_literal_2043916[p4_array_index_2047299_comb] ^ p3_literal_2043914[p4_array_index_2047316_comb] ^ p3_literal_2043912[p4_array_index_2047301_comb] ^ p3_literal_2043910[p4_array_index_2047318_comb] ^ p4_array_index_2047303_comb;
  assign p4_array_index_2047410_comb = p3_literal_2043916[p4_res7__454_comb];
  assign p4_array_index_2047411_comb = p3_literal_2043918[p4_res7__452_comb];
  assign p4_array_index_2047412_comb = p3_literal_2043920[p4_res7__450_comb];
  assign p4_res7__462_comb = p3_literal_2043910[p4_res7__460_comb] ^ p3_literal_2043912[p4_res7__458_comb] ^ p3_literal_2043914[p4_res7__456_comb] ^ p4_array_index_2047410_comb ^ p4_array_index_2047411_comb ^ p4_array_index_2047412_comb ^ p4_res7__448_comb ^ p3_literal_2043923[p4_array_index_2047294_comb] ^ p4_array_index_2047295_comb ^ p4_array_index_2047360_comb ^ p4_array_index_2047331_comb ^ p3_literal_2043916[p4_array_index_2047298_comb] ^ p3_literal_2043914[p4_array_index_2047299_comb] ^ p3_literal_2043912[p4_array_index_2047316_comb] ^ p3_literal_2043910[p4_array_index_2047301_comb] ^ p4_array_index_2047318_comb;
  assign p4_array_index_2047423_comb = p3_literal_2043918[p4_res7__454_comb];
  assign p4_array_index_2047424_comb = p3_literal_2043920[p4_res7__452_comb];
  assign p4_res7__464_comb = p3_literal_2043910[p4_res7__462_comb] ^ p3_literal_2043912[p4_res7__460_comb] ^ p3_literal_2043914[p4_res7__458_comb] ^ p3_literal_2043916[p4_res7__456_comb] ^ p4_array_index_2047423_comb ^ p4_array_index_2047424_comb ^ p4_res7__450_comb ^ p3_literal_2043923[p4_res7__448_comb] ^ p4_array_index_2047294_comb ^ p4_array_index_2047374_comb ^ p4_array_index_2047345_comb ^ p4_array_index_2047313_comb ^ p3_literal_2043914[p4_array_index_2047298_comb] ^ p3_literal_2043912[p4_array_index_2047299_comb] ^ p3_literal_2043910[p4_array_index_2047316_comb] ^ p4_array_index_2047301_comb;
  assign p4_array_index_2047434_comb = p3_literal_2043918[p4_res7__456_comb];
  assign p4_array_index_2047435_comb = p3_literal_2043920[p4_res7__454_comb];
  assign p4_res7__466_comb = p3_literal_2043910[p4_res7__464_comb] ^ p3_literal_2043912[p4_res7__462_comb] ^ p3_literal_2043914[p4_res7__460_comb] ^ p3_literal_2043916[p4_res7__458_comb] ^ p4_array_index_2047434_comb ^ p4_array_index_2047435_comb ^ p4_res7__452_comb ^ p3_literal_2043923[p4_res7__450_comb] ^ p4_res7__448_comb ^ p4_array_index_2047387_comb ^ p4_array_index_2047359_comb ^ p4_array_index_2047330_comb ^ p3_literal_2043914[p4_array_index_2047297_comb] ^ p3_literal_2043912[p4_array_index_2047298_comb] ^ p3_literal_2043910[p4_array_index_2047299_comb] ^ p4_array_index_2047316_comb;
  assign p4_array_index_2047446_comb = p3_literal_2043920[p4_res7__456_comb];
  assign p4_res7__468_comb = p3_literal_2043910[p4_res7__466_comb] ^ p3_literal_2043912[p4_res7__464_comb] ^ p3_literal_2043914[p4_res7__462_comb] ^ p3_literal_2043916[p4_res7__460_comb] ^ p3_literal_2043918[p4_res7__458_comb] ^ p4_array_index_2047446_comb ^ p4_res7__454_comb ^ p3_literal_2043923[p4_res7__452_comb] ^ p4_res7__450_comb ^ p4_array_index_2047400_comb ^ p4_array_index_2047373_comb ^ p4_array_index_2047344_comb ^ p4_array_index_2047312_comb ^ p3_literal_2043912[p4_array_index_2047297_comb] ^ p3_literal_2043910[p4_array_index_2047298_comb] ^ p4_array_index_2047299_comb;
  assign p4_array_index_2047456_comb = p3_literal_2043920[p4_res7__458_comb];
  assign p4_res7__470_comb = p3_literal_2043910[p4_res7__468_comb] ^ p3_literal_2043912[p4_res7__466_comb] ^ p3_literal_2043914[p4_res7__464_comb] ^ p3_literal_2043916[p4_res7__462_comb] ^ p3_literal_2043918[p4_res7__460_comb] ^ p4_array_index_2047456_comb ^ p4_res7__456_comb ^ p3_literal_2043923[p4_res7__454_comb] ^ p4_res7__452_comb ^ p4_array_index_2047412_comb ^ p4_array_index_2047386_comb ^ p4_array_index_2047358_comb ^ p4_array_index_2047329_comb ^ p3_literal_2043912[p4_array_index_2047296_comb] ^ p3_literal_2043910[p4_array_index_2047297_comb] ^ p4_array_index_2047298_comb;
  assign p4_res7__472_comb = p3_literal_2043910[p4_res7__470_comb] ^ p3_literal_2043912[p4_res7__468_comb] ^ p3_literal_2043914[p4_res7__466_comb] ^ p3_literal_2043916[p4_res7__464_comb] ^ p3_literal_2043918[p4_res7__462_comb] ^ p3_literal_2043920[p4_res7__460_comb] ^ p4_res7__458_comb ^ p3_literal_2043923[p4_res7__456_comb] ^ p4_res7__454_comb ^ p4_array_index_2047424_comb ^ p4_array_index_2047399_comb ^ p4_array_index_2047372_comb ^ p4_array_index_2047343_comb ^ p4_array_index_2047311_comb ^ p3_literal_2043910[p4_array_index_2047296_comb] ^ p4_array_index_2047297_comb;
  assign p4_res7__474_comb = p3_literal_2043910[p4_res7__472_comb] ^ p3_literal_2043912[p4_res7__470_comb] ^ p3_literal_2043914[p4_res7__468_comb] ^ p3_literal_2043916[p4_res7__466_comb] ^ p3_literal_2043918[p4_res7__464_comb] ^ p3_literal_2043920[p4_res7__462_comb] ^ p4_res7__460_comb ^ p3_literal_2043923[p4_res7__458_comb] ^ p4_res7__456_comb ^ p4_array_index_2047435_comb ^ p4_array_index_2047411_comb ^ p4_array_index_2047385_comb ^ p4_array_index_2047357_comb ^ p4_array_index_2047328_comb ^ p3_literal_2043910[p4_array_index_2047295_comb] ^ p4_array_index_2047296_comb;
  assign p4_res7__476_comb = p3_literal_2043910[p4_res7__474_comb] ^ p3_literal_2043912[p4_res7__472_comb] ^ p3_literal_2043914[p4_res7__470_comb] ^ p3_literal_2043916[p4_res7__468_comb] ^ p3_literal_2043918[p4_res7__466_comb] ^ p3_literal_2043920[p4_res7__464_comb] ^ p4_res7__462_comb ^ p3_literal_2043923[p4_res7__460_comb] ^ p4_res7__458_comb ^ p4_array_index_2047446_comb ^ p4_array_index_2047423_comb ^ p4_array_index_2047398_comb ^ p4_array_index_2047371_comb ^ p4_array_index_2047342_comb ^ p4_array_index_2047310_comb ^ p4_array_index_2047295_comb;
  assign p4_res7__478_comb = p3_literal_2043910[p4_res7__476_comb] ^ p3_literal_2043912[p4_res7__474_comb] ^ p3_literal_2043914[p4_res7__472_comb] ^ p3_literal_2043916[p4_res7__470_comb] ^ p3_literal_2043918[p4_res7__468_comb] ^ p3_literal_2043920[p4_res7__466_comb] ^ p4_res7__464_comb ^ p3_literal_2043923[p4_res7__462_comb] ^ p4_res7__460_comb ^ p4_array_index_2047456_comb ^ p4_array_index_2047434_comb ^ p4_array_index_2047410_comb ^ p4_array_index_2047384_comb ^ p4_array_index_2047356_comb ^ p4_array_index_2047327_comb ^ p4_array_index_2047294_comb;
  assign p4_res__14_comb = {p4_res7__478_comb, p4_res7__476_comb, p4_res7__474_comb, p4_res7__472_comb, p4_res7__470_comb, p4_res7__468_comb, p4_res7__466_comb, p4_res7__464_comb, p4_res7__462_comb, p4_res7__460_comb, p4_res7__458_comb, p4_res7__456_comb, p4_res7__454_comb, p4_res7__452_comb, p4_res7__450_comb, p4_res7__448_comb};
  assign p4_k5_comb = p4_res__14_comb ^ p3_xor_2046948;
  assign p4_addedKey__47_comb = p4_k5_comb ^ 128'h2fb2_6c2c_0f0a_acd1_9935_81c3_4e97_5410;
  assign p4_array_index_2047512_comb = p3_literal_2043896[p4_addedKey__47_comb[127:120]];
  assign p4_array_index_2047513_comb = p3_literal_2043896[p4_addedKey__47_comb[119:112]];
  assign p4_array_index_2047514_comb = p3_literal_2043896[p4_addedKey__47_comb[111:104]];
  assign p4_array_index_2047515_comb = p3_literal_2043896[p4_addedKey__47_comb[103:96]];
  assign p4_array_index_2047516_comb = p3_literal_2043896[p4_addedKey__47_comb[95:88]];
  assign p4_array_index_2047517_comb = p3_literal_2043896[p4_addedKey__47_comb[87:80]];
  assign p4_array_index_2047519_comb = p3_literal_2043896[p4_addedKey__47_comb[71:64]];
  assign p4_array_index_2047521_comb = p3_literal_2043896[p4_addedKey__47_comb[55:48]];
  assign p4_array_index_2047522_comb = p3_literal_2043896[p4_addedKey__47_comb[47:40]];
  assign p4_array_index_2047523_comb = p3_literal_2043896[p4_addedKey__47_comb[39:32]];
  assign p4_array_index_2047524_comb = p3_literal_2043896[p4_addedKey__47_comb[31:24]];
  assign p4_array_index_2047525_comb = p3_literal_2043896[p4_addedKey__47_comb[23:16]];
  assign p4_array_index_2047526_comb = p3_literal_2043896[p4_addedKey__47_comb[15:8]];
  assign p4_array_index_2047528_comb = p3_literal_2043910[p4_array_index_2047512_comb];
  assign p4_array_index_2047529_comb = p3_literal_2043912[p4_array_index_2047513_comb];
  assign p4_array_index_2047530_comb = p3_literal_2043914[p4_array_index_2047514_comb];
  assign p4_array_index_2047531_comb = p3_literal_2043916[p4_array_index_2047515_comb];
  assign p4_array_index_2047532_comb = p3_literal_2043918[p4_array_index_2047516_comb];
  assign p4_array_index_2047533_comb = p3_literal_2043920[p4_array_index_2047517_comb];
  assign p4_array_index_2047534_comb = p3_literal_2043896[p4_addedKey__47_comb[79:72]];
  assign p4_array_index_2047536_comb = p3_literal_2043896[p4_addedKey__47_comb[63:56]];
  assign p4_res7__480_comb = p4_array_index_2047528_comb ^ p4_array_index_2047529_comb ^ p4_array_index_2047530_comb ^ p4_array_index_2047531_comb ^ p4_array_index_2047532_comb ^ p4_array_index_2047533_comb ^ p4_array_index_2047534_comb ^ p3_literal_2043923[p4_array_index_2047519_comb] ^ p4_array_index_2047536_comb ^ p3_literal_2043920[p4_array_index_2047521_comb] ^ p3_literal_2043918[p4_array_index_2047522_comb] ^ p3_literal_2043916[p4_array_index_2047523_comb] ^ p3_literal_2043914[p4_array_index_2047524_comb] ^ p3_literal_2043912[p4_array_index_2047525_comb] ^ p3_literal_2043910[p4_array_index_2047526_comb] ^ p3_literal_2043896[p4_addedKey__47_comb[7:0]];
  assign p4_array_index_2047545_comb = p3_literal_2043910[p4_res7__480_comb];
  assign p4_array_index_2047546_comb = p3_literal_2043912[p4_array_index_2047512_comb];
  assign p4_array_index_2047547_comb = p3_literal_2043914[p4_array_index_2047513_comb];
  assign p4_array_index_2047548_comb = p3_literal_2043916[p4_array_index_2047514_comb];
  assign p4_array_index_2047549_comb = p3_literal_2043918[p4_array_index_2047515_comb];
  assign p4_array_index_2047550_comb = p3_literal_2043920[p4_array_index_2047516_comb];
  assign p4_res7__482_comb = p4_array_index_2047545_comb ^ p4_array_index_2047546_comb ^ p4_array_index_2047547_comb ^ p4_array_index_2047548_comb ^ p4_array_index_2047549_comb ^ p4_array_index_2047550_comb ^ p4_array_index_2047517_comb ^ p3_literal_2043923[p4_array_index_2047534_comb] ^ p4_array_index_2047519_comb ^ p3_literal_2043920[p4_array_index_2047536_comb] ^ p3_literal_2043918[p4_array_index_2047521_comb] ^ p3_literal_2043916[p4_array_index_2047522_comb] ^ p3_literal_2043914[p4_array_index_2047523_comb] ^ p3_literal_2043912[p4_array_index_2047524_comb] ^ p3_literal_2043910[p4_array_index_2047525_comb] ^ p4_array_index_2047526_comb;
  assign p4_array_index_2047560_comb = p3_literal_2043912[p4_res7__480_comb];
  assign p4_array_index_2047561_comb = p3_literal_2043914[p4_array_index_2047512_comb];
  assign p4_array_index_2047562_comb = p3_literal_2043916[p4_array_index_2047513_comb];
  assign p4_array_index_2047563_comb = p3_literal_2043918[p4_array_index_2047514_comb];
  assign p4_array_index_2047564_comb = p3_literal_2043920[p4_array_index_2047515_comb];
  assign p4_res7__484_comb = p3_literal_2043910[p4_res7__482_comb] ^ p4_array_index_2047560_comb ^ p4_array_index_2047561_comb ^ p4_array_index_2047562_comb ^ p4_array_index_2047563_comb ^ p4_array_index_2047564_comb ^ p4_array_index_2047516_comb ^ p3_literal_2043923[p4_array_index_2047517_comb] ^ p4_array_index_2047534_comb ^ p3_literal_2043920[p4_array_index_2047519_comb] ^ p3_literal_2043918[p4_array_index_2047536_comb] ^ p3_literal_2043916[p4_array_index_2047521_comb] ^ p3_literal_2043914[p4_array_index_2047522_comb] ^ p3_literal_2043912[p4_array_index_2047523_comb] ^ p3_literal_2043910[p4_array_index_2047524_comb] ^ p4_array_index_2047525_comb;
  assign p4_array_index_2047574_comb = p3_literal_2043912[p4_res7__482_comb];
  assign p4_array_index_2047575_comb = p3_literal_2043914[p4_res7__480_comb];
  assign p4_array_index_2047576_comb = p3_literal_2043916[p4_array_index_2047512_comb];
  assign p4_array_index_2047577_comb = p3_literal_2043918[p4_array_index_2047513_comb];
  assign p4_array_index_2047578_comb = p3_literal_2043920[p4_array_index_2047514_comb];
  assign p4_res7__486_comb = p3_literal_2043910[p4_res7__484_comb] ^ p4_array_index_2047574_comb ^ p4_array_index_2047575_comb ^ p4_array_index_2047576_comb ^ p4_array_index_2047577_comb ^ p4_array_index_2047578_comb ^ p4_array_index_2047515_comb ^ p3_literal_2043923[p4_array_index_2047516_comb] ^ p4_array_index_2047517_comb ^ p3_literal_2043920[p4_array_index_2047534_comb] ^ p3_literal_2043918[p4_array_index_2047519_comb] ^ p3_literal_2043916[p4_array_index_2047536_comb] ^ p3_literal_2043914[p4_array_index_2047521_comb] ^ p3_literal_2043912[p4_array_index_2047522_comb] ^ p3_literal_2043910[p4_array_index_2047523_comb] ^ p4_array_index_2047524_comb;
  assign p4_array_index_2047589_comb = p3_literal_2043914[p4_res7__482_comb];
  assign p4_array_index_2047590_comb = p3_literal_2043916[p4_res7__480_comb];
  assign p4_array_index_2047591_comb = p3_literal_2043918[p4_array_index_2047512_comb];
  assign p4_array_index_2047592_comb = p3_literal_2043920[p4_array_index_2047513_comb];
  assign p4_res7__488_comb = p3_literal_2043910[p4_res7__486_comb] ^ p3_literal_2043912[p4_res7__484_comb] ^ p4_array_index_2047589_comb ^ p4_array_index_2047590_comb ^ p4_array_index_2047591_comb ^ p4_array_index_2047592_comb ^ p4_array_index_2047514_comb ^ p3_literal_2043923[p4_array_index_2047515_comb] ^ p4_array_index_2047516_comb ^ p4_array_index_2047533_comb ^ p3_literal_2043918[p4_array_index_2047534_comb] ^ p3_literal_2043916[p4_array_index_2047519_comb] ^ p3_literal_2043914[p4_array_index_2047536_comb] ^ p3_literal_2043912[p4_array_index_2047521_comb] ^ p3_literal_2043910[p4_array_index_2047522_comb] ^ p4_array_index_2047523_comb;
  assign p4_array_index_2047602_comb = p3_literal_2043914[p4_res7__484_comb];
  assign p4_array_index_2047603_comb = p3_literal_2043916[p4_res7__482_comb];
  assign p4_array_index_2047604_comb = p3_literal_2043918[p4_res7__480_comb];
  assign p4_array_index_2047605_comb = p3_literal_2043920[p4_array_index_2047512_comb];
  assign p4_res7__490_comb = p3_literal_2043910[p4_res7__488_comb] ^ p3_literal_2043912[p4_res7__486_comb] ^ p4_array_index_2047602_comb ^ p4_array_index_2047603_comb ^ p4_array_index_2047604_comb ^ p4_array_index_2047605_comb ^ p4_array_index_2047513_comb ^ p3_literal_2043923[p4_array_index_2047514_comb] ^ p4_array_index_2047515_comb ^ p4_array_index_2047550_comb ^ p3_literal_2043918[p4_array_index_2047517_comb] ^ p3_literal_2043916[p4_array_index_2047534_comb] ^ p3_literal_2043914[p4_array_index_2047519_comb] ^ p3_literal_2043912[p4_array_index_2047536_comb] ^ p3_literal_2043910[p4_array_index_2047521_comb] ^ p4_array_index_2047522_comb;
  assign p4_array_index_2047616_comb = p3_literal_2043916[p4_res7__484_comb];
  assign p4_array_index_2047617_comb = p3_literal_2043918[p4_res7__482_comb];
  assign p4_array_index_2047618_comb = p3_literal_2043920[p4_res7__480_comb];
  assign p4_res7__492_comb = p3_literal_2043910[p4_res7__490_comb] ^ p3_literal_2043912[p4_res7__488_comb] ^ p3_literal_2043914[p4_res7__486_comb] ^ p4_array_index_2047616_comb ^ p4_array_index_2047617_comb ^ p4_array_index_2047618_comb ^ p4_array_index_2047512_comb ^ p3_literal_2043923[p4_array_index_2047513_comb] ^ p4_array_index_2047514_comb ^ p4_array_index_2047564_comb ^ p4_array_index_2047532_comb ^ p3_literal_2043916[p4_array_index_2047517_comb] ^ p3_literal_2043914[p4_array_index_2047534_comb] ^ p3_literal_2043912[p4_array_index_2047519_comb] ^ p3_literal_2043910[p4_array_index_2047536_comb] ^ p4_array_index_2047521_comb;
  assign p4_array_index_2047628_comb = p3_literal_2043916[p4_res7__486_comb];
  assign p4_array_index_2047629_comb = p3_literal_2043918[p4_res7__484_comb];
  assign p4_array_index_2047630_comb = p3_literal_2043920[p4_res7__482_comb];
  assign p4_res7__494_comb = p3_literal_2043910[p4_res7__492_comb] ^ p3_literal_2043912[p4_res7__490_comb] ^ p3_literal_2043914[p4_res7__488_comb] ^ p4_array_index_2047628_comb ^ p4_array_index_2047629_comb ^ p4_array_index_2047630_comb ^ p4_res7__480_comb ^ p3_literal_2043923[p4_array_index_2047512_comb] ^ p4_array_index_2047513_comb ^ p4_array_index_2047578_comb ^ p4_array_index_2047549_comb ^ p3_literal_2043916[p4_array_index_2047516_comb] ^ p3_literal_2043914[p4_array_index_2047517_comb] ^ p3_literal_2043912[p4_array_index_2047534_comb] ^ p3_literal_2043910[p4_array_index_2047519_comb] ^ p4_array_index_2047536_comb;
  assign p4_array_index_2047641_comb = p3_literal_2043918[p4_res7__486_comb];
  assign p4_array_index_2047642_comb = p3_literal_2043920[p4_res7__484_comb];
  assign p4_res7__496_comb = p3_literal_2043910[p4_res7__494_comb] ^ p3_literal_2043912[p4_res7__492_comb] ^ p3_literal_2043914[p4_res7__490_comb] ^ p3_literal_2043916[p4_res7__488_comb] ^ p4_array_index_2047641_comb ^ p4_array_index_2047642_comb ^ p4_res7__482_comb ^ p3_literal_2043923[p4_res7__480_comb] ^ p4_array_index_2047512_comb ^ p4_array_index_2047592_comb ^ p4_array_index_2047563_comb ^ p4_array_index_2047531_comb ^ p3_literal_2043914[p4_array_index_2047516_comb] ^ p3_literal_2043912[p4_array_index_2047517_comb] ^ p3_literal_2043910[p4_array_index_2047534_comb] ^ p4_array_index_2047519_comb;
  assign p4_array_index_2047652_comb = p3_literal_2043918[p4_res7__488_comb];
  assign p4_array_index_2047653_comb = p3_literal_2043920[p4_res7__486_comb];
  assign p4_res7__498_comb = p3_literal_2043910[p4_res7__496_comb] ^ p3_literal_2043912[p4_res7__494_comb] ^ p3_literal_2043914[p4_res7__492_comb] ^ p3_literal_2043916[p4_res7__490_comb] ^ p4_array_index_2047652_comb ^ p4_array_index_2047653_comb ^ p4_res7__484_comb ^ p3_literal_2043923[p4_res7__482_comb] ^ p4_res7__480_comb ^ p4_array_index_2047605_comb ^ p4_array_index_2047577_comb ^ p4_array_index_2047548_comb ^ p3_literal_2043914[p4_array_index_2047515_comb] ^ p3_literal_2043912[p4_array_index_2047516_comb] ^ p3_literal_2043910[p4_array_index_2047517_comb] ^ p4_array_index_2047534_comb;
  assign p4_array_index_2047664_comb = p3_literal_2043920[p4_res7__488_comb];
  assign p4_res7__500_comb = p3_literal_2043910[p4_res7__498_comb] ^ p3_literal_2043912[p4_res7__496_comb] ^ p3_literal_2043914[p4_res7__494_comb] ^ p3_literal_2043916[p4_res7__492_comb] ^ p3_literal_2043918[p4_res7__490_comb] ^ p4_array_index_2047664_comb ^ p4_res7__486_comb ^ p3_literal_2043923[p4_res7__484_comb] ^ p4_res7__482_comb ^ p4_array_index_2047618_comb ^ p4_array_index_2047591_comb ^ p4_array_index_2047562_comb ^ p4_array_index_2047530_comb ^ p3_literal_2043912[p4_array_index_2047515_comb] ^ p3_literal_2043910[p4_array_index_2047516_comb] ^ p4_array_index_2047517_comb;
  assign p4_array_index_2047674_comb = p3_literal_2043920[p4_res7__490_comb];
  assign p4_res7__502_comb = p3_literal_2043910[p4_res7__500_comb] ^ p3_literal_2043912[p4_res7__498_comb] ^ p3_literal_2043914[p4_res7__496_comb] ^ p3_literal_2043916[p4_res7__494_comb] ^ p3_literal_2043918[p4_res7__492_comb] ^ p4_array_index_2047674_comb ^ p4_res7__488_comb ^ p3_literal_2043923[p4_res7__486_comb] ^ p4_res7__484_comb ^ p4_array_index_2047630_comb ^ p4_array_index_2047604_comb ^ p4_array_index_2047576_comb ^ p4_array_index_2047547_comb ^ p3_literal_2043912[p4_array_index_2047514_comb] ^ p3_literal_2043910[p4_array_index_2047515_comb] ^ p4_array_index_2047516_comb;
  assign p4_res7__504_comb = p3_literal_2043910[p4_res7__502_comb] ^ p3_literal_2043912[p4_res7__500_comb] ^ p3_literal_2043914[p4_res7__498_comb] ^ p3_literal_2043916[p4_res7__496_comb] ^ p3_literal_2043918[p4_res7__494_comb] ^ p3_literal_2043920[p4_res7__492_comb] ^ p4_res7__490_comb ^ p3_literal_2043923[p4_res7__488_comb] ^ p4_res7__486_comb ^ p4_array_index_2047642_comb ^ p4_array_index_2047617_comb ^ p4_array_index_2047590_comb ^ p4_array_index_2047561_comb ^ p4_array_index_2047529_comb ^ p3_literal_2043910[p4_array_index_2047514_comb] ^ p4_array_index_2047515_comb;
  assign p4_res7__506_comb = p3_literal_2043910[p4_res7__504_comb] ^ p3_literal_2043912[p4_res7__502_comb] ^ p3_literal_2043914[p4_res7__500_comb] ^ p3_literal_2043916[p4_res7__498_comb] ^ p3_literal_2043918[p4_res7__496_comb] ^ p3_literal_2043920[p4_res7__494_comb] ^ p4_res7__492_comb ^ p3_literal_2043923[p4_res7__490_comb] ^ p4_res7__488_comb ^ p4_array_index_2047653_comb ^ p4_array_index_2047629_comb ^ p4_array_index_2047603_comb ^ p4_array_index_2047575_comb ^ p4_array_index_2047546_comb ^ p3_literal_2043910[p4_array_index_2047513_comb] ^ p4_array_index_2047514_comb;
  assign p4_res7__508_comb = p3_literal_2043910[p4_res7__506_comb] ^ p3_literal_2043912[p4_res7__504_comb] ^ p3_literal_2043914[p4_res7__502_comb] ^ p3_literal_2043916[p4_res7__500_comb] ^ p3_literal_2043918[p4_res7__498_comb] ^ p3_literal_2043920[p4_res7__496_comb] ^ p4_res7__494_comb ^ p3_literal_2043923[p4_res7__492_comb] ^ p4_res7__490_comb ^ p4_array_index_2047664_comb ^ p4_array_index_2047641_comb ^ p4_array_index_2047616_comb ^ p4_array_index_2047589_comb ^ p4_array_index_2047560_comb ^ p4_array_index_2047528_comb ^ p4_array_index_2047513_comb;
  assign p4_res7__510_comb = p3_literal_2043910[p4_res7__508_comb] ^ p3_literal_2043912[p4_res7__506_comb] ^ p3_literal_2043914[p4_res7__504_comb] ^ p3_literal_2043916[p4_res7__502_comb] ^ p3_literal_2043918[p4_res7__500_comb] ^ p3_literal_2043920[p4_res7__498_comb] ^ p4_res7__496_comb ^ p3_literal_2043923[p4_res7__494_comb] ^ p4_res7__492_comb ^ p4_array_index_2047674_comb ^ p4_array_index_2047652_comb ^ p4_array_index_2047628_comb ^ p4_array_index_2047602_comb ^ p4_array_index_2047574_comb ^ p4_array_index_2047545_comb ^ p4_array_index_2047512_comb;
  assign p4_res__15_comb = {p4_res7__510_comb, p4_res7__508_comb, p4_res7__506_comb, p4_res7__504_comb, p4_res7__502_comb, p4_res7__500_comb, p4_res7__498_comb, p4_res7__496_comb, p4_res7__494_comb, p4_res7__492_comb, p4_res7__490_comb, p4_res7__488_comb, p4_res7__486_comb, p4_res7__484_comb, p4_res7__482_comb, p4_res7__480_comb};
  assign p4_k4_comb = p4_res__15_comb ^ p4_xor_2047278_comb;
  assign p4_addedKey__48_comb = p4_k4_comb ^ 128'h4110_1a5e_6342_d669_c412_3cd3_9313_c011;
  assign p4_array_index_2047730_comb = p3_literal_2043896[p4_addedKey__48_comb[127:120]];
  assign p4_array_index_2047731_comb = p3_literal_2043896[p4_addedKey__48_comb[119:112]];
  assign p4_array_index_2047732_comb = p3_literal_2043896[p4_addedKey__48_comb[111:104]];
  assign p4_array_index_2047733_comb = p3_literal_2043896[p4_addedKey__48_comb[103:96]];
  assign p4_array_index_2047734_comb = p3_literal_2043896[p4_addedKey__48_comb[95:88]];
  assign p4_array_index_2047735_comb = p3_literal_2043896[p4_addedKey__48_comb[87:80]];
  assign p4_array_index_2047737_comb = p3_literal_2043896[p4_addedKey__48_comb[71:64]];
  assign p4_array_index_2047739_comb = p3_literal_2043896[p4_addedKey__48_comb[55:48]];
  assign p4_array_index_2047740_comb = p3_literal_2043896[p4_addedKey__48_comb[47:40]];
  assign p4_array_index_2047741_comb = p3_literal_2043896[p4_addedKey__48_comb[39:32]];
  assign p4_array_index_2047742_comb = p3_literal_2043896[p4_addedKey__48_comb[31:24]];
  assign p4_array_index_2047743_comb = p3_literal_2043896[p4_addedKey__48_comb[23:16]];
  assign p4_array_index_2047744_comb = p3_literal_2043896[p4_addedKey__48_comb[15:8]];
  assign p4_array_index_2047746_comb = p3_literal_2043910[p4_array_index_2047730_comb];
  assign p4_array_index_2047747_comb = p3_literal_2043912[p4_array_index_2047731_comb];
  assign p4_array_index_2047748_comb = p3_literal_2043914[p4_array_index_2047732_comb];
  assign p4_array_index_2047749_comb = p3_literal_2043916[p4_array_index_2047733_comb];
  assign p4_array_index_2047750_comb = p3_literal_2043918[p4_array_index_2047734_comb];
  assign p4_array_index_2047751_comb = p3_literal_2043920[p4_array_index_2047735_comb];
  assign p4_array_index_2047752_comb = p3_literal_2043896[p4_addedKey__48_comb[79:72]];
  assign p4_array_index_2047754_comb = p3_literal_2043896[p4_addedKey__48_comb[63:56]];
  assign p4_res7__512_comb = p4_array_index_2047746_comb ^ p4_array_index_2047747_comb ^ p4_array_index_2047748_comb ^ p4_array_index_2047749_comb ^ p4_array_index_2047750_comb ^ p4_array_index_2047751_comb ^ p4_array_index_2047752_comb ^ p3_literal_2043923[p4_array_index_2047737_comb] ^ p4_array_index_2047754_comb ^ p3_literal_2043920[p4_array_index_2047739_comb] ^ p3_literal_2043918[p4_array_index_2047740_comb] ^ p3_literal_2043916[p4_array_index_2047741_comb] ^ p3_literal_2043914[p4_array_index_2047742_comb] ^ p3_literal_2043912[p4_array_index_2047743_comb] ^ p3_literal_2043910[p4_array_index_2047744_comb] ^ p3_literal_2043896[p4_addedKey__48_comb[7:0]];
  assign p4_array_index_2047763_comb = p3_literal_2043910[p4_res7__512_comb];
  assign p4_array_index_2047764_comb = p3_literal_2043912[p4_array_index_2047730_comb];
  assign p4_array_index_2047765_comb = p3_literal_2043914[p4_array_index_2047731_comb];
  assign p4_array_index_2047766_comb = p3_literal_2043916[p4_array_index_2047732_comb];
  assign p4_array_index_2047767_comb = p3_literal_2043918[p4_array_index_2047733_comb];
  assign p4_array_index_2047768_comb = p3_literal_2043920[p4_array_index_2047734_comb];
  assign p4_res7__514_comb = p4_array_index_2047763_comb ^ p4_array_index_2047764_comb ^ p4_array_index_2047765_comb ^ p4_array_index_2047766_comb ^ p4_array_index_2047767_comb ^ p4_array_index_2047768_comb ^ p4_array_index_2047735_comb ^ p3_literal_2043923[p4_array_index_2047752_comb] ^ p4_array_index_2047737_comb ^ p3_literal_2043920[p4_array_index_2047754_comb] ^ p3_literal_2043918[p4_array_index_2047739_comb] ^ p3_literal_2043916[p4_array_index_2047740_comb] ^ p3_literal_2043914[p4_array_index_2047741_comb] ^ p3_literal_2043912[p4_array_index_2047742_comb] ^ p3_literal_2043910[p4_array_index_2047743_comb] ^ p4_array_index_2047744_comb;
  assign p4_array_index_2047778_comb = p3_literal_2043912[p4_res7__512_comb];
  assign p4_array_index_2047779_comb = p3_literal_2043914[p4_array_index_2047730_comb];
  assign p4_array_index_2047780_comb = p3_literal_2043916[p4_array_index_2047731_comb];
  assign p4_array_index_2047781_comb = p3_literal_2043918[p4_array_index_2047732_comb];
  assign p4_array_index_2047782_comb = p3_literal_2043920[p4_array_index_2047733_comb];
  assign p4_res7__516_comb = p3_literal_2043910[p4_res7__514_comb] ^ p4_array_index_2047778_comb ^ p4_array_index_2047779_comb ^ p4_array_index_2047780_comb ^ p4_array_index_2047781_comb ^ p4_array_index_2047782_comb ^ p4_array_index_2047734_comb ^ p3_literal_2043923[p4_array_index_2047735_comb] ^ p4_array_index_2047752_comb ^ p3_literal_2043920[p4_array_index_2047737_comb] ^ p3_literal_2043918[p4_array_index_2047754_comb] ^ p3_literal_2043916[p4_array_index_2047739_comb] ^ p3_literal_2043914[p4_array_index_2047740_comb] ^ p3_literal_2043912[p4_array_index_2047741_comb] ^ p3_literal_2043910[p4_array_index_2047742_comb] ^ p4_array_index_2047743_comb;
  assign p4_array_index_2047792_comb = p3_literal_2043912[p4_res7__514_comb];
  assign p4_array_index_2047793_comb = p3_literal_2043914[p4_res7__512_comb];
  assign p4_array_index_2047794_comb = p3_literal_2043916[p4_array_index_2047730_comb];
  assign p4_array_index_2047795_comb = p3_literal_2043918[p4_array_index_2047731_comb];
  assign p4_array_index_2047796_comb = p3_literal_2043920[p4_array_index_2047732_comb];
  assign p4_res7__518_comb = p3_literal_2043910[p4_res7__516_comb] ^ p4_array_index_2047792_comb ^ p4_array_index_2047793_comb ^ p4_array_index_2047794_comb ^ p4_array_index_2047795_comb ^ p4_array_index_2047796_comb ^ p4_array_index_2047733_comb ^ p3_literal_2043923[p4_array_index_2047734_comb] ^ p4_array_index_2047735_comb ^ p3_literal_2043920[p4_array_index_2047752_comb] ^ p3_literal_2043918[p4_array_index_2047737_comb] ^ p3_literal_2043916[p4_array_index_2047754_comb] ^ p3_literal_2043914[p4_array_index_2047739_comb] ^ p3_literal_2043912[p4_array_index_2047740_comb] ^ p3_literal_2043910[p4_array_index_2047741_comb] ^ p4_array_index_2047742_comb;
  assign p4_array_index_2047807_comb = p3_literal_2043914[p4_res7__514_comb];
  assign p4_array_index_2047808_comb = p3_literal_2043916[p4_res7__512_comb];
  assign p4_array_index_2047809_comb = p3_literal_2043918[p4_array_index_2047730_comb];
  assign p4_array_index_2047810_comb = p3_literal_2043920[p4_array_index_2047731_comb];
  assign p4_res7__520_comb = p3_literal_2043910[p4_res7__518_comb] ^ p3_literal_2043912[p4_res7__516_comb] ^ p4_array_index_2047807_comb ^ p4_array_index_2047808_comb ^ p4_array_index_2047809_comb ^ p4_array_index_2047810_comb ^ p4_array_index_2047732_comb ^ p3_literal_2043923[p4_array_index_2047733_comb] ^ p4_array_index_2047734_comb ^ p4_array_index_2047751_comb ^ p3_literal_2043918[p4_array_index_2047752_comb] ^ p3_literal_2043916[p4_array_index_2047737_comb] ^ p3_literal_2043914[p4_array_index_2047754_comb] ^ p3_literal_2043912[p4_array_index_2047739_comb] ^ p3_literal_2043910[p4_array_index_2047740_comb] ^ p4_array_index_2047741_comb;
  assign p4_array_index_2047820_comb = p3_literal_2043914[p4_res7__516_comb];
  assign p4_array_index_2047821_comb = p3_literal_2043916[p4_res7__514_comb];
  assign p4_array_index_2047822_comb = p3_literal_2043918[p4_res7__512_comb];
  assign p4_array_index_2047823_comb = p3_literal_2043920[p4_array_index_2047730_comb];
  assign p4_res7__522_comb = p3_literal_2043910[p4_res7__520_comb] ^ p3_literal_2043912[p4_res7__518_comb] ^ p4_array_index_2047820_comb ^ p4_array_index_2047821_comb ^ p4_array_index_2047822_comb ^ p4_array_index_2047823_comb ^ p4_array_index_2047731_comb ^ p3_literal_2043923[p4_array_index_2047732_comb] ^ p4_array_index_2047733_comb ^ p4_array_index_2047768_comb ^ p3_literal_2043918[p4_array_index_2047735_comb] ^ p3_literal_2043916[p4_array_index_2047752_comb] ^ p3_literal_2043914[p4_array_index_2047737_comb] ^ p3_literal_2043912[p4_array_index_2047754_comb] ^ p3_literal_2043910[p4_array_index_2047739_comb] ^ p4_array_index_2047740_comb;
  assign p4_array_index_2047834_comb = p3_literal_2043916[p4_res7__516_comb];
  assign p4_array_index_2047835_comb = p3_literal_2043918[p4_res7__514_comb];
  assign p4_array_index_2047836_comb = p3_literal_2043920[p4_res7__512_comb];
  assign p4_res7__524_comb = p3_literal_2043910[p4_res7__522_comb] ^ p3_literal_2043912[p4_res7__520_comb] ^ p3_literal_2043914[p4_res7__518_comb] ^ p4_array_index_2047834_comb ^ p4_array_index_2047835_comb ^ p4_array_index_2047836_comb ^ p4_array_index_2047730_comb ^ p3_literal_2043923[p4_array_index_2047731_comb] ^ p4_array_index_2047732_comb ^ p4_array_index_2047782_comb ^ p4_array_index_2047750_comb ^ p3_literal_2043916[p4_array_index_2047735_comb] ^ p3_literal_2043914[p4_array_index_2047752_comb] ^ p3_literal_2043912[p4_array_index_2047737_comb] ^ p3_literal_2043910[p4_array_index_2047754_comb] ^ p4_array_index_2047739_comb;
  assign p4_array_index_2047846_comb = p3_literal_2043916[p4_res7__518_comb];
  assign p4_array_index_2047847_comb = p3_literal_2043918[p4_res7__516_comb];
  assign p4_array_index_2047848_comb = p3_literal_2043920[p4_res7__514_comb];
  assign p4_res7__526_comb = p3_literal_2043910[p4_res7__524_comb] ^ p3_literal_2043912[p4_res7__522_comb] ^ p3_literal_2043914[p4_res7__520_comb] ^ p4_array_index_2047846_comb ^ p4_array_index_2047847_comb ^ p4_array_index_2047848_comb ^ p4_res7__512_comb ^ p3_literal_2043923[p4_array_index_2047730_comb] ^ p4_array_index_2047731_comb ^ p4_array_index_2047796_comb ^ p4_array_index_2047767_comb ^ p3_literal_2043916[p4_array_index_2047734_comb] ^ p3_literal_2043914[p4_array_index_2047735_comb] ^ p3_literal_2043912[p4_array_index_2047752_comb] ^ p3_literal_2043910[p4_array_index_2047737_comb] ^ p4_array_index_2047754_comb;
  assign p4_array_index_2047859_comb = p3_literal_2043918[p4_res7__518_comb];
  assign p4_array_index_2047860_comb = p3_literal_2043920[p4_res7__516_comb];
  assign p4_res7__528_comb = p3_literal_2043910[p4_res7__526_comb] ^ p3_literal_2043912[p4_res7__524_comb] ^ p3_literal_2043914[p4_res7__522_comb] ^ p3_literal_2043916[p4_res7__520_comb] ^ p4_array_index_2047859_comb ^ p4_array_index_2047860_comb ^ p4_res7__514_comb ^ p3_literal_2043923[p4_res7__512_comb] ^ p4_array_index_2047730_comb ^ p4_array_index_2047810_comb ^ p4_array_index_2047781_comb ^ p4_array_index_2047749_comb ^ p3_literal_2043914[p4_array_index_2047734_comb] ^ p3_literal_2043912[p4_array_index_2047735_comb] ^ p3_literal_2043910[p4_array_index_2047752_comb] ^ p4_array_index_2047737_comb;
  assign p4_array_index_2047870_comb = p3_literal_2043918[p4_res7__520_comb];
  assign p4_array_index_2047871_comb = p3_literal_2043920[p4_res7__518_comb];
  assign p4_res7__530_comb = p3_literal_2043910[p4_res7__528_comb] ^ p3_literal_2043912[p4_res7__526_comb] ^ p3_literal_2043914[p4_res7__524_comb] ^ p3_literal_2043916[p4_res7__522_comb] ^ p4_array_index_2047870_comb ^ p4_array_index_2047871_comb ^ p4_res7__516_comb ^ p3_literal_2043923[p4_res7__514_comb] ^ p4_res7__512_comb ^ p4_array_index_2047823_comb ^ p4_array_index_2047795_comb ^ p4_array_index_2047766_comb ^ p3_literal_2043914[p4_array_index_2047733_comb] ^ p3_literal_2043912[p4_array_index_2047734_comb] ^ p3_literal_2043910[p4_array_index_2047735_comb] ^ p4_array_index_2047752_comb;
  assign p4_array_index_2047882_comb = p3_literal_2043920[p4_res7__520_comb];
  assign p4_res7__532_comb = p3_literal_2043910[p4_res7__530_comb] ^ p3_literal_2043912[p4_res7__528_comb] ^ p3_literal_2043914[p4_res7__526_comb] ^ p3_literal_2043916[p4_res7__524_comb] ^ p3_literal_2043918[p4_res7__522_comb] ^ p4_array_index_2047882_comb ^ p4_res7__518_comb ^ p3_literal_2043923[p4_res7__516_comb] ^ p4_res7__514_comb ^ p4_array_index_2047836_comb ^ p4_array_index_2047809_comb ^ p4_array_index_2047780_comb ^ p4_array_index_2047748_comb ^ p3_literal_2043912[p4_array_index_2047733_comb] ^ p3_literal_2043910[p4_array_index_2047734_comb] ^ p4_array_index_2047735_comb;
  assign p4_array_index_2047892_comb = p3_literal_2043920[p4_res7__522_comb];
  assign p4_res7__534_comb = p3_literal_2043910[p4_res7__532_comb] ^ p3_literal_2043912[p4_res7__530_comb] ^ p3_literal_2043914[p4_res7__528_comb] ^ p3_literal_2043916[p4_res7__526_comb] ^ p3_literal_2043918[p4_res7__524_comb] ^ p4_array_index_2047892_comb ^ p4_res7__520_comb ^ p3_literal_2043923[p4_res7__518_comb] ^ p4_res7__516_comb ^ p4_array_index_2047848_comb ^ p4_array_index_2047822_comb ^ p4_array_index_2047794_comb ^ p4_array_index_2047765_comb ^ p3_literal_2043912[p4_array_index_2047732_comb] ^ p3_literal_2043910[p4_array_index_2047733_comb] ^ p4_array_index_2047734_comb;
  assign p4_res7__536_comb = p3_literal_2043910[p4_res7__534_comb] ^ p3_literal_2043912[p4_res7__532_comb] ^ p3_literal_2043914[p4_res7__530_comb] ^ p3_literal_2043916[p4_res7__528_comb] ^ p3_literal_2043918[p4_res7__526_comb] ^ p3_literal_2043920[p4_res7__524_comb] ^ p4_res7__522_comb ^ p3_literal_2043923[p4_res7__520_comb] ^ p4_res7__518_comb ^ p4_array_index_2047860_comb ^ p4_array_index_2047835_comb ^ p4_array_index_2047808_comb ^ p4_array_index_2047779_comb ^ p4_array_index_2047747_comb ^ p3_literal_2043910[p4_array_index_2047732_comb] ^ p4_array_index_2047733_comb;
  assign p4_res7__538_comb = p3_literal_2043910[p4_res7__536_comb] ^ p3_literal_2043912[p4_res7__534_comb] ^ p3_literal_2043914[p4_res7__532_comb] ^ p3_literal_2043916[p4_res7__530_comb] ^ p3_literal_2043918[p4_res7__528_comb] ^ p3_literal_2043920[p4_res7__526_comb] ^ p4_res7__524_comb ^ p3_literal_2043923[p4_res7__522_comb] ^ p4_res7__520_comb ^ p4_array_index_2047871_comb ^ p4_array_index_2047847_comb ^ p4_array_index_2047821_comb ^ p4_array_index_2047793_comb ^ p4_array_index_2047764_comb ^ p3_literal_2043910[p4_array_index_2047731_comb] ^ p4_array_index_2047732_comb;
  assign p4_res7__540_comb = p3_literal_2043910[p4_res7__538_comb] ^ p3_literal_2043912[p4_res7__536_comb] ^ p3_literal_2043914[p4_res7__534_comb] ^ p3_literal_2043916[p4_res7__532_comb] ^ p3_literal_2043918[p4_res7__530_comb] ^ p3_literal_2043920[p4_res7__528_comb] ^ p4_res7__526_comb ^ p3_literal_2043923[p4_res7__524_comb] ^ p4_res7__522_comb ^ p4_array_index_2047882_comb ^ p4_array_index_2047859_comb ^ p4_array_index_2047834_comb ^ p4_array_index_2047807_comb ^ p4_array_index_2047778_comb ^ p4_array_index_2047746_comb ^ p4_array_index_2047731_comb;
  assign p4_res7__542_comb = p3_literal_2043910[p4_res7__540_comb] ^ p3_literal_2043912[p4_res7__538_comb] ^ p3_literal_2043914[p4_res7__536_comb] ^ p3_literal_2043916[p4_res7__534_comb] ^ p3_literal_2043918[p4_res7__532_comb] ^ p3_literal_2043920[p4_res7__530_comb] ^ p4_res7__528_comb ^ p3_literal_2043923[p4_res7__526_comb] ^ p4_res7__524_comb ^ p4_array_index_2047892_comb ^ p4_array_index_2047870_comb ^ p4_array_index_2047846_comb ^ p4_array_index_2047820_comb ^ p4_array_index_2047792_comb ^ p4_array_index_2047763_comb ^ p4_array_index_2047730_comb;
  assign p4_res__16_comb = {p4_res7__542_comb, p4_res7__540_comb, p4_res7__538_comb, p4_res7__536_comb, p4_res7__534_comb, p4_res7__532_comb, p4_res7__530_comb, p4_res7__528_comb, p4_res7__526_comb, p4_res7__524_comb, p4_res7__522_comb, p4_res7__520_comb, p4_res7__518_comb, p4_res7__516_comb, p4_res7__514_comb, p4_res7__512_comb};
  assign p4_xor_2047932_comb = p4_res__16_comb ^ p4_k5_comb;
  assign p4_addedKey__49_comb = p4_xor_2047932_comb ^ 128'hf335_80c8_d79a_5862_237b_38e3_375c_bf12;
  assign p4_array_index_2047948_comb = p3_literal_2043896[p4_addedKey__49_comb[127:120]];
  assign p4_array_index_2047949_comb = p3_literal_2043896[p4_addedKey__49_comb[119:112]];
  assign p4_array_index_2047950_comb = p3_literal_2043896[p4_addedKey__49_comb[111:104]];
  assign p4_array_index_2047951_comb = p3_literal_2043896[p4_addedKey__49_comb[103:96]];
  assign p4_array_index_2047952_comb = p3_literal_2043896[p4_addedKey__49_comb[95:88]];
  assign p4_array_index_2047953_comb = p3_literal_2043896[p4_addedKey__49_comb[87:80]];
  assign p4_array_index_2047955_comb = p3_literal_2043896[p4_addedKey__49_comb[71:64]];
  assign p4_array_index_2047957_comb = p3_literal_2043896[p4_addedKey__49_comb[55:48]];
  assign p4_array_index_2047958_comb = p3_literal_2043896[p4_addedKey__49_comb[47:40]];
  assign p4_array_index_2047959_comb = p3_literal_2043896[p4_addedKey__49_comb[39:32]];
  assign p4_array_index_2047960_comb = p3_literal_2043896[p4_addedKey__49_comb[31:24]];
  assign p4_array_index_2047961_comb = p3_literal_2043896[p4_addedKey__49_comb[23:16]];
  assign p4_array_index_2047962_comb = p3_literal_2043896[p4_addedKey__49_comb[15:8]];
  assign p4_array_index_2047964_comb = p3_literal_2043910[p4_array_index_2047948_comb];
  assign p4_array_index_2047965_comb = p3_literal_2043912[p4_array_index_2047949_comb];
  assign p4_array_index_2047966_comb = p3_literal_2043914[p4_array_index_2047950_comb];
  assign p4_array_index_2047967_comb = p3_literal_2043916[p4_array_index_2047951_comb];
  assign p4_array_index_2047968_comb = p3_literal_2043918[p4_array_index_2047952_comb];
  assign p4_array_index_2047969_comb = p3_literal_2043920[p4_array_index_2047953_comb];
  assign p4_array_index_2047970_comb = p3_literal_2043896[p4_addedKey__49_comb[79:72]];
  assign p4_array_index_2047972_comb = p3_literal_2043896[p4_addedKey__49_comb[63:56]];
  assign p4_res7__544_comb = p4_array_index_2047964_comb ^ p4_array_index_2047965_comb ^ p4_array_index_2047966_comb ^ p4_array_index_2047967_comb ^ p4_array_index_2047968_comb ^ p4_array_index_2047969_comb ^ p4_array_index_2047970_comb ^ p3_literal_2043923[p4_array_index_2047955_comb] ^ p4_array_index_2047972_comb ^ p3_literal_2043920[p4_array_index_2047957_comb] ^ p3_literal_2043918[p4_array_index_2047958_comb] ^ p3_literal_2043916[p4_array_index_2047959_comb] ^ p3_literal_2043914[p4_array_index_2047960_comb] ^ p3_literal_2043912[p4_array_index_2047961_comb] ^ p3_literal_2043910[p4_array_index_2047962_comb] ^ p3_literal_2043896[p4_addedKey__49_comb[7:0]];
  assign p4_array_index_2047981_comb = p3_literal_2043910[p4_res7__544_comb];
  assign p4_array_index_2047982_comb = p3_literal_2043912[p4_array_index_2047948_comb];
  assign p4_array_index_2047983_comb = p3_literal_2043914[p4_array_index_2047949_comb];
  assign p4_array_index_2047984_comb = p3_literal_2043916[p4_array_index_2047950_comb];
  assign p4_array_index_2047985_comb = p3_literal_2043918[p4_array_index_2047951_comb];
  assign p4_array_index_2047986_comb = p3_literal_2043920[p4_array_index_2047952_comb];
  assign p4_res7__546_comb = p4_array_index_2047981_comb ^ p4_array_index_2047982_comb ^ p4_array_index_2047983_comb ^ p4_array_index_2047984_comb ^ p4_array_index_2047985_comb ^ p4_array_index_2047986_comb ^ p4_array_index_2047953_comb ^ p3_literal_2043923[p4_array_index_2047970_comb] ^ p4_array_index_2047955_comb ^ p3_literal_2043920[p4_array_index_2047972_comb] ^ p3_literal_2043918[p4_array_index_2047957_comb] ^ p3_literal_2043916[p4_array_index_2047958_comb] ^ p3_literal_2043914[p4_array_index_2047959_comb] ^ p3_literal_2043912[p4_array_index_2047960_comb] ^ p3_literal_2043910[p4_array_index_2047961_comb] ^ p4_array_index_2047962_comb;
  assign p4_array_index_2047996_comb = p3_literal_2043912[p4_res7__544_comb];
  assign p4_array_index_2047997_comb = p3_literal_2043914[p4_array_index_2047948_comb];
  assign p4_array_index_2047998_comb = p3_literal_2043916[p4_array_index_2047949_comb];
  assign p4_array_index_2047999_comb = p3_literal_2043918[p4_array_index_2047950_comb];
  assign p4_array_index_2048000_comb = p3_literal_2043920[p4_array_index_2047951_comb];
  assign p4_res7__548_comb = p3_literal_2043910[p4_res7__546_comb] ^ p4_array_index_2047996_comb ^ p4_array_index_2047997_comb ^ p4_array_index_2047998_comb ^ p4_array_index_2047999_comb ^ p4_array_index_2048000_comb ^ p4_array_index_2047952_comb ^ p3_literal_2043923[p4_array_index_2047953_comb] ^ p4_array_index_2047970_comb ^ p3_literal_2043920[p4_array_index_2047955_comb] ^ p3_literal_2043918[p4_array_index_2047972_comb] ^ p3_literal_2043916[p4_array_index_2047957_comb] ^ p3_literal_2043914[p4_array_index_2047958_comb] ^ p3_literal_2043912[p4_array_index_2047959_comb] ^ p3_literal_2043910[p4_array_index_2047960_comb] ^ p4_array_index_2047961_comb;
  assign p4_array_index_2048010_comb = p3_literal_2043912[p4_res7__546_comb];
  assign p4_array_index_2048011_comb = p3_literal_2043914[p4_res7__544_comb];
  assign p4_array_index_2048012_comb = p3_literal_2043916[p4_array_index_2047948_comb];
  assign p4_array_index_2048013_comb = p3_literal_2043918[p4_array_index_2047949_comb];
  assign p4_array_index_2048014_comb = p3_literal_2043920[p4_array_index_2047950_comb];
  assign p4_res7__550_comb = p3_literal_2043910[p4_res7__548_comb] ^ p4_array_index_2048010_comb ^ p4_array_index_2048011_comb ^ p4_array_index_2048012_comb ^ p4_array_index_2048013_comb ^ p4_array_index_2048014_comb ^ p4_array_index_2047951_comb ^ p3_literal_2043923[p4_array_index_2047952_comb] ^ p4_array_index_2047953_comb ^ p3_literal_2043920[p4_array_index_2047970_comb] ^ p3_literal_2043918[p4_array_index_2047955_comb] ^ p3_literal_2043916[p4_array_index_2047972_comb] ^ p3_literal_2043914[p4_array_index_2047957_comb] ^ p3_literal_2043912[p4_array_index_2047958_comb] ^ p3_literal_2043910[p4_array_index_2047959_comb] ^ p4_array_index_2047960_comb;
  assign p4_array_index_2048025_comb = p3_literal_2043914[p4_res7__546_comb];
  assign p4_array_index_2048026_comb = p3_literal_2043916[p4_res7__544_comb];
  assign p4_array_index_2048027_comb = p3_literal_2043918[p4_array_index_2047948_comb];
  assign p4_array_index_2048028_comb = p3_literal_2043920[p4_array_index_2047949_comb];
  assign p4_res7__552_comb = p3_literal_2043910[p4_res7__550_comb] ^ p3_literal_2043912[p4_res7__548_comb] ^ p4_array_index_2048025_comb ^ p4_array_index_2048026_comb ^ p4_array_index_2048027_comb ^ p4_array_index_2048028_comb ^ p4_array_index_2047950_comb ^ p3_literal_2043923[p4_array_index_2047951_comb] ^ p4_array_index_2047952_comb ^ p4_array_index_2047969_comb ^ p3_literal_2043918[p4_array_index_2047970_comb] ^ p3_literal_2043916[p4_array_index_2047955_comb] ^ p3_literal_2043914[p4_array_index_2047972_comb] ^ p3_literal_2043912[p4_array_index_2047957_comb] ^ p3_literal_2043910[p4_array_index_2047958_comb] ^ p4_array_index_2047959_comb;
  assign p4_array_index_2048038_comb = p3_literal_2043914[p4_res7__548_comb];
  assign p4_array_index_2048039_comb = p3_literal_2043916[p4_res7__546_comb];
  assign p4_array_index_2048040_comb = p3_literal_2043918[p4_res7__544_comb];
  assign p4_array_index_2048041_comb = p3_literal_2043920[p4_array_index_2047948_comb];
  assign p4_res7__554_comb = p3_literal_2043910[p4_res7__552_comb] ^ p3_literal_2043912[p4_res7__550_comb] ^ p4_array_index_2048038_comb ^ p4_array_index_2048039_comb ^ p4_array_index_2048040_comb ^ p4_array_index_2048041_comb ^ p4_array_index_2047949_comb ^ p3_literal_2043923[p4_array_index_2047950_comb] ^ p4_array_index_2047951_comb ^ p4_array_index_2047986_comb ^ p3_literal_2043918[p4_array_index_2047953_comb] ^ p3_literal_2043916[p4_array_index_2047970_comb] ^ p3_literal_2043914[p4_array_index_2047955_comb] ^ p3_literal_2043912[p4_array_index_2047972_comb] ^ p3_literal_2043910[p4_array_index_2047957_comb] ^ p4_array_index_2047958_comb;
  assign p4_array_index_2048052_comb = p3_literal_2043916[p4_res7__548_comb];
  assign p4_array_index_2048053_comb = p3_literal_2043918[p4_res7__546_comb];
  assign p4_array_index_2048054_comb = p3_literal_2043920[p4_res7__544_comb];
  assign p4_res7__556_comb = p3_literal_2043910[p4_res7__554_comb] ^ p3_literal_2043912[p4_res7__552_comb] ^ p3_literal_2043914[p4_res7__550_comb] ^ p4_array_index_2048052_comb ^ p4_array_index_2048053_comb ^ p4_array_index_2048054_comb ^ p4_array_index_2047948_comb ^ p3_literal_2043923[p4_array_index_2047949_comb] ^ p4_array_index_2047950_comb ^ p4_array_index_2048000_comb ^ p4_array_index_2047968_comb ^ p3_literal_2043916[p4_array_index_2047953_comb] ^ p3_literal_2043914[p4_array_index_2047970_comb] ^ p3_literal_2043912[p4_array_index_2047955_comb] ^ p3_literal_2043910[p4_array_index_2047972_comb] ^ p4_array_index_2047957_comb;
  assign p4_array_index_2048064_comb = p3_literal_2043916[p4_res7__550_comb];
  assign p4_array_index_2048065_comb = p3_literal_2043918[p4_res7__548_comb];
  assign p4_array_index_2048066_comb = p3_literal_2043920[p4_res7__546_comb];
  assign p4_res7__558_comb = p3_literal_2043910[p4_res7__556_comb] ^ p3_literal_2043912[p4_res7__554_comb] ^ p3_literal_2043914[p4_res7__552_comb] ^ p4_array_index_2048064_comb ^ p4_array_index_2048065_comb ^ p4_array_index_2048066_comb ^ p4_res7__544_comb ^ p3_literal_2043923[p4_array_index_2047948_comb] ^ p4_array_index_2047949_comb ^ p4_array_index_2048014_comb ^ p4_array_index_2047985_comb ^ p3_literal_2043916[p4_array_index_2047952_comb] ^ p3_literal_2043914[p4_array_index_2047953_comb] ^ p3_literal_2043912[p4_array_index_2047970_comb] ^ p3_literal_2043910[p4_array_index_2047955_comb] ^ p4_array_index_2047972_comb;
  assign p4_array_index_2048077_comb = p3_literal_2043918[p4_res7__550_comb];
  assign p4_array_index_2048078_comb = p3_literal_2043920[p4_res7__548_comb];
  assign p4_res7__560_comb = p3_literal_2043910[p4_res7__558_comb] ^ p3_literal_2043912[p4_res7__556_comb] ^ p3_literal_2043914[p4_res7__554_comb] ^ p3_literal_2043916[p4_res7__552_comb] ^ p4_array_index_2048077_comb ^ p4_array_index_2048078_comb ^ p4_res7__546_comb ^ p3_literal_2043923[p4_res7__544_comb] ^ p4_array_index_2047948_comb ^ p4_array_index_2048028_comb ^ p4_array_index_2047999_comb ^ p4_array_index_2047967_comb ^ p3_literal_2043914[p4_array_index_2047952_comb] ^ p3_literal_2043912[p4_array_index_2047953_comb] ^ p3_literal_2043910[p4_array_index_2047970_comb] ^ p4_array_index_2047955_comb;
  assign p4_array_index_2048088_comb = p3_literal_2043918[p4_res7__552_comb];
  assign p4_array_index_2048089_comb = p3_literal_2043920[p4_res7__550_comb];
  assign p4_res7__562_comb = p3_literal_2043910[p4_res7__560_comb] ^ p3_literal_2043912[p4_res7__558_comb] ^ p3_literal_2043914[p4_res7__556_comb] ^ p3_literal_2043916[p4_res7__554_comb] ^ p4_array_index_2048088_comb ^ p4_array_index_2048089_comb ^ p4_res7__548_comb ^ p3_literal_2043923[p4_res7__546_comb] ^ p4_res7__544_comb ^ p4_array_index_2048041_comb ^ p4_array_index_2048013_comb ^ p4_array_index_2047984_comb ^ p3_literal_2043914[p4_array_index_2047951_comb] ^ p3_literal_2043912[p4_array_index_2047952_comb] ^ p3_literal_2043910[p4_array_index_2047953_comb] ^ p4_array_index_2047970_comb;
  assign p4_array_index_2048100_comb = p3_literal_2043920[p4_res7__552_comb];
  assign p4_res7__564_comb = p3_literal_2043910[p4_res7__562_comb] ^ p3_literal_2043912[p4_res7__560_comb] ^ p3_literal_2043914[p4_res7__558_comb] ^ p3_literal_2043916[p4_res7__556_comb] ^ p3_literal_2043918[p4_res7__554_comb] ^ p4_array_index_2048100_comb ^ p4_res7__550_comb ^ p3_literal_2043923[p4_res7__548_comb] ^ p4_res7__546_comb ^ p4_array_index_2048054_comb ^ p4_array_index_2048027_comb ^ p4_array_index_2047998_comb ^ p4_array_index_2047966_comb ^ p3_literal_2043912[p4_array_index_2047951_comb] ^ p3_literal_2043910[p4_array_index_2047952_comb] ^ p4_array_index_2047953_comb;
  assign p4_array_index_2048110_comb = p3_literal_2043920[p4_res7__554_comb];
  assign p4_res7__566_comb = p3_literal_2043910[p4_res7__564_comb] ^ p3_literal_2043912[p4_res7__562_comb] ^ p3_literal_2043914[p4_res7__560_comb] ^ p3_literal_2043916[p4_res7__558_comb] ^ p3_literal_2043918[p4_res7__556_comb] ^ p4_array_index_2048110_comb ^ p4_res7__552_comb ^ p3_literal_2043923[p4_res7__550_comb] ^ p4_res7__548_comb ^ p4_array_index_2048066_comb ^ p4_array_index_2048040_comb ^ p4_array_index_2048012_comb ^ p4_array_index_2047983_comb ^ p3_literal_2043912[p4_array_index_2047950_comb] ^ p3_literal_2043910[p4_array_index_2047951_comb] ^ p4_array_index_2047952_comb;
  assign p4_array_index_2048115_comb = p3_literal_2043910[p4_res7__566_comb];
  assign p4_array_index_2048116_comb = p3_literal_2043912[p4_res7__564_comb];
  assign p4_array_index_2048117_comb = p3_literal_2043914[p4_res7__562_comb];
  assign p4_array_index_2048118_comb = p3_literal_2043916[p4_res7__560_comb];
  assign p4_array_index_2048119_comb = p3_literal_2043918[p4_res7__558_comb];
  assign p4_array_index_2048120_comb = p3_literal_2043920[p4_res7__556_comb];
  assign p4_array_index_2048121_comb = p3_literal_2043923[p4_res7__552_comb];
  assign p4_array_index_2048122_comb = p3_literal_2043910[p4_array_index_2047950_comb];

  // Registers for pipe stage 4:
  reg [127:0] p4_encoded;
  reg [127:0] p4_bit_slice_2043893;
  reg [127:0] p4_bit_slice_2044119;
  reg [127:0] p4_k3;
  reg [127:0] p4_k2;
  reg [127:0] p4_k5;
  reg [127:0] p4_k4;
  reg [127:0] p4_xor_2047932;
  reg [7:0] p4_array_index_2047948;
  reg [7:0] p4_array_index_2047949;
  reg [7:0] p4_array_index_2047950;
  reg [7:0] p4_array_index_2047951;
  reg [7:0] p4_array_index_2047964;
  reg [7:0] p4_array_index_2047965;
  reg [7:0] p4_res7__544;
  reg [7:0] p4_array_index_2047981;
  reg [7:0] p4_array_index_2047982;
  reg [7:0] p4_res7__546;
  reg [7:0] p4_array_index_2047996;
  reg [7:0] p4_array_index_2047997;
  reg [7:0] p4_res7__548;
  reg [7:0] p4_array_index_2048010;
  reg [7:0] p4_array_index_2048011;
  reg [7:0] p4_res7__550;
  reg [7:0] p4_array_index_2048025;
  reg [7:0] p4_array_index_2048026;
  reg [7:0] p4_res7__552;
  reg [7:0] p4_array_index_2048038;
  reg [7:0] p4_array_index_2048039;
  reg [7:0] p4_res7__554;
  reg [7:0] p4_array_index_2048052;
  reg [7:0] p4_array_index_2048053;
  reg [7:0] p4_res7__556;
  reg [7:0] p4_array_index_2048064;
  reg [7:0] p4_array_index_2048065;
  reg [7:0] p4_res7__558;
  reg [7:0] p4_array_index_2048077;
  reg [7:0] p4_array_index_2048078;
  reg [7:0] p4_res7__560;
  reg [7:0] p4_array_index_2048088;
  reg [7:0] p4_array_index_2048089;
  reg [7:0] p4_res7__562;
  reg [7:0] p4_array_index_2048100;
  reg [7:0] p4_res7__564;
  reg [7:0] p4_array_index_2048110;
  reg [7:0] p4_res7__566;
  reg [7:0] p4_array_index_2048115;
  reg [7:0] p4_array_index_2048116;
  reg [7:0] p4_array_index_2048117;
  reg [7:0] p4_array_index_2048118;
  reg [7:0] p4_array_index_2048119;
  reg [7:0] p4_array_index_2048120;
  reg [7:0] p4_array_index_2048121;
  reg [7:0] p4_array_index_2048122;
  reg [7:0] p5_literal_2043896[256];
  reg [7:0] p5_literal_2043910[256];
  reg [7:0] p5_literal_2043912[256];
  reg [7:0] p5_literal_2043914[256];
  reg [7:0] p5_literal_2043916[256];
  reg [7:0] p5_literal_2043918[256];
  reg [7:0] p5_literal_2043920[256];
  reg [7:0] p5_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p4_encoded <= p3_encoded;
    p4_bit_slice_2043893 <= p3_bit_slice_2043893;
    p4_bit_slice_2044119 <= p3_bit_slice_2044119;
    p4_k3 <= p3_k3;
    p4_k2 <= p3_k2;
    p4_k5 <= p4_k5_comb;
    p4_k4 <= p4_k4_comb;
    p4_xor_2047932 <= p4_xor_2047932_comb;
    p4_array_index_2047948 <= p4_array_index_2047948_comb;
    p4_array_index_2047949 <= p4_array_index_2047949_comb;
    p4_array_index_2047950 <= p4_array_index_2047950_comb;
    p4_array_index_2047951 <= p4_array_index_2047951_comb;
    p4_array_index_2047964 <= p4_array_index_2047964_comb;
    p4_array_index_2047965 <= p4_array_index_2047965_comb;
    p4_res7__544 <= p4_res7__544_comb;
    p4_array_index_2047981 <= p4_array_index_2047981_comb;
    p4_array_index_2047982 <= p4_array_index_2047982_comb;
    p4_res7__546 <= p4_res7__546_comb;
    p4_array_index_2047996 <= p4_array_index_2047996_comb;
    p4_array_index_2047997 <= p4_array_index_2047997_comb;
    p4_res7__548 <= p4_res7__548_comb;
    p4_array_index_2048010 <= p4_array_index_2048010_comb;
    p4_array_index_2048011 <= p4_array_index_2048011_comb;
    p4_res7__550 <= p4_res7__550_comb;
    p4_array_index_2048025 <= p4_array_index_2048025_comb;
    p4_array_index_2048026 <= p4_array_index_2048026_comb;
    p4_res7__552 <= p4_res7__552_comb;
    p4_array_index_2048038 <= p4_array_index_2048038_comb;
    p4_array_index_2048039 <= p4_array_index_2048039_comb;
    p4_res7__554 <= p4_res7__554_comb;
    p4_array_index_2048052 <= p4_array_index_2048052_comb;
    p4_array_index_2048053 <= p4_array_index_2048053_comb;
    p4_res7__556 <= p4_res7__556_comb;
    p4_array_index_2048064 <= p4_array_index_2048064_comb;
    p4_array_index_2048065 <= p4_array_index_2048065_comb;
    p4_res7__558 <= p4_res7__558_comb;
    p4_array_index_2048077 <= p4_array_index_2048077_comb;
    p4_array_index_2048078 <= p4_array_index_2048078_comb;
    p4_res7__560 <= p4_res7__560_comb;
    p4_array_index_2048088 <= p4_array_index_2048088_comb;
    p4_array_index_2048089 <= p4_array_index_2048089_comb;
    p4_res7__562 <= p4_res7__562_comb;
    p4_array_index_2048100 <= p4_array_index_2048100_comb;
    p4_res7__564 <= p4_res7__564_comb;
    p4_array_index_2048110 <= p4_array_index_2048110_comb;
    p4_res7__566 <= p4_res7__566_comb;
    p4_array_index_2048115 <= p4_array_index_2048115_comb;
    p4_array_index_2048116 <= p4_array_index_2048116_comb;
    p4_array_index_2048117 <= p4_array_index_2048117_comb;
    p4_array_index_2048118 <= p4_array_index_2048118_comb;
    p4_array_index_2048119 <= p4_array_index_2048119_comb;
    p4_array_index_2048120 <= p4_array_index_2048120_comb;
    p4_array_index_2048121 <= p4_array_index_2048121_comb;
    p4_array_index_2048122 <= p4_array_index_2048122_comb;
    p5_literal_2043896 <= p4_literal_2043896;
    p5_literal_2043910 <= p4_literal_2043910;
    p5_literal_2043912 <= p4_literal_2043912;
    p5_literal_2043914 <= p4_literal_2043914;
    p5_literal_2043916 <= p4_literal_2043916;
    p5_literal_2043918 <= p4_literal_2043918;
    p5_literal_2043920 <= p4_literal_2043920;
    p5_literal_2043923 <= p4_literal_2043923;
  end

  // ===== Pipe stage 5:
  wire [7:0] p5_res7__568_comb;
  wire [7:0] p5_res7__570_comb;
  wire [7:0] p5_res7__572_comb;
  wire [7:0] p5_res7__574_comb;
  wire [127:0] p5_res__17_comb;
  wire [127:0] p5_xor_2048274_comb;
  wire [127:0] p5_addedKey__50_comb;
  wire [7:0] p5_array_index_2048290_comb;
  wire [7:0] p5_array_index_2048291_comb;
  wire [7:0] p5_array_index_2048292_comb;
  wire [7:0] p5_array_index_2048293_comb;
  wire [7:0] p5_array_index_2048294_comb;
  wire [7:0] p5_array_index_2048295_comb;
  wire [7:0] p5_array_index_2048297_comb;
  wire [7:0] p5_array_index_2048299_comb;
  wire [7:0] p5_array_index_2048300_comb;
  wire [7:0] p5_array_index_2048301_comb;
  wire [7:0] p5_array_index_2048302_comb;
  wire [7:0] p5_array_index_2048303_comb;
  wire [7:0] p5_array_index_2048304_comb;
  wire [7:0] p5_array_index_2048306_comb;
  wire [7:0] p5_array_index_2048307_comb;
  wire [7:0] p5_array_index_2048308_comb;
  wire [7:0] p5_array_index_2048309_comb;
  wire [7:0] p5_array_index_2048310_comb;
  wire [7:0] p5_array_index_2048311_comb;
  wire [7:0] p5_array_index_2048312_comb;
  wire [7:0] p5_array_index_2048314_comb;
  wire [7:0] p5_res7__576_comb;
  wire [7:0] p5_array_index_2048323_comb;
  wire [7:0] p5_array_index_2048324_comb;
  wire [7:0] p5_array_index_2048325_comb;
  wire [7:0] p5_array_index_2048326_comb;
  wire [7:0] p5_array_index_2048327_comb;
  wire [7:0] p5_array_index_2048328_comb;
  wire [7:0] p5_res7__578_comb;
  wire [7:0] p5_array_index_2048338_comb;
  wire [7:0] p5_array_index_2048339_comb;
  wire [7:0] p5_array_index_2048340_comb;
  wire [7:0] p5_array_index_2048341_comb;
  wire [7:0] p5_array_index_2048342_comb;
  wire [7:0] p5_res7__580_comb;
  wire [7:0] p5_array_index_2048352_comb;
  wire [7:0] p5_array_index_2048353_comb;
  wire [7:0] p5_array_index_2048354_comb;
  wire [7:0] p5_array_index_2048355_comb;
  wire [7:0] p5_array_index_2048356_comb;
  wire [7:0] p5_res7__582_comb;
  wire [7:0] p5_array_index_2048367_comb;
  wire [7:0] p5_array_index_2048368_comb;
  wire [7:0] p5_array_index_2048369_comb;
  wire [7:0] p5_array_index_2048370_comb;
  wire [7:0] p5_res7__584_comb;
  wire [7:0] p5_array_index_2048380_comb;
  wire [7:0] p5_array_index_2048381_comb;
  wire [7:0] p5_array_index_2048382_comb;
  wire [7:0] p5_array_index_2048383_comb;
  wire [7:0] p5_res7__586_comb;
  wire [7:0] p5_array_index_2048394_comb;
  wire [7:0] p5_array_index_2048395_comb;
  wire [7:0] p5_array_index_2048396_comb;
  wire [7:0] p5_res7__588_comb;
  wire [7:0] p5_array_index_2048406_comb;
  wire [7:0] p5_array_index_2048407_comb;
  wire [7:0] p5_array_index_2048408_comb;
  wire [7:0] p5_res7__590_comb;
  wire [7:0] p5_array_index_2048419_comb;
  wire [7:0] p5_array_index_2048420_comb;
  wire [7:0] p5_res7__592_comb;
  wire [7:0] p5_array_index_2048430_comb;
  wire [7:0] p5_array_index_2048431_comb;
  wire [7:0] p5_res7__594_comb;
  wire [7:0] p5_array_index_2048442_comb;
  wire [7:0] p5_res7__596_comb;
  wire [7:0] p5_array_index_2048452_comb;
  wire [7:0] p5_res7__598_comb;
  wire [7:0] p5_res7__600_comb;
  wire [7:0] p5_res7__602_comb;
  wire [7:0] p5_res7__604_comb;
  wire [7:0] p5_res7__606_comb;
  wire [127:0] p5_res__18_comb;
  wire [127:0] p5_xor_2048492_comb;
  wire [127:0] p5_addedKey__51_comb;
  wire [7:0] p5_array_index_2048508_comb;
  wire [7:0] p5_array_index_2048509_comb;
  wire [7:0] p5_array_index_2048510_comb;
  wire [7:0] p5_array_index_2048511_comb;
  wire [7:0] p5_array_index_2048512_comb;
  wire [7:0] p5_array_index_2048513_comb;
  wire [7:0] p5_array_index_2048515_comb;
  wire [7:0] p5_array_index_2048517_comb;
  wire [7:0] p5_array_index_2048518_comb;
  wire [7:0] p5_array_index_2048519_comb;
  wire [7:0] p5_array_index_2048520_comb;
  wire [7:0] p5_array_index_2048521_comb;
  wire [7:0] p5_array_index_2048522_comb;
  wire [7:0] p5_array_index_2048524_comb;
  wire [7:0] p5_array_index_2048525_comb;
  wire [7:0] p5_array_index_2048526_comb;
  wire [7:0] p5_array_index_2048527_comb;
  wire [7:0] p5_array_index_2048528_comb;
  wire [7:0] p5_array_index_2048529_comb;
  wire [7:0] p5_array_index_2048530_comb;
  wire [7:0] p5_array_index_2048532_comb;
  wire [7:0] p5_res7__608_comb;
  wire [7:0] p5_array_index_2048541_comb;
  wire [7:0] p5_array_index_2048542_comb;
  wire [7:0] p5_array_index_2048543_comb;
  wire [7:0] p5_array_index_2048544_comb;
  wire [7:0] p5_array_index_2048545_comb;
  wire [7:0] p5_array_index_2048546_comb;
  wire [7:0] p5_res7__610_comb;
  wire [7:0] p5_array_index_2048556_comb;
  wire [7:0] p5_array_index_2048557_comb;
  wire [7:0] p5_array_index_2048558_comb;
  wire [7:0] p5_array_index_2048559_comb;
  wire [7:0] p5_array_index_2048560_comb;
  wire [7:0] p5_res7__612_comb;
  wire [7:0] p5_array_index_2048570_comb;
  wire [7:0] p5_array_index_2048571_comb;
  wire [7:0] p5_array_index_2048572_comb;
  wire [7:0] p5_array_index_2048573_comb;
  wire [7:0] p5_array_index_2048574_comb;
  wire [7:0] p5_res7__614_comb;
  wire [7:0] p5_array_index_2048585_comb;
  wire [7:0] p5_array_index_2048586_comb;
  wire [7:0] p5_array_index_2048587_comb;
  wire [7:0] p5_array_index_2048588_comb;
  wire [7:0] p5_res7__616_comb;
  wire [7:0] p5_array_index_2048598_comb;
  wire [7:0] p5_array_index_2048599_comb;
  wire [7:0] p5_array_index_2048600_comb;
  wire [7:0] p5_array_index_2048601_comb;
  wire [7:0] p5_res7__618_comb;
  wire [7:0] p5_array_index_2048612_comb;
  wire [7:0] p5_array_index_2048613_comb;
  wire [7:0] p5_array_index_2048614_comb;
  wire [7:0] p5_res7__620_comb;
  wire [7:0] p5_array_index_2048624_comb;
  wire [7:0] p5_array_index_2048625_comb;
  wire [7:0] p5_array_index_2048626_comb;
  wire [7:0] p5_res7__622_comb;
  wire [7:0] p5_array_index_2048637_comb;
  wire [7:0] p5_array_index_2048638_comb;
  wire [7:0] p5_res7__624_comb;
  wire [7:0] p5_array_index_2048648_comb;
  wire [7:0] p5_array_index_2048649_comb;
  wire [7:0] p5_res7__626_comb;
  wire [7:0] p5_array_index_2048660_comb;
  wire [7:0] p5_res7__628_comb;
  wire [7:0] p5_array_index_2048670_comb;
  wire [7:0] p5_res7__630_comb;
  wire [7:0] p5_res7__632_comb;
  wire [7:0] p5_res7__634_comb;
  wire [7:0] p5_res7__636_comb;
  wire [7:0] p5_res7__638_comb;
  wire [127:0] p5_res__19_comb;
  wire [127:0] p5_xor_2048710_comb;
  wire [127:0] p5_addedKey__52_comb;
  wire [7:0] p5_array_index_2048726_comb;
  wire [7:0] p5_array_index_2048727_comb;
  wire [7:0] p5_array_index_2048728_comb;
  wire [7:0] p5_array_index_2048729_comb;
  wire [7:0] p5_array_index_2048730_comb;
  wire [7:0] p5_array_index_2048731_comb;
  wire [7:0] p5_array_index_2048733_comb;
  wire [7:0] p5_array_index_2048735_comb;
  wire [7:0] p5_array_index_2048736_comb;
  wire [7:0] p5_array_index_2048737_comb;
  wire [7:0] p5_array_index_2048738_comb;
  wire [7:0] p5_array_index_2048739_comb;
  wire [7:0] p5_array_index_2048740_comb;
  wire [7:0] p5_array_index_2048742_comb;
  wire [7:0] p5_array_index_2048743_comb;
  wire [7:0] p5_array_index_2048744_comb;
  wire [7:0] p5_array_index_2048745_comb;
  wire [7:0] p5_array_index_2048746_comb;
  wire [7:0] p5_array_index_2048747_comb;
  wire [7:0] p5_array_index_2048748_comb;
  wire [7:0] p5_array_index_2048750_comb;
  wire [7:0] p5_res7__640_comb;
  wire [7:0] p5_array_index_2048759_comb;
  wire [7:0] p5_array_index_2048760_comb;
  wire [7:0] p5_array_index_2048761_comb;
  wire [7:0] p5_array_index_2048762_comb;
  wire [7:0] p5_array_index_2048763_comb;
  wire [7:0] p5_array_index_2048764_comb;
  wire [7:0] p5_res7__642_comb;
  wire [7:0] p5_array_index_2048774_comb;
  wire [7:0] p5_array_index_2048775_comb;
  wire [7:0] p5_array_index_2048776_comb;
  wire [7:0] p5_array_index_2048777_comb;
  wire [7:0] p5_array_index_2048778_comb;
  wire [7:0] p5_res7__644_comb;
  wire [7:0] p5_array_index_2048788_comb;
  wire [7:0] p5_array_index_2048789_comb;
  wire [7:0] p5_array_index_2048790_comb;
  wire [7:0] p5_array_index_2048791_comb;
  wire [7:0] p5_array_index_2048792_comb;
  wire [7:0] p5_res7__646_comb;
  wire [7:0] p5_array_index_2048803_comb;
  wire [7:0] p5_array_index_2048804_comb;
  wire [7:0] p5_array_index_2048805_comb;
  wire [7:0] p5_array_index_2048806_comb;
  wire [7:0] p5_res7__648_comb;
  wire [7:0] p5_array_index_2048816_comb;
  wire [7:0] p5_array_index_2048817_comb;
  wire [7:0] p5_array_index_2048818_comb;
  wire [7:0] p5_array_index_2048819_comb;
  wire [7:0] p5_res7__650_comb;
  wire [7:0] p5_array_index_2048830_comb;
  wire [7:0] p5_array_index_2048831_comb;
  wire [7:0] p5_array_index_2048832_comb;
  wire [7:0] p5_res7__652_comb;
  wire [7:0] p5_array_index_2048842_comb;
  wire [7:0] p5_array_index_2048843_comb;
  wire [7:0] p5_array_index_2048844_comb;
  wire [7:0] p5_res7__654_comb;
  wire [7:0] p5_array_index_2048855_comb;
  wire [7:0] p5_array_index_2048856_comb;
  wire [7:0] p5_res7__656_comb;
  wire [7:0] p5_array_index_2048866_comb;
  wire [7:0] p5_array_index_2048867_comb;
  wire [7:0] p5_res7__658_comb;
  wire [7:0] p5_array_index_2048878_comb;
  wire [7:0] p5_res7__660_comb;
  wire [7:0] p5_array_index_2048888_comb;
  wire [7:0] p5_res7__662_comb;
  wire [7:0] p5_res7__664_comb;
  wire [7:0] p5_res7__666_comb;
  wire [7:0] p5_res7__668_comb;
  wire [7:0] p5_res7__670_comb;
  wire [127:0] p5_res__20_comb;
  wire [127:0] p5_xor_2048928_comb;
  wire [127:0] p5_addedKey__53_comb;
  wire [7:0] p5_array_index_2048944_comb;
  wire [7:0] p5_array_index_2048945_comb;
  wire [7:0] p5_array_index_2048946_comb;
  wire [7:0] p5_array_index_2048947_comb;
  wire [7:0] p5_array_index_2048948_comb;
  wire [7:0] p5_array_index_2048949_comb;
  wire [7:0] p5_array_index_2048951_comb;
  wire [7:0] p5_array_index_2048953_comb;
  wire [7:0] p5_array_index_2048954_comb;
  wire [7:0] p5_array_index_2048955_comb;
  wire [7:0] p5_array_index_2048956_comb;
  wire [7:0] p5_array_index_2048957_comb;
  wire [7:0] p5_array_index_2048958_comb;
  wire [7:0] p5_array_index_2048960_comb;
  wire [7:0] p5_array_index_2048961_comb;
  wire [7:0] p5_array_index_2048962_comb;
  wire [7:0] p5_array_index_2048963_comb;
  wire [7:0] p5_array_index_2048964_comb;
  wire [7:0] p5_array_index_2048965_comb;
  wire [7:0] p5_array_index_2048966_comb;
  wire [7:0] p5_array_index_2048968_comb;
  wire [7:0] p5_res7__672_comb;
  wire [7:0] p5_array_index_2048977_comb;
  wire [7:0] p5_array_index_2048978_comb;
  wire [7:0] p5_array_index_2048979_comb;
  wire [7:0] p5_array_index_2048980_comb;
  wire [7:0] p5_array_index_2048981_comb;
  wire [7:0] p5_array_index_2048982_comb;
  wire [7:0] p5_res7__674_comb;
  wire [7:0] p5_array_index_2048992_comb;
  wire [7:0] p5_array_index_2048993_comb;
  wire [7:0] p5_array_index_2048994_comb;
  wire [7:0] p5_array_index_2048995_comb;
  wire [7:0] p5_array_index_2048996_comb;
  wire [7:0] p5_res7__676_comb;
  wire [7:0] p5_array_index_2049006_comb;
  wire [7:0] p5_array_index_2049007_comb;
  wire [7:0] p5_array_index_2049008_comb;
  wire [7:0] p5_array_index_2049009_comb;
  wire [7:0] p5_array_index_2049010_comb;
  wire [7:0] p5_res7__678_comb;
  wire [7:0] p5_array_index_2049021_comb;
  wire [7:0] p5_array_index_2049022_comb;
  wire [7:0] p5_array_index_2049023_comb;
  wire [7:0] p5_array_index_2049024_comb;
  wire [7:0] p5_res7__680_comb;
  wire [7:0] p5_array_index_2049034_comb;
  wire [7:0] p5_array_index_2049035_comb;
  wire [7:0] p5_array_index_2049036_comb;
  wire [7:0] p5_array_index_2049037_comb;
  wire [7:0] p5_res7__682_comb;
  wire [7:0] p5_array_index_2049048_comb;
  wire [7:0] p5_array_index_2049049_comb;
  wire [7:0] p5_array_index_2049050_comb;
  wire [7:0] p5_res7__684_comb;
  wire [7:0] p5_array_index_2049060_comb;
  wire [7:0] p5_array_index_2049061_comb;
  wire [7:0] p5_array_index_2049062_comb;
  wire [7:0] p5_res7__686_comb;
  wire [7:0] p5_array_index_2049073_comb;
  wire [7:0] p5_array_index_2049074_comb;
  wire [7:0] p5_res7__688_comb;
  wire [7:0] p5_array_index_2049084_comb;
  wire [7:0] p5_array_index_2049085_comb;
  wire [7:0] p5_res7__690_comb;
  wire [7:0] p5_array_index_2049096_comb;
  wire [7:0] p5_res7__692_comb;
  wire [7:0] p5_array_index_2049106_comb;
  wire [7:0] p5_res7__694_comb;
  wire [7:0] p5_res7__696_comb;
  wire [7:0] p5_res7__698_comb;
  wire [7:0] p5_res7__700_comb;
  wire [7:0] p5_res7__702_comb;
  wire [127:0] p5_res__21_comb;
  wire [127:0] p5_xor_2049146_comb;
  wire [127:0] p5_addedKey__54_comb;
  wire [7:0] p5_array_index_2049162_comb;
  wire [7:0] p5_array_index_2049163_comb;
  wire [7:0] p5_array_index_2049164_comb;
  wire [7:0] p5_array_index_2049165_comb;
  wire [7:0] p5_array_index_2049166_comb;
  wire [7:0] p5_array_index_2049167_comb;
  wire [7:0] p5_array_index_2049169_comb;
  wire [7:0] p5_array_index_2049171_comb;
  wire [7:0] p5_array_index_2049172_comb;
  wire [7:0] p5_array_index_2049173_comb;
  wire [7:0] p5_array_index_2049174_comb;
  wire [7:0] p5_array_index_2049175_comb;
  wire [7:0] p5_array_index_2049176_comb;
  wire [7:0] p5_array_index_2049178_comb;
  wire [7:0] p5_array_index_2049179_comb;
  wire [7:0] p5_array_index_2049180_comb;
  wire [7:0] p5_array_index_2049181_comb;
  wire [7:0] p5_array_index_2049182_comb;
  wire [7:0] p5_array_index_2049183_comb;
  wire [7:0] p5_array_index_2049184_comb;
  wire [7:0] p5_array_index_2049186_comb;
  wire [7:0] p5_res7__704_comb;
  wire [7:0] p5_array_index_2049195_comb;
  wire [7:0] p5_array_index_2049196_comb;
  wire [7:0] p5_array_index_2049197_comb;
  wire [7:0] p5_array_index_2049198_comb;
  wire [7:0] p5_array_index_2049199_comb;
  wire [7:0] p5_array_index_2049200_comb;
  wire [7:0] p5_res7__706_comb;
  wire [7:0] p5_array_index_2049210_comb;
  wire [7:0] p5_array_index_2049211_comb;
  wire [7:0] p5_array_index_2049212_comb;
  wire [7:0] p5_array_index_2049213_comb;
  wire [7:0] p5_array_index_2049214_comb;
  wire [7:0] p5_res7__708_comb;
  assign p5_res7__568_comb = p4_array_index_2048115 ^ p4_array_index_2048116 ^ p4_array_index_2048117 ^ p4_array_index_2048118 ^ p4_array_index_2048119 ^ p4_array_index_2048120 ^ p4_res7__554 ^ p4_array_index_2048121 ^ p4_res7__550 ^ p4_array_index_2048078 ^ p4_array_index_2048053 ^ p4_array_index_2048026 ^ p4_array_index_2047997 ^ p4_array_index_2047965 ^ p4_array_index_2048122 ^ p4_array_index_2047951;
  assign p5_res7__570_comb = p4_literal_2043910[p5_res7__568_comb] ^ p4_literal_2043912[p4_res7__566] ^ p4_literal_2043914[p4_res7__564] ^ p4_literal_2043916[p4_res7__562] ^ p4_literal_2043918[p4_res7__560] ^ p4_literal_2043920[p4_res7__558] ^ p4_res7__556 ^ p4_literal_2043923[p4_res7__554] ^ p4_res7__552 ^ p4_array_index_2048089 ^ p4_array_index_2048065 ^ p4_array_index_2048039 ^ p4_array_index_2048011 ^ p4_array_index_2047982 ^ p4_literal_2043910[p4_array_index_2047949] ^ p4_array_index_2047950;
  assign p5_res7__572_comb = p4_literal_2043910[p5_res7__570_comb] ^ p4_literal_2043912[p5_res7__568_comb] ^ p4_literal_2043914[p4_res7__566] ^ p4_literal_2043916[p4_res7__564] ^ p4_literal_2043918[p4_res7__562] ^ p4_literal_2043920[p4_res7__560] ^ p4_res7__558 ^ p4_literal_2043923[p4_res7__556] ^ p4_res7__554 ^ p4_array_index_2048100 ^ p4_array_index_2048077 ^ p4_array_index_2048052 ^ p4_array_index_2048025 ^ p4_array_index_2047996 ^ p4_array_index_2047964 ^ p4_array_index_2047949;
  assign p5_res7__574_comb = p4_literal_2043910[p5_res7__572_comb] ^ p4_literal_2043912[p5_res7__570_comb] ^ p4_literal_2043914[p5_res7__568_comb] ^ p4_literal_2043916[p4_res7__566] ^ p4_literal_2043918[p4_res7__564] ^ p4_literal_2043920[p4_res7__562] ^ p4_res7__560 ^ p4_literal_2043923[p4_res7__558] ^ p4_res7__556 ^ p4_array_index_2048110 ^ p4_array_index_2048088 ^ p4_array_index_2048064 ^ p4_array_index_2048038 ^ p4_array_index_2048010 ^ p4_array_index_2047981 ^ p4_array_index_2047948;
  assign p5_res__17_comb = {p5_res7__574_comb, p5_res7__572_comb, p5_res7__570_comb, p5_res7__568_comb, p4_res7__566, p4_res7__564, p4_res7__562, p4_res7__560, p4_res7__558, p4_res7__556, p4_res7__554, p4_res7__552, p4_res7__550, p4_res7__548, p4_res7__546, p4_res7__544};
  assign p5_xor_2048274_comb = p5_res__17_comb ^ p4_k4;
  assign p5_addedKey__50_comb = p5_xor_2048274_comb ^ 128'h9d97_f6ba_bbd2_22da_7e5c_85f3_ead8_2b13;
  assign p5_array_index_2048290_comb = p4_literal_2043896[p5_addedKey__50_comb[127:120]];
  assign p5_array_index_2048291_comb = p4_literal_2043896[p5_addedKey__50_comb[119:112]];
  assign p5_array_index_2048292_comb = p4_literal_2043896[p5_addedKey__50_comb[111:104]];
  assign p5_array_index_2048293_comb = p4_literal_2043896[p5_addedKey__50_comb[103:96]];
  assign p5_array_index_2048294_comb = p4_literal_2043896[p5_addedKey__50_comb[95:88]];
  assign p5_array_index_2048295_comb = p4_literal_2043896[p5_addedKey__50_comb[87:80]];
  assign p5_array_index_2048297_comb = p4_literal_2043896[p5_addedKey__50_comb[71:64]];
  assign p5_array_index_2048299_comb = p4_literal_2043896[p5_addedKey__50_comb[55:48]];
  assign p5_array_index_2048300_comb = p4_literal_2043896[p5_addedKey__50_comb[47:40]];
  assign p5_array_index_2048301_comb = p4_literal_2043896[p5_addedKey__50_comb[39:32]];
  assign p5_array_index_2048302_comb = p4_literal_2043896[p5_addedKey__50_comb[31:24]];
  assign p5_array_index_2048303_comb = p4_literal_2043896[p5_addedKey__50_comb[23:16]];
  assign p5_array_index_2048304_comb = p4_literal_2043896[p5_addedKey__50_comb[15:8]];
  assign p5_array_index_2048306_comb = p4_literal_2043910[p5_array_index_2048290_comb];
  assign p5_array_index_2048307_comb = p4_literal_2043912[p5_array_index_2048291_comb];
  assign p5_array_index_2048308_comb = p4_literal_2043914[p5_array_index_2048292_comb];
  assign p5_array_index_2048309_comb = p4_literal_2043916[p5_array_index_2048293_comb];
  assign p5_array_index_2048310_comb = p4_literal_2043918[p5_array_index_2048294_comb];
  assign p5_array_index_2048311_comb = p4_literal_2043920[p5_array_index_2048295_comb];
  assign p5_array_index_2048312_comb = p4_literal_2043896[p5_addedKey__50_comb[79:72]];
  assign p5_array_index_2048314_comb = p4_literal_2043896[p5_addedKey__50_comb[63:56]];
  assign p5_res7__576_comb = p5_array_index_2048306_comb ^ p5_array_index_2048307_comb ^ p5_array_index_2048308_comb ^ p5_array_index_2048309_comb ^ p5_array_index_2048310_comb ^ p5_array_index_2048311_comb ^ p5_array_index_2048312_comb ^ p4_literal_2043923[p5_array_index_2048297_comb] ^ p5_array_index_2048314_comb ^ p4_literal_2043920[p5_array_index_2048299_comb] ^ p4_literal_2043918[p5_array_index_2048300_comb] ^ p4_literal_2043916[p5_array_index_2048301_comb] ^ p4_literal_2043914[p5_array_index_2048302_comb] ^ p4_literal_2043912[p5_array_index_2048303_comb] ^ p4_literal_2043910[p5_array_index_2048304_comb] ^ p4_literal_2043896[p5_addedKey__50_comb[7:0]];
  assign p5_array_index_2048323_comb = p4_literal_2043910[p5_res7__576_comb];
  assign p5_array_index_2048324_comb = p4_literal_2043912[p5_array_index_2048290_comb];
  assign p5_array_index_2048325_comb = p4_literal_2043914[p5_array_index_2048291_comb];
  assign p5_array_index_2048326_comb = p4_literal_2043916[p5_array_index_2048292_comb];
  assign p5_array_index_2048327_comb = p4_literal_2043918[p5_array_index_2048293_comb];
  assign p5_array_index_2048328_comb = p4_literal_2043920[p5_array_index_2048294_comb];
  assign p5_res7__578_comb = p5_array_index_2048323_comb ^ p5_array_index_2048324_comb ^ p5_array_index_2048325_comb ^ p5_array_index_2048326_comb ^ p5_array_index_2048327_comb ^ p5_array_index_2048328_comb ^ p5_array_index_2048295_comb ^ p4_literal_2043923[p5_array_index_2048312_comb] ^ p5_array_index_2048297_comb ^ p4_literal_2043920[p5_array_index_2048314_comb] ^ p4_literal_2043918[p5_array_index_2048299_comb] ^ p4_literal_2043916[p5_array_index_2048300_comb] ^ p4_literal_2043914[p5_array_index_2048301_comb] ^ p4_literal_2043912[p5_array_index_2048302_comb] ^ p4_literal_2043910[p5_array_index_2048303_comb] ^ p5_array_index_2048304_comb;
  assign p5_array_index_2048338_comb = p4_literal_2043912[p5_res7__576_comb];
  assign p5_array_index_2048339_comb = p4_literal_2043914[p5_array_index_2048290_comb];
  assign p5_array_index_2048340_comb = p4_literal_2043916[p5_array_index_2048291_comb];
  assign p5_array_index_2048341_comb = p4_literal_2043918[p5_array_index_2048292_comb];
  assign p5_array_index_2048342_comb = p4_literal_2043920[p5_array_index_2048293_comb];
  assign p5_res7__580_comb = p4_literal_2043910[p5_res7__578_comb] ^ p5_array_index_2048338_comb ^ p5_array_index_2048339_comb ^ p5_array_index_2048340_comb ^ p5_array_index_2048341_comb ^ p5_array_index_2048342_comb ^ p5_array_index_2048294_comb ^ p4_literal_2043923[p5_array_index_2048295_comb] ^ p5_array_index_2048312_comb ^ p4_literal_2043920[p5_array_index_2048297_comb] ^ p4_literal_2043918[p5_array_index_2048314_comb] ^ p4_literal_2043916[p5_array_index_2048299_comb] ^ p4_literal_2043914[p5_array_index_2048300_comb] ^ p4_literal_2043912[p5_array_index_2048301_comb] ^ p4_literal_2043910[p5_array_index_2048302_comb] ^ p5_array_index_2048303_comb;
  assign p5_array_index_2048352_comb = p4_literal_2043912[p5_res7__578_comb];
  assign p5_array_index_2048353_comb = p4_literal_2043914[p5_res7__576_comb];
  assign p5_array_index_2048354_comb = p4_literal_2043916[p5_array_index_2048290_comb];
  assign p5_array_index_2048355_comb = p4_literal_2043918[p5_array_index_2048291_comb];
  assign p5_array_index_2048356_comb = p4_literal_2043920[p5_array_index_2048292_comb];
  assign p5_res7__582_comb = p4_literal_2043910[p5_res7__580_comb] ^ p5_array_index_2048352_comb ^ p5_array_index_2048353_comb ^ p5_array_index_2048354_comb ^ p5_array_index_2048355_comb ^ p5_array_index_2048356_comb ^ p5_array_index_2048293_comb ^ p4_literal_2043923[p5_array_index_2048294_comb] ^ p5_array_index_2048295_comb ^ p4_literal_2043920[p5_array_index_2048312_comb] ^ p4_literal_2043918[p5_array_index_2048297_comb] ^ p4_literal_2043916[p5_array_index_2048314_comb] ^ p4_literal_2043914[p5_array_index_2048299_comb] ^ p4_literal_2043912[p5_array_index_2048300_comb] ^ p4_literal_2043910[p5_array_index_2048301_comb] ^ p5_array_index_2048302_comb;
  assign p5_array_index_2048367_comb = p4_literal_2043914[p5_res7__578_comb];
  assign p5_array_index_2048368_comb = p4_literal_2043916[p5_res7__576_comb];
  assign p5_array_index_2048369_comb = p4_literal_2043918[p5_array_index_2048290_comb];
  assign p5_array_index_2048370_comb = p4_literal_2043920[p5_array_index_2048291_comb];
  assign p5_res7__584_comb = p4_literal_2043910[p5_res7__582_comb] ^ p4_literal_2043912[p5_res7__580_comb] ^ p5_array_index_2048367_comb ^ p5_array_index_2048368_comb ^ p5_array_index_2048369_comb ^ p5_array_index_2048370_comb ^ p5_array_index_2048292_comb ^ p4_literal_2043923[p5_array_index_2048293_comb] ^ p5_array_index_2048294_comb ^ p5_array_index_2048311_comb ^ p4_literal_2043918[p5_array_index_2048312_comb] ^ p4_literal_2043916[p5_array_index_2048297_comb] ^ p4_literal_2043914[p5_array_index_2048314_comb] ^ p4_literal_2043912[p5_array_index_2048299_comb] ^ p4_literal_2043910[p5_array_index_2048300_comb] ^ p5_array_index_2048301_comb;
  assign p5_array_index_2048380_comb = p4_literal_2043914[p5_res7__580_comb];
  assign p5_array_index_2048381_comb = p4_literal_2043916[p5_res7__578_comb];
  assign p5_array_index_2048382_comb = p4_literal_2043918[p5_res7__576_comb];
  assign p5_array_index_2048383_comb = p4_literal_2043920[p5_array_index_2048290_comb];
  assign p5_res7__586_comb = p4_literal_2043910[p5_res7__584_comb] ^ p4_literal_2043912[p5_res7__582_comb] ^ p5_array_index_2048380_comb ^ p5_array_index_2048381_comb ^ p5_array_index_2048382_comb ^ p5_array_index_2048383_comb ^ p5_array_index_2048291_comb ^ p4_literal_2043923[p5_array_index_2048292_comb] ^ p5_array_index_2048293_comb ^ p5_array_index_2048328_comb ^ p4_literal_2043918[p5_array_index_2048295_comb] ^ p4_literal_2043916[p5_array_index_2048312_comb] ^ p4_literal_2043914[p5_array_index_2048297_comb] ^ p4_literal_2043912[p5_array_index_2048314_comb] ^ p4_literal_2043910[p5_array_index_2048299_comb] ^ p5_array_index_2048300_comb;
  assign p5_array_index_2048394_comb = p4_literal_2043916[p5_res7__580_comb];
  assign p5_array_index_2048395_comb = p4_literal_2043918[p5_res7__578_comb];
  assign p5_array_index_2048396_comb = p4_literal_2043920[p5_res7__576_comb];
  assign p5_res7__588_comb = p4_literal_2043910[p5_res7__586_comb] ^ p4_literal_2043912[p5_res7__584_comb] ^ p4_literal_2043914[p5_res7__582_comb] ^ p5_array_index_2048394_comb ^ p5_array_index_2048395_comb ^ p5_array_index_2048396_comb ^ p5_array_index_2048290_comb ^ p4_literal_2043923[p5_array_index_2048291_comb] ^ p5_array_index_2048292_comb ^ p5_array_index_2048342_comb ^ p5_array_index_2048310_comb ^ p4_literal_2043916[p5_array_index_2048295_comb] ^ p4_literal_2043914[p5_array_index_2048312_comb] ^ p4_literal_2043912[p5_array_index_2048297_comb] ^ p4_literal_2043910[p5_array_index_2048314_comb] ^ p5_array_index_2048299_comb;
  assign p5_array_index_2048406_comb = p4_literal_2043916[p5_res7__582_comb];
  assign p5_array_index_2048407_comb = p4_literal_2043918[p5_res7__580_comb];
  assign p5_array_index_2048408_comb = p4_literal_2043920[p5_res7__578_comb];
  assign p5_res7__590_comb = p4_literal_2043910[p5_res7__588_comb] ^ p4_literal_2043912[p5_res7__586_comb] ^ p4_literal_2043914[p5_res7__584_comb] ^ p5_array_index_2048406_comb ^ p5_array_index_2048407_comb ^ p5_array_index_2048408_comb ^ p5_res7__576_comb ^ p4_literal_2043923[p5_array_index_2048290_comb] ^ p5_array_index_2048291_comb ^ p5_array_index_2048356_comb ^ p5_array_index_2048327_comb ^ p4_literal_2043916[p5_array_index_2048294_comb] ^ p4_literal_2043914[p5_array_index_2048295_comb] ^ p4_literal_2043912[p5_array_index_2048312_comb] ^ p4_literal_2043910[p5_array_index_2048297_comb] ^ p5_array_index_2048314_comb;
  assign p5_array_index_2048419_comb = p4_literal_2043918[p5_res7__582_comb];
  assign p5_array_index_2048420_comb = p4_literal_2043920[p5_res7__580_comb];
  assign p5_res7__592_comb = p4_literal_2043910[p5_res7__590_comb] ^ p4_literal_2043912[p5_res7__588_comb] ^ p4_literal_2043914[p5_res7__586_comb] ^ p4_literal_2043916[p5_res7__584_comb] ^ p5_array_index_2048419_comb ^ p5_array_index_2048420_comb ^ p5_res7__578_comb ^ p4_literal_2043923[p5_res7__576_comb] ^ p5_array_index_2048290_comb ^ p5_array_index_2048370_comb ^ p5_array_index_2048341_comb ^ p5_array_index_2048309_comb ^ p4_literal_2043914[p5_array_index_2048294_comb] ^ p4_literal_2043912[p5_array_index_2048295_comb] ^ p4_literal_2043910[p5_array_index_2048312_comb] ^ p5_array_index_2048297_comb;
  assign p5_array_index_2048430_comb = p4_literal_2043918[p5_res7__584_comb];
  assign p5_array_index_2048431_comb = p4_literal_2043920[p5_res7__582_comb];
  assign p5_res7__594_comb = p4_literal_2043910[p5_res7__592_comb] ^ p4_literal_2043912[p5_res7__590_comb] ^ p4_literal_2043914[p5_res7__588_comb] ^ p4_literal_2043916[p5_res7__586_comb] ^ p5_array_index_2048430_comb ^ p5_array_index_2048431_comb ^ p5_res7__580_comb ^ p4_literal_2043923[p5_res7__578_comb] ^ p5_res7__576_comb ^ p5_array_index_2048383_comb ^ p5_array_index_2048355_comb ^ p5_array_index_2048326_comb ^ p4_literal_2043914[p5_array_index_2048293_comb] ^ p4_literal_2043912[p5_array_index_2048294_comb] ^ p4_literal_2043910[p5_array_index_2048295_comb] ^ p5_array_index_2048312_comb;
  assign p5_array_index_2048442_comb = p4_literal_2043920[p5_res7__584_comb];
  assign p5_res7__596_comb = p4_literal_2043910[p5_res7__594_comb] ^ p4_literal_2043912[p5_res7__592_comb] ^ p4_literal_2043914[p5_res7__590_comb] ^ p4_literal_2043916[p5_res7__588_comb] ^ p4_literal_2043918[p5_res7__586_comb] ^ p5_array_index_2048442_comb ^ p5_res7__582_comb ^ p4_literal_2043923[p5_res7__580_comb] ^ p5_res7__578_comb ^ p5_array_index_2048396_comb ^ p5_array_index_2048369_comb ^ p5_array_index_2048340_comb ^ p5_array_index_2048308_comb ^ p4_literal_2043912[p5_array_index_2048293_comb] ^ p4_literal_2043910[p5_array_index_2048294_comb] ^ p5_array_index_2048295_comb;
  assign p5_array_index_2048452_comb = p4_literal_2043920[p5_res7__586_comb];
  assign p5_res7__598_comb = p4_literal_2043910[p5_res7__596_comb] ^ p4_literal_2043912[p5_res7__594_comb] ^ p4_literal_2043914[p5_res7__592_comb] ^ p4_literal_2043916[p5_res7__590_comb] ^ p4_literal_2043918[p5_res7__588_comb] ^ p5_array_index_2048452_comb ^ p5_res7__584_comb ^ p4_literal_2043923[p5_res7__582_comb] ^ p5_res7__580_comb ^ p5_array_index_2048408_comb ^ p5_array_index_2048382_comb ^ p5_array_index_2048354_comb ^ p5_array_index_2048325_comb ^ p4_literal_2043912[p5_array_index_2048292_comb] ^ p4_literal_2043910[p5_array_index_2048293_comb] ^ p5_array_index_2048294_comb;
  assign p5_res7__600_comb = p4_literal_2043910[p5_res7__598_comb] ^ p4_literal_2043912[p5_res7__596_comb] ^ p4_literal_2043914[p5_res7__594_comb] ^ p4_literal_2043916[p5_res7__592_comb] ^ p4_literal_2043918[p5_res7__590_comb] ^ p4_literal_2043920[p5_res7__588_comb] ^ p5_res7__586_comb ^ p4_literal_2043923[p5_res7__584_comb] ^ p5_res7__582_comb ^ p5_array_index_2048420_comb ^ p5_array_index_2048395_comb ^ p5_array_index_2048368_comb ^ p5_array_index_2048339_comb ^ p5_array_index_2048307_comb ^ p4_literal_2043910[p5_array_index_2048292_comb] ^ p5_array_index_2048293_comb;
  assign p5_res7__602_comb = p4_literal_2043910[p5_res7__600_comb] ^ p4_literal_2043912[p5_res7__598_comb] ^ p4_literal_2043914[p5_res7__596_comb] ^ p4_literal_2043916[p5_res7__594_comb] ^ p4_literal_2043918[p5_res7__592_comb] ^ p4_literal_2043920[p5_res7__590_comb] ^ p5_res7__588_comb ^ p4_literal_2043923[p5_res7__586_comb] ^ p5_res7__584_comb ^ p5_array_index_2048431_comb ^ p5_array_index_2048407_comb ^ p5_array_index_2048381_comb ^ p5_array_index_2048353_comb ^ p5_array_index_2048324_comb ^ p4_literal_2043910[p5_array_index_2048291_comb] ^ p5_array_index_2048292_comb;
  assign p5_res7__604_comb = p4_literal_2043910[p5_res7__602_comb] ^ p4_literal_2043912[p5_res7__600_comb] ^ p4_literal_2043914[p5_res7__598_comb] ^ p4_literal_2043916[p5_res7__596_comb] ^ p4_literal_2043918[p5_res7__594_comb] ^ p4_literal_2043920[p5_res7__592_comb] ^ p5_res7__590_comb ^ p4_literal_2043923[p5_res7__588_comb] ^ p5_res7__586_comb ^ p5_array_index_2048442_comb ^ p5_array_index_2048419_comb ^ p5_array_index_2048394_comb ^ p5_array_index_2048367_comb ^ p5_array_index_2048338_comb ^ p5_array_index_2048306_comb ^ p5_array_index_2048291_comb;
  assign p5_res7__606_comb = p4_literal_2043910[p5_res7__604_comb] ^ p4_literal_2043912[p5_res7__602_comb] ^ p4_literal_2043914[p5_res7__600_comb] ^ p4_literal_2043916[p5_res7__598_comb] ^ p4_literal_2043918[p5_res7__596_comb] ^ p4_literal_2043920[p5_res7__594_comb] ^ p5_res7__592_comb ^ p4_literal_2043923[p5_res7__590_comb] ^ p5_res7__588_comb ^ p5_array_index_2048452_comb ^ p5_array_index_2048430_comb ^ p5_array_index_2048406_comb ^ p5_array_index_2048380_comb ^ p5_array_index_2048352_comb ^ p5_array_index_2048323_comb ^ p5_array_index_2048290_comb;
  assign p5_res__18_comb = {p5_res7__606_comb, p5_res7__604_comb, p5_res7__602_comb, p5_res7__600_comb, p5_res7__598_comb, p5_res7__596_comb, p5_res7__594_comb, p5_res7__592_comb, p5_res7__590_comb, p5_res7__588_comb, p5_res7__586_comb, p5_res7__584_comb, p5_res7__582_comb, p5_res7__580_comb, p5_res7__578_comb, p5_res7__576_comb};
  assign p5_xor_2048492_comb = p5_res__18_comb ^ p4_xor_2047932;
  assign p5_addedKey__51_comb = p5_xor_2048492_comb ^ 128'h547f_7727_7ce9_8774_2ea9_3083_bcc2_4114;
  assign p5_array_index_2048508_comb = p4_literal_2043896[p5_addedKey__51_comb[127:120]];
  assign p5_array_index_2048509_comb = p4_literal_2043896[p5_addedKey__51_comb[119:112]];
  assign p5_array_index_2048510_comb = p4_literal_2043896[p5_addedKey__51_comb[111:104]];
  assign p5_array_index_2048511_comb = p4_literal_2043896[p5_addedKey__51_comb[103:96]];
  assign p5_array_index_2048512_comb = p4_literal_2043896[p5_addedKey__51_comb[95:88]];
  assign p5_array_index_2048513_comb = p4_literal_2043896[p5_addedKey__51_comb[87:80]];
  assign p5_array_index_2048515_comb = p4_literal_2043896[p5_addedKey__51_comb[71:64]];
  assign p5_array_index_2048517_comb = p4_literal_2043896[p5_addedKey__51_comb[55:48]];
  assign p5_array_index_2048518_comb = p4_literal_2043896[p5_addedKey__51_comb[47:40]];
  assign p5_array_index_2048519_comb = p4_literal_2043896[p5_addedKey__51_comb[39:32]];
  assign p5_array_index_2048520_comb = p4_literal_2043896[p5_addedKey__51_comb[31:24]];
  assign p5_array_index_2048521_comb = p4_literal_2043896[p5_addedKey__51_comb[23:16]];
  assign p5_array_index_2048522_comb = p4_literal_2043896[p5_addedKey__51_comb[15:8]];
  assign p5_array_index_2048524_comb = p4_literal_2043910[p5_array_index_2048508_comb];
  assign p5_array_index_2048525_comb = p4_literal_2043912[p5_array_index_2048509_comb];
  assign p5_array_index_2048526_comb = p4_literal_2043914[p5_array_index_2048510_comb];
  assign p5_array_index_2048527_comb = p4_literal_2043916[p5_array_index_2048511_comb];
  assign p5_array_index_2048528_comb = p4_literal_2043918[p5_array_index_2048512_comb];
  assign p5_array_index_2048529_comb = p4_literal_2043920[p5_array_index_2048513_comb];
  assign p5_array_index_2048530_comb = p4_literal_2043896[p5_addedKey__51_comb[79:72]];
  assign p5_array_index_2048532_comb = p4_literal_2043896[p5_addedKey__51_comb[63:56]];
  assign p5_res7__608_comb = p5_array_index_2048524_comb ^ p5_array_index_2048525_comb ^ p5_array_index_2048526_comb ^ p5_array_index_2048527_comb ^ p5_array_index_2048528_comb ^ p5_array_index_2048529_comb ^ p5_array_index_2048530_comb ^ p4_literal_2043923[p5_array_index_2048515_comb] ^ p5_array_index_2048532_comb ^ p4_literal_2043920[p5_array_index_2048517_comb] ^ p4_literal_2043918[p5_array_index_2048518_comb] ^ p4_literal_2043916[p5_array_index_2048519_comb] ^ p4_literal_2043914[p5_array_index_2048520_comb] ^ p4_literal_2043912[p5_array_index_2048521_comb] ^ p4_literal_2043910[p5_array_index_2048522_comb] ^ p4_literal_2043896[p5_addedKey__51_comb[7:0]];
  assign p5_array_index_2048541_comb = p4_literal_2043910[p5_res7__608_comb];
  assign p5_array_index_2048542_comb = p4_literal_2043912[p5_array_index_2048508_comb];
  assign p5_array_index_2048543_comb = p4_literal_2043914[p5_array_index_2048509_comb];
  assign p5_array_index_2048544_comb = p4_literal_2043916[p5_array_index_2048510_comb];
  assign p5_array_index_2048545_comb = p4_literal_2043918[p5_array_index_2048511_comb];
  assign p5_array_index_2048546_comb = p4_literal_2043920[p5_array_index_2048512_comb];
  assign p5_res7__610_comb = p5_array_index_2048541_comb ^ p5_array_index_2048542_comb ^ p5_array_index_2048543_comb ^ p5_array_index_2048544_comb ^ p5_array_index_2048545_comb ^ p5_array_index_2048546_comb ^ p5_array_index_2048513_comb ^ p4_literal_2043923[p5_array_index_2048530_comb] ^ p5_array_index_2048515_comb ^ p4_literal_2043920[p5_array_index_2048532_comb] ^ p4_literal_2043918[p5_array_index_2048517_comb] ^ p4_literal_2043916[p5_array_index_2048518_comb] ^ p4_literal_2043914[p5_array_index_2048519_comb] ^ p4_literal_2043912[p5_array_index_2048520_comb] ^ p4_literal_2043910[p5_array_index_2048521_comb] ^ p5_array_index_2048522_comb;
  assign p5_array_index_2048556_comb = p4_literal_2043912[p5_res7__608_comb];
  assign p5_array_index_2048557_comb = p4_literal_2043914[p5_array_index_2048508_comb];
  assign p5_array_index_2048558_comb = p4_literal_2043916[p5_array_index_2048509_comb];
  assign p5_array_index_2048559_comb = p4_literal_2043918[p5_array_index_2048510_comb];
  assign p5_array_index_2048560_comb = p4_literal_2043920[p5_array_index_2048511_comb];
  assign p5_res7__612_comb = p4_literal_2043910[p5_res7__610_comb] ^ p5_array_index_2048556_comb ^ p5_array_index_2048557_comb ^ p5_array_index_2048558_comb ^ p5_array_index_2048559_comb ^ p5_array_index_2048560_comb ^ p5_array_index_2048512_comb ^ p4_literal_2043923[p5_array_index_2048513_comb] ^ p5_array_index_2048530_comb ^ p4_literal_2043920[p5_array_index_2048515_comb] ^ p4_literal_2043918[p5_array_index_2048532_comb] ^ p4_literal_2043916[p5_array_index_2048517_comb] ^ p4_literal_2043914[p5_array_index_2048518_comb] ^ p4_literal_2043912[p5_array_index_2048519_comb] ^ p4_literal_2043910[p5_array_index_2048520_comb] ^ p5_array_index_2048521_comb;
  assign p5_array_index_2048570_comb = p4_literal_2043912[p5_res7__610_comb];
  assign p5_array_index_2048571_comb = p4_literal_2043914[p5_res7__608_comb];
  assign p5_array_index_2048572_comb = p4_literal_2043916[p5_array_index_2048508_comb];
  assign p5_array_index_2048573_comb = p4_literal_2043918[p5_array_index_2048509_comb];
  assign p5_array_index_2048574_comb = p4_literal_2043920[p5_array_index_2048510_comb];
  assign p5_res7__614_comb = p4_literal_2043910[p5_res7__612_comb] ^ p5_array_index_2048570_comb ^ p5_array_index_2048571_comb ^ p5_array_index_2048572_comb ^ p5_array_index_2048573_comb ^ p5_array_index_2048574_comb ^ p5_array_index_2048511_comb ^ p4_literal_2043923[p5_array_index_2048512_comb] ^ p5_array_index_2048513_comb ^ p4_literal_2043920[p5_array_index_2048530_comb] ^ p4_literal_2043918[p5_array_index_2048515_comb] ^ p4_literal_2043916[p5_array_index_2048532_comb] ^ p4_literal_2043914[p5_array_index_2048517_comb] ^ p4_literal_2043912[p5_array_index_2048518_comb] ^ p4_literal_2043910[p5_array_index_2048519_comb] ^ p5_array_index_2048520_comb;
  assign p5_array_index_2048585_comb = p4_literal_2043914[p5_res7__610_comb];
  assign p5_array_index_2048586_comb = p4_literal_2043916[p5_res7__608_comb];
  assign p5_array_index_2048587_comb = p4_literal_2043918[p5_array_index_2048508_comb];
  assign p5_array_index_2048588_comb = p4_literal_2043920[p5_array_index_2048509_comb];
  assign p5_res7__616_comb = p4_literal_2043910[p5_res7__614_comb] ^ p4_literal_2043912[p5_res7__612_comb] ^ p5_array_index_2048585_comb ^ p5_array_index_2048586_comb ^ p5_array_index_2048587_comb ^ p5_array_index_2048588_comb ^ p5_array_index_2048510_comb ^ p4_literal_2043923[p5_array_index_2048511_comb] ^ p5_array_index_2048512_comb ^ p5_array_index_2048529_comb ^ p4_literal_2043918[p5_array_index_2048530_comb] ^ p4_literal_2043916[p5_array_index_2048515_comb] ^ p4_literal_2043914[p5_array_index_2048532_comb] ^ p4_literal_2043912[p5_array_index_2048517_comb] ^ p4_literal_2043910[p5_array_index_2048518_comb] ^ p5_array_index_2048519_comb;
  assign p5_array_index_2048598_comb = p4_literal_2043914[p5_res7__612_comb];
  assign p5_array_index_2048599_comb = p4_literal_2043916[p5_res7__610_comb];
  assign p5_array_index_2048600_comb = p4_literal_2043918[p5_res7__608_comb];
  assign p5_array_index_2048601_comb = p4_literal_2043920[p5_array_index_2048508_comb];
  assign p5_res7__618_comb = p4_literal_2043910[p5_res7__616_comb] ^ p4_literal_2043912[p5_res7__614_comb] ^ p5_array_index_2048598_comb ^ p5_array_index_2048599_comb ^ p5_array_index_2048600_comb ^ p5_array_index_2048601_comb ^ p5_array_index_2048509_comb ^ p4_literal_2043923[p5_array_index_2048510_comb] ^ p5_array_index_2048511_comb ^ p5_array_index_2048546_comb ^ p4_literal_2043918[p5_array_index_2048513_comb] ^ p4_literal_2043916[p5_array_index_2048530_comb] ^ p4_literal_2043914[p5_array_index_2048515_comb] ^ p4_literal_2043912[p5_array_index_2048532_comb] ^ p4_literal_2043910[p5_array_index_2048517_comb] ^ p5_array_index_2048518_comb;
  assign p5_array_index_2048612_comb = p4_literal_2043916[p5_res7__612_comb];
  assign p5_array_index_2048613_comb = p4_literal_2043918[p5_res7__610_comb];
  assign p5_array_index_2048614_comb = p4_literal_2043920[p5_res7__608_comb];
  assign p5_res7__620_comb = p4_literal_2043910[p5_res7__618_comb] ^ p4_literal_2043912[p5_res7__616_comb] ^ p4_literal_2043914[p5_res7__614_comb] ^ p5_array_index_2048612_comb ^ p5_array_index_2048613_comb ^ p5_array_index_2048614_comb ^ p5_array_index_2048508_comb ^ p4_literal_2043923[p5_array_index_2048509_comb] ^ p5_array_index_2048510_comb ^ p5_array_index_2048560_comb ^ p5_array_index_2048528_comb ^ p4_literal_2043916[p5_array_index_2048513_comb] ^ p4_literal_2043914[p5_array_index_2048530_comb] ^ p4_literal_2043912[p5_array_index_2048515_comb] ^ p4_literal_2043910[p5_array_index_2048532_comb] ^ p5_array_index_2048517_comb;
  assign p5_array_index_2048624_comb = p4_literal_2043916[p5_res7__614_comb];
  assign p5_array_index_2048625_comb = p4_literal_2043918[p5_res7__612_comb];
  assign p5_array_index_2048626_comb = p4_literal_2043920[p5_res7__610_comb];
  assign p5_res7__622_comb = p4_literal_2043910[p5_res7__620_comb] ^ p4_literal_2043912[p5_res7__618_comb] ^ p4_literal_2043914[p5_res7__616_comb] ^ p5_array_index_2048624_comb ^ p5_array_index_2048625_comb ^ p5_array_index_2048626_comb ^ p5_res7__608_comb ^ p4_literal_2043923[p5_array_index_2048508_comb] ^ p5_array_index_2048509_comb ^ p5_array_index_2048574_comb ^ p5_array_index_2048545_comb ^ p4_literal_2043916[p5_array_index_2048512_comb] ^ p4_literal_2043914[p5_array_index_2048513_comb] ^ p4_literal_2043912[p5_array_index_2048530_comb] ^ p4_literal_2043910[p5_array_index_2048515_comb] ^ p5_array_index_2048532_comb;
  assign p5_array_index_2048637_comb = p4_literal_2043918[p5_res7__614_comb];
  assign p5_array_index_2048638_comb = p4_literal_2043920[p5_res7__612_comb];
  assign p5_res7__624_comb = p4_literal_2043910[p5_res7__622_comb] ^ p4_literal_2043912[p5_res7__620_comb] ^ p4_literal_2043914[p5_res7__618_comb] ^ p4_literal_2043916[p5_res7__616_comb] ^ p5_array_index_2048637_comb ^ p5_array_index_2048638_comb ^ p5_res7__610_comb ^ p4_literal_2043923[p5_res7__608_comb] ^ p5_array_index_2048508_comb ^ p5_array_index_2048588_comb ^ p5_array_index_2048559_comb ^ p5_array_index_2048527_comb ^ p4_literal_2043914[p5_array_index_2048512_comb] ^ p4_literal_2043912[p5_array_index_2048513_comb] ^ p4_literal_2043910[p5_array_index_2048530_comb] ^ p5_array_index_2048515_comb;
  assign p5_array_index_2048648_comb = p4_literal_2043918[p5_res7__616_comb];
  assign p5_array_index_2048649_comb = p4_literal_2043920[p5_res7__614_comb];
  assign p5_res7__626_comb = p4_literal_2043910[p5_res7__624_comb] ^ p4_literal_2043912[p5_res7__622_comb] ^ p4_literal_2043914[p5_res7__620_comb] ^ p4_literal_2043916[p5_res7__618_comb] ^ p5_array_index_2048648_comb ^ p5_array_index_2048649_comb ^ p5_res7__612_comb ^ p4_literal_2043923[p5_res7__610_comb] ^ p5_res7__608_comb ^ p5_array_index_2048601_comb ^ p5_array_index_2048573_comb ^ p5_array_index_2048544_comb ^ p4_literal_2043914[p5_array_index_2048511_comb] ^ p4_literal_2043912[p5_array_index_2048512_comb] ^ p4_literal_2043910[p5_array_index_2048513_comb] ^ p5_array_index_2048530_comb;
  assign p5_array_index_2048660_comb = p4_literal_2043920[p5_res7__616_comb];
  assign p5_res7__628_comb = p4_literal_2043910[p5_res7__626_comb] ^ p4_literal_2043912[p5_res7__624_comb] ^ p4_literal_2043914[p5_res7__622_comb] ^ p4_literal_2043916[p5_res7__620_comb] ^ p4_literal_2043918[p5_res7__618_comb] ^ p5_array_index_2048660_comb ^ p5_res7__614_comb ^ p4_literal_2043923[p5_res7__612_comb] ^ p5_res7__610_comb ^ p5_array_index_2048614_comb ^ p5_array_index_2048587_comb ^ p5_array_index_2048558_comb ^ p5_array_index_2048526_comb ^ p4_literal_2043912[p5_array_index_2048511_comb] ^ p4_literal_2043910[p5_array_index_2048512_comb] ^ p5_array_index_2048513_comb;
  assign p5_array_index_2048670_comb = p4_literal_2043920[p5_res7__618_comb];
  assign p5_res7__630_comb = p4_literal_2043910[p5_res7__628_comb] ^ p4_literal_2043912[p5_res7__626_comb] ^ p4_literal_2043914[p5_res7__624_comb] ^ p4_literal_2043916[p5_res7__622_comb] ^ p4_literal_2043918[p5_res7__620_comb] ^ p5_array_index_2048670_comb ^ p5_res7__616_comb ^ p4_literal_2043923[p5_res7__614_comb] ^ p5_res7__612_comb ^ p5_array_index_2048626_comb ^ p5_array_index_2048600_comb ^ p5_array_index_2048572_comb ^ p5_array_index_2048543_comb ^ p4_literal_2043912[p5_array_index_2048510_comb] ^ p4_literal_2043910[p5_array_index_2048511_comb] ^ p5_array_index_2048512_comb;
  assign p5_res7__632_comb = p4_literal_2043910[p5_res7__630_comb] ^ p4_literal_2043912[p5_res7__628_comb] ^ p4_literal_2043914[p5_res7__626_comb] ^ p4_literal_2043916[p5_res7__624_comb] ^ p4_literal_2043918[p5_res7__622_comb] ^ p4_literal_2043920[p5_res7__620_comb] ^ p5_res7__618_comb ^ p4_literal_2043923[p5_res7__616_comb] ^ p5_res7__614_comb ^ p5_array_index_2048638_comb ^ p5_array_index_2048613_comb ^ p5_array_index_2048586_comb ^ p5_array_index_2048557_comb ^ p5_array_index_2048525_comb ^ p4_literal_2043910[p5_array_index_2048510_comb] ^ p5_array_index_2048511_comb;
  assign p5_res7__634_comb = p4_literal_2043910[p5_res7__632_comb] ^ p4_literal_2043912[p5_res7__630_comb] ^ p4_literal_2043914[p5_res7__628_comb] ^ p4_literal_2043916[p5_res7__626_comb] ^ p4_literal_2043918[p5_res7__624_comb] ^ p4_literal_2043920[p5_res7__622_comb] ^ p5_res7__620_comb ^ p4_literal_2043923[p5_res7__618_comb] ^ p5_res7__616_comb ^ p5_array_index_2048649_comb ^ p5_array_index_2048625_comb ^ p5_array_index_2048599_comb ^ p5_array_index_2048571_comb ^ p5_array_index_2048542_comb ^ p4_literal_2043910[p5_array_index_2048509_comb] ^ p5_array_index_2048510_comb;
  assign p5_res7__636_comb = p4_literal_2043910[p5_res7__634_comb] ^ p4_literal_2043912[p5_res7__632_comb] ^ p4_literal_2043914[p5_res7__630_comb] ^ p4_literal_2043916[p5_res7__628_comb] ^ p4_literal_2043918[p5_res7__626_comb] ^ p4_literal_2043920[p5_res7__624_comb] ^ p5_res7__622_comb ^ p4_literal_2043923[p5_res7__620_comb] ^ p5_res7__618_comb ^ p5_array_index_2048660_comb ^ p5_array_index_2048637_comb ^ p5_array_index_2048612_comb ^ p5_array_index_2048585_comb ^ p5_array_index_2048556_comb ^ p5_array_index_2048524_comb ^ p5_array_index_2048509_comb;
  assign p5_res7__638_comb = p4_literal_2043910[p5_res7__636_comb] ^ p4_literal_2043912[p5_res7__634_comb] ^ p4_literal_2043914[p5_res7__632_comb] ^ p4_literal_2043916[p5_res7__630_comb] ^ p4_literal_2043918[p5_res7__628_comb] ^ p4_literal_2043920[p5_res7__626_comb] ^ p5_res7__624_comb ^ p4_literal_2043923[p5_res7__622_comb] ^ p5_res7__620_comb ^ p5_array_index_2048670_comb ^ p5_array_index_2048648_comb ^ p5_array_index_2048624_comb ^ p5_array_index_2048598_comb ^ p5_array_index_2048570_comb ^ p5_array_index_2048541_comb ^ p5_array_index_2048508_comb;
  assign p5_res__19_comb = {p5_res7__638_comb, p5_res7__636_comb, p5_res7__634_comb, p5_res7__632_comb, p5_res7__630_comb, p5_res7__628_comb, p5_res7__626_comb, p5_res7__624_comb, p5_res7__622_comb, p5_res7__620_comb, p5_res7__618_comb, p5_res7__616_comb, p5_res7__614_comb, p5_res7__612_comb, p5_res7__610_comb, p5_res7__608_comb};
  assign p5_xor_2048710_comb = p5_res__19_comb ^ p5_xor_2048274_comb;
  assign p5_addedKey__52_comb = p5_xor_2048710_comb ^ 128'h3add_0155_10a1_fdcc_738e_8d93_6146_d515;
  assign p5_array_index_2048726_comb = p4_literal_2043896[p5_addedKey__52_comb[127:120]];
  assign p5_array_index_2048727_comb = p4_literal_2043896[p5_addedKey__52_comb[119:112]];
  assign p5_array_index_2048728_comb = p4_literal_2043896[p5_addedKey__52_comb[111:104]];
  assign p5_array_index_2048729_comb = p4_literal_2043896[p5_addedKey__52_comb[103:96]];
  assign p5_array_index_2048730_comb = p4_literal_2043896[p5_addedKey__52_comb[95:88]];
  assign p5_array_index_2048731_comb = p4_literal_2043896[p5_addedKey__52_comb[87:80]];
  assign p5_array_index_2048733_comb = p4_literal_2043896[p5_addedKey__52_comb[71:64]];
  assign p5_array_index_2048735_comb = p4_literal_2043896[p5_addedKey__52_comb[55:48]];
  assign p5_array_index_2048736_comb = p4_literal_2043896[p5_addedKey__52_comb[47:40]];
  assign p5_array_index_2048737_comb = p4_literal_2043896[p5_addedKey__52_comb[39:32]];
  assign p5_array_index_2048738_comb = p4_literal_2043896[p5_addedKey__52_comb[31:24]];
  assign p5_array_index_2048739_comb = p4_literal_2043896[p5_addedKey__52_comb[23:16]];
  assign p5_array_index_2048740_comb = p4_literal_2043896[p5_addedKey__52_comb[15:8]];
  assign p5_array_index_2048742_comb = p4_literal_2043910[p5_array_index_2048726_comb];
  assign p5_array_index_2048743_comb = p4_literal_2043912[p5_array_index_2048727_comb];
  assign p5_array_index_2048744_comb = p4_literal_2043914[p5_array_index_2048728_comb];
  assign p5_array_index_2048745_comb = p4_literal_2043916[p5_array_index_2048729_comb];
  assign p5_array_index_2048746_comb = p4_literal_2043918[p5_array_index_2048730_comb];
  assign p5_array_index_2048747_comb = p4_literal_2043920[p5_array_index_2048731_comb];
  assign p5_array_index_2048748_comb = p4_literal_2043896[p5_addedKey__52_comb[79:72]];
  assign p5_array_index_2048750_comb = p4_literal_2043896[p5_addedKey__52_comb[63:56]];
  assign p5_res7__640_comb = p5_array_index_2048742_comb ^ p5_array_index_2048743_comb ^ p5_array_index_2048744_comb ^ p5_array_index_2048745_comb ^ p5_array_index_2048746_comb ^ p5_array_index_2048747_comb ^ p5_array_index_2048748_comb ^ p4_literal_2043923[p5_array_index_2048733_comb] ^ p5_array_index_2048750_comb ^ p4_literal_2043920[p5_array_index_2048735_comb] ^ p4_literal_2043918[p5_array_index_2048736_comb] ^ p4_literal_2043916[p5_array_index_2048737_comb] ^ p4_literal_2043914[p5_array_index_2048738_comb] ^ p4_literal_2043912[p5_array_index_2048739_comb] ^ p4_literal_2043910[p5_array_index_2048740_comb] ^ p4_literal_2043896[p5_addedKey__52_comb[7:0]];
  assign p5_array_index_2048759_comb = p4_literal_2043910[p5_res7__640_comb];
  assign p5_array_index_2048760_comb = p4_literal_2043912[p5_array_index_2048726_comb];
  assign p5_array_index_2048761_comb = p4_literal_2043914[p5_array_index_2048727_comb];
  assign p5_array_index_2048762_comb = p4_literal_2043916[p5_array_index_2048728_comb];
  assign p5_array_index_2048763_comb = p4_literal_2043918[p5_array_index_2048729_comb];
  assign p5_array_index_2048764_comb = p4_literal_2043920[p5_array_index_2048730_comb];
  assign p5_res7__642_comb = p5_array_index_2048759_comb ^ p5_array_index_2048760_comb ^ p5_array_index_2048761_comb ^ p5_array_index_2048762_comb ^ p5_array_index_2048763_comb ^ p5_array_index_2048764_comb ^ p5_array_index_2048731_comb ^ p4_literal_2043923[p5_array_index_2048748_comb] ^ p5_array_index_2048733_comb ^ p4_literal_2043920[p5_array_index_2048750_comb] ^ p4_literal_2043918[p5_array_index_2048735_comb] ^ p4_literal_2043916[p5_array_index_2048736_comb] ^ p4_literal_2043914[p5_array_index_2048737_comb] ^ p4_literal_2043912[p5_array_index_2048738_comb] ^ p4_literal_2043910[p5_array_index_2048739_comb] ^ p5_array_index_2048740_comb;
  assign p5_array_index_2048774_comb = p4_literal_2043912[p5_res7__640_comb];
  assign p5_array_index_2048775_comb = p4_literal_2043914[p5_array_index_2048726_comb];
  assign p5_array_index_2048776_comb = p4_literal_2043916[p5_array_index_2048727_comb];
  assign p5_array_index_2048777_comb = p4_literal_2043918[p5_array_index_2048728_comb];
  assign p5_array_index_2048778_comb = p4_literal_2043920[p5_array_index_2048729_comb];
  assign p5_res7__644_comb = p4_literal_2043910[p5_res7__642_comb] ^ p5_array_index_2048774_comb ^ p5_array_index_2048775_comb ^ p5_array_index_2048776_comb ^ p5_array_index_2048777_comb ^ p5_array_index_2048778_comb ^ p5_array_index_2048730_comb ^ p4_literal_2043923[p5_array_index_2048731_comb] ^ p5_array_index_2048748_comb ^ p4_literal_2043920[p5_array_index_2048733_comb] ^ p4_literal_2043918[p5_array_index_2048750_comb] ^ p4_literal_2043916[p5_array_index_2048735_comb] ^ p4_literal_2043914[p5_array_index_2048736_comb] ^ p4_literal_2043912[p5_array_index_2048737_comb] ^ p4_literal_2043910[p5_array_index_2048738_comb] ^ p5_array_index_2048739_comb;
  assign p5_array_index_2048788_comb = p4_literal_2043912[p5_res7__642_comb];
  assign p5_array_index_2048789_comb = p4_literal_2043914[p5_res7__640_comb];
  assign p5_array_index_2048790_comb = p4_literal_2043916[p5_array_index_2048726_comb];
  assign p5_array_index_2048791_comb = p4_literal_2043918[p5_array_index_2048727_comb];
  assign p5_array_index_2048792_comb = p4_literal_2043920[p5_array_index_2048728_comb];
  assign p5_res7__646_comb = p4_literal_2043910[p5_res7__644_comb] ^ p5_array_index_2048788_comb ^ p5_array_index_2048789_comb ^ p5_array_index_2048790_comb ^ p5_array_index_2048791_comb ^ p5_array_index_2048792_comb ^ p5_array_index_2048729_comb ^ p4_literal_2043923[p5_array_index_2048730_comb] ^ p5_array_index_2048731_comb ^ p4_literal_2043920[p5_array_index_2048748_comb] ^ p4_literal_2043918[p5_array_index_2048733_comb] ^ p4_literal_2043916[p5_array_index_2048750_comb] ^ p4_literal_2043914[p5_array_index_2048735_comb] ^ p4_literal_2043912[p5_array_index_2048736_comb] ^ p4_literal_2043910[p5_array_index_2048737_comb] ^ p5_array_index_2048738_comb;
  assign p5_array_index_2048803_comb = p4_literal_2043914[p5_res7__642_comb];
  assign p5_array_index_2048804_comb = p4_literal_2043916[p5_res7__640_comb];
  assign p5_array_index_2048805_comb = p4_literal_2043918[p5_array_index_2048726_comb];
  assign p5_array_index_2048806_comb = p4_literal_2043920[p5_array_index_2048727_comb];
  assign p5_res7__648_comb = p4_literal_2043910[p5_res7__646_comb] ^ p4_literal_2043912[p5_res7__644_comb] ^ p5_array_index_2048803_comb ^ p5_array_index_2048804_comb ^ p5_array_index_2048805_comb ^ p5_array_index_2048806_comb ^ p5_array_index_2048728_comb ^ p4_literal_2043923[p5_array_index_2048729_comb] ^ p5_array_index_2048730_comb ^ p5_array_index_2048747_comb ^ p4_literal_2043918[p5_array_index_2048748_comb] ^ p4_literal_2043916[p5_array_index_2048733_comb] ^ p4_literal_2043914[p5_array_index_2048750_comb] ^ p4_literal_2043912[p5_array_index_2048735_comb] ^ p4_literal_2043910[p5_array_index_2048736_comb] ^ p5_array_index_2048737_comb;
  assign p5_array_index_2048816_comb = p4_literal_2043914[p5_res7__644_comb];
  assign p5_array_index_2048817_comb = p4_literal_2043916[p5_res7__642_comb];
  assign p5_array_index_2048818_comb = p4_literal_2043918[p5_res7__640_comb];
  assign p5_array_index_2048819_comb = p4_literal_2043920[p5_array_index_2048726_comb];
  assign p5_res7__650_comb = p4_literal_2043910[p5_res7__648_comb] ^ p4_literal_2043912[p5_res7__646_comb] ^ p5_array_index_2048816_comb ^ p5_array_index_2048817_comb ^ p5_array_index_2048818_comb ^ p5_array_index_2048819_comb ^ p5_array_index_2048727_comb ^ p4_literal_2043923[p5_array_index_2048728_comb] ^ p5_array_index_2048729_comb ^ p5_array_index_2048764_comb ^ p4_literal_2043918[p5_array_index_2048731_comb] ^ p4_literal_2043916[p5_array_index_2048748_comb] ^ p4_literal_2043914[p5_array_index_2048733_comb] ^ p4_literal_2043912[p5_array_index_2048750_comb] ^ p4_literal_2043910[p5_array_index_2048735_comb] ^ p5_array_index_2048736_comb;
  assign p5_array_index_2048830_comb = p4_literal_2043916[p5_res7__644_comb];
  assign p5_array_index_2048831_comb = p4_literal_2043918[p5_res7__642_comb];
  assign p5_array_index_2048832_comb = p4_literal_2043920[p5_res7__640_comb];
  assign p5_res7__652_comb = p4_literal_2043910[p5_res7__650_comb] ^ p4_literal_2043912[p5_res7__648_comb] ^ p4_literal_2043914[p5_res7__646_comb] ^ p5_array_index_2048830_comb ^ p5_array_index_2048831_comb ^ p5_array_index_2048832_comb ^ p5_array_index_2048726_comb ^ p4_literal_2043923[p5_array_index_2048727_comb] ^ p5_array_index_2048728_comb ^ p5_array_index_2048778_comb ^ p5_array_index_2048746_comb ^ p4_literal_2043916[p5_array_index_2048731_comb] ^ p4_literal_2043914[p5_array_index_2048748_comb] ^ p4_literal_2043912[p5_array_index_2048733_comb] ^ p4_literal_2043910[p5_array_index_2048750_comb] ^ p5_array_index_2048735_comb;
  assign p5_array_index_2048842_comb = p4_literal_2043916[p5_res7__646_comb];
  assign p5_array_index_2048843_comb = p4_literal_2043918[p5_res7__644_comb];
  assign p5_array_index_2048844_comb = p4_literal_2043920[p5_res7__642_comb];
  assign p5_res7__654_comb = p4_literal_2043910[p5_res7__652_comb] ^ p4_literal_2043912[p5_res7__650_comb] ^ p4_literal_2043914[p5_res7__648_comb] ^ p5_array_index_2048842_comb ^ p5_array_index_2048843_comb ^ p5_array_index_2048844_comb ^ p5_res7__640_comb ^ p4_literal_2043923[p5_array_index_2048726_comb] ^ p5_array_index_2048727_comb ^ p5_array_index_2048792_comb ^ p5_array_index_2048763_comb ^ p4_literal_2043916[p5_array_index_2048730_comb] ^ p4_literal_2043914[p5_array_index_2048731_comb] ^ p4_literal_2043912[p5_array_index_2048748_comb] ^ p4_literal_2043910[p5_array_index_2048733_comb] ^ p5_array_index_2048750_comb;
  assign p5_array_index_2048855_comb = p4_literal_2043918[p5_res7__646_comb];
  assign p5_array_index_2048856_comb = p4_literal_2043920[p5_res7__644_comb];
  assign p5_res7__656_comb = p4_literal_2043910[p5_res7__654_comb] ^ p4_literal_2043912[p5_res7__652_comb] ^ p4_literal_2043914[p5_res7__650_comb] ^ p4_literal_2043916[p5_res7__648_comb] ^ p5_array_index_2048855_comb ^ p5_array_index_2048856_comb ^ p5_res7__642_comb ^ p4_literal_2043923[p5_res7__640_comb] ^ p5_array_index_2048726_comb ^ p5_array_index_2048806_comb ^ p5_array_index_2048777_comb ^ p5_array_index_2048745_comb ^ p4_literal_2043914[p5_array_index_2048730_comb] ^ p4_literal_2043912[p5_array_index_2048731_comb] ^ p4_literal_2043910[p5_array_index_2048748_comb] ^ p5_array_index_2048733_comb;
  assign p5_array_index_2048866_comb = p4_literal_2043918[p5_res7__648_comb];
  assign p5_array_index_2048867_comb = p4_literal_2043920[p5_res7__646_comb];
  assign p5_res7__658_comb = p4_literal_2043910[p5_res7__656_comb] ^ p4_literal_2043912[p5_res7__654_comb] ^ p4_literal_2043914[p5_res7__652_comb] ^ p4_literal_2043916[p5_res7__650_comb] ^ p5_array_index_2048866_comb ^ p5_array_index_2048867_comb ^ p5_res7__644_comb ^ p4_literal_2043923[p5_res7__642_comb] ^ p5_res7__640_comb ^ p5_array_index_2048819_comb ^ p5_array_index_2048791_comb ^ p5_array_index_2048762_comb ^ p4_literal_2043914[p5_array_index_2048729_comb] ^ p4_literal_2043912[p5_array_index_2048730_comb] ^ p4_literal_2043910[p5_array_index_2048731_comb] ^ p5_array_index_2048748_comb;
  assign p5_array_index_2048878_comb = p4_literal_2043920[p5_res7__648_comb];
  assign p5_res7__660_comb = p4_literal_2043910[p5_res7__658_comb] ^ p4_literal_2043912[p5_res7__656_comb] ^ p4_literal_2043914[p5_res7__654_comb] ^ p4_literal_2043916[p5_res7__652_comb] ^ p4_literal_2043918[p5_res7__650_comb] ^ p5_array_index_2048878_comb ^ p5_res7__646_comb ^ p4_literal_2043923[p5_res7__644_comb] ^ p5_res7__642_comb ^ p5_array_index_2048832_comb ^ p5_array_index_2048805_comb ^ p5_array_index_2048776_comb ^ p5_array_index_2048744_comb ^ p4_literal_2043912[p5_array_index_2048729_comb] ^ p4_literal_2043910[p5_array_index_2048730_comb] ^ p5_array_index_2048731_comb;
  assign p5_array_index_2048888_comb = p4_literal_2043920[p5_res7__650_comb];
  assign p5_res7__662_comb = p4_literal_2043910[p5_res7__660_comb] ^ p4_literal_2043912[p5_res7__658_comb] ^ p4_literal_2043914[p5_res7__656_comb] ^ p4_literal_2043916[p5_res7__654_comb] ^ p4_literal_2043918[p5_res7__652_comb] ^ p5_array_index_2048888_comb ^ p5_res7__648_comb ^ p4_literal_2043923[p5_res7__646_comb] ^ p5_res7__644_comb ^ p5_array_index_2048844_comb ^ p5_array_index_2048818_comb ^ p5_array_index_2048790_comb ^ p5_array_index_2048761_comb ^ p4_literal_2043912[p5_array_index_2048728_comb] ^ p4_literal_2043910[p5_array_index_2048729_comb] ^ p5_array_index_2048730_comb;
  assign p5_res7__664_comb = p4_literal_2043910[p5_res7__662_comb] ^ p4_literal_2043912[p5_res7__660_comb] ^ p4_literal_2043914[p5_res7__658_comb] ^ p4_literal_2043916[p5_res7__656_comb] ^ p4_literal_2043918[p5_res7__654_comb] ^ p4_literal_2043920[p5_res7__652_comb] ^ p5_res7__650_comb ^ p4_literal_2043923[p5_res7__648_comb] ^ p5_res7__646_comb ^ p5_array_index_2048856_comb ^ p5_array_index_2048831_comb ^ p5_array_index_2048804_comb ^ p5_array_index_2048775_comb ^ p5_array_index_2048743_comb ^ p4_literal_2043910[p5_array_index_2048728_comb] ^ p5_array_index_2048729_comb;
  assign p5_res7__666_comb = p4_literal_2043910[p5_res7__664_comb] ^ p4_literal_2043912[p5_res7__662_comb] ^ p4_literal_2043914[p5_res7__660_comb] ^ p4_literal_2043916[p5_res7__658_comb] ^ p4_literal_2043918[p5_res7__656_comb] ^ p4_literal_2043920[p5_res7__654_comb] ^ p5_res7__652_comb ^ p4_literal_2043923[p5_res7__650_comb] ^ p5_res7__648_comb ^ p5_array_index_2048867_comb ^ p5_array_index_2048843_comb ^ p5_array_index_2048817_comb ^ p5_array_index_2048789_comb ^ p5_array_index_2048760_comb ^ p4_literal_2043910[p5_array_index_2048727_comb] ^ p5_array_index_2048728_comb;
  assign p5_res7__668_comb = p4_literal_2043910[p5_res7__666_comb] ^ p4_literal_2043912[p5_res7__664_comb] ^ p4_literal_2043914[p5_res7__662_comb] ^ p4_literal_2043916[p5_res7__660_comb] ^ p4_literal_2043918[p5_res7__658_comb] ^ p4_literal_2043920[p5_res7__656_comb] ^ p5_res7__654_comb ^ p4_literal_2043923[p5_res7__652_comb] ^ p5_res7__650_comb ^ p5_array_index_2048878_comb ^ p5_array_index_2048855_comb ^ p5_array_index_2048830_comb ^ p5_array_index_2048803_comb ^ p5_array_index_2048774_comb ^ p5_array_index_2048742_comb ^ p5_array_index_2048727_comb;
  assign p5_res7__670_comb = p4_literal_2043910[p5_res7__668_comb] ^ p4_literal_2043912[p5_res7__666_comb] ^ p4_literal_2043914[p5_res7__664_comb] ^ p4_literal_2043916[p5_res7__662_comb] ^ p4_literal_2043918[p5_res7__660_comb] ^ p4_literal_2043920[p5_res7__658_comb] ^ p5_res7__656_comb ^ p4_literal_2043923[p5_res7__654_comb] ^ p5_res7__652_comb ^ p5_array_index_2048888_comb ^ p5_array_index_2048866_comb ^ p5_array_index_2048842_comb ^ p5_array_index_2048816_comb ^ p5_array_index_2048788_comb ^ p5_array_index_2048759_comb ^ p5_array_index_2048726_comb;
  assign p5_res__20_comb = {p5_res7__670_comb, p5_res7__668_comb, p5_res7__666_comb, p5_res7__664_comb, p5_res7__662_comb, p5_res7__660_comb, p5_res7__658_comb, p5_res7__656_comb, p5_res7__654_comb, p5_res7__652_comb, p5_res7__650_comb, p5_res7__648_comb, p5_res7__646_comb, p5_res7__644_comb, p5_res7__642_comb, p5_res7__640_comb};
  assign p5_xor_2048928_comb = p5_res__20_comb ^ p5_xor_2048492_comb;
  assign p5_addedKey__53_comb = p5_xor_2048928_comb ^ 128'h88f8_9bc3_a479_73c7_94e7_89a3_c509_aa16;
  assign p5_array_index_2048944_comb = p4_literal_2043896[p5_addedKey__53_comb[127:120]];
  assign p5_array_index_2048945_comb = p4_literal_2043896[p5_addedKey__53_comb[119:112]];
  assign p5_array_index_2048946_comb = p4_literal_2043896[p5_addedKey__53_comb[111:104]];
  assign p5_array_index_2048947_comb = p4_literal_2043896[p5_addedKey__53_comb[103:96]];
  assign p5_array_index_2048948_comb = p4_literal_2043896[p5_addedKey__53_comb[95:88]];
  assign p5_array_index_2048949_comb = p4_literal_2043896[p5_addedKey__53_comb[87:80]];
  assign p5_array_index_2048951_comb = p4_literal_2043896[p5_addedKey__53_comb[71:64]];
  assign p5_array_index_2048953_comb = p4_literal_2043896[p5_addedKey__53_comb[55:48]];
  assign p5_array_index_2048954_comb = p4_literal_2043896[p5_addedKey__53_comb[47:40]];
  assign p5_array_index_2048955_comb = p4_literal_2043896[p5_addedKey__53_comb[39:32]];
  assign p5_array_index_2048956_comb = p4_literal_2043896[p5_addedKey__53_comb[31:24]];
  assign p5_array_index_2048957_comb = p4_literal_2043896[p5_addedKey__53_comb[23:16]];
  assign p5_array_index_2048958_comb = p4_literal_2043896[p5_addedKey__53_comb[15:8]];
  assign p5_array_index_2048960_comb = p4_literal_2043910[p5_array_index_2048944_comb];
  assign p5_array_index_2048961_comb = p4_literal_2043912[p5_array_index_2048945_comb];
  assign p5_array_index_2048962_comb = p4_literal_2043914[p5_array_index_2048946_comb];
  assign p5_array_index_2048963_comb = p4_literal_2043916[p5_array_index_2048947_comb];
  assign p5_array_index_2048964_comb = p4_literal_2043918[p5_array_index_2048948_comb];
  assign p5_array_index_2048965_comb = p4_literal_2043920[p5_array_index_2048949_comb];
  assign p5_array_index_2048966_comb = p4_literal_2043896[p5_addedKey__53_comb[79:72]];
  assign p5_array_index_2048968_comb = p4_literal_2043896[p5_addedKey__53_comb[63:56]];
  assign p5_res7__672_comb = p5_array_index_2048960_comb ^ p5_array_index_2048961_comb ^ p5_array_index_2048962_comb ^ p5_array_index_2048963_comb ^ p5_array_index_2048964_comb ^ p5_array_index_2048965_comb ^ p5_array_index_2048966_comb ^ p4_literal_2043923[p5_array_index_2048951_comb] ^ p5_array_index_2048968_comb ^ p4_literal_2043920[p5_array_index_2048953_comb] ^ p4_literal_2043918[p5_array_index_2048954_comb] ^ p4_literal_2043916[p5_array_index_2048955_comb] ^ p4_literal_2043914[p5_array_index_2048956_comb] ^ p4_literal_2043912[p5_array_index_2048957_comb] ^ p4_literal_2043910[p5_array_index_2048958_comb] ^ p4_literal_2043896[p5_addedKey__53_comb[7:0]];
  assign p5_array_index_2048977_comb = p4_literal_2043910[p5_res7__672_comb];
  assign p5_array_index_2048978_comb = p4_literal_2043912[p5_array_index_2048944_comb];
  assign p5_array_index_2048979_comb = p4_literal_2043914[p5_array_index_2048945_comb];
  assign p5_array_index_2048980_comb = p4_literal_2043916[p5_array_index_2048946_comb];
  assign p5_array_index_2048981_comb = p4_literal_2043918[p5_array_index_2048947_comb];
  assign p5_array_index_2048982_comb = p4_literal_2043920[p5_array_index_2048948_comb];
  assign p5_res7__674_comb = p5_array_index_2048977_comb ^ p5_array_index_2048978_comb ^ p5_array_index_2048979_comb ^ p5_array_index_2048980_comb ^ p5_array_index_2048981_comb ^ p5_array_index_2048982_comb ^ p5_array_index_2048949_comb ^ p4_literal_2043923[p5_array_index_2048966_comb] ^ p5_array_index_2048951_comb ^ p4_literal_2043920[p5_array_index_2048968_comb] ^ p4_literal_2043918[p5_array_index_2048953_comb] ^ p4_literal_2043916[p5_array_index_2048954_comb] ^ p4_literal_2043914[p5_array_index_2048955_comb] ^ p4_literal_2043912[p5_array_index_2048956_comb] ^ p4_literal_2043910[p5_array_index_2048957_comb] ^ p5_array_index_2048958_comb;
  assign p5_array_index_2048992_comb = p4_literal_2043912[p5_res7__672_comb];
  assign p5_array_index_2048993_comb = p4_literal_2043914[p5_array_index_2048944_comb];
  assign p5_array_index_2048994_comb = p4_literal_2043916[p5_array_index_2048945_comb];
  assign p5_array_index_2048995_comb = p4_literal_2043918[p5_array_index_2048946_comb];
  assign p5_array_index_2048996_comb = p4_literal_2043920[p5_array_index_2048947_comb];
  assign p5_res7__676_comb = p4_literal_2043910[p5_res7__674_comb] ^ p5_array_index_2048992_comb ^ p5_array_index_2048993_comb ^ p5_array_index_2048994_comb ^ p5_array_index_2048995_comb ^ p5_array_index_2048996_comb ^ p5_array_index_2048948_comb ^ p4_literal_2043923[p5_array_index_2048949_comb] ^ p5_array_index_2048966_comb ^ p4_literal_2043920[p5_array_index_2048951_comb] ^ p4_literal_2043918[p5_array_index_2048968_comb] ^ p4_literal_2043916[p5_array_index_2048953_comb] ^ p4_literal_2043914[p5_array_index_2048954_comb] ^ p4_literal_2043912[p5_array_index_2048955_comb] ^ p4_literal_2043910[p5_array_index_2048956_comb] ^ p5_array_index_2048957_comb;
  assign p5_array_index_2049006_comb = p4_literal_2043912[p5_res7__674_comb];
  assign p5_array_index_2049007_comb = p4_literal_2043914[p5_res7__672_comb];
  assign p5_array_index_2049008_comb = p4_literal_2043916[p5_array_index_2048944_comb];
  assign p5_array_index_2049009_comb = p4_literal_2043918[p5_array_index_2048945_comb];
  assign p5_array_index_2049010_comb = p4_literal_2043920[p5_array_index_2048946_comb];
  assign p5_res7__678_comb = p4_literal_2043910[p5_res7__676_comb] ^ p5_array_index_2049006_comb ^ p5_array_index_2049007_comb ^ p5_array_index_2049008_comb ^ p5_array_index_2049009_comb ^ p5_array_index_2049010_comb ^ p5_array_index_2048947_comb ^ p4_literal_2043923[p5_array_index_2048948_comb] ^ p5_array_index_2048949_comb ^ p4_literal_2043920[p5_array_index_2048966_comb] ^ p4_literal_2043918[p5_array_index_2048951_comb] ^ p4_literal_2043916[p5_array_index_2048968_comb] ^ p4_literal_2043914[p5_array_index_2048953_comb] ^ p4_literal_2043912[p5_array_index_2048954_comb] ^ p4_literal_2043910[p5_array_index_2048955_comb] ^ p5_array_index_2048956_comb;
  assign p5_array_index_2049021_comb = p4_literal_2043914[p5_res7__674_comb];
  assign p5_array_index_2049022_comb = p4_literal_2043916[p5_res7__672_comb];
  assign p5_array_index_2049023_comb = p4_literal_2043918[p5_array_index_2048944_comb];
  assign p5_array_index_2049024_comb = p4_literal_2043920[p5_array_index_2048945_comb];
  assign p5_res7__680_comb = p4_literal_2043910[p5_res7__678_comb] ^ p4_literal_2043912[p5_res7__676_comb] ^ p5_array_index_2049021_comb ^ p5_array_index_2049022_comb ^ p5_array_index_2049023_comb ^ p5_array_index_2049024_comb ^ p5_array_index_2048946_comb ^ p4_literal_2043923[p5_array_index_2048947_comb] ^ p5_array_index_2048948_comb ^ p5_array_index_2048965_comb ^ p4_literal_2043918[p5_array_index_2048966_comb] ^ p4_literal_2043916[p5_array_index_2048951_comb] ^ p4_literal_2043914[p5_array_index_2048968_comb] ^ p4_literal_2043912[p5_array_index_2048953_comb] ^ p4_literal_2043910[p5_array_index_2048954_comb] ^ p5_array_index_2048955_comb;
  assign p5_array_index_2049034_comb = p4_literal_2043914[p5_res7__676_comb];
  assign p5_array_index_2049035_comb = p4_literal_2043916[p5_res7__674_comb];
  assign p5_array_index_2049036_comb = p4_literal_2043918[p5_res7__672_comb];
  assign p5_array_index_2049037_comb = p4_literal_2043920[p5_array_index_2048944_comb];
  assign p5_res7__682_comb = p4_literal_2043910[p5_res7__680_comb] ^ p4_literal_2043912[p5_res7__678_comb] ^ p5_array_index_2049034_comb ^ p5_array_index_2049035_comb ^ p5_array_index_2049036_comb ^ p5_array_index_2049037_comb ^ p5_array_index_2048945_comb ^ p4_literal_2043923[p5_array_index_2048946_comb] ^ p5_array_index_2048947_comb ^ p5_array_index_2048982_comb ^ p4_literal_2043918[p5_array_index_2048949_comb] ^ p4_literal_2043916[p5_array_index_2048966_comb] ^ p4_literal_2043914[p5_array_index_2048951_comb] ^ p4_literal_2043912[p5_array_index_2048968_comb] ^ p4_literal_2043910[p5_array_index_2048953_comb] ^ p5_array_index_2048954_comb;
  assign p5_array_index_2049048_comb = p4_literal_2043916[p5_res7__676_comb];
  assign p5_array_index_2049049_comb = p4_literal_2043918[p5_res7__674_comb];
  assign p5_array_index_2049050_comb = p4_literal_2043920[p5_res7__672_comb];
  assign p5_res7__684_comb = p4_literal_2043910[p5_res7__682_comb] ^ p4_literal_2043912[p5_res7__680_comb] ^ p4_literal_2043914[p5_res7__678_comb] ^ p5_array_index_2049048_comb ^ p5_array_index_2049049_comb ^ p5_array_index_2049050_comb ^ p5_array_index_2048944_comb ^ p4_literal_2043923[p5_array_index_2048945_comb] ^ p5_array_index_2048946_comb ^ p5_array_index_2048996_comb ^ p5_array_index_2048964_comb ^ p4_literal_2043916[p5_array_index_2048949_comb] ^ p4_literal_2043914[p5_array_index_2048966_comb] ^ p4_literal_2043912[p5_array_index_2048951_comb] ^ p4_literal_2043910[p5_array_index_2048968_comb] ^ p5_array_index_2048953_comb;
  assign p5_array_index_2049060_comb = p4_literal_2043916[p5_res7__678_comb];
  assign p5_array_index_2049061_comb = p4_literal_2043918[p5_res7__676_comb];
  assign p5_array_index_2049062_comb = p4_literal_2043920[p5_res7__674_comb];
  assign p5_res7__686_comb = p4_literal_2043910[p5_res7__684_comb] ^ p4_literal_2043912[p5_res7__682_comb] ^ p4_literal_2043914[p5_res7__680_comb] ^ p5_array_index_2049060_comb ^ p5_array_index_2049061_comb ^ p5_array_index_2049062_comb ^ p5_res7__672_comb ^ p4_literal_2043923[p5_array_index_2048944_comb] ^ p5_array_index_2048945_comb ^ p5_array_index_2049010_comb ^ p5_array_index_2048981_comb ^ p4_literal_2043916[p5_array_index_2048948_comb] ^ p4_literal_2043914[p5_array_index_2048949_comb] ^ p4_literal_2043912[p5_array_index_2048966_comb] ^ p4_literal_2043910[p5_array_index_2048951_comb] ^ p5_array_index_2048968_comb;
  assign p5_array_index_2049073_comb = p4_literal_2043918[p5_res7__678_comb];
  assign p5_array_index_2049074_comb = p4_literal_2043920[p5_res7__676_comb];
  assign p5_res7__688_comb = p4_literal_2043910[p5_res7__686_comb] ^ p4_literal_2043912[p5_res7__684_comb] ^ p4_literal_2043914[p5_res7__682_comb] ^ p4_literal_2043916[p5_res7__680_comb] ^ p5_array_index_2049073_comb ^ p5_array_index_2049074_comb ^ p5_res7__674_comb ^ p4_literal_2043923[p5_res7__672_comb] ^ p5_array_index_2048944_comb ^ p5_array_index_2049024_comb ^ p5_array_index_2048995_comb ^ p5_array_index_2048963_comb ^ p4_literal_2043914[p5_array_index_2048948_comb] ^ p4_literal_2043912[p5_array_index_2048949_comb] ^ p4_literal_2043910[p5_array_index_2048966_comb] ^ p5_array_index_2048951_comb;
  assign p5_array_index_2049084_comb = p4_literal_2043918[p5_res7__680_comb];
  assign p5_array_index_2049085_comb = p4_literal_2043920[p5_res7__678_comb];
  assign p5_res7__690_comb = p4_literal_2043910[p5_res7__688_comb] ^ p4_literal_2043912[p5_res7__686_comb] ^ p4_literal_2043914[p5_res7__684_comb] ^ p4_literal_2043916[p5_res7__682_comb] ^ p5_array_index_2049084_comb ^ p5_array_index_2049085_comb ^ p5_res7__676_comb ^ p4_literal_2043923[p5_res7__674_comb] ^ p5_res7__672_comb ^ p5_array_index_2049037_comb ^ p5_array_index_2049009_comb ^ p5_array_index_2048980_comb ^ p4_literal_2043914[p5_array_index_2048947_comb] ^ p4_literal_2043912[p5_array_index_2048948_comb] ^ p4_literal_2043910[p5_array_index_2048949_comb] ^ p5_array_index_2048966_comb;
  assign p5_array_index_2049096_comb = p4_literal_2043920[p5_res7__680_comb];
  assign p5_res7__692_comb = p4_literal_2043910[p5_res7__690_comb] ^ p4_literal_2043912[p5_res7__688_comb] ^ p4_literal_2043914[p5_res7__686_comb] ^ p4_literal_2043916[p5_res7__684_comb] ^ p4_literal_2043918[p5_res7__682_comb] ^ p5_array_index_2049096_comb ^ p5_res7__678_comb ^ p4_literal_2043923[p5_res7__676_comb] ^ p5_res7__674_comb ^ p5_array_index_2049050_comb ^ p5_array_index_2049023_comb ^ p5_array_index_2048994_comb ^ p5_array_index_2048962_comb ^ p4_literal_2043912[p5_array_index_2048947_comb] ^ p4_literal_2043910[p5_array_index_2048948_comb] ^ p5_array_index_2048949_comb;
  assign p5_array_index_2049106_comb = p4_literal_2043920[p5_res7__682_comb];
  assign p5_res7__694_comb = p4_literal_2043910[p5_res7__692_comb] ^ p4_literal_2043912[p5_res7__690_comb] ^ p4_literal_2043914[p5_res7__688_comb] ^ p4_literal_2043916[p5_res7__686_comb] ^ p4_literal_2043918[p5_res7__684_comb] ^ p5_array_index_2049106_comb ^ p5_res7__680_comb ^ p4_literal_2043923[p5_res7__678_comb] ^ p5_res7__676_comb ^ p5_array_index_2049062_comb ^ p5_array_index_2049036_comb ^ p5_array_index_2049008_comb ^ p5_array_index_2048979_comb ^ p4_literal_2043912[p5_array_index_2048946_comb] ^ p4_literal_2043910[p5_array_index_2048947_comb] ^ p5_array_index_2048948_comb;
  assign p5_res7__696_comb = p4_literal_2043910[p5_res7__694_comb] ^ p4_literal_2043912[p5_res7__692_comb] ^ p4_literal_2043914[p5_res7__690_comb] ^ p4_literal_2043916[p5_res7__688_comb] ^ p4_literal_2043918[p5_res7__686_comb] ^ p4_literal_2043920[p5_res7__684_comb] ^ p5_res7__682_comb ^ p4_literal_2043923[p5_res7__680_comb] ^ p5_res7__678_comb ^ p5_array_index_2049074_comb ^ p5_array_index_2049049_comb ^ p5_array_index_2049022_comb ^ p5_array_index_2048993_comb ^ p5_array_index_2048961_comb ^ p4_literal_2043910[p5_array_index_2048946_comb] ^ p5_array_index_2048947_comb;
  assign p5_res7__698_comb = p4_literal_2043910[p5_res7__696_comb] ^ p4_literal_2043912[p5_res7__694_comb] ^ p4_literal_2043914[p5_res7__692_comb] ^ p4_literal_2043916[p5_res7__690_comb] ^ p4_literal_2043918[p5_res7__688_comb] ^ p4_literal_2043920[p5_res7__686_comb] ^ p5_res7__684_comb ^ p4_literal_2043923[p5_res7__682_comb] ^ p5_res7__680_comb ^ p5_array_index_2049085_comb ^ p5_array_index_2049061_comb ^ p5_array_index_2049035_comb ^ p5_array_index_2049007_comb ^ p5_array_index_2048978_comb ^ p4_literal_2043910[p5_array_index_2048945_comb] ^ p5_array_index_2048946_comb;
  assign p5_res7__700_comb = p4_literal_2043910[p5_res7__698_comb] ^ p4_literal_2043912[p5_res7__696_comb] ^ p4_literal_2043914[p5_res7__694_comb] ^ p4_literal_2043916[p5_res7__692_comb] ^ p4_literal_2043918[p5_res7__690_comb] ^ p4_literal_2043920[p5_res7__688_comb] ^ p5_res7__686_comb ^ p4_literal_2043923[p5_res7__684_comb] ^ p5_res7__682_comb ^ p5_array_index_2049096_comb ^ p5_array_index_2049073_comb ^ p5_array_index_2049048_comb ^ p5_array_index_2049021_comb ^ p5_array_index_2048992_comb ^ p5_array_index_2048960_comb ^ p5_array_index_2048945_comb;
  assign p5_res7__702_comb = p4_literal_2043910[p5_res7__700_comb] ^ p4_literal_2043912[p5_res7__698_comb] ^ p4_literal_2043914[p5_res7__696_comb] ^ p4_literal_2043916[p5_res7__694_comb] ^ p4_literal_2043918[p5_res7__692_comb] ^ p4_literal_2043920[p5_res7__690_comb] ^ p5_res7__688_comb ^ p4_literal_2043923[p5_res7__686_comb] ^ p5_res7__684_comb ^ p5_array_index_2049106_comb ^ p5_array_index_2049084_comb ^ p5_array_index_2049060_comb ^ p5_array_index_2049034_comb ^ p5_array_index_2049006_comb ^ p5_array_index_2048977_comb ^ p5_array_index_2048944_comb;
  assign p5_res__21_comb = {p5_res7__702_comb, p5_res7__700_comb, p5_res7__698_comb, p5_res7__696_comb, p5_res7__694_comb, p5_res7__692_comb, p5_res7__690_comb, p5_res7__688_comb, p5_res7__686_comb, p5_res7__684_comb, p5_res7__682_comb, p5_res7__680_comb, p5_res7__678_comb, p5_res7__676_comb, p5_res7__674_comb, p5_res7__672_comb};
  assign p5_xor_2049146_comb = p5_res__21_comb ^ p5_xor_2048710_comb;
  assign p5_addedKey__54_comb = p5_xor_2049146_comb ^ 128'he65a_edb1_c831_097f_c9c0_34b3_188d_3e17;
  assign p5_array_index_2049162_comb = p4_literal_2043896[p5_addedKey__54_comb[127:120]];
  assign p5_array_index_2049163_comb = p4_literal_2043896[p5_addedKey__54_comb[119:112]];
  assign p5_array_index_2049164_comb = p4_literal_2043896[p5_addedKey__54_comb[111:104]];
  assign p5_array_index_2049165_comb = p4_literal_2043896[p5_addedKey__54_comb[103:96]];
  assign p5_array_index_2049166_comb = p4_literal_2043896[p5_addedKey__54_comb[95:88]];
  assign p5_array_index_2049167_comb = p4_literal_2043896[p5_addedKey__54_comb[87:80]];
  assign p5_array_index_2049169_comb = p4_literal_2043896[p5_addedKey__54_comb[71:64]];
  assign p5_array_index_2049171_comb = p4_literal_2043896[p5_addedKey__54_comb[55:48]];
  assign p5_array_index_2049172_comb = p4_literal_2043896[p5_addedKey__54_comb[47:40]];
  assign p5_array_index_2049173_comb = p4_literal_2043896[p5_addedKey__54_comb[39:32]];
  assign p5_array_index_2049174_comb = p4_literal_2043896[p5_addedKey__54_comb[31:24]];
  assign p5_array_index_2049175_comb = p4_literal_2043896[p5_addedKey__54_comb[23:16]];
  assign p5_array_index_2049176_comb = p4_literal_2043896[p5_addedKey__54_comb[15:8]];
  assign p5_array_index_2049178_comb = p4_literal_2043910[p5_array_index_2049162_comb];
  assign p5_array_index_2049179_comb = p4_literal_2043912[p5_array_index_2049163_comb];
  assign p5_array_index_2049180_comb = p4_literal_2043914[p5_array_index_2049164_comb];
  assign p5_array_index_2049181_comb = p4_literal_2043916[p5_array_index_2049165_comb];
  assign p5_array_index_2049182_comb = p4_literal_2043918[p5_array_index_2049166_comb];
  assign p5_array_index_2049183_comb = p4_literal_2043920[p5_array_index_2049167_comb];
  assign p5_array_index_2049184_comb = p4_literal_2043896[p5_addedKey__54_comb[79:72]];
  assign p5_array_index_2049186_comb = p4_literal_2043896[p5_addedKey__54_comb[63:56]];
  assign p5_res7__704_comb = p5_array_index_2049178_comb ^ p5_array_index_2049179_comb ^ p5_array_index_2049180_comb ^ p5_array_index_2049181_comb ^ p5_array_index_2049182_comb ^ p5_array_index_2049183_comb ^ p5_array_index_2049184_comb ^ p4_literal_2043923[p5_array_index_2049169_comb] ^ p5_array_index_2049186_comb ^ p4_literal_2043920[p5_array_index_2049171_comb] ^ p4_literal_2043918[p5_array_index_2049172_comb] ^ p4_literal_2043916[p5_array_index_2049173_comb] ^ p4_literal_2043914[p5_array_index_2049174_comb] ^ p4_literal_2043912[p5_array_index_2049175_comb] ^ p4_literal_2043910[p5_array_index_2049176_comb] ^ p4_literal_2043896[p5_addedKey__54_comb[7:0]];
  assign p5_array_index_2049195_comb = p4_literal_2043910[p5_res7__704_comb];
  assign p5_array_index_2049196_comb = p4_literal_2043912[p5_array_index_2049162_comb];
  assign p5_array_index_2049197_comb = p4_literal_2043914[p5_array_index_2049163_comb];
  assign p5_array_index_2049198_comb = p4_literal_2043916[p5_array_index_2049164_comb];
  assign p5_array_index_2049199_comb = p4_literal_2043918[p5_array_index_2049165_comb];
  assign p5_array_index_2049200_comb = p4_literal_2043920[p5_array_index_2049166_comb];
  assign p5_res7__706_comb = p5_array_index_2049195_comb ^ p5_array_index_2049196_comb ^ p5_array_index_2049197_comb ^ p5_array_index_2049198_comb ^ p5_array_index_2049199_comb ^ p5_array_index_2049200_comb ^ p5_array_index_2049167_comb ^ p4_literal_2043923[p5_array_index_2049184_comb] ^ p5_array_index_2049169_comb ^ p4_literal_2043920[p5_array_index_2049186_comb] ^ p4_literal_2043918[p5_array_index_2049171_comb] ^ p4_literal_2043916[p5_array_index_2049172_comb] ^ p4_literal_2043914[p5_array_index_2049173_comb] ^ p4_literal_2043912[p5_array_index_2049174_comb] ^ p4_literal_2043910[p5_array_index_2049175_comb] ^ p5_array_index_2049176_comb;
  assign p5_array_index_2049210_comb = p4_literal_2043912[p5_res7__704_comb];
  assign p5_array_index_2049211_comb = p4_literal_2043914[p5_array_index_2049162_comb];
  assign p5_array_index_2049212_comb = p4_literal_2043916[p5_array_index_2049163_comb];
  assign p5_array_index_2049213_comb = p4_literal_2043918[p5_array_index_2049164_comb];
  assign p5_array_index_2049214_comb = p4_literal_2043920[p5_array_index_2049165_comb];
  assign p5_res7__708_comb = p4_literal_2043910[p5_res7__706_comb] ^ p5_array_index_2049210_comb ^ p5_array_index_2049211_comb ^ p5_array_index_2049212_comb ^ p5_array_index_2049213_comb ^ p5_array_index_2049214_comb ^ p5_array_index_2049166_comb ^ p4_literal_2043923[p5_array_index_2049167_comb] ^ p5_array_index_2049184_comb ^ p4_literal_2043920[p5_array_index_2049169_comb] ^ p4_literal_2043918[p5_array_index_2049186_comb] ^ p4_literal_2043916[p5_array_index_2049171_comb] ^ p4_literal_2043914[p5_array_index_2049172_comb] ^ p4_literal_2043912[p5_array_index_2049173_comb] ^ p4_literal_2043910[p5_array_index_2049174_comb] ^ p5_array_index_2049175_comb;

  // Registers for pipe stage 5:
  reg [127:0] p5_encoded;
  reg [127:0] p5_bit_slice_2043893;
  reg [127:0] p5_bit_slice_2044119;
  reg [127:0] p5_k3;
  reg [127:0] p5_k2;
  reg [127:0] p5_k5;
  reg [127:0] p5_k4;
  reg [127:0] p5_xor_2048928;
  reg [127:0] p5_xor_2049146;
  reg [7:0] p5_array_index_2049162;
  reg [7:0] p5_array_index_2049163;
  reg [7:0] p5_array_index_2049164;
  reg [7:0] p5_array_index_2049165;
  reg [7:0] p5_array_index_2049166;
  reg [7:0] p5_array_index_2049167;
  reg [7:0] p5_array_index_2049169;
  reg [7:0] p5_array_index_2049171;
  reg [7:0] p5_array_index_2049172;
  reg [7:0] p5_array_index_2049173;
  reg [7:0] p5_array_index_2049174;
  reg [7:0] p5_array_index_2049178;
  reg [7:0] p5_array_index_2049179;
  reg [7:0] p5_array_index_2049180;
  reg [7:0] p5_array_index_2049181;
  reg [7:0] p5_array_index_2049182;
  reg [7:0] p5_array_index_2049183;
  reg [7:0] p5_array_index_2049184;
  reg [7:0] p5_array_index_2049186;
  reg [7:0] p5_res7__704;
  reg [7:0] p5_array_index_2049195;
  reg [7:0] p5_array_index_2049196;
  reg [7:0] p5_array_index_2049197;
  reg [7:0] p5_array_index_2049198;
  reg [7:0] p5_array_index_2049199;
  reg [7:0] p5_array_index_2049200;
  reg [7:0] p5_res7__706;
  reg [7:0] p5_array_index_2049210;
  reg [7:0] p5_array_index_2049211;
  reg [7:0] p5_array_index_2049212;
  reg [7:0] p5_array_index_2049213;
  reg [7:0] p5_array_index_2049214;
  reg [7:0] p5_res7__708;
  reg [7:0] p6_literal_2043896[256];
  reg [7:0] p6_literal_2043910[256];
  reg [7:0] p6_literal_2043912[256];
  reg [7:0] p6_literal_2043914[256];
  reg [7:0] p6_literal_2043916[256];
  reg [7:0] p6_literal_2043918[256];
  reg [7:0] p6_literal_2043920[256];
  reg [7:0] p6_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p5_encoded <= p4_encoded;
    p5_bit_slice_2043893 <= p4_bit_slice_2043893;
    p5_bit_slice_2044119 <= p4_bit_slice_2044119;
    p5_k3 <= p4_k3;
    p5_k2 <= p4_k2;
    p5_k5 <= p4_k5;
    p5_k4 <= p4_k4;
    p5_xor_2048928 <= p5_xor_2048928_comb;
    p5_xor_2049146 <= p5_xor_2049146_comb;
    p5_array_index_2049162 <= p5_array_index_2049162_comb;
    p5_array_index_2049163 <= p5_array_index_2049163_comb;
    p5_array_index_2049164 <= p5_array_index_2049164_comb;
    p5_array_index_2049165 <= p5_array_index_2049165_comb;
    p5_array_index_2049166 <= p5_array_index_2049166_comb;
    p5_array_index_2049167 <= p5_array_index_2049167_comb;
    p5_array_index_2049169 <= p5_array_index_2049169_comb;
    p5_array_index_2049171 <= p5_array_index_2049171_comb;
    p5_array_index_2049172 <= p5_array_index_2049172_comb;
    p5_array_index_2049173 <= p5_array_index_2049173_comb;
    p5_array_index_2049174 <= p5_array_index_2049174_comb;
    p5_array_index_2049178 <= p5_array_index_2049178_comb;
    p5_array_index_2049179 <= p5_array_index_2049179_comb;
    p5_array_index_2049180 <= p5_array_index_2049180_comb;
    p5_array_index_2049181 <= p5_array_index_2049181_comb;
    p5_array_index_2049182 <= p5_array_index_2049182_comb;
    p5_array_index_2049183 <= p5_array_index_2049183_comb;
    p5_array_index_2049184 <= p5_array_index_2049184_comb;
    p5_array_index_2049186 <= p5_array_index_2049186_comb;
    p5_res7__704 <= p5_res7__704_comb;
    p5_array_index_2049195 <= p5_array_index_2049195_comb;
    p5_array_index_2049196 <= p5_array_index_2049196_comb;
    p5_array_index_2049197 <= p5_array_index_2049197_comb;
    p5_array_index_2049198 <= p5_array_index_2049198_comb;
    p5_array_index_2049199 <= p5_array_index_2049199_comb;
    p5_array_index_2049200 <= p5_array_index_2049200_comb;
    p5_res7__706 <= p5_res7__706_comb;
    p5_array_index_2049210 <= p5_array_index_2049210_comb;
    p5_array_index_2049211 <= p5_array_index_2049211_comb;
    p5_array_index_2049212 <= p5_array_index_2049212_comb;
    p5_array_index_2049213 <= p5_array_index_2049213_comb;
    p5_array_index_2049214 <= p5_array_index_2049214_comb;
    p5_res7__708 <= p5_res7__708_comb;
    p6_literal_2043896 <= p5_literal_2043896;
    p6_literal_2043910 <= p5_literal_2043910;
    p6_literal_2043912 <= p5_literal_2043912;
    p6_literal_2043914 <= p5_literal_2043914;
    p6_literal_2043916 <= p5_literal_2043916;
    p6_literal_2043918 <= p5_literal_2043918;
    p6_literal_2043920 <= p5_literal_2043920;
    p6_literal_2043923 <= p5_literal_2043923;
  end

  // ===== Pipe stage 6:
  wire [7:0] p6_array_index_2049324_comb;
  wire [7:0] p6_array_index_2049325_comb;
  wire [7:0] p6_array_index_2049326_comb;
  wire [7:0] p6_array_index_2049327_comb;
  wire [7:0] p6_array_index_2049328_comb;
  wire [7:0] p6_res7__710_comb;
  wire [7:0] p6_array_index_2049339_comb;
  wire [7:0] p6_array_index_2049340_comb;
  wire [7:0] p6_array_index_2049341_comb;
  wire [7:0] p6_array_index_2049342_comb;
  wire [7:0] p6_res7__712_comb;
  wire [7:0] p6_array_index_2049352_comb;
  wire [7:0] p6_array_index_2049353_comb;
  wire [7:0] p6_array_index_2049354_comb;
  wire [7:0] p6_array_index_2049355_comb;
  wire [7:0] p6_res7__714_comb;
  wire [7:0] p6_array_index_2049366_comb;
  wire [7:0] p6_array_index_2049367_comb;
  wire [7:0] p6_array_index_2049368_comb;
  wire [7:0] p6_res7__716_comb;
  wire [7:0] p6_array_index_2049378_comb;
  wire [7:0] p6_array_index_2049379_comb;
  wire [7:0] p6_array_index_2049380_comb;
  wire [7:0] p6_res7__718_comb;
  wire [7:0] p6_array_index_2049391_comb;
  wire [7:0] p6_array_index_2049392_comb;
  wire [7:0] p6_res7__720_comb;
  wire [7:0] p6_array_index_2049402_comb;
  wire [7:0] p6_array_index_2049403_comb;
  wire [7:0] p6_res7__722_comb;
  wire [7:0] p6_array_index_2049414_comb;
  wire [7:0] p6_res7__724_comb;
  wire [7:0] p6_array_index_2049424_comb;
  wire [7:0] p6_res7__726_comb;
  wire [7:0] p6_res7__728_comb;
  wire [7:0] p6_res7__730_comb;
  wire [7:0] p6_res7__732_comb;
  wire [7:0] p6_res7__734_comb;
  wire [127:0] p6_res__22_comb;
  wire [127:0] p6_k7_comb;
  wire [127:0] p6_addedKey__55_comb;
  wire [7:0] p6_array_index_2049480_comb;
  wire [7:0] p6_array_index_2049481_comb;
  wire [7:0] p6_array_index_2049482_comb;
  wire [7:0] p6_array_index_2049483_comb;
  wire [7:0] p6_array_index_2049484_comb;
  wire [7:0] p6_array_index_2049485_comb;
  wire [7:0] p6_array_index_2049487_comb;
  wire [7:0] p6_array_index_2049489_comb;
  wire [7:0] p6_array_index_2049490_comb;
  wire [7:0] p6_array_index_2049491_comb;
  wire [7:0] p6_array_index_2049492_comb;
  wire [7:0] p6_array_index_2049493_comb;
  wire [7:0] p6_array_index_2049494_comb;
  wire [7:0] p6_array_index_2049496_comb;
  wire [7:0] p6_array_index_2049497_comb;
  wire [7:0] p6_array_index_2049498_comb;
  wire [7:0] p6_array_index_2049499_comb;
  wire [7:0] p6_array_index_2049500_comb;
  wire [7:0] p6_array_index_2049501_comb;
  wire [7:0] p6_array_index_2049502_comb;
  wire [7:0] p6_array_index_2049504_comb;
  wire [7:0] p6_res7__736_comb;
  wire [7:0] p6_array_index_2049513_comb;
  wire [7:0] p6_array_index_2049514_comb;
  wire [7:0] p6_array_index_2049515_comb;
  wire [7:0] p6_array_index_2049516_comb;
  wire [7:0] p6_array_index_2049517_comb;
  wire [7:0] p6_array_index_2049518_comb;
  wire [7:0] p6_res7__738_comb;
  wire [7:0] p6_array_index_2049528_comb;
  wire [7:0] p6_array_index_2049529_comb;
  wire [7:0] p6_array_index_2049530_comb;
  wire [7:0] p6_array_index_2049531_comb;
  wire [7:0] p6_array_index_2049532_comb;
  wire [7:0] p6_res7__740_comb;
  wire [7:0] p6_array_index_2049542_comb;
  wire [7:0] p6_array_index_2049543_comb;
  wire [7:0] p6_array_index_2049544_comb;
  wire [7:0] p6_array_index_2049545_comb;
  wire [7:0] p6_array_index_2049546_comb;
  wire [7:0] p6_res7__742_comb;
  wire [7:0] p6_array_index_2049557_comb;
  wire [7:0] p6_array_index_2049558_comb;
  wire [7:0] p6_array_index_2049559_comb;
  wire [7:0] p6_array_index_2049560_comb;
  wire [7:0] p6_res7__744_comb;
  wire [7:0] p6_array_index_2049570_comb;
  wire [7:0] p6_array_index_2049571_comb;
  wire [7:0] p6_array_index_2049572_comb;
  wire [7:0] p6_array_index_2049573_comb;
  wire [7:0] p6_res7__746_comb;
  wire [7:0] p6_array_index_2049584_comb;
  wire [7:0] p6_array_index_2049585_comb;
  wire [7:0] p6_array_index_2049586_comb;
  wire [7:0] p6_res7__748_comb;
  wire [7:0] p6_array_index_2049596_comb;
  wire [7:0] p6_array_index_2049597_comb;
  wire [7:0] p6_array_index_2049598_comb;
  wire [7:0] p6_res7__750_comb;
  wire [7:0] p6_array_index_2049609_comb;
  wire [7:0] p6_array_index_2049610_comb;
  wire [7:0] p6_res7__752_comb;
  wire [7:0] p6_array_index_2049620_comb;
  wire [7:0] p6_array_index_2049621_comb;
  wire [7:0] p6_res7__754_comb;
  wire [7:0] p6_array_index_2049632_comb;
  wire [7:0] p6_res7__756_comb;
  wire [7:0] p6_array_index_2049642_comb;
  wire [7:0] p6_res7__758_comb;
  wire [7:0] p6_res7__760_comb;
  wire [7:0] p6_res7__762_comb;
  wire [7:0] p6_res7__764_comb;
  wire [7:0] p6_res7__766_comb;
  wire [127:0] p6_res__23_comb;
  wire [127:0] p6_k6_comb;
  wire [127:0] p6_addedKey__56_comb;
  wire [7:0] p6_array_index_2049698_comb;
  wire [7:0] p6_array_index_2049699_comb;
  wire [7:0] p6_array_index_2049700_comb;
  wire [7:0] p6_array_index_2049701_comb;
  wire [7:0] p6_array_index_2049702_comb;
  wire [7:0] p6_array_index_2049703_comb;
  wire [7:0] p6_array_index_2049705_comb;
  wire [7:0] p6_array_index_2049707_comb;
  wire [7:0] p6_array_index_2049708_comb;
  wire [7:0] p6_array_index_2049709_comb;
  wire [7:0] p6_array_index_2049710_comb;
  wire [7:0] p6_array_index_2049711_comb;
  wire [7:0] p6_array_index_2049712_comb;
  wire [7:0] p6_array_index_2049714_comb;
  wire [7:0] p6_array_index_2049715_comb;
  wire [7:0] p6_array_index_2049716_comb;
  wire [7:0] p6_array_index_2049717_comb;
  wire [7:0] p6_array_index_2049718_comb;
  wire [7:0] p6_array_index_2049719_comb;
  wire [7:0] p6_array_index_2049720_comb;
  wire [7:0] p6_array_index_2049722_comb;
  wire [7:0] p6_res7__768_comb;
  wire [7:0] p6_array_index_2049731_comb;
  wire [7:0] p6_array_index_2049732_comb;
  wire [7:0] p6_array_index_2049733_comb;
  wire [7:0] p6_array_index_2049734_comb;
  wire [7:0] p6_array_index_2049735_comb;
  wire [7:0] p6_array_index_2049736_comb;
  wire [7:0] p6_res7__770_comb;
  wire [7:0] p6_array_index_2049746_comb;
  wire [7:0] p6_array_index_2049747_comb;
  wire [7:0] p6_array_index_2049748_comb;
  wire [7:0] p6_array_index_2049749_comb;
  wire [7:0] p6_array_index_2049750_comb;
  wire [7:0] p6_res7__772_comb;
  wire [7:0] p6_array_index_2049760_comb;
  wire [7:0] p6_array_index_2049761_comb;
  wire [7:0] p6_array_index_2049762_comb;
  wire [7:0] p6_array_index_2049763_comb;
  wire [7:0] p6_array_index_2049764_comb;
  wire [7:0] p6_res7__774_comb;
  wire [7:0] p6_array_index_2049775_comb;
  wire [7:0] p6_array_index_2049776_comb;
  wire [7:0] p6_array_index_2049777_comb;
  wire [7:0] p6_array_index_2049778_comb;
  wire [7:0] p6_res7__776_comb;
  wire [7:0] p6_array_index_2049788_comb;
  wire [7:0] p6_array_index_2049789_comb;
  wire [7:0] p6_array_index_2049790_comb;
  wire [7:0] p6_array_index_2049791_comb;
  wire [7:0] p6_res7__778_comb;
  wire [7:0] p6_array_index_2049802_comb;
  wire [7:0] p6_array_index_2049803_comb;
  wire [7:0] p6_array_index_2049804_comb;
  wire [7:0] p6_res7__780_comb;
  wire [7:0] p6_array_index_2049814_comb;
  wire [7:0] p6_array_index_2049815_comb;
  wire [7:0] p6_array_index_2049816_comb;
  wire [7:0] p6_res7__782_comb;
  wire [7:0] p6_array_index_2049827_comb;
  wire [7:0] p6_array_index_2049828_comb;
  wire [7:0] p6_res7__784_comb;
  wire [7:0] p6_array_index_2049838_comb;
  wire [7:0] p6_array_index_2049839_comb;
  wire [7:0] p6_res7__786_comb;
  wire [7:0] p6_array_index_2049850_comb;
  wire [7:0] p6_res7__788_comb;
  wire [7:0] p6_array_index_2049860_comb;
  wire [7:0] p6_res7__790_comb;
  wire [7:0] p6_res7__792_comb;
  wire [7:0] p6_res7__794_comb;
  wire [7:0] p6_res7__796_comb;
  wire [7:0] p6_res7__798_comb;
  wire [127:0] p6_res__24_comb;
  wire [127:0] p6_xor_2049900_comb;
  wire [127:0] p6_addedKey__57_comb;
  wire [7:0] p6_array_index_2049916_comb;
  wire [7:0] p6_array_index_2049917_comb;
  wire [7:0] p6_array_index_2049918_comb;
  wire [7:0] p6_array_index_2049919_comb;
  wire [7:0] p6_array_index_2049920_comb;
  wire [7:0] p6_array_index_2049921_comb;
  wire [7:0] p6_array_index_2049923_comb;
  wire [7:0] p6_array_index_2049925_comb;
  wire [7:0] p6_array_index_2049926_comb;
  wire [7:0] p6_array_index_2049927_comb;
  wire [7:0] p6_array_index_2049928_comb;
  wire [7:0] p6_array_index_2049929_comb;
  wire [7:0] p6_array_index_2049930_comb;
  wire [7:0] p6_array_index_2049932_comb;
  wire [7:0] p6_array_index_2049933_comb;
  wire [7:0] p6_array_index_2049934_comb;
  wire [7:0] p6_array_index_2049935_comb;
  wire [7:0] p6_array_index_2049936_comb;
  wire [7:0] p6_array_index_2049937_comb;
  wire [7:0] p6_array_index_2049938_comb;
  wire [7:0] p6_array_index_2049940_comb;
  wire [7:0] p6_res7__800_comb;
  wire [7:0] p6_array_index_2049949_comb;
  wire [7:0] p6_array_index_2049950_comb;
  wire [7:0] p6_array_index_2049951_comb;
  wire [7:0] p6_array_index_2049952_comb;
  wire [7:0] p6_array_index_2049953_comb;
  wire [7:0] p6_array_index_2049954_comb;
  wire [7:0] p6_res7__802_comb;
  wire [7:0] p6_array_index_2049964_comb;
  wire [7:0] p6_array_index_2049965_comb;
  wire [7:0] p6_array_index_2049966_comb;
  wire [7:0] p6_array_index_2049967_comb;
  wire [7:0] p6_array_index_2049968_comb;
  wire [7:0] p6_res7__804_comb;
  wire [7:0] p6_array_index_2049978_comb;
  wire [7:0] p6_array_index_2049979_comb;
  wire [7:0] p6_array_index_2049980_comb;
  wire [7:0] p6_array_index_2049981_comb;
  wire [7:0] p6_array_index_2049982_comb;
  wire [7:0] p6_res7__806_comb;
  wire [7:0] p6_array_index_2049993_comb;
  wire [7:0] p6_array_index_2049994_comb;
  wire [7:0] p6_array_index_2049995_comb;
  wire [7:0] p6_array_index_2049996_comb;
  wire [7:0] p6_res7__808_comb;
  wire [7:0] p6_array_index_2050006_comb;
  wire [7:0] p6_array_index_2050007_comb;
  wire [7:0] p6_array_index_2050008_comb;
  wire [7:0] p6_array_index_2050009_comb;
  wire [7:0] p6_res7__810_comb;
  wire [7:0] p6_array_index_2050020_comb;
  wire [7:0] p6_array_index_2050021_comb;
  wire [7:0] p6_array_index_2050022_comb;
  wire [7:0] p6_res7__812_comb;
  wire [7:0] p6_array_index_2050032_comb;
  wire [7:0] p6_array_index_2050033_comb;
  wire [7:0] p6_array_index_2050034_comb;
  wire [7:0] p6_res7__814_comb;
  wire [7:0] p6_array_index_2050045_comb;
  wire [7:0] p6_array_index_2050046_comb;
  wire [7:0] p6_res7__816_comb;
  wire [7:0] p6_array_index_2050056_comb;
  wire [7:0] p6_array_index_2050057_comb;
  wire [7:0] p6_res7__818_comb;
  wire [7:0] p6_array_index_2050068_comb;
  wire [7:0] p6_res7__820_comb;
  wire [7:0] p6_array_index_2050078_comb;
  wire [7:0] p6_res7__822_comb;
  wire [7:0] p6_res7__824_comb;
  wire [7:0] p6_res7__826_comb;
  wire [7:0] p6_res7__828_comb;
  wire [7:0] p6_res7__830_comb;
  wire [127:0] p6_res__25_comb;
  wire [127:0] p6_xor_2050118_comb;
  wire [127:0] p6_addedKey__58_comb;
  wire [7:0] p6_array_index_2050134_comb;
  wire [7:0] p6_array_index_2050135_comb;
  wire [7:0] p6_array_index_2050136_comb;
  wire [7:0] p6_array_index_2050137_comb;
  wire [7:0] p6_array_index_2050138_comb;
  wire [7:0] p6_array_index_2050139_comb;
  wire [7:0] p6_array_index_2050141_comb;
  wire [7:0] p6_array_index_2050143_comb;
  wire [7:0] p6_array_index_2050144_comb;
  wire [7:0] p6_array_index_2050145_comb;
  wire [7:0] p6_array_index_2050146_comb;
  wire [7:0] p6_array_index_2050147_comb;
  wire [7:0] p6_array_index_2050148_comb;
  wire [7:0] p6_array_index_2050150_comb;
  wire [7:0] p6_array_index_2050151_comb;
  wire [7:0] p6_array_index_2050152_comb;
  wire [7:0] p6_array_index_2050153_comb;
  wire [7:0] p6_array_index_2050154_comb;
  wire [7:0] p6_array_index_2050155_comb;
  wire [7:0] p6_array_index_2050156_comb;
  wire [7:0] p6_array_index_2050158_comb;
  wire [7:0] p6_res7__832_comb;
  wire [7:0] p6_array_index_2050167_comb;
  wire [7:0] p6_array_index_2050168_comb;
  wire [7:0] p6_array_index_2050169_comb;
  wire [7:0] p6_array_index_2050170_comb;
  wire [7:0] p6_array_index_2050171_comb;
  wire [7:0] p6_array_index_2050172_comb;
  wire [7:0] p6_res7__834_comb;
  wire [7:0] p6_array_index_2050182_comb;
  wire [7:0] p6_array_index_2050183_comb;
  wire [7:0] p6_array_index_2050184_comb;
  wire [7:0] p6_array_index_2050185_comb;
  wire [7:0] p6_array_index_2050186_comb;
  wire [7:0] p6_res7__836_comb;
  wire [7:0] p6_array_index_2050196_comb;
  wire [7:0] p6_array_index_2050197_comb;
  wire [7:0] p6_array_index_2050198_comb;
  wire [7:0] p6_array_index_2050199_comb;
  wire [7:0] p6_array_index_2050200_comb;
  wire [7:0] p6_res7__838_comb;
  wire [7:0] p6_array_index_2050211_comb;
  wire [7:0] p6_array_index_2050212_comb;
  wire [7:0] p6_array_index_2050213_comb;
  wire [7:0] p6_array_index_2050214_comb;
  wire [7:0] p6_res7__840_comb;
  wire [7:0] p6_array_index_2050224_comb;
  wire [7:0] p6_array_index_2050225_comb;
  wire [7:0] p6_array_index_2050226_comb;
  wire [7:0] p6_array_index_2050227_comb;
  wire [7:0] p6_res7__842_comb;
  wire [7:0] p6_array_index_2050238_comb;
  wire [7:0] p6_array_index_2050239_comb;
  wire [7:0] p6_array_index_2050240_comb;
  wire [7:0] p6_res7__844_comb;
  wire [7:0] p6_array_index_2050250_comb;
  wire [7:0] p6_array_index_2050251_comb;
  wire [7:0] p6_array_index_2050252_comb;
  wire [7:0] p6_res7__846_comb;
  wire [7:0] p6_array_index_2050263_comb;
  wire [7:0] p6_array_index_2050264_comb;
  wire [7:0] p6_res7__848_comb;
  wire [7:0] p6_array_index_2050274_comb;
  wire [7:0] p6_array_index_2050275_comb;
  wire [7:0] p6_res7__850_comb;
  wire [7:0] p6_array_index_2050281_comb;
  wire [7:0] p6_array_index_2050282_comb;
  wire [7:0] p6_array_index_2050283_comb;
  wire [7:0] p6_array_index_2050284_comb;
  wire [7:0] p6_array_index_2050285_comb;
  wire [7:0] p6_array_index_2050286_comb;
  wire [7:0] p6_array_index_2050287_comb;
  wire [7:0] p6_array_index_2050288_comb;
  wire [7:0] p6_array_index_2050289_comb;
  assign p6_array_index_2049324_comb = p5_literal_2043912[p5_res7__706];
  assign p6_array_index_2049325_comb = p5_literal_2043914[p5_res7__704];
  assign p6_array_index_2049326_comb = p5_literal_2043916[p5_array_index_2049162];
  assign p6_array_index_2049327_comb = p5_literal_2043918[p5_array_index_2049163];
  assign p6_array_index_2049328_comb = p5_literal_2043920[p5_array_index_2049164];
  assign p6_res7__710_comb = p5_literal_2043910[p5_res7__708] ^ p6_array_index_2049324_comb ^ p6_array_index_2049325_comb ^ p6_array_index_2049326_comb ^ p6_array_index_2049327_comb ^ p6_array_index_2049328_comb ^ p5_array_index_2049165 ^ p5_literal_2043923[p5_array_index_2049166] ^ p5_array_index_2049167 ^ p5_literal_2043920[p5_array_index_2049184] ^ p5_literal_2043918[p5_array_index_2049169] ^ p5_literal_2043916[p5_array_index_2049186] ^ p5_literal_2043914[p5_array_index_2049171] ^ p5_literal_2043912[p5_array_index_2049172] ^ p5_literal_2043910[p5_array_index_2049173] ^ p5_array_index_2049174;
  assign p6_array_index_2049339_comb = p5_literal_2043914[p5_res7__706];
  assign p6_array_index_2049340_comb = p5_literal_2043916[p5_res7__704];
  assign p6_array_index_2049341_comb = p5_literal_2043918[p5_array_index_2049162];
  assign p6_array_index_2049342_comb = p5_literal_2043920[p5_array_index_2049163];
  assign p6_res7__712_comb = p5_literal_2043910[p6_res7__710_comb] ^ p5_literal_2043912[p5_res7__708] ^ p6_array_index_2049339_comb ^ p6_array_index_2049340_comb ^ p6_array_index_2049341_comb ^ p6_array_index_2049342_comb ^ p5_array_index_2049164 ^ p5_literal_2043923[p5_array_index_2049165] ^ p5_array_index_2049166 ^ p5_array_index_2049183 ^ p5_literal_2043918[p5_array_index_2049184] ^ p5_literal_2043916[p5_array_index_2049169] ^ p5_literal_2043914[p5_array_index_2049186] ^ p5_literal_2043912[p5_array_index_2049171] ^ p5_literal_2043910[p5_array_index_2049172] ^ p5_array_index_2049173;
  assign p6_array_index_2049352_comb = p5_literal_2043914[p5_res7__708];
  assign p6_array_index_2049353_comb = p5_literal_2043916[p5_res7__706];
  assign p6_array_index_2049354_comb = p5_literal_2043918[p5_res7__704];
  assign p6_array_index_2049355_comb = p5_literal_2043920[p5_array_index_2049162];
  assign p6_res7__714_comb = p5_literal_2043910[p6_res7__712_comb] ^ p5_literal_2043912[p6_res7__710_comb] ^ p6_array_index_2049352_comb ^ p6_array_index_2049353_comb ^ p6_array_index_2049354_comb ^ p6_array_index_2049355_comb ^ p5_array_index_2049163 ^ p5_literal_2043923[p5_array_index_2049164] ^ p5_array_index_2049165 ^ p5_array_index_2049200 ^ p5_literal_2043918[p5_array_index_2049167] ^ p5_literal_2043916[p5_array_index_2049184] ^ p5_literal_2043914[p5_array_index_2049169] ^ p5_literal_2043912[p5_array_index_2049186] ^ p5_literal_2043910[p5_array_index_2049171] ^ p5_array_index_2049172;
  assign p6_array_index_2049366_comb = p5_literal_2043916[p5_res7__708];
  assign p6_array_index_2049367_comb = p5_literal_2043918[p5_res7__706];
  assign p6_array_index_2049368_comb = p5_literal_2043920[p5_res7__704];
  assign p6_res7__716_comb = p5_literal_2043910[p6_res7__714_comb] ^ p5_literal_2043912[p6_res7__712_comb] ^ p5_literal_2043914[p6_res7__710_comb] ^ p6_array_index_2049366_comb ^ p6_array_index_2049367_comb ^ p6_array_index_2049368_comb ^ p5_array_index_2049162 ^ p5_literal_2043923[p5_array_index_2049163] ^ p5_array_index_2049164 ^ p5_array_index_2049214 ^ p5_array_index_2049182 ^ p5_literal_2043916[p5_array_index_2049167] ^ p5_literal_2043914[p5_array_index_2049184] ^ p5_literal_2043912[p5_array_index_2049169] ^ p5_literal_2043910[p5_array_index_2049186] ^ p5_array_index_2049171;
  assign p6_array_index_2049378_comb = p5_literal_2043916[p6_res7__710_comb];
  assign p6_array_index_2049379_comb = p5_literal_2043918[p5_res7__708];
  assign p6_array_index_2049380_comb = p5_literal_2043920[p5_res7__706];
  assign p6_res7__718_comb = p5_literal_2043910[p6_res7__716_comb] ^ p5_literal_2043912[p6_res7__714_comb] ^ p5_literal_2043914[p6_res7__712_comb] ^ p6_array_index_2049378_comb ^ p6_array_index_2049379_comb ^ p6_array_index_2049380_comb ^ p5_res7__704 ^ p5_literal_2043923[p5_array_index_2049162] ^ p5_array_index_2049163 ^ p6_array_index_2049328_comb ^ p5_array_index_2049199 ^ p5_literal_2043916[p5_array_index_2049166] ^ p5_literal_2043914[p5_array_index_2049167] ^ p5_literal_2043912[p5_array_index_2049184] ^ p5_literal_2043910[p5_array_index_2049169] ^ p5_array_index_2049186;
  assign p6_array_index_2049391_comb = p5_literal_2043918[p6_res7__710_comb];
  assign p6_array_index_2049392_comb = p5_literal_2043920[p5_res7__708];
  assign p6_res7__720_comb = p5_literal_2043910[p6_res7__718_comb] ^ p5_literal_2043912[p6_res7__716_comb] ^ p5_literal_2043914[p6_res7__714_comb] ^ p5_literal_2043916[p6_res7__712_comb] ^ p6_array_index_2049391_comb ^ p6_array_index_2049392_comb ^ p5_res7__706 ^ p5_literal_2043923[p5_res7__704] ^ p5_array_index_2049162 ^ p6_array_index_2049342_comb ^ p5_array_index_2049213 ^ p5_array_index_2049181 ^ p5_literal_2043914[p5_array_index_2049166] ^ p5_literal_2043912[p5_array_index_2049167] ^ p5_literal_2043910[p5_array_index_2049184] ^ p5_array_index_2049169;
  assign p6_array_index_2049402_comb = p5_literal_2043918[p6_res7__712_comb];
  assign p6_array_index_2049403_comb = p5_literal_2043920[p6_res7__710_comb];
  assign p6_res7__722_comb = p5_literal_2043910[p6_res7__720_comb] ^ p5_literal_2043912[p6_res7__718_comb] ^ p5_literal_2043914[p6_res7__716_comb] ^ p5_literal_2043916[p6_res7__714_comb] ^ p6_array_index_2049402_comb ^ p6_array_index_2049403_comb ^ p5_res7__708 ^ p5_literal_2043923[p5_res7__706] ^ p5_res7__704 ^ p6_array_index_2049355_comb ^ p6_array_index_2049327_comb ^ p5_array_index_2049198 ^ p5_literal_2043914[p5_array_index_2049165] ^ p5_literal_2043912[p5_array_index_2049166] ^ p5_literal_2043910[p5_array_index_2049167] ^ p5_array_index_2049184;
  assign p6_array_index_2049414_comb = p5_literal_2043920[p6_res7__712_comb];
  assign p6_res7__724_comb = p5_literal_2043910[p6_res7__722_comb] ^ p5_literal_2043912[p6_res7__720_comb] ^ p5_literal_2043914[p6_res7__718_comb] ^ p5_literal_2043916[p6_res7__716_comb] ^ p5_literal_2043918[p6_res7__714_comb] ^ p6_array_index_2049414_comb ^ p6_res7__710_comb ^ p5_literal_2043923[p5_res7__708] ^ p5_res7__706 ^ p6_array_index_2049368_comb ^ p6_array_index_2049341_comb ^ p5_array_index_2049212 ^ p5_array_index_2049180 ^ p5_literal_2043912[p5_array_index_2049165] ^ p5_literal_2043910[p5_array_index_2049166] ^ p5_array_index_2049167;
  assign p6_array_index_2049424_comb = p5_literal_2043920[p6_res7__714_comb];
  assign p6_res7__726_comb = p5_literal_2043910[p6_res7__724_comb] ^ p5_literal_2043912[p6_res7__722_comb] ^ p5_literal_2043914[p6_res7__720_comb] ^ p5_literal_2043916[p6_res7__718_comb] ^ p5_literal_2043918[p6_res7__716_comb] ^ p6_array_index_2049424_comb ^ p6_res7__712_comb ^ p5_literal_2043923[p6_res7__710_comb] ^ p5_res7__708 ^ p6_array_index_2049380_comb ^ p6_array_index_2049354_comb ^ p6_array_index_2049326_comb ^ p5_array_index_2049197 ^ p5_literal_2043912[p5_array_index_2049164] ^ p5_literal_2043910[p5_array_index_2049165] ^ p5_array_index_2049166;
  assign p6_res7__728_comb = p5_literal_2043910[p6_res7__726_comb] ^ p5_literal_2043912[p6_res7__724_comb] ^ p5_literal_2043914[p6_res7__722_comb] ^ p5_literal_2043916[p6_res7__720_comb] ^ p5_literal_2043918[p6_res7__718_comb] ^ p5_literal_2043920[p6_res7__716_comb] ^ p6_res7__714_comb ^ p5_literal_2043923[p6_res7__712_comb] ^ p6_res7__710_comb ^ p6_array_index_2049392_comb ^ p6_array_index_2049367_comb ^ p6_array_index_2049340_comb ^ p5_array_index_2049211 ^ p5_array_index_2049179 ^ p5_literal_2043910[p5_array_index_2049164] ^ p5_array_index_2049165;
  assign p6_res7__730_comb = p5_literal_2043910[p6_res7__728_comb] ^ p5_literal_2043912[p6_res7__726_comb] ^ p5_literal_2043914[p6_res7__724_comb] ^ p5_literal_2043916[p6_res7__722_comb] ^ p5_literal_2043918[p6_res7__720_comb] ^ p5_literal_2043920[p6_res7__718_comb] ^ p6_res7__716_comb ^ p5_literal_2043923[p6_res7__714_comb] ^ p6_res7__712_comb ^ p6_array_index_2049403_comb ^ p6_array_index_2049379_comb ^ p6_array_index_2049353_comb ^ p6_array_index_2049325_comb ^ p5_array_index_2049196 ^ p5_literal_2043910[p5_array_index_2049163] ^ p5_array_index_2049164;
  assign p6_res7__732_comb = p5_literal_2043910[p6_res7__730_comb] ^ p5_literal_2043912[p6_res7__728_comb] ^ p5_literal_2043914[p6_res7__726_comb] ^ p5_literal_2043916[p6_res7__724_comb] ^ p5_literal_2043918[p6_res7__722_comb] ^ p5_literal_2043920[p6_res7__720_comb] ^ p6_res7__718_comb ^ p5_literal_2043923[p6_res7__716_comb] ^ p6_res7__714_comb ^ p6_array_index_2049414_comb ^ p6_array_index_2049391_comb ^ p6_array_index_2049366_comb ^ p6_array_index_2049339_comb ^ p5_array_index_2049210 ^ p5_array_index_2049178 ^ p5_array_index_2049163;
  assign p6_res7__734_comb = p5_literal_2043910[p6_res7__732_comb] ^ p5_literal_2043912[p6_res7__730_comb] ^ p5_literal_2043914[p6_res7__728_comb] ^ p5_literal_2043916[p6_res7__726_comb] ^ p5_literal_2043918[p6_res7__724_comb] ^ p5_literal_2043920[p6_res7__722_comb] ^ p6_res7__720_comb ^ p5_literal_2043923[p6_res7__718_comb] ^ p6_res7__716_comb ^ p6_array_index_2049424_comb ^ p6_array_index_2049402_comb ^ p6_array_index_2049378_comb ^ p6_array_index_2049352_comb ^ p6_array_index_2049324_comb ^ p5_array_index_2049195 ^ p5_array_index_2049162;
  assign p6_res__22_comb = {p6_res7__734_comb, p6_res7__732_comb, p6_res7__730_comb, p6_res7__728_comb, p6_res7__726_comb, p6_res7__724_comb, p6_res7__722_comb, p6_res7__720_comb, p6_res7__718_comb, p6_res7__716_comb, p6_res7__714_comb, p6_res7__712_comb, p6_res7__710_comb, p5_res7__708, p5_res7__706, p5_res7__704};
  assign p6_k7_comb = p6_res__22_comb ^ p5_xor_2048928;
  assign p6_addedKey__55_comb = p6_k7_comb ^ 128'hd9eb_5a3a_e90f_fa58_34ce_2043_693d_7e18;
  assign p6_array_index_2049480_comb = p5_literal_2043896[p6_addedKey__55_comb[127:120]];
  assign p6_array_index_2049481_comb = p5_literal_2043896[p6_addedKey__55_comb[119:112]];
  assign p6_array_index_2049482_comb = p5_literal_2043896[p6_addedKey__55_comb[111:104]];
  assign p6_array_index_2049483_comb = p5_literal_2043896[p6_addedKey__55_comb[103:96]];
  assign p6_array_index_2049484_comb = p5_literal_2043896[p6_addedKey__55_comb[95:88]];
  assign p6_array_index_2049485_comb = p5_literal_2043896[p6_addedKey__55_comb[87:80]];
  assign p6_array_index_2049487_comb = p5_literal_2043896[p6_addedKey__55_comb[71:64]];
  assign p6_array_index_2049489_comb = p5_literal_2043896[p6_addedKey__55_comb[55:48]];
  assign p6_array_index_2049490_comb = p5_literal_2043896[p6_addedKey__55_comb[47:40]];
  assign p6_array_index_2049491_comb = p5_literal_2043896[p6_addedKey__55_comb[39:32]];
  assign p6_array_index_2049492_comb = p5_literal_2043896[p6_addedKey__55_comb[31:24]];
  assign p6_array_index_2049493_comb = p5_literal_2043896[p6_addedKey__55_comb[23:16]];
  assign p6_array_index_2049494_comb = p5_literal_2043896[p6_addedKey__55_comb[15:8]];
  assign p6_array_index_2049496_comb = p5_literal_2043910[p6_array_index_2049480_comb];
  assign p6_array_index_2049497_comb = p5_literal_2043912[p6_array_index_2049481_comb];
  assign p6_array_index_2049498_comb = p5_literal_2043914[p6_array_index_2049482_comb];
  assign p6_array_index_2049499_comb = p5_literal_2043916[p6_array_index_2049483_comb];
  assign p6_array_index_2049500_comb = p5_literal_2043918[p6_array_index_2049484_comb];
  assign p6_array_index_2049501_comb = p5_literal_2043920[p6_array_index_2049485_comb];
  assign p6_array_index_2049502_comb = p5_literal_2043896[p6_addedKey__55_comb[79:72]];
  assign p6_array_index_2049504_comb = p5_literal_2043896[p6_addedKey__55_comb[63:56]];
  assign p6_res7__736_comb = p6_array_index_2049496_comb ^ p6_array_index_2049497_comb ^ p6_array_index_2049498_comb ^ p6_array_index_2049499_comb ^ p6_array_index_2049500_comb ^ p6_array_index_2049501_comb ^ p6_array_index_2049502_comb ^ p5_literal_2043923[p6_array_index_2049487_comb] ^ p6_array_index_2049504_comb ^ p5_literal_2043920[p6_array_index_2049489_comb] ^ p5_literal_2043918[p6_array_index_2049490_comb] ^ p5_literal_2043916[p6_array_index_2049491_comb] ^ p5_literal_2043914[p6_array_index_2049492_comb] ^ p5_literal_2043912[p6_array_index_2049493_comb] ^ p5_literal_2043910[p6_array_index_2049494_comb] ^ p5_literal_2043896[p6_addedKey__55_comb[7:0]];
  assign p6_array_index_2049513_comb = p5_literal_2043910[p6_res7__736_comb];
  assign p6_array_index_2049514_comb = p5_literal_2043912[p6_array_index_2049480_comb];
  assign p6_array_index_2049515_comb = p5_literal_2043914[p6_array_index_2049481_comb];
  assign p6_array_index_2049516_comb = p5_literal_2043916[p6_array_index_2049482_comb];
  assign p6_array_index_2049517_comb = p5_literal_2043918[p6_array_index_2049483_comb];
  assign p6_array_index_2049518_comb = p5_literal_2043920[p6_array_index_2049484_comb];
  assign p6_res7__738_comb = p6_array_index_2049513_comb ^ p6_array_index_2049514_comb ^ p6_array_index_2049515_comb ^ p6_array_index_2049516_comb ^ p6_array_index_2049517_comb ^ p6_array_index_2049518_comb ^ p6_array_index_2049485_comb ^ p5_literal_2043923[p6_array_index_2049502_comb] ^ p6_array_index_2049487_comb ^ p5_literal_2043920[p6_array_index_2049504_comb] ^ p5_literal_2043918[p6_array_index_2049489_comb] ^ p5_literal_2043916[p6_array_index_2049490_comb] ^ p5_literal_2043914[p6_array_index_2049491_comb] ^ p5_literal_2043912[p6_array_index_2049492_comb] ^ p5_literal_2043910[p6_array_index_2049493_comb] ^ p6_array_index_2049494_comb;
  assign p6_array_index_2049528_comb = p5_literal_2043912[p6_res7__736_comb];
  assign p6_array_index_2049529_comb = p5_literal_2043914[p6_array_index_2049480_comb];
  assign p6_array_index_2049530_comb = p5_literal_2043916[p6_array_index_2049481_comb];
  assign p6_array_index_2049531_comb = p5_literal_2043918[p6_array_index_2049482_comb];
  assign p6_array_index_2049532_comb = p5_literal_2043920[p6_array_index_2049483_comb];
  assign p6_res7__740_comb = p5_literal_2043910[p6_res7__738_comb] ^ p6_array_index_2049528_comb ^ p6_array_index_2049529_comb ^ p6_array_index_2049530_comb ^ p6_array_index_2049531_comb ^ p6_array_index_2049532_comb ^ p6_array_index_2049484_comb ^ p5_literal_2043923[p6_array_index_2049485_comb] ^ p6_array_index_2049502_comb ^ p5_literal_2043920[p6_array_index_2049487_comb] ^ p5_literal_2043918[p6_array_index_2049504_comb] ^ p5_literal_2043916[p6_array_index_2049489_comb] ^ p5_literal_2043914[p6_array_index_2049490_comb] ^ p5_literal_2043912[p6_array_index_2049491_comb] ^ p5_literal_2043910[p6_array_index_2049492_comb] ^ p6_array_index_2049493_comb;
  assign p6_array_index_2049542_comb = p5_literal_2043912[p6_res7__738_comb];
  assign p6_array_index_2049543_comb = p5_literal_2043914[p6_res7__736_comb];
  assign p6_array_index_2049544_comb = p5_literal_2043916[p6_array_index_2049480_comb];
  assign p6_array_index_2049545_comb = p5_literal_2043918[p6_array_index_2049481_comb];
  assign p6_array_index_2049546_comb = p5_literal_2043920[p6_array_index_2049482_comb];
  assign p6_res7__742_comb = p5_literal_2043910[p6_res7__740_comb] ^ p6_array_index_2049542_comb ^ p6_array_index_2049543_comb ^ p6_array_index_2049544_comb ^ p6_array_index_2049545_comb ^ p6_array_index_2049546_comb ^ p6_array_index_2049483_comb ^ p5_literal_2043923[p6_array_index_2049484_comb] ^ p6_array_index_2049485_comb ^ p5_literal_2043920[p6_array_index_2049502_comb] ^ p5_literal_2043918[p6_array_index_2049487_comb] ^ p5_literal_2043916[p6_array_index_2049504_comb] ^ p5_literal_2043914[p6_array_index_2049489_comb] ^ p5_literal_2043912[p6_array_index_2049490_comb] ^ p5_literal_2043910[p6_array_index_2049491_comb] ^ p6_array_index_2049492_comb;
  assign p6_array_index_2049557_comb = p5_literal_2043914[p6_res7__738_comb];
  assign p6_array_index_2049558_comb = p5_literal_2043916[p6_res7__736_comb];
  assign p6_array_index_2049559_comb = p5_literal_2043918[p6_array_index_2049480_comb];
  assign p6_array_index_2049560_comb = p5_literal_2043920[p6_array_index_2049481_comb];
  assign p6_res7__744_comb = p5_literal_2043910[p6_res7__742_comb] ^ p5_literal_2043912[p6_res7__740_comb] ^ p6_array_index_2049557_comb ^ p6_array_index_2049558_comb ^ p6_array_index_2049559_comb ^ p6_array_index_2049560_comb ^ p6_array_index_2049482_comb ^ p5_literal_2043923[p6_array_index_2049483_comb] ^ p6_array_index_2049484_comb ^ p6_array_index_2049501_comb ^ p5_literal_2043918[p6_array_index_2049502_comb] ^ p5_literal_2043916[p6_array_index_2049487_comb] ^ p5_literal_2043914[p6_array_index_2049504_comb] ^ p5_literal_2043912[p6_array_index_2049489_comb] ^ p5_literal_2043910[p6_array_index_2049490_comb] ^ p6_array_index_2049491_comb;
  assign p6_array_index_2049570_comb = p5_literal_2043914[p6_res7__740_comb];
  assign p6_array_index_2049571_comb = p5_literal_2043916[p6_res7__738_comb];
  assign p6_array_index_2049572_comb = p5_literal_2043918[p6_res7__736_comb];
  assign p6_array_index_2049573_comb = p5_literal_2043920[p6_array_index_2049480_comb];
  assign p6_res7__746_comb = p5_literal_2043910[p6_res7__744_comb] ^ p5_literal_2043912[p6_res7__742_comb] ^ p6_array_index_2049570_comb ^ p6_array_index_2049571_comb ^ p6_array_index_2049572_comb ^ p6_array_index_2049573_comb ^ p6_array_index_2049481_comb ^ p5_literal_2043923[p6_array_index_2049482_comb] ^ p6_array_index_2049483_comb ^ p6_array_index_2049518_comb ^ p5_literal_2043918[p6_array_index_2049485_comb] ^ p5_literal_2043916[p6_array_index_2049502_comb] ^ p5_literal_2043914[p6_array_index_2049487_comb] ^ p5_literal_2043912[p6_array_index_2049504_comb] ^ p5_literal_2043910[p6_array_index_2049489_comb] ^ p6_array_index_2049490_comb;
  assign p6_array_index_2049584_comb = p5_literal_2043916[p6_res7__740_comb];
  assign p6_array_index_2049585_comb = p5_literal_2043918[p6_res7__738_comb];
  assign p6_array_index_2049586_comb = p5_literal_2043920[p6_res7__736_comb];
  assign p6_res7__748_comb = p5_literal_2043910[p6_res7__746_comb] ^ p5_literal_2043912[p6_res7__744_comb] ^ p5_literal_2043914[p6_res7__742_comb] ^ p6_array_index_2049584_comb ^ p6_array_index_2049585_comb ^ p6_array_index_2049586_comb ^ p6_array_index_2049480_comb ^ p5_literal_2043923[p6_array_index_2049481_comb] ^ p6_array_index_2049482_comb ^ p6_array_index_2049532_comb ^ p6_array_index_2049500_comb ^ p5_literal_2043916[p6_array_index_2049485_comb] ^ p5_literal_2043914[p6_array_index_2049502_comb] ^ p5_literal_2043912[p6_array_index_2049487_comb] ^ p5_literal_2043910[p6_array_index_2049504_comb] ^ p6_array_index_2049489_comb;
  assign p6_array_index_2049596_comb = p5_literal_2043916[p6_res7__742_comb];
  assign p6_array_index_2049597_comb = p5_literal_2043918[p6_res7__740_comb];
  assign p6_array_index_2049598_comb = p5_literal_2043920[p6_res7__738_comb];
  assign p6_res7__750_comb = p5_literal_2043910[p6_res7__748_comb] ^ p5_literal_2043912[p6_res7__746_comb] ^ p5_literal_2043914[p6_res7__744_comb] ^ p6_array_index_2049596_comb ^ p6_array_index_2049597_comb ^ p6_array_index_2049598_comb ^ p6_res7__736_comb ^ p5_literal_2043923[p6_array_index_2049480_comb] ^ p6_array_index_2049481_comb ^ p6_array_index_2049546_comb ^ p6_array_index_2049517_comb ^ p5_literal_2043916[p6_array_index_2049484_comb] ^ p5_literal_2043914[p6_array_index_2049485_comb] ^ p5_literal_2043912[p6_array_index_2049502_comb] ^ p5_literal_2043910[p6_array_index_2049487_comb] ^ p6_array_index_2049504_comb;
  assign p6_array_index_2049609_comb = p5_literal_2043918[p6_res7__742_comb];
  assign p6_array_index_2049610_comb = p5_literal_2043920[p6_res7__740_comb];
  assign p6_res7__752_comb = p5_literal_2043910[p6_res7__750_comb] ^ p5_literal_2043912[p6_res7__748_comb] ^ p5_literal_2043914[p6_res7__746_comb] ^ p5_literal_2043916[p6_res7__744_comb] ^ p6_array_index_2049609_comb ^ p6_array_index_2049610_comb ^ p6_res7__738_comb ^ p5_literal_2043923[p6_res7__736_comb] ^ p6_array_index_2049480_comb ^ p6_array_index_2049560_comb ^ p6_array_index_2049531_comb ^ p6_array_index_2049499_comb ^ p5_literal_2043914[p6_array_index_2049484_comb] ^ p5_literal_2043912[p6_array_index_2049485_comb] ^ p5_literal_2043910[p6_array_index_2049502_comb] ^ p6_array_index_2049487_comb;
  assign p6_array_index_2049620_comb = p5_literal_2043918[p6_res7__744_comb];
  assign p6_array_index_2049621_comb = p5_literal_2043920[p6_res7__742_comb];
  assign p6_res7__754_comb = p5_literal_2043910[p6_res7__752_comb] ^ p5_literal_2043912[p6_res7__750_comb] ^ p5_literal_2043914[p6_res7__748_comb] ^ p5_literal_2043916[p6_res7__746_comb] ^ p6_array_index_2049620_comb ^ p6_array_index_2049621_comb ^ p6_res7__740_comb ^ p5_literal_2043923[p6_res7__738_comb] ^ p6_res7__736_comb ^ p6_array_index_2049573_comb ^ p6_array_index_2049545_comb ^ p6_array_index_2049516_comb ^ p5_literal_2043914[p6_array_index_2049483_comb] ^ p5_literal_2043912[p6_array_index_2049484_comb] ^ p5_literal_2043910[p6_array_index_2049485_comb] ^ p6_array_index_2049502_comb;
  assign p6_array_index_2049632_comb = p5_literal_2043920[p6_res7__744_comb];
  assign p6_res7__756_comb = p5_literal_2043910[p6_res7__754_comb] ^ p5_literal_2043912[p6_res7__752_comb] ^ p5_literal_2043914[p6_res7__750_comb] ^ p5_literal_2043916[p6_res7__748_comb] ^ p5_literal_2043918[p6_res7__746_comb] ^ p6_array_index_2049632_comb ^ p6_res7__742_comb ^ p5_literal_2043923[p6_res7__740_comb] ^ p6_res7__738_comb ^ p6_array_index_2049586_comb ^ p6_array_index_2049559_comb ^ p6_array_index_2049530_comb ^ p6_array_index_2049498_comb ^ p5_literal_2043912[p6_array_index_2049483_comb] ^ p5_literal_2043910[p6_array_index_2049484_comb] ^ p6_array_index_2049485_comb;
  assign p6_array_index_2049642_comb = p5_literal_2043920[p6_res7__746_comb];
  assign p6_res7__758_comb = p5_literal_2043910[p6_res7__756_comb] ^ p5_literal_2043912[p6_res7__754_comb] ^ p5_literal_2043914[p6_res7__752_comb] ^ p5_literal_2043916[p6_res7__750_comb] ^ p5_literal_2043918[p6_res7__748_comb] ^ p6_array_index_2049642_comb ^ p6_res7__744_comb ^ p5_literal_2043923[p6_res7__742_comb] ^ p6_res7__740_comb ^ p6_array_index_2049598_comb ^ p6_array_index_2049572_comb ^ p6_array_index_2049544_comb ^ p6_array_index_2049515_comb ^ p5_literal_2043912[p6_array_index_2049482_comb] ^ p5_literal_2043910[p6_array_index_2049483_comb] ^ p6_array_index_2049484_comb;
  assign p6_res7__760_comb = p5_literal_2043910[p6_res7__758_comb] ^ p5_literal_2043912[p6_res7__756_comb] ^ p5_literal_2043914[p6_res7__754_comb] ^ p5_literal_2043916[p6_res7__752_comb] ^ p5_literal_2043918[p6_res7__750_comb] ^ p5_literal_2043920[p6_res7__748_comb] ^ p6_res7__746_comb ^ p5_literal_2043923[p6_res7__744_comb] ^ p6_res7__742_comb ^ p6_array_index_2049610_comb ^ p6_array_index_2049585_comb ^ p6_array_index_2049558_comb ^ p6_array_index_2049529_comb ^ p6_array_index_2049497_comb ^ p5_literal_2043910[p6_array_index_2049482_comb] ^ p6_array_index_2049483_comb;
  assign p6_res7__762_comb = p5_literal_2043910[p6_res7__760_comb] ^ p5_literal_2043912[p6_res7__758_comb] ^ p5_literal_2043914[p6_res7__756_comb] ^ p5_literal_2043916[p6_res7__754_comb] ^ p5_literal_2043918[p6_res7__752_comb] ^ p5_literal_2043920[p6_res7__750_comb] ^ p6_res7__748_comb ^ p5_literal_2043923[p6_res7__746_comb] ^ p6_res7__744_comb ^ p6_array_index_2049621_comb ^ p6_array_index_2049597_comb ^ p6_array_index_2049571_comb ^ p6_array_index_2049543_comb ^ p6_array_index_2049514_comb ^ p5_literal_2043910[p6_array_index_2049481_comb] ^ p6_array_index_2049482_comb;
  assign p6_res7__764_comb = p5_literal_2043910[p6_res7__762_comb] ^ p5_literal_2043912[p6_res7__760_comb] ^ p5_literal_2043914[p6_res7__758_comb] ^ p5_literal_2043916[p6_res7__756_comb] ^ p5_literal_2043918[p6_res7__754_comb] ^ p5_literal_2043920[p6_res7__752_comb] ^ p6_res7__750_comb ^ p5_literal_2043923[p6_res7__748_comb] ^ p6_res7__746_comb ^ p6_array_index_2049632_comb ^ p6_array_index_2049609_comb ^ p6_array_index_2049584_comb ^ p6_array_index_2049557_comb ^ p6_array_index_2049528_comb ^ p6_array_index_2049496_comb ^ p6_array_index_2049481_comb;
  assign p6_res7__766_comb = p5_literal_2043910[p6_res7__764_comb] ^ p5_literal_2043912[p6_res7__762_comb] ^ p5_literal_2043914[p6_res7__760_comb] ^ p5_literal_2043916[p6_res7__758_comb] ^ p5_literal_2043918[p6_res7__756_comb] ^ p5_literal_2043920[p6_res7__754_comb] ^ p6_res7__752_comb ^ p5_literal_2043923[p6_res7__750_comb] ^ p6_res7__748_comb ^ p6_array_index_2049642_comb ^ p6_array_index_2049620_comb ^ p6_array_index_2049596_comb ^ p6_array_index_2049570_comb ^ p6_array_index_2049542_comb ^ p6_array_index_2049513_comb ^ p6_array_index_2049480_comb;
  assign p6_res__23_comb = {p6_res7__766_comb, p6_res7__764_comb, p6_res7__762_comb, p6_res7__760_comb, p6_res7__758_comb, p6_res7__756_comb, p6_res7__754_comb, p6_res7__752_comb, p6_res7__750_comb, p6_res7__748_comb, p6_res7__746_comb, p6_res7__744_comb, p6_res7__742_comb, p6_res7__740_comb, p6_res7__738_comb, p6_res7__736_comb};
  assign p6_k6_comb = p6_res__23_comb ^ p5_xor_2049146;
  assign p6_addedKey__56_comb = p6_k6_comb ^ 128'hb749_2c48_8547_80e0_69e9_9d53_b4b9_ea19;
  assign p6_array_index_2049698_comb = p5_literal_2043896[p6_addedKey__56_comb[127:120]];
  assign p6_array_index_2049699_comb = p5_literal_2043896[p6_addedKey__56_comb[119:112]];
  assign p6_array_index_2049700_comb = p5_literal_2043896[p6_addedKey__56_comb[111:104]];
  assign p6_array_index_2049701_comb = p5_literal_2043896[p6_addedKey__56_comb[103:96]];
  assign p6_array_index_2049702_comb = p5_literal_2043896[p6_addedKey__56_comb[95:88]];
  assign p6_array_index_2049703_comb = p5_literal_2043896[p6_addedKey__56_comb[87:80]];
  assign p6_array_index_2049705_comb = p5_literal_2043896[p6_addedKey__56_comb[71:64]];
  assign p6_array_index_2049707_comb = p5_literal_2043896[p6_addedKey__56_comb[55:48]];
  assign p6_array_index_2049708_comb = p5_literal_2043896[p6_addedKey__56_comb[47:40]];
  assign p6_array_index_2049709_comb = p5_literal_2043896[p6_addedKey__56_comb[39:32]];
  assign p6_array_index_2049710_comb = p5_literal_2043896[p6_addedKey__56_comb[31:24]];
  assign p6_array_index_2049711_comb = p5_literal_2043896[p6_addedKey__56_comb[23:16]];
  assign p6_array_index_2049712_comb = p5_literal_2043896[p6_addedKey__56_comb[15:8]];
  assign p6_array_index_2049714_comb = p5_literal_2043910[p6_array_index_2049698_comb];
  assign p6_array_index_2049715_comb = p5_literal_2043912[p6_array_index_2049699_comb];
  assign p6_array_index_2049716_comb = p5_literal_2043914[p6_array_index_2049700_comb];
  assign p6_array_index_2049717_comb = p5_literal_2043916[p6_array_index_2049701_comb];
  assign p6_array_index_2049718_comb = p5_literal_2043918[p6_array_index_2049702_comb];
  assign p6_array_index_2049719_comb = p5_literal_2043920[p6_array_index_2049703_comb];
  assign p6_array_index_2049720_comb = p5_literal_2043896[p6_addedKey__56_comb[79:72]];
  assign p6_array_index_2049722_comb = p5_literal_2043896[p6_addedKey__56_comb[63:56]];
  assign p6_res7__768_comb = p6_array_index_2049714_comb ^ p6_array_index_2049715_comb ^ p6_array_index_2049716_comb ^ p6_array_index_2049717_comb ^ p6_array_index_2049718_comb ^ p6_array_index_2049719_comb ^ p6_array_index_2049720_comb ^ p5_literal_2043923[p6_array_index_2049705_comb] ^ p6_array_index_2049722_comb ^ p5_literal_2043920[p6_array_index_2049707_comb] ^ p5_literal_2043918[p6_array_index_2049708_comb] ^ p5_literal_2043916[p6_array_index_2049709_comb] ^ p5_literal_2043914[p6_array_index_2049710_comb] ^ p5_literal_2043912[p6_array_index_2049711_comb] ^ p5_literal_2043910[p6_array_index_2049712_comb] ^ p5_literal_2043896[p6_addedKey__56_comb[7:0]];
  assign p6_array_index_2049731_comb = p5_literal_2043910[p6_res7__768_comb];
  assign p6_array_index_2049732_comb = p5_literal_2043912[p6_array_index_2049698_comb];
  assign p6_array_index_2049733_comb = p5_literal_2043914[p6_array_index_2049699_comb];
  assign p6_array_index_2049734_comb = p5_literal_2043916[p6_array_index_2049700_comb];
  assign p6_array_index_2049735_comb = p5_literal_2043918[p6_array_index_2049701_comb];
  assign p6_array_index_2049736_comb = p5_literal_2043920[p6_array_index_2049702_comb];
  assign p6_res7__770_comb = p6_array_index_2049731_comb ^ p6_array_index_2049732_comb ^ p6_array_index_2049733_comb ^ p6_array_index_2049734_comb ^ p6_array_index_2049735_comb ^ p6_array_index_2049736_comb ^ p6_array_index_2049703_comb ^ p5_literal_2043923[p6_array_index_2049720_comb] ^ p6_array_index_2049705_comb ^ p5_literal_2043920[p6_array_index_2049722_comb] ^ p5_literal_2043918[p6_array_index_2049707_comb] ^ p5_literal_2043916[p6_array_index_2049708_comb] ^ p5_literal_2043914[p6_array_index_2049709_comb] ^ p5_literal_2043912[p6_array_index_2049710_comb] ^ p5_literal_2043910[p6_array_index_2049711_comb] ^ p6_array_index_2049712_comb;
  assign p6_array_index_2049746_comb = p5_literal_2043912[p6_res7__768_comb];
  assign p6_array_index_2049747_comb = p5_literal_2043914[p6_array_index_2049698_comb];
  assign p6_array_index_2049748_comb = p5_literal_2043916[p6_array_index_2049699_comb];
  assign p6_array_index_2049749_comb = p5_literal_2043918[p6_array_index_2049700_comb];
  assign p6_array_index_2049750_comb = p5_literal_2043920[p6_array_index_2049701_comb];
  assign p6_res7__772_comb = p5_literal_2043910[p6_res7__770_comb] ^ p6_array_index_2049746_comb ^ p6_array_index_2049747_comb ^ p6_array_index_2049748_comb ^ p6_array_index_2049749_comb ^ p6_array_index_2049750_comb ^ p6_array_index_2049702_comb ^ p5_literal_2043923[p6_array_index_2049703_comb] ^ p6_array_index_2049720_comb ^ p5_literal_2043920[p6_array_index_2049705_comb] ^ p5_literal_2043918[p6_array_index_2049722_comb] ^ p5_literal_2043916[p6_array_index_2049707_comb] ^ p5_literal_2043914[p6_array_index_2049708_comb] ^ p5_literal_2043912[p6_array_index_2049709_comb] ^ p5_literal_2043910[p6_array_index_2049710_comb] ^ p6_array_index_2049711_comb;
  assign p6_array_index_2049760_comb = p5_literal_2043912[p6_res7__770_comb];
  assign p6_array_index_2049761_comb = p5_literal_2043914[p6_res7__768_comb];
  assign p6_array_index_2049762_comb = p5_literal_2043916[p6_array_index_2049698_comb];
  assign p6_array_index_2049763_comb = p5_literal_2043918[p6_array_index_2049699_comb];
  assign p6_array_index_2049764_comb = p5_literal_2043920[p6_array_index_2049700_comb];
  assign p6_res7__774_comb = p5_literal_2043910[p6_res7__772_comb] ^ p6_array_index_2049760_comb ^ p6_array_index_2049761_comb ^ p6_array_index_2049762_comb ^ p6_array_index_2049763_comb ^ p6_array_index_2049764_comb ^ p6_array_index_2049701_comb ^ p5_literal_2043923[p6_array_index_2049702_comb] ^ p6_array_index_2049703_comb ^ p5_literal_2043920[p6_array_index_2049720_comb] ^ p5_literal_2043918[p6_array_index_2049705_comb] ^ p5_literal_2043916[p6_array_index_2049722_comb] ^ p5_literal_2043914[p6_array_index_2049707_comb] ^ p5_literal_2043912[p6_array_index_2049708_comb] ^ p5_literal_2043910[p6_array_index_2049709_comb] ^ p6_array_index_2049710_comb;
  assign p6_array_index_2049775_comb = p5_literal_2043914[p6_res7__770_comb];
  assign p6_array_index_2049776_comb = p5_literal_2043916[p6_res7__768_comb];
  assign p6_array_index_2049777_comb = p5_literal_2043918[p6_array_index_2049698_comb];
  assign p6_array_index_2049778_comb = p5_literal_2043920[p6_array_index_2049699_comb];
  assign p6_res7__776_comb = p5_literal_2043910[p6_res7__774_comb] ^ p5_literal_2043912[p6_res7__772_comb] ^ p6_array_index_2049775_comb ^ p6_array_index_2049776_comb ^ p6_array_index_2049777_comb ^ p6_array_index_2049778_comb ^ p6_array_index_2049700_comb ^ p5_literal_2043923[p6_array_index_2049701_comb] ^ p6_array_index_2049702_comb ^ p6_array_index_2049719_comb ^ p5_literal_2043918[p6_array_index_2049720_comb] ^ p5_literal_2043916[p6_array_index_2049705_comb] ^ p5_literal_2043914[p6_array_index_2049722_comb] ^ p5_literal_2043912[p6_array_index_2049707_comb] ^ p5_literal_2043910[p6_array_index_2049708_comb] ^ p6_array_index_2049709_comb;
  assign p6_array_index_2049788_comb = p5_literal_2043914[p6_res7__772_comb];
  assign p6_array_index_2049789_comb = p5_literal_2043916[p6_res7__770_comb];
  assign p6_array_index_2049790_comb = p5_literal_2043918[p6_res7__768_comb];
  assign p6_array_index_2049791_comb = p5_literal_2043920[p6_array_index_2049698_comb];
  assign p6_res7__778_comb = p5_literal_2043910[p6_res7__776_comb] ^ p5_literal_2043912[p6_res7__774_comb] ^ p6_array_index_2049788_comb ^ p6_array_index_2049789_comb ^ p6_array_index_2049790_comb ^ p6_array_index_2049791_comb ^ p6_array_index_2049699_comb ^ p5_literal_2043923[p6_array_index_2049700_comb] ^ p6_array_index_2049701_comb ^ p6_array_index_2049736_comb ^ p5_literal_2043918[p6_array_index_2049703_comb] ^ p5_literal_2043916[p6_array_index_2049720_comb] ^ p5_literal_2043914[p6_array_index_2049705_comb] ^ p5_literal_2043912[p6_array_index_2049722_comb] ^ p5_literal_2043910[p6_array_index_2049707_comb] ^ p6_array_index_2049708_comb;
  assign p6_array_index_2049802_comb = p5_literal_2043916[p6_res7__772_comb];
  assign p6_array_index_2049803_comb = p5_literal_2043918[p6_res7__770_comb];
  assign p6_array_index_2049804_comb = p5_literal_2043920[p6_res7__768_comb];
  assign p6_res7__780_comb = p5_literal_2043910[p6_res7__778_comb] ^ p5_literal_2043912[p6_res7__776_comb] ^ p5_literal_2043914[p6_res7__774_comb] ^ p6_array_index_2049802_comb ^ p6_array_index_2049803_comb ^ p6_array_index_2049804_comb ^ p6_array_index_2049698_comb ^ p5_literal_2043923[p6_array_index_2049699_comb] ^ p6_array_index_2049700_comb ^ p6_array_index_2049750_comb ^ p6_array_index_2049718_comb ^ p5_literal_2043916[p6_array_index_2049703_comb] ^ p5_literal_2043914[p6_array_index_2049720_comb] ^ p5_literal_2043912[p6_array_index_2049705_comb] ^ p5_literal_2043910[p6_array_index_2049722_comb] ^ p6_array_index_2049707_comb;
  assign p6_array_index_2049814_comb = p5_literal_2043916[p6_res7__774_comb];
  assign p6_array_index_2049815_comb = p5_literal_2043918[p6_res7__772_comb];
  assign p6_array_index_2049816_comb = p5_literal_2043920[p6_res7__770_comb];
  assign p6_res7__782_comb = p5_literal_2043910[p6_res7__780_comb] ^ p5_literal_2043912[p6_res7__778_comb] ^ p5_literal_2043914[p6_res7__776_comb] ^ p6_array_index_2049814_comb ^ p6_array_index_2049815_comb ^ p6_array_index_2049816_comb ^ p6_res7__768_comb ^ p5_literal_2043923[p6_array_index_2049698_comb] ^ p6_array_index_2049699_comb ^ p6_array_index_2049764_comb ^ p6_array_index_2049735_comb ^ p5_literal_2043916[p6_array_index_2049702_comb] ^ p5_literal_2043914[p6_array_index_2049703_comb] ^ p5_literal_2043912[p6_array_index_2049720_comb] ^ p5_literal_2043910[p6_array_index_2049705_comb] ^ p6_array_index_2049722_comb;
  assign p6_array_index_2049827_comb = p5_literal_2043918[p6_res7__774_comb];
  assign p6_array_index_2049828_comb = p5_literal_2043920[p6_res7__772_comb];
  assign p6_res7__784_comb = p5_literal_2043910[p6_res7__782_comb] ^ p5_literal_2043912[p6_res7__780_comb] ^ p5_literal_2043914[p6_res7__778_comb] ^ p5_literal_2043916[p6_res7__776_comb] ^ p6_array_index_2049827_comb ^ p6_array_index_2049828_comb ^ p6_res7__770_comb ^ p5_literal_2043923[p6_res7__768_comb] ^ p6_array_index_2049698_comb ^ p6_array_index_2049778_comb ^ p6_array_index_2049749_comb ^ p6_array_index_2049717_comb ^ p5_literal_2043914[p6_array_index_2049702_comb] ^ p5_literal_2043912[p6_array_index_2049703_comb] ^ p5_literal_2043910[p6_array_index_2049720_comb] ^ p6_array_index_2049705_comb;
  assign p6_array_index_2049838_comb = p5_literal_2043918[p6_res7__776_comb];
  assign p6_array_index_2049839_comb = p5_literal_2043920[p6_res7__774_comb];
  assign p6_res7__786_comb = p5_literal_2043910[p6_res7__784_comb] ^ p5_literal_2043912[p6_res7__782_comb] ^ p5_literal_2043914[p6_res7__780_comb] ^ p5_literal_2043916[p6_res7__778_comb] ^ p6_array_index_2049838_comb ^ p6_array_index_2049839_comb ^ p6_res7__772_comb ^ p5_literal_2043923[p6_res7__770_comb] ^ p6_res7__768_comb ^ p6_array_index_2049791_comb ^ p6_array_index_2049763_comb ^ p6_array_index_2049734_comb ^ p5_literal_2043914[p6_array_index_2049701_comb] ^ p5_literal_2043912[p6_array_index_2049702_comb] ^ p5_literal_2043910[p6_array_index_2049703_comb] ^ p6_array_index_2049720_comb;
  assign p6_array_index_2049850_comb = p5_literal_2043920[p6_res7__776_comb];
  assign p6_res7__788_comb = p5_literal_2043910[p6_res7__786_comb] ^ p5_literal_2043912[p6_res7__784_comb] ^ p5_literal_2043914[p6_res7__782_comb] ^ p5_literal_2043916[p6_res7__780_comb] ^ p5_literal_2043918[p6_res7__778_comb] ^ p6_array_index_2049850_comb ^ p6_res7__774_comb ^ p5_literal_2043923[p6_res7__772_comb] ^ p6_res7__770_comb ^ p6_array_index_2049804_comb ^ p6_array_index_2049777_comb ^ p6_array_index_2049748_comb ^ p6_array_index_2049716_comb ^ p5_literal_2043912[p6_array_index_2049701_comb] ^ p5_literal_2043910[p6_array_index_2049702_comb] ^ p6_array_index_2049703_comb;
  assign p6_array_index_2049860_comb = p5_literal_2043920[p6_res7__778_comb];
  assign p6_res7__790_comb = p5_literal_2043910[p6_res7__788_comb] ^ p5_literal_2043912[p6_res7__786_comb] ^ p5_literal_2043914[p6_res7__784_comb] ^ p5_literal_2043916[p6_res7__782_comb] ^ p5_literal_2043918[p6_res7__780_comb] ^ p6_array_index_2049860_comb ^ p6_res7__776_comb ^ p5_literal_2043923[p6_res7__774_comb] ^ p6_res7__772_comb ^ p6_array_index_2049816_comb ^ p6_array_index_2049790_comb ^ p6_array_index_2049762_comb ^ p6_array_index_2049733_comb ^ p5_literal_2043912[p6_array_index_2049700_comb] ^ p5_literal_2043910[p6_array_index_2049701_comb] ^ p6_array_index_2049702_comb;
  assign p6_res7__792_comb = p5_literal_2043910[p6_res7__790_comb] ^ p5_literal_2043912[p6_res7__788_comb] ^ p5_literal_2043914[p6_res7__786_comb] ^ p5_literal_2043916[p6_res7__784_comb] ^ p5_literal_2043918[p6_res7__782_comb] ^ p5_literal_2043920[p6_res7__780_comb] ^ p6_res7__778_comb ^ p5_literal_2043923[p6_res7__776_comb] ^ p6_res7__774_comb ^ p6_array_index_2049828_comb ^ p6_array_index_2049803_comb ^ p6_array_index_2049776_comb ^ p6_array_index_2049747_comb ^ p6_array_index_2049715_comb ^ p5_literal_2043910[p6_array_index_2049700_comb] ^ p6_array_index_2049701_comb;
  assign p6_res7__794_comb = p5_literal_2043910[p6_res7__792_comb] ^ p5_literal_2043912[p6_res7__790_comb] ^ p5_literal_2043914[p6_res7__788_comb] ^ p5_literal_2043916[p6_res7__786_comb] ^ p5_literal_2043918[p6_res7__784_comb] ^ p5_literal_2043920[p6_res7__782_comb] ^ p6_res7__780_comb ^ p5_literal_2043923[p6_res7__778_comb] ^ p6_res7__776_comb ^ p6_array_index_2049839_comb ^ p6_array_index_2049815_comb ^ p6_array_index_2049789_comb ^ p6_array_index_2049761_comb ^ p6_array_index_2049732_comb ^ p5_literal_2043910[p6_array_index_2049699_comb] ^ p6_array_index_2049700_comb;
  assign p6_res7__796_comb = p5_literal_2043910[p6_res7__794_comb] ^ p5_literal_2043912[p6_res7__792_comb] ^ p5_literal_2043914[p6_res7__790_comb] ^ p5_literal_2043916[p6_res7__788_comb] ^ p5_literal_2043918[p6_res7__786_comb] ^ p5_literal_2043920[p6_res7__784_comb] ^ p6_res7__782_comb ^ p5_literal_2043923[p6_res7__780_comb] ^ p6_res7__778_comb ^ p6_array_index_2049850_comb ^ p6_array_index_2049827_comb ^ p6_array_index_2049802_comb ^ p6_array_index_2049775_comb ^ p6_array_index_2049746_comb ^ p6_array_index_2049714_comb ^ p6_array_index_2049699_comb;
  assign p6_res7__798_comb = p5_literal_2043910[p6_res7__796_comb] ^ p5_literal_2043912[p6_res7__794_comb] ^ p5_literal_2043914[p6_res7__792_comb] ^ p5_literal_2043916[p6_res7__790_comb] ^ p5_literal_2043918[p6_res7__788_comb] ^ p5_literal_2043920[p6_res7__786_comb] ^ p6_res7__784_comb ^ p5_literal_2043923[p6_res7__782_comb] ^ p6_res7__780_comb ^ p6_array_index_2049860_comb ^ p6_array_index_2049838_comb ^ p6_array_index_2049814_comb ^ p6_array_index_2049788_comb ^ p6_array_index_2049760_comb ^ p6_array_index_2049731_comb ^ p6_array_index_2049698_comb;
  assign p6_res__24_comb = {p6_res7__798_comb, p6_res7__796_comb, p6_res7__794_comb, p6_res7__792_comb, p6_res7__790_comb, p6_res7__788_comb, p6_res7__786_comb, p6_res7__784_comb, p6_res7__782_comb, p6_res7__780_comb, p6_res7__778_comb, p6_res7__776_comb, p6_res7__774_comb, p6_res7__772_comb, p6_res7__770_comb, p6_res7__768_comb};
  assign p6_xor_2049900_comb = p6_res__24_comb ^ p6_k7_comb;
  assign p6_addedKey__57_comb = p6_xor_2049900_comb ^ 128'h056c_b6de_319f_0eeb_8e80_9963_10f6_951a;
  assign p6_array_index_2049916_comb = p5_literal_2043896[p6_addedKey__57_comb[127:120]];
  assign p6_array_index_2049917_comb = p5_literal_2043896[p6_addedKey__57_comb[119:112]];
  assign p6_array_index_2049918_comb = p5_literal_2043896[p6_addedKey__57_comb[111:104]];
  assign p6_array_index_2049919_comb = p5_literal_2043896[p6_addedKey__57_comb[103:96]];
  assign p6_array_index_2049920_comb = p5_literal_2043896[p6_addedKey__57_comb[95:88]];
  assign p6_array_index_2049921_comb = p5_literal_2043896[p6_addedKey__57_comb[87:80]];
  assign p6_array_index_2049923_comb = p5_literal_2043896[p6_addedKey__57_comb[71:64]];
  assign p6_array_index_2049925_comb = p5_literal_2043896[p6_addedKey__57_comb[55:48]];
  assign p6_array_index_2049926_comb = p5_literal_2043896[p6_addedKey__57_comb[47:40]];
  assign p6_array_index_2049927_comb = p5_literal_2043896[p6_addedKey__57_comb[39:32]];
  assign p6_array_index_2049928_comb = p5_literal_2043896[p6_addedKey__57_comb[31:24]];
  assign p6_array_index_2049929_comb = p5_literal_2043896[p6_addedKey__57_comb[23:16]];
  assign p6_array_index_2049930_comb = p5_literal_2043896[p6_addedKey__57_comb[15:8]];
  assign p6_array_index_2049932_comb = p5_literal_2043910[p6_array_index_2049916_comb];
  assign p6_array_index_2049933_comb = p5_literal_2043912[p6_array_index_2049917_comb];
  assign p6_array_index_2049934_comb = p5_literal_2043914[p6_array_index_2049918_comb];
  assign p6_array_index_2049935_comb = p5_literal_2043916[p6_array_index_2049919_comb];
  assign p6_array_index_2049936_comb = p5_literal_2043918[p6_array_index_2049920_comb];
  assign p6_array_index_2049937_comb = p5_literal_2043920[p6_array_index_2049921_comb];
  assign p6_array_index_2049938_comb = p5_literal_2043896[p6_addedKey__57_comb[79:72]];
  assign p6_array_index_2049940_comb = p5_literal_2043896[p6_addedKey__57_comb[63:56]];
  assign p6_res7__800_comb = p6_array_index_2049932_comb ^ p6_array_index_2049933_comb ^ p6_array_index_2049934_comb ^ p6_array_index_2049935_comb ^ p6_array_index_2049936_comb ^ p6_array_index_2049937_comb ^ p6_array_index_2049938_comb ^ p5_literal_2043923[p6_array_index_2049923_comb] ^ p6_array_index_2049940_comb ^ p5_literal_2043920[p6_array_index_2049925_comb] ^ p5_literal_2043918[p6_array_index_2049926_comb] ^ p5_literal_2043916[p6_array_index_2049927_comb] ^ p5_literal_2043914[p6_array_index_2049928_comb] ^ p5_literal_2043912[p6_array_index_2049929_comb] ^ p5_literal_2043910[p6_array_index_2049930_comb] ^ p5_literal_2043896[p6_addedKey__57_comb[7:0]];
  assign p6_array_index_2049949_comb = p5_literal_2043910[p6_res7__800_comb];
  assign p6_array_index_2049950_comb = p5_literal_2043912[p6_array_index_2049916_comb];
  assign p6_array_index_2049951_comb = p5_literal_2043914[p6_array_index_2049917_comb];
  assign p6_array_index_2049952_comb = p5_literal_2043916[p6_array_index_2049918_comb];
  assign p6_array_index_2049953_comb = p5_literal_2043918[p6_array_index_2049919_comb];
  assign p6_array_index_2049954_comb = p5_literal_2043920[p6_array_index_2049920_comb];
  assign p6_res7__802_comb = p6_array_index_2049949_comb ^ p6_array_index_2049950_comb ^ p6_array_index_2049951_comb ^ p6_array_index_2049952_comb ^ p6_array_index_2049953_comb ^ p6_array_index_2049954_comb ^ p6_array_index_2049921_comb ^ p5_literal_2043923[p6_array_index_2049938_comb] ^ p6_array_index_2049923_comb ^ p5_literal_2043920[p6_array_index_2049940_comb] ^ p5_literal_2043918[p6_array_index_2049925_comb] ^ p5_literal_2043916[p6_array_index_2049926_comb] ^ p5_literal_2043914[p6_array_index_2049927_comb] ^ p5_literal_2043912[p6_array_index_2049928_comb] ^ p5_literal_2043910[p6_array_index_2049929_comb] ^ p6_array_index_2049930_comb;
  assign p6_array_index_2049964_comb = p5_literal_2043912[p6_res7__800_comb];
  assign p6_array_index_2049965_comb = p5_literal_2043914[p6_array_index_2049916_comb];
  assign p6_array_index_2049966_comb = p5_literal_2043916[p6_array_index_2049917_comb];
  assign p6_array_index_2049967_comb = p5_literal_2043918[p6_array_index_2049918_comb];
  assign p6_array_index_2049968_comb = p5_literal_2043920[p6_array_index_2049919_comb];
  assign p6_res7__804_comb = p5_literal_2043910[p6_res7__802_comb] ^ p6_array_index_2049964_comb ^ p6_array_index_2049965_comb ^ p6_array_index_2049966_comb ^ p6_array_index_2049967_comb ^ p6_array_index_2049968_comb ^ p6_array_index_2049920_comb ^ p5_literal_2043923[p6_array_index_2049921_comb] ^ p6_array_index_2049938_comb ^ p5_literal_2043920[p6_array_index_2049923_comb] ^ p5_literal_2043918[p6_array_index_2049940_comb] ^ p5_literal_2043916[p6_array_index_2049925_comb] ^ p5_literal_2043914[p6_array_index_2049926_comb] ^ p5_literal_2043912[p6_array_index_2049927_comb] ^ p5_literal_2043910[p6_array_index_2049928_comb] ^ p6_array_index_2049929_comb;
  assign p6_array_index_2049978_comb = p5_literal_2043912[p6_res7__802_comb];
  assign p6_array_index_2049979_comb = p5_literal_2043914[p6_res7__800_comb];
  assign p6_array_index_2049980_comb = p5_literal_2043916[p6_array_index_2049916_comb];
  assign p6_array_index_2049981_comb = p5_literal_2043918[p6_array_index_2049917_comb];
  assign p6_array_index_2049982_comb = p5_literal_2043920[p6_array_index_2049918_comb];
  assign p6_res7__806_comb = p5_literal_2043910[p6_res7__804_comb] ^ p6_array_index_2049978_comb ^ p6_array_index_2049979_comb ^ p6_array_index_2049980_comb ^ p6_array_index_2049981_comb ^ p6_array_index_2049982_comb ^ p6_array_index_2049919_comb ^ p5_literal_2043923[p6_array_index_2049920_comb] ^ p6_array_index_2049921_comb ^ p5_literal_2043920[p6_array_index_2049938_comb] ^ p5_literal_2043918[p6_array_index_2049923_comb] ^ p5_literal_2043916[p6_array_index_2049940_comb] ^ p5_literal_2043914[p6_array_index_2049925_comb] ^ p5_literal_2043912[p6_array_index_2049926_comb] ^ p5_literal_2043910[p6_array_index_2049927_comb] ^ p6_array_index_2049928_comb;
  assign p6_array_index_2049993_comb = p5_literal_2043914[p6_res7__802_comb];
  assign p6_array_index_2049994_comb = p5_literal_2043916[p6_res7__800_comb];
  assign p6_array_index_2049995_comb = p5_literal_2043918[p6_array_index_2049916_comb];
  assign p6_array_index_2049996_comb = p5_literal_2043920[p6_array_index_2049917_comb];
  assign p6_res7__808_comb = p5_literal_2043910[p6_res7__806_comb] ^ p5_literal_2043912[p6_res7__804_comb] ^ p6_array_index_2049993_comb ^ p6_array_index_2049994_comb ^ p6_array_index_2049995_comb ^ p6_array_index_2049996_comb ^ p6_array_index_2049918_comb ^ p5_literal_2043923[p6_array_index_2049919_comb] ^ p6_array_index_2049920_comb ^ p6_array_index_2049937_comb ^ p5_literal_2043918[p6_array_index_2049938_comb] ^ p5_literal_2043916[p6_array_index_2049923_comb] ^ p5_literal_2043914[p6_array_index_2049940_comb] ^ p5_literal_2043912[p6_array_index_2049925_comb] ^ p5_literal_2043910[p6_array_index_2049926_comb] ^ p6_array_index_2049927_comb;
  assign p6_array_index_2050006_comb = p5_literal_2043914[p6_res7__804_comb];
  assign p6_array_index_2050007_comb = p5_literal_2043916[p6_res7__802_comb];
  assign p6_array_index_2050008_comb = p5_literal_2043918[p6_res7__800_comb];
  assign p6_array_index_2050009_comb = p5_literal_2043920[p6_array_index_2049916_comb];
  assign p6_res7__810_comb = p5_literal_2043910[p6_res7__808_comb] ^ p5_literal_2043912[p6_res7__806_comb] ^ p6_array_index_2050006_comb ^ p6_array_index_2050007_comb ^ p6_array_index_2050008_comb ^ p6_array_index_2050009_comb ^ p6_array_index_2049917_comb ^ p5_literal_2043923[p6_array_index_2049918_comb] ^ p6_array_index_2049919_comb ^ p6_array_index_2049954_comb ^ p5_literal_2043918[p6_array_index_2049921_comb] ^ p5_literal_2043916[p6_array_index_2049938_comb] ^ p5_literal_2043914[p6_array_index_2049923_comb] ^ p5_literal_2043912[p6_array_index_2049940_comb] ^ p5_literal_2043910[p6_array_index_2049925_comb] ^ p6_array_index_2049926_comb;
  assign p6_array_index_2050020_comb = p5_literal_2043916[p6_res7__804_comb];
  assign p6_array_index_2050021_comb = p5_literal_2043918[p6_res7__802_comb];
  assign p6_array_index_2050022_comb = p5_literal_2043920[p6_res7__800_comb];
  assign p6_res7__812_comb = p5_literal_2043910[p6_res7__810_comb] ^ p5_literal_2043912[p6_res7__808_comb] ^ p5_literal_2043914[p6_res7__806_comb] ^ p6_array_index_2050020_comb ^ p6_array_index_2050021_comb ^ p6_array_index_2050022_comb ^ p6_array_index_2049916_comb ^ p5_literal_2043923[p6_array_index_2049917_comb] ^ p6_array_index_2049918_comb ^ p6_array_index_2049968_comb ^ p6_array_index_2049936_comb ^ p5_literal_2043916[p6_array_index_2049921_comb] ^ p5_literal_2043914[p6_array_index_2049938_comb] ^ p5_literal_2043912[p6_array_index_2049923_comb] ^ p5_literal_2043910[p6_array_index_2049940_comb] ^ p6_array_index_2049925_comb;
  assign p6_array_index_2050032_comb = p5_literal_2043916[p6_res7__806_comb];
  assign p6_array_index_2050033_comb = p5_literal_2043918[p6_res7__804_comb];
  assign p6_array_index_2050034_comb = p5_literal_2043920[p6_res7__802_comb];
  assign p6_res7__814_comb = p5_literal_2043910[p6_res7__812_comb] ^ p5_literal_2043912[p6_res7__810_comb] ^ p5_literal_2043914[p6_res7__808_comb] ^ p6_array_index_2050032_comb ^ p6_array_index_2050033_comb ^ p6_array_index_2050034_comb ^ p6_res7__800_comb ^ p5_literal_2043923[p6_array_index_2049916_comb] ^ p6_array_index_2049917_comb ^ p6_array_index_2049982_comb ^ p6_array_index_2049953_comb ^ p5_literal_2043916[p6_array_index_2049920_comb] ^ p5_literal_2043914[p6_array_index_2049921_comb] ^ p5_literal_2043912[p6_array_index_2049938_comb] ^ p5_literal_2043910[p6_array_index_2049923_comb] ^ p6_array_index_2049940_comb;
  assign p6_array_index_2050045_comb = p5_literal_2043918[p6_res7__806_comb];
  assign p6_array_index_2050046_comb = p5_literal_2043920[p6_res7__804_comb];
  assign p6_res7__816_comb = p5_literal_2043910[p6_res7__814_comb] ^ p5_literal_2043912[p6_res7__812_comb] ^ p5_literal_2043914[p6_res7__810_comb] ^ p5_literal_2043916[p6_res7__808_comb] ^ p6_array_index_2050045_comb ^ p6_array_index_2050046_comb ^ p6_res7__802_comb ^ p5_literal_2043923[p6_res7__800_comb] ^ p6_array_index_2049916_comb ^ p6_array_index_2049996_comb ^ p6_array_index_2049967_comb ^ p6_array_index_2049935_comb ^ p5_literal_2043914[p6_array_index_2049920_comb] ^ p5_literal_2043912[p6_array_index_2049921_comb] ^ p5_literal_2043910[p6_array_index_2049938_comb] ^ p6_array_index_2049923_comb;
  assign p6_array_index_2050056_comb = p5_literal_2043918[p6_res7__808_comb];
  assign p6_array_index_2050057_comb = p5_literal_2043920[p6_res7__806_comb];
  assign p6_res7__818_comb = p5_literal_2043910[p6_res7__816_comb] ^ p5_literal_2043912[p6_res7__814_comb] ^ p5_literal_2043914[p6_res7__812_comb] ^ p5_literal_2043916[p6_res7__810_comb] ^ p6_array_index_2050056_comb ^ p6_array_index_2050057_comb ^ p6_res7__804_comb ^ p5_literal_2043923[p6_res7__802_comb] ^ p6_res7__800_comb ^ p6_array_index_2050009_comb ^ p6_array_index_2049981_comb ^ p6_array_index_2049952_comb ^ p5_literal_2043914[p6_array_index_2049919_comb] ^ p5_literal_2043912[p6_array_index_2049920_comb] ^ p5_literal_2043910[p6_array_index_2049921_comb] ^ p6_array_index_2049938_comb;
  assign p6_array_index_2050068_comb = p5_literal_2043920[p6_res7__808_comb];
  assign p6_res7__820_comb = p5_literal_2043910[p6_res7__818_comb] ^ p5_literal_2043912[p6_res7__816_comb] ^ p5_literal_2043914[p6_res7__814_comb] ^ p5_literal_2043916[p6_res7__812_comb] ^ p5_literal_2043918[p6_res7__810_comb] ^ p6_array_index_2050068_comb ^ p6_res7__806_comb ^ p5_literal_2043923[p6_res7__804_comb] ^ p6_res7__802_comb ^ p6_array_index_2050022_comb ^ p6_array_index_2049995_comb ^ p6_array_index_2049966_comb ^ p6_array_index_2049934_comb ^ p5_literal_2043912[p6_array_index_2049919_comb] ^ p5_literal_2043910[p6_array_index_2049920_comb] ^ p6_array_index_2049921_comb;
  assign p6_array_index_2050078_comb = p5_literal_2043920[p6_res7__810_comb];
  assign p6_res7__822_comb = p5_literal_2043910[p6_res7__820_comb] ^ p5_literal_2043912[p6_res7__818_comb] ^ p5_literal_2043914[p6_res7__816_comb] ^ p5_literal_2043916[p6_res7__814_comb] ^ p5_literal_2043918[p6_res7__812_comb] ^ p6_array_index_2050078_comb ^ p6_res7__808_comb ^ p5_literal_2043923[p6_res7__806_comb] ^ p6_res7__804_comb ^ p6_array_index_2050034_comb ^ p6_array_index_2050008_comb ^ p6_array_index_2049980_comb ^ p6_array_index_2049951_comb ^ p5_literal_2043912[p6_array_index_2049918_comb] ^ p5_literal_2043910[p6_array_index_2049919_comb] ^ p6_array_index_2049920_comb;
  assign p6_res7__824_comb = p5_literal_2043910[p6_res7__822_comb] ^ p5_literal_2043912[p6_res7__820_comb] ^ p5_literal_2043914[p6_res7__818_comb] ^ p5_literal_2043916[p6_res7__816_comb] ^ p5_literal_2043918[p6_res7__814_comb] ^ p5_literal_2043920[p6_res7__812_comb] ^ p6_res7__810_comb ^ p5_literal_2043923[p6_res7__808_comb] ^ p6_res7__806_comb ^ p6_array_index_2050046_comb ^ p6_array_index_2050021_comb ^ p6_array_index_2049994_comb ^ p6_array_index_2049965_comb ^ p6_array_index_2049933_comb ^ p5_literal_2043910[p6_array_index_2049918_comb] ^ p6_array_index_2049919_comb;
  assign p6_res7__826_comb = p5_literal_2043910[p6_res7__824_comb] ^ p5_literal_2043912[p6_res7__822_comb] ^ p5_literal_2043914[p6_res7__820_comb] ^ p5_literal_2043916[p6_res7__818_comb] ^ p5_literal_2043918[p6_res7__816_comb] ^ p5_literal_2043920[p6_res7__814_comb] ^ p6_res7__812_comb ^ p5_literal_2043923[p6_res7__810_comb] ^ p6_res7__808_comb ^ p6_array_index_2050057_comb ^ p6_array_index_2050033_comb ^ p6_array_index_2050007_comb ^ p6_array_index_2049979_comb ^ p6_array_index_2049950_comb ^ p5_literal_2043910[p6_array_index_2049917_comb] ^ p6_array_index_2049918_comb;
  assign p6_res7__828_comb = p5_literal_2043910[p6_res7__826_comb] ^ p5_literal_2043912[p6_res7__824_comb] ^ p5_literal_2043914[p6_res7__822_comb] ^ p5_literal_2043916[p6_res7__820_comb] ^ p5_literal_2043918[p6_res7__818_comb] ^ p5_literal_2043920[p6_res7__816_comb] ^ p6_res7__814_comb ^ p5_literal_2043923[p6_res7__812_comb] ^ p6_res7__810_comb ^ p6_array_index_2050068_comb ^ p6_array_index_2050045_comb ^ p6_array_index_2050020_comb ^ p6_array_index_2049993_comb ^ p6_array_index_2049964_comb ^ p6_array_index_2049932_comb ^ p6_array_index_2049917_comb;
  assign p6_res7__830_comb = p5_literal_2043910[p6_res7__828_comb] ^ p5_literal_2043912[p6_res7__826_comb] ^ p5_literal_2043914[p6_res7__824_comb] ^ p5_literal_2043916[p6_res7__822_comb] ^ p5_literal_2043918[p6_res7__820_comb] ^ p5_literal_2043920[p6_res7__818_comb] ^ p6_res7__816_comb ^ p5_literal_2043923[p6_res7__814_comb] ^ p6_res7__812_comb ^ p6_array_index_2050078_comb ^ p6_array_index_2050056_comb ^ p6_array_index_2050032_comb ^ p6_array_index_2050006_comb ^ p6_array_index_2049978_comb ^ p6_array_index_2049949_comb ^ p6_array_index_2049916_comb;
  assign p6_res__25_comb = {p6_res7__830_comb, p6_res7__828_comb, p6_res7__826_comb, p6_res7__824_comb, p6_res7__822_comb, p6_res7__820_comb, p6_res7__818_comb, p6_res7__816_comb, p6_res7__814_comb, p6_res7__812_comb, p6_res7__810_comb, p6_res7__808_comb, p6_res7__806_comb, p6_res7__804_comb, p6_res7__802_comb, p6_res7__800_comb};
  assign p6_xor_2050118_comb = p6_res__25_comb ^ p6_k6_comb;
  assign p6_addedKey__58_comb = p6_xor_2050118_comb ^ 128'h6bce_c0ac_5dd7_7453_d3a7_2473_cd72_011b;
  assign p6_array_index_2050134_comb = p5_literal_2043896[p6_addedKey__58_comb[127:120]];
  assign p6_array_index_2050135_comb = p5_literal_2043896[p6_addedKey__58_comb[119:112]];
  assign p6_array_index_2050136_comb = p5_literal_2043896[p6_addedKey__58_comb[111:104]];
  assign p6_array_index_2050137_comb = p5_literal_2043896[p6_addedKey__58_comb[103:96]];
  assign p6_array_index_2050138_comb = p5_literal_2043896[p6_addedKey__58_comb[95:88]];
  assign p6_array_index_2050139_comb = p5_literal_2043896[p6_addedKey__58_comb[87:80]];
  assign p6_array_index_2050141_comb = p5_literal_2043896[p6_addedKey__58_comb[71:64]];
  assign p6_array_index_2050143_comb = p5_literal_2043896[p6_addedKey__58_comb[55:48]];
  assign p6_array_index_2050144_comb = p5_literal_2043896[p6_addedKey__58_comb[47:40]];
  assign p6_array_index_2050145_comb = p5_literal_2043896[p6_addedKey__58_comb[39:32]];
  assign p6_array_index_2050146_comb = p5_literal_2043896[p6_addedKey__58_comb[31:24]];
  assign p6_array_index_2050147_comb = p5_literal_2043896[p6_addedKey__58_comb[23:16]];
  assign p6_array_index_2050148_comb = p5_literal_2043896[p6_addedKey__58_comb[15:8]];
  assign p6_array_index_2050150_comb = p5_literal_2043910[p6_array_index_2050134_comb];
  assign p6_array_index_2050151_comb = p5_literal_2043912[p6_array_index_2050135_comb];
  assign p6_array_index_2050152_comb = p5_literal_2043914[p6_array_index_2050136_comb];
  assign p6_array_index_2050153_comb = p5_literal_2043916[p6_array_index_2050137_comb];
  assign p6_array_index_2050154_comb = p5_literal_2043918[p6_array_index_2050138_comb];
  assign p6_array_index_2050155_comb = p5_literal_2043920[p6_array_index_2050139_comb];
  assign p6_array_index_2050156_comb = p5_literal_2043896[p6_addedKey__58_comb[79:72]];
  assign p6_array_index_2050158_comb = p5_literal_2043896[p6_addedKey__58_comb[63:56]];
  assign p6_res7__832_comb = p6_array_index_2050150_comb ^ p6_array_index_2050151_comb ^ p6_array_index_2050152_comb ^ p6_array_index_2050153_comb ^ p6_array_index_2050154_comb ^ p6_array_index_2050155_comb ^ p6_array_index_2050156_comb ^ p5_literal_2043923[p6_array_index_2050141_comb] ^ p6_array_index_2050158_comb ^ p5_literal_2043920[p6_array_index_2050143_comb] ^ p5_literal_2043918[p6_array_index_2050144_comb] ^ p5_literal_2043916[p6_array_index_2050145_comb] ^ p5_literal_2043914[p6_array_index_2050146_comb] ^ p5_literal_2043912[p6_array_index_2050147_comb] ^ p5_literal_2043910[p6_array_index_2050148_comb] ^ p5_literal_2043896[p6_addedKey__58_comb[7:0]];
  assign p6_array_index_2050167_comb = p5_literal_2043910[p6_res7__832_comb];
  assign p6_array_index_2050168_comb = p5_literal_2043912[p6_array_index_2050134_comb];
  assign p6_array_index_2050169_comb = p5_literal_2043914[p6_array_index_2050135_comb];
  assign p6_array_index_2050170_comb = p5_literal_2043916[p6_array_index_2050136_comb];
  assign p6_array_index_2050171_comb = p5_literal_2043918[p6_array_index_2050137_comb];
  assign p6_array_index_2050172_comb = p5_literal_2043920[p6_array_index_2050138_comb];
  assign p6_res7__834_comb = p6_array_index_2050167_comb ^ p6_array_index_2050168_comb ^ p6_array_index_2050169_comb ^ p6_array_index_2050170_comb ^ p6_array_index_2050171_comb ^ p6_array_index_2050172_comb ^ p6_array_index_2050139_comb ^ p5_literal_2043923[p6_array_index_2050156_comb] ^ p6_array_index_2050141_comb ^ p5_literal_2043920[p6_array_index_2050158_comb] ^ p5_literal_2043918[p6_array_index_2050143_comb] ^ p5_literal_2043916[p6_array_index_2050144_comb] ^ p5_literal_2043914[p6_array_index_2050145_comb] ^ p5_literal_2043912[p6_array_index_2050146_comb] ^ p5_literal_2043910[p6_array_index_2050147_comb] ^ p6_array_index_2050148_comb;
  assign p6_array_index_2050182_comb = p5_literal_2043912[p6_res7__832_comb];
  assign p6_array_index_2050183_comb = p5_literal_2043914[p6_array_index_2050134_comb];
  assign p6_array_index_2050184_comb = p5_literal_2043916[p6_array_index_2050135_comb];
  assign p6_array_index_2050185_comb = p5_literal_2043918[p6_array_index_2050136_comb];
  assign p6_array_index_2050186_comb = p5_literal_2043920[p6_array_index_2050137_comb];
  assign p6_res7__836_comb = p5_literal_2043910[p6_res7__834_comb] ^ p6_array_index_2050182_comb ^ p6_array_index_2050183_comb ^ p6_array_index_2050184_comb ^ p6_array_index_2050185_comb ^ p6_array_index_2050186_comb ^ p6_array_index_2050138_comb ^ p5_literal_2043923[p6_array_index_2050139_comb] ^ p6_array_index_2050156_comb ^ p5_literal_2043920[p6_array_index_2050141_comb] ^ p5_literal_2043918[p6_array_index_2050158_comb] ^ p5_literal_2043916[p6_array_index_2050143_comb] ^ p5_literal_2043914[p6_array_index_2050144_comb] ^ p5_literal_2043912[p6_array_index_2050145_comb] ^ p5_literal_2043910[p6_array_index_2050146_comb] ^ p6_array_index_2050147_comb;
  assign p6_array_index_2050196_comb = p5_literal_2043912[p6_res7__834_comb];
  assign p6_array_index_2050197_comb = p5_literal_2043914[p6_res7__832_comb];
  assign p6_array_index_2050198_comb = p5_literal_2043916[p6_array_index_2050134_comb];
  assign p6_array_index_2050199_comb = p5_literal_2043918[p6_array_index_2050135_comb];
  assign p6_array_index_2050200_comb = p5_literal_2043920[p6_array_index_2050136_comb];
  assign p6_res7__838_comb = p5_literal_2043910[p6_res7__836_comb] ^ p6_array_index_2050196_comb ^ p6_array_index_2050197_comb ^ p6_array_index_2050198_comb ^ p6_array_index_2050199_comb ^ p6_array_index_2050200_comb ^ p6_array_index_2050137_comb ^ p5_literal_2043923[p6_array_index_2050138_comb] ^ p6_array_index_2050139_comb ^ p5_literal_2043920[p6_array_index_2050156_comb] ^ p5_literal_2043918[p6_array_index_2050141_comb] ^ p5_literal_2043916[p6_array_index_2050158_comb] ^ p5_literal_2043914[p6_array_index_2050143_comb] ^ p5_literal_2043912[p6_array_index_2050144_comb] ^ p5_literal_2043910[p6_array_index_2050145_comb] ^ p6_array_index_2050146_comb;
  assign p6_array_index_2050211_comb = p5_literal_2043914[p6_res7__834_comb];
  assign p6_array_index_2050212_comb = p5_literal_2043916[p6_res7__832_comb];
  assign p6_array_index_2050213_comb = p5_literal_2043918[p6_array_index_2050134_comb];
  assign p6_array_index_2050214_comb = p5_literal_2043920[p6_array_index_2050135_comb];
  assign p6_res7__840_comb = p5_literal_2043910[p6_res7__838_comb] ^ p5_literal_2043912[p6_res7__836_comb] ^ p6_array_index_2050211_comb ^ p6_array_index_2050212_comb ^ p6_array_index_2050213_comb ^ p6_array_index_2050214_comb ^ p6_array_index_2050136_comb ^ p5_literal_2043923[p6_array_index_2050137_comb] ^ p6_array_index_2050138_comb ^ p6_array_index_2050155_comb ^ p5_literal_2043918[p6_array_index_2050156_comb] ^ p5_literal_2043916[p6_array_index_2050141_comb] ^ p5_literal_2043914[p6_array_index_2050158_comb] ^ p5_literal_2043912[p6_array_index_2050143_comb] ^ p5_literal_2043910[p6_array_index_2050144_comb] ^ p6_array_index_2050145_comb;
  assign p6_array_index_2050224_comb = p5_literal_2043914[p6_res7__836_comb];
  assign p6_array_index_2050225_comb = p5_literal_2043916[p6_res7__834_comb];
  assign p6_array_index_2050226_comb = p5_literal_2043918[p6_res7__832_comb];
  assign p6_array_index_2050227_comb = p5_literal_2043920[p6_array_index_2050134_comb];
  assign p6_res7__842_comb = p5_literal_2043910[p6_res7__840_comb] ^ p5_literal_2043912[p6_res7__838_comb] ^ p6_array_index_2050224_comb ^ p6_array_index_2050225_comb ^ p6_array_index_2050226_comb ^ p6_array_index_2050227_comb ^ p6_array_index_2050135_comb ^ p5_literal_2043923[p6_array_index_2050136_comb] ^ p6_array_index_2050137_comb ^ p6_array_index_2050172_comb ^ p5_literal_2043918[p6_array_index_2050139_comb] ^ p5_literal_2043916[p6_array_index_2050156_comb] ^ p5_literal_2043914[p6_array_index_2050141_comb] ^ p5_literal_2043912[p6_array_index_2050158_comb] ^ p5_literal_2043910[p6_array_index_2050143_comb] ^ p6_array_index_2050144_comb;
  assign p6_array_index_2050238_comb = p5_literal_2043916[p6_res7__836_comb];
  assign p6_array_index_2050239_comb = p5_literal_2043918[p6_res7__834_comb];
  assign p6_array_index_2050240_comb = p5_literal_2043920[p6_res7__832_comb];
  assign p6_res7__844_comb = p5_literal_2043910[p6_res7__842_comb] ^ p5_literal_2043912[p6_res7__840_comb] ^ p5_literal_2043914[p6_res7__838_comb] ^ p6_array_index_2050238_comb ^ p6_array_index_2050239_comb ^ p6_array_index_2050240_comb ^ p6_array_index_2050134_comb ^ p5_literal_2043923[p6_array_index_2050135_comb] ^ p6_array_index_2050136_comb ^ p6_array_index_2050186_comb ^ p6_array_index_2050154_comb ^ p5_literal_2043916[p6_array_index_2050139_comb] ^ p5_literal_2043914[p6_array_index_2050156_comb] ^ p5_literal_2043912[p6_array_index_2050141_comb] ^ p5_literal_2043910[p6_array_index_2050158_comb] ^ p6_array_index_2050143_comb;
  assign p6_array_index_2050250_comb = p5_literal_2043916[p6_res7__838_comb];
  assign p6_array_index_2050251_comb = p5_literal_2043918[p6_res7__836_comb];
  assign p6_array_index_2050252_comb = p5_literal_2043920[p6_res7__834_comb];
  assign p6_res7__846_comb = p5_literal_2043910[p6_res7__844_comb] ^ p5_literal_2043912[p6_res7__842_comb] ^ p5_literal_2043914[p6_res7__840_comb] ^ p6_array_index_2050250_comb ^ p6_array_index_2050251_comb ^ p6_array_index_2050252_comb ^ p6_res7__832_comb ^ p5_literal_2043923[p6_array_index_2050134_comb] ^ p6_array_index_2050135_comb ^ p6_array_index_2050200_comb ^ p6_array_index_2050171_comb ^ p5_literal_2043916[p6_array_index_2050138_comb] ^ p5_literal_2043914[p6_array_index_2050139_comb] ^ p5_literal_2043912[p6_array_index_2050156_comb] ^ p5_literal_2043910[p6_array_index_2050141_comb] ^ p6_array_index_2050158_comb;
  assign p6_array_index_2050263_comb = p5_literal_2043918[p6_res7__838_comb];
  assign p6_array_index_2050264_comb = p5_literal_2043920[p6_res7__836_comb];
  assign p6_res7__848_comb = p5_literal_2043910[p6_res7__846_comb] ^ p5_literal_2043912[p6_res7__844_comb] ^ p5_literal_2043914[p6_res7__842_comb] ^ p5_literal_2043916[p6_res7__840_comb] ^ p6_array_index_2050263_comb ^ p6_array_index_2050264_comb ^ p6_res7__834_comb ^ p5_literal_2043923[p6_res7__832_comb] ^ p6_array_index_2050134_comb ^ p6_array_index_2050214_comb ^ p6_array_index_2050185_comb ^ p6_array_index_2050153_comb ^ p5_literal_2043914[p6_array_index_2050138_comb] ^ p5_literal_2043912[p6_array_index_2050139_comb] ^ p5_literal_2043910[p6_array_index_2050156_comb] ^ p6_array_index_2050141_comb;
  assign p6_array_index_2050274_comb = p5_literal_2043918[p6_res7__840_comb];
  assign p6_array_index_2050275_comb = p5_literal_2043920[p6_res7__838_comb];
  assign p6_res7__850_comb = p5_literal_2043910[p6_res7__848_comb] ^ p5_literal_2043912[p6_res7__846_comb] ^ p5_literal_2043914[p6_res7__844_comb] ^ p5_literal_2043916[p6_res7__842_comb] ^ p6_array_index_2050274_comb ^ p6_array_index_2050275_comb ^ p6_res7__836_comb ^ p5_literal_2043923[p6_res7__834_comb] ^ p6_res7__832_comb ^ p6_array_index_2050227_comb ^ p6_array_index_2050199_comb ^ p6_array_index_2050170_comb ^ p5_literal_2043914[p6_array_index_2050137_comb] ^ p5_literal_2043912[p6_array_index_2050138_comb] ^ p5_literal_2043910[p6_array_index_2050139_comb] ^ p6_array_index_2050156_comb;
  assign p6_array_index_2050281_comb = p5_literal_2043910[p6_res7__850_comb];
  assign p6_array_index_2050282_comb = p5_literal_2043912[p6_res7__848_comb];
  assign p6_array_index_2050283_comb = p5_literal_2043914[p6_res7__846_comb];
  assign p6_array_index_2050284_comb = p5_literal_2043916[p6_res7__844_comb];
  assign p6_array_index_2050285_comb = p5_literal_2043918[p6_res7__842_comb];
  assign p6_array_index_2050286_comb = p5_literal_2043920[p6_res7__840_comb];
  assign p6_array_index_2050287_comb = p5_literal_2043923[p6_res7__836_comb];
  assign p6_array_index_2050288_comb = p5_literal_2043912[p6_array_index_2050137_comb];
  assign p6_array_index_2050289_comb = p5_literal_2043910[p6_array_index_2050138_comb];

  // Registers for pipe stage 6:
  reg [127:0] p6_encoded;
  reg [127:0] p6_bit_slice_2043893;
  reg [127:0] p6_bit_slice_2044119;
  reg [127:0] p6_k3;
  reg [127:0] p6_k2;
  reg [127:0] p6_k5;
  reg [127:0] p6_k4;
  reg [127:0] p6_k7;
  reg [127:0] p6_k6;
  reg [127:0] p6_xor_2049900;
  reg [127:0] p6_xor_2050118;
  reg [7:0] p6_array_index_2050134;
  reg [7:0] p6_array_index_2050135;
  reg [7:0] p6_array_index_2050136;
  reg [7:0] p6_array_index_2050137;
  reg [7:0] p6_array_index_2050138;
  reg [7:0] p6_array_index_2050139;
  reg [7:0] p6_array_index_2050150;
  reg [7:0] p6_array_index_2050151;
  reg [7:0] p6_array_index_2050152;
  reg [7:0] p6_res7__832;
  reg [7:0] p6_array_index_2050167;
  reg [7:0] p6_array_index_2050168;
  reg [7:0] p6_array_index_2050169;
  reg [7:0] p6_res7__834;
  reg [7:0] p6_array_index_2050182;
  reg [7:0] p6_array_index_2050183;
  reg [7:0] p6_array_index_2050184;
  reg [7:0] p6_res7__836;
  reg [7:0] p6_array_index_2050196;
  reg [7:0] p6_array_index_2050197;
  reg [7:0] p6_array_index_2050198;
  reg [7:0] p6_res7__838;
  reg [7:0] p6_array_index_2050211;
  reg [7:0] p6_array_index_2050212;
  reg [7:0] p6_array_index_2050213;
  reg [7:0] p6_res7__840;
  reg [7:0] p6_array_index_2050224;
  reg [7:0] p6_array_index_2050225;
  reg [7:0] p6_array_index_2050226;
  reg [7:0] p6_res7__842;
  reg [7:0] p6_array_index_2050238;
  reg [7:0] p6_array_index_2050239;
  reg [7:0] p6_array_index_2050240;
  reg [7:0] p6_res7__844;
  reg [7:0] p6_array_index_2050250;
  reg [7:0] p6_array_index_2050251;
  reg [7:0] p6_array_index_2050252;
  reg [7:0] p6_res7__846;
  reg [7:0] p6_array_index_2050263;
  reg [7:0] p6_array_index_2050264;
  reg [7:0] p6_res7__848;
  reg [7:0] p6_array_index_2050274;
  reg [7:0] p6_array_index_2050275;
  reg [7:0] p6_res7__850;
  reg [7:0] p6_array_index_2050281;
  reg [7:0] p6_array_index_2050282;
  reg [7:0] p6_array_index_2050283;
  reg [7:0] p6_array_index_2050284;
  reg [7:0] p6_array_index_2050285;
  reg [7:0] p6_array_index_2050286;
  reg [7:0] p6_array_index_2050287;
  reg [7:0] p6_array_index_2050288;
  reg [7:0] p6_array_index_2050289;
  reg [7:0] p7_literal_2043910[256];
  reg [7:0] p7_literal_2043912[256];
  reg [7:0] p7_literal_2043914[256];
  reg [7:0] p7_literal_2043916[256];
  reg [7:0] p7_literal_2043918[256];
  reg [7:0] p7_literal_2043920[256];
  reg [7:0] p7_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p6_encoded <= p5_encoded;
    p6_bit_slice_2043893 <= p5_bit_slice_2043893;
    p6_bit_slice_2044119 <= p5_bit_slice_2044119;
    p6_k3 <= p5_k3;
    p6_k2 <= p5_k2;
    p6_k5 <= p5_k5;
    p6_k4 <= p5_k4;
    p6_k7 <= p6_k7_comb;
    p6_k6 <= p6_k6_comb;
    p6_xor_2049900 <= p6_xor_2049900_comb;
    p6_xor_2050118 <= p6_xor_2050118_comb;
    p6_array_index_2050134 <= p6_array_index_2050134_comb;
    p6_array_index_2050135 <= p6_array_index_2050135_comb;
    p6_array_index_2050136 <= p6_array_index_2050136_comb;
    p6_array_index_2050137 <= p6_array_index_2050137_comb;
    p6_array_index_2050138 <= p6_array_index_2050138_comb;
    p6_array_index_2050139 <= p6_array_index_2050139_comb;
    p6_array_index_2050150 <= p6_array_index_2050150_comb;
    p6_array_index_2050151 <= p6_array_index_2050151_comb;
    p6_array_index_2050152 <= p6_array_index_2050152_comb;
    p6_res7__832 <= p6_res7__832_comb;
    p6_array_index_2050167 <= p6_array_index_2050167_comb;
    p6_array_index_2050168 <= p6_array_index_2050168_comb;
    p6_array_index_2050169 <= p6_array_index_2050169_comb;
    p6_res7__834 <= p6_res7__834_comb;
    p6_array_index_2050182 <= p6_array_index_2050182_comb;
    p6_array_index_2050183 <= p6_array_index_2050183_comb;
    p6_array_index_2050184 <= p6_array_index_2050184_comb;
    p6_res7__836 <= p6_res7__836_comb;
    p6_array_index_2050196 <= p6_array_index_2050196_comb;
    p6_array_index_2050197 <= p6_array_index_2050197_comb;
    p6_array_index_2050198 <= p6_array_index_2050198_comb;
    p6_res7__838 <= p6_res7__838_comb;
    p6_array_index_2050211 <= p6_array_index_2050211_comb;
    p6_array_index_2050212 <= p6_array_index_2050212_comb;
    p6_array_index_2050213 <= p6_array_index_2050213_comb;
    p6_res7__840 <= p6_res7__840_comb;
    p6_array_index_2050224 <= p6_array_index_2050224_comb;
    p6_array_index_2050225 <= p6_array_index_2050225_comb;
    p6_array_index_2050226 <= p6_array_index_2050226_comb;
    p6_res7__842 <= p6_res7__842_comb;
    p6_array_index_2050238 <= p6_array_index_2050238_comb;
    p6_array_index_2050239 <= p6_array_index_2050239_comb;
    p6_array_index_2050240 <= p6_array_index_2050240_comb;
    p6_res7__844 <= p6_res7__844_comb;
    p6_array_index_2050250 <= p6_array_index_2050250_comb;
    p6_array_index_2050251 <= p6_array_index_2050251_comb;
    p6_array_index_2050252 <= p6_array_index_2050252_comb;
    p6_res7__846 <= p6_res7__846_comb;
    p6_array_index_2050263 <= p6_array_index_2050263_comb;
    p6_array_index_2050264 <= p6_array_index_2050264_comb;
    p6_res7__848 <= p6_res7__848_comb;
    p6_array_index_2050274 <= p6_array_index_2050274_comb;
    p6_array_index_2050275 <= p6_array_index_2050275_comb;
    p6_res7__850 <= p6_res7__850_comb;
    p6_array_index_2050281 <= p6_array_index_2050281_comb;
    p6_array_index_2050282 <= p6_array_index_2050282_comb;
    p6_array_index_2050283 <= p6_array_index_2050283_comb;
    p6_array_index_2050284 <= p6_array_index_2050284_comb;
    p6_array_index_2050285 <= p6_array_index_2050285_comb;
    p6_array_index_2050286 <= p6_array_index_2050286_comb;
    p6_array_index_2050287 <= p6_array_index_2050287_comb;
    p6_array_index_2050288 <= p6_array_index_2050288_comb;
    p6_array_index_2050289 <= p6_array_index_2050289_comb;
    p7_literal_2043910 <= p6_literal_2043910;
    p7_literal_2043912 <= p6_literal_2043912;
    p7_literal_2043914 <= p6_literal_2043914;
    p7_literal_2043916 <= p6_literal_2043916;
    p7_literal_2043918 <= p6_literal_2043918;
    p7_literal_2043920 <= p6_literal_2043920;
    p7_literal_2043923 <= p6_literal_2043923;
  end

  // ===== Pipe stage 7:
  wire [7:0] p7_res7__852_comb;
  wire [7:0] p7_array_index_2050440_comb;
  wire [7:0] p7_res7__854_comb;
  wire [7:0] p7_res7__856_comb;
  wire [7:0] p7_res7__858_comb;
  wire [7:0] p7_res7__860_comb;
  wire [7:0] p7_res7__862_comb;
  wire [127:0] p7_res__26_comb;
  wire [127:0] p7_xor_2050480_comb;
  wire [127:0] p7_addedKey__59_comb;
  wire [7:0] p7_array_index_2050496_comb;
  wire [7:0] p7_array_index_2050497_comb;
  wire [7:0] p7_array_index_2050498_comb;
  wire [7:0] p7_array_index_2050499_comb;
  wire [7:0] p7_array_index_2050500_comb;
  wire [7:0] p7_array_index_2050501_comb;
  wire [7:0] p7_array_index_2050503_comb;
  wire [7:0] p7_array_index_2050505_comb;
  wire [7:0] p7_array_index_2050506_comb;
  wire [7:0] p7_array_index_2050507_comb;
  wire [7:0] p7_array_index_2050508_comb;
  wire [7:0] p7_array_index_2050509_comb;
  wire [7:0] p7_array_index_2050510_comb;
  wire [7:0] p7_array_index_2050512_comb;
  wire [7:0] p7_array_index_2050513_comb;
  wire [7:0] p7_array_index_2050514_comb;
  wire [7:0] p7_array_index_2050515_comb;
  wire [7:0] p7_array_index_2050516_comb;
  wire [7:0] p7_array_index_2050517_comb;
  wire [7:0] p7_array_index_2050518_comb;
  wire [7:0] p7_array_index_2050520_comb;
  wire [7:0] p7_res7__864_comb;
  wire [7:0] p7_array_index_2050529_comb;
  wire [7:0] p7_array_index_2050530_comb;
  wire [7:0] p7_array_index_2050531_comb;
  wire [7:0] p7_array_index_2050532_comb;
  wire [7:0] p7_array_index_2050533_comb;
  wire [7:0] p7_array_index_2050534_comb;
  wire [7:0] p7_res7__866_comb;
  wire [7:0] p7_array_index_2050544_comb;
  wire [7:0] p7_array_index_2050545_comb;
  wire [7:0] p7_array_index_2050546_comb;
  wire [7:0] p7_array_index_2050547_comb;
  wire [7:0] p7_array_index_2050548_comb;
  wire [7:0] p7_res7__868_comb;
  wire [7:0] p7_array_index_2050558_comb;
  wire [7:0] p7_array_index_2050559_comb;
  wire [7:0] p7_array_index_2050560_comb;
  wire [7:0] p7_array_index_2050561_comb;
  wire [7:0] p7_array_index_2050562_comb;
  wire [7:0] p7_res7__870_comb;
  wire [7:0] p7_array_index_2050573_comb;
  wire [7:0] p7_array_index_2050574_comb;
  wire [7:0] p7_array_index_2050575_comb;
  wire [7:0] p7_array_index_2050576_comb;
  wire [7:0] p7_res7__872_comb;
  wire [7:0] p7_array_index_2050586_comb;
  wire [7:0] p7_array_index_2050587_comb;
  wire [7:0] p7_array_index_2050588_comb;
  wire [7:0] p7_array_index_2050589_comb;
  wire [7:0] p7_res7__874_comb;
  wire [7:0] p7_array_index_2050600_comb;
  wire [7:0] p7_array_index_2050601_comb;
  wire [7:0] p7_array_index_2050602_comb;
  wire [7:0] p7_res7__876_comb;
  wire [7:0] p7_array_index_2050612_comb;
  wire [7:0] p7_array_index_2050613_comb;
  wire [7:0] p7_array_index_2050614_comb;
  wire [7:0] p7_res7__878_comb;
  wire [7:0] p7_array_index_2050625_comb;
  wire [7:0] p7_array_index_2050626_comb;
  wire [7:0] p7_res7__880_comb;
  wire [7:0] p7_array_index_2050636_comb;
  wire [7:0] p7_array_index_2050637_comb;
  wire [7:0] p7_res7__882_comb;
  wire [7:0] p7_array_index_2050648_comb;
  wire [7:0] p7_res7__884_comb;
  wire [7:0] p7_array_index_2050658_comb;
  wire [7:0] p7_res7__886_comb;
  wire [7:0] p7_res7__888_comb;
  wire [7:0] p7_res7__890_comb;
  wire [7:0] p7_res7__892_comb;
  wire [7:0] p7_res7__894_comb;
  wire [127:0] p7_res__27_comb;
  wire [127:0] p7_xor_2050698_comb;
  wire [127:0] p7_addedKey__60_comb;
  wire [7:0] p7_array_index_2050714_comb;
  wire [7:0] p7_array_index_2050715_comb;
  wire [7:0] p7_array_index_2050716_comb;
  wire [7:0] p7_array_index_2050717_comb;
  wire [7:0] p7_array_index_2050718_comb;
  wire [7:0] p7_array_index_2050719_comb;
  wire [7:0] p7_array_index_2050721_comb;
  wire [7:0] p7_array_index_2050723_comb;
  wire [7:0] p7_array_index_2050724_comb;
  wire [7:0] p7_array_index_2050725_comb;
  wire [7:0] p7_array_index_2050726_comb;
  wire [7:0] p7_array_index_2050727_comb;
  wire [7:0] p7_array_index_2050728_comb;
  wire [7:0] p7_array_index_2050730_comb;
  wire [7:0] p7_array_index_2050731_comb;
  wire [7:0] p7_array_index_2050732_comb;
  wire [7:0] p7_array_index_2050733_comb;
  wire [7:0] p7_array_index_2050734_comb;
  wire [7:0] p7_array_index_2050735_comb;
  wire [7:0] p7_array_index_2050736_comb;
  wire [7:0] p7_array_index_2050738_comb;
  wire [7:0] p7_res7__896_comb;
  wire [7:0] p7_array_index_2050747_comb;
  wire [7:0] p7_array_index_2050748_comb;
  wire [7:0] p7_array_index_2050749_comb;
  wire [7:0] p7_array_index_2050750_comb;
  wire [7:0] p7_array_index_2050751_comb;
  wire [7:0] p7_array_index_2050752_comb;
  wire [7:0] p7_res7__898_comb;
  wire [7:0] p7_array_index_2050762_comb;
  wire [7:0] p7_array_index_2050763_comb;
  wire [7:0] p7_array_index_2050764_comb;
  wire [7:0] p7_array_index_2050765_comb;
  wire [7:0] p7_array_index_2050766_comb;
  wire [7:0] p7_res7__900_comb;
  wire [7:0] p7_array_index_2050776_comb;
  wire [7:0] p7_array_index_2050777_comb;
  wire [7:0] p7_array_index_2050778_comb;
  wire [7:0] p7_array_index_2050779_comb;
  wire [7:0] p7_array_index_2050780_comb;
  wire [7:0] p7_res7__902_comb;
  wire [7:0] p7_array_index_2050791_comb;
  wire [7:0] p7_array_index_2050792_comb;
  wire [7:0] p7_array_index_2050793_comb;
  wire [7:0] p7_array_index_2050794_comb;
  wire [7:0] p7_res7__904_comb;
  wire [7:0] p7_array_index_2050804_comb;
  wire [7:0] p7_array_index_2050805_comb;
  wire [7:0] p7_array_index_2050806_comb;
  wire [7:0] p7_array_index_2050807_comb;
  wire [7:0] p7_res7__906_comb;
  wire [7:0] p7_array_index_2050818_comb;
  wire [7:0] p7_array_index_2050819_comb;
  wire [7:0] p7_array_index_2050820_comb;
  wire [7:0] p7_res7__908_comb;
  wire [7:0] p7_array_index_2050830_comb;
  wire [7:0] p7_array_index_2050831_comb;
  wire [7:0] p7_array_index_2050832_comb;
  wire [7:0] p7_res7__910_comb;
  wire [7:0] p7_array_index_2050843_comb;
  wire [7:0] p7_array_index_2050844_comb;
  wire [7:0] p7_res7__912_comb;
  wire [7:0] p7_array_index_2050854_comb;
  wire [7:0] p7_array_index_2050855_comb;
  wire [7:0] p7_res7__914_comb;
  wire [7:0] p7_array_index_2050866_comb;
  wire [7:0] p7_res7__916_comb;
  wire [7:0] p7_array_index_2050876_comb;
  wire [7:0] p7_res7__918_comb;
  wire [7:0] p7_res7__920_comb;
  wire [7:0] p7_res7__922_comb;
  wire [7:0] p7_res7__924_comb;
  wire [7:0] p7_res7__926_comb;
  wire [127:0] p7_res__28_comb;
  wire [127:0] p7_xor_2050916_comb;
  wire [127:0] p7_addedKey__61_comb;
  wire [7:0] p7_array_index_2050932_comb;
  wire [7:0] p7_array_index_2050933_comb;
  wire [7:0] p7_array_index_2050934_comb;
  wire [7:0] p7_array_index_2050935_comb;
  wire [7:0] p7_array_index_2050936_comb;
  wire [7:0] p7_array_index_2050937_comb;
  wire [7:0] p7_array_index_2050939_comb;
  wire [7:0] p7_array_index_2050941_comb;
  wire [7:0] p7_array_index_2050942_comb;
  wire [7:0] p7_array_index_2050943_comb;
  wire [7:0] p7_array_index_2050944_comb;
  wire [7:0] p7_array_index_2050945_comb;
  wire [7:0] p7_array_index_2050946_comb;
  wire [7:0] p7_array_index_2050948_comb;
  wire [7:0] p7_array_index_2050949_comb;
  wire [7:0] p7_array_index_2050950_comb;
  wire [7:0] p7_array_index_2050951_comb;
  wire [7:0] p7_array_index_2050952_comb;
  wire [7:0] p7_array_index_2050953_comb;
  wire [7:0] p7_array_index_2050954_comb;
  wire [7:0] p7_array_index_2050956_comb;
  wire [7:0] p7_res7__928_comb;
  wire [7:0] p7_array_index_2050965_comb;
  wire [7:0] p7_array_index_2050966_comb;
  wire [7:0] p7_array_index_2050967_comb;
  wire [7:0] p7_array_index_2050968_comb;
  wire [7:0] p7_array_index_2050969_comb;
  wire [7:0] p7_array_index_2050970_comb;
  wire [7:0] p7_res7__930_comb;
  wire [7:0] p7_array_index_2050980_comb;
  wire [7:0] p7_array_index_2050981_comb;
  wire [7:0] p7_array_index_2050982_comb;
  wire [7:0] p7_array_index_2050983_comb;
  wire [7:0] p7_array_index_2050984_comb;
  wire [7:0] p7_res7__932_comb;
  wire [7:0] p7_array_index_2050994_comb;
  wire [7:0] p7_array_index_2050995_comb;
  wire [7:0] p7_array_index_2050996_comb;
  wire [7:0] p7_array_index_2050997_comb;
  wire [7:0] p7_array_index_2050998_comb;
  wire [7:0] p7_res7__934_comb;
  wire [7:0] p7_array_index_2051009_comb;
  wire [7:0] p7_array_index_2051010_comb;
  wire [7:0] p7_array_index_2051011_comb;
  wire [7:0] p7_array_index_2051012_comb;
  wire [7:0] p7_res7__936_comb;
  wire [7:0] p7_array_index_2051022_comb;
  wire [7:0] p7_array_index_2051023_comb;
  wire [7:0] p7_array_index_2051024_comb;
  wire [7:0] p7_array_index_2051025_comb;
  wire [7:0] p7_res7__938_comb;
  wire [7:0] p7_array_index_2051036_comb;
  wire [7:0] p7_array_index_2051037_comb;
  wire [7:0] p7_array_index_2051038_comb;
  wire [7:0] p7_res7__940_comb;
  wire [7:0] p7_array_index_2051048_comb;
  wire [7:0] p7_array_index_2051049_comb;
  wire [7:0] p7_array_index_2051050_comb;
  wire [7:0] p7_res7__942_comb;
  wire [7:0] p7_array_index_2051061_comb;
  wire [7:0] p7_array_index_2051062_comb;
  wire [7:0] p7_res7__944_comb;
  wire [7:0] p7_array_index_2051072_comb;
  wire [7:0] p7_array_index_2051073_comb;
  wire [7:0] p7_res7__946_comb;
  wire [7:0] p7_array_index_2051084_comb;
  wire [7:0] p7_res7__948_comb;
  wire [7:0] p7_array_index_2051094_comb;
  wire [7:0] p7_res7__950_comb;
  wire [7:0] p7_res7__952_comb;
  wire [7:0] p7_res7__954_comb;
  wire [7:0] p7_res7__956_comb;
  wire [7:0] p7_res7__958_comb;
  wire [127:0] p7_res__29_comb;
  wire [127:0] p7_xor_2051134_comb;
  wire [127:0] p7_addedKey__62_comb;
  wire [7:0] p7_array_index_2051150_comb;
  wire [7:0] p7_array_index_2051151_comb;
  wire [7:0] p7_array_index_2051152_comb;
  wire [7:0] p7_array_index_2051153_comb;
  wire [7:0] p7_array_index_2051154_comb;
  wire [7:0] p7_array_index_2051155_comb;
  wire [7:0] p7_array_index_2051157_comb;
  wire [7:0] p7_array_index_2051159_comb;
  wire [7:0] p7_array_index_2051160_comb;
  wire [7:0] p7_array_index_2051161_comb;
  wire [7:0] p7_array_index_2051162_comb;
  wire [7:0] p7_array_index_2051163_comb;
  wire [7:0] p7_array_index_2051164_comb;
  wire [7:0] p7_array_index_2051166_comb;
  wire [7:0] p7_array_index_2051167_comb;
  wire [7:0] p7_array_index_2051168_comb;
  wire [7:0] p7_array_index_2051169_comb;
  wire [7:0] p7_array_index_2051170_comb;
  wire [7:0] p7_array_index_2051171_comb;
  wire [7:0] p7_array_index_2051172_comb;
  wire [7:0] p7_array_index_2051174_comb;
  wire [7:0] p7_res7__960_comb;
  wire [7:0] p7_array_index_2051183_comb;
  wire [7:0] p7_array_index_2051184_comb;
  wire [7:0] p7_array_index_2051185_comb;
  wire [7:0] p7_array_index_2051186_comb;
  wire [7:0] p7_array_index_2051187_comb;
  wire [7:0] p7_array_index_2051188_comb;
  wire [7:0] p7_res7__962_comb;
  wire [7:0] p7_array_index_2051198_comb;
  wire [7:0] p7_array_index_2051199_comb;
  wire [7:0] p7_array_index_2051200_comb;
  wire [7:0] p7_array_index_2051201_comb;
  wire [7:0] p7_array_index_2051202_comb;
  wire [7:0] p7_res7__964_comb;
  wire [7:0] p7_array_index_2051212_comb;
  wire [7:0] p7_array_index_2051213_comb;
  wire [7:0] p7_array_index_2051214_comb;
  wire [7:0] p7_array_index_2051215_comb;
  wire [7:0] p7_array_index_2051216_comb;
  wire [7:0] p7_res7__966_comb;
  wire [7:0] p7_array_index_2051227_comb;
  wire [7:0] p7_array_index_2051228_comb;
  wire [7:0] p7_array_index_2051229_comb;
  wire [7:0] p7_array_index_2051230_comb;
  wire [7:0] p7_res7__968_comb;
  wire [7:0] p7_array_index_2051240_comb;
  wire [7:0] p7_array_index_2051241_comb;
  wire [7:0] p7_array_index_2051242_comb;
  wire [7:0] p7_array_index_2051243_comb;
  wire [7:0] p7_res7__970_comb;
  wire [7:0] p7_array_index_2051254_comb;
  wire [7:0] p7_array_index_2051255_comb;
  wire [7:0] p7_array_index_2051256_comb;
  wire [7:0] p7_res7__972_comb;
  wire [7:0] p7_array_index_2051266_comb;
  wire [7:0] p7_array_index_2051267_comb;
  wire [7:0] p7_array_index_2051268_comb;
  wire [7:0] p7_res7__974_comb;
  wire [7:0] p7_array_index_2051279_comb;
  wire [7:0] p7_array_index_2051280_comb;
  wire [7:0] p7_res7__976_comb;
  wire [7:0] p7_array_index_2051290_comb;
  wire [7:0] p7_array_index_2051291_comb;
  wire [7:0] p7_res7__978_comb;
  wire [7:0] p7_array_index_2051302_comb;
  wire [7:0] p7_res7__980_comb;
  wire [7:0] p7_array_index_2051312_comb;
  wire [7:0] p7_res7__982_comb;
  wire [7:0] p7_res7__984_comb;
  wire [7:0] p7_res7__986_comb;
  wire [7:0] p7_res7__988_comb;
  wire [7:0] p7_res7__990_comb;
  wire [127:0] p7_res__30_comb;
  wire [127:0] p7_k9_comb;
  wire [127:0] p7_xor_2051355_comb;
  wire [127:0] p7_addedKey__63_comb;
  wire [7:0] p7_bit_slice_2051370_comb;
  wire [7:0] p7_bit_slice_2051371_comb;
  wire [7:0] p7_bit_slice_2051372_comb;
  wire [7:0] p7_bit_slice_2051373_comb;
  wire [7:0] p7_bit_slice_2051374_comb;
  wire [7:0] p7_bit_slice_2051375_comb;
  wire [7:0] p7_bit_slice_2051376_comb;
  wire [7:0] p7_bit_slice_2051377_comb;
  wire [7:0] p7_bit_slice_2051378_comb;
  wire [7:0] p7_bit_slice_2051379_comb;
  wire [7:0] p7_bit_slice_2051380_comb;
  wire [7:0] p7_bit_slice_2051381_comb;
  wire [7:0] p7_bit_slice_2051404_comb;
  wire [7:0] p7_bit_slice_2051406_comb;
  wire [7:0] p7_array_index_2051407_comb;
  wire [7:0] p7_array_index_2051408_comb;
  wire [7:0] p7_array_index_2051409_comb;
  wire [7:0] p7_array_index_2051410_comb;
  wire [7:0] p7_array_index_2051411_comb;
  wire [7:0] p7_array_index_2051412_comb;
  wire [7:0] p7_array_index_2051382_comb;
  wire [7:0] p7_array_index_2051383_comb;
  wire [7:0] p7_array_index_2051384_comb;
  wire [7:0] p7_array_index_2051385_comb;
  wire [7:0] p7_array_index_2051386_comb;
  wire [7:0] p7_array_index_2051387_comb;
  wire [7:0] p7_array_index_2051389_comb;
  wire [7:0] p7_array_index_2051391_comb;
  wire [7:0] p7_array_index_2051392_comb;
  wire [7:0] p7_array_index_2051393_comb;
  wire [7:0] p7_array_index_2051394_comb;
  wire [7:0] p7_array_index_2051395_comb;
  wire [7:0] p7_array_index_2051396_comb;
  wire [7:0] p7_res7__1025_comb;
  wire [7:0] p7_array_index_2051414_comb;
  wire [7:0] p7_array_index_2051415_comb;
  wire [7:0] p7_array_index_2051416_comb;
  wire [7:0] p7_array_index_2051417_comb;
  wire [7:0] p7_array_index_2051418_comb;
  wire [7:0] p7_array_index_2051419_comb;
  wire [7:0] p7_array_index_2051420_comb;
  wire [7:0] p7_array_index_2051422_comb;
  wire [7:0] p7_array_index_2051439_comb;
  wire [7:0] p7_array_index_2051440_comb;
  wire [7:0] p7_array_index_2051441_comb;
  wire [7:0] p7_array_index_2051442_comb;
  wire [7:0] p7_array_index_2051443_comb;
  wire [7:0] p7_array_index_2051444_comb;
  wire [7:0] p7_res7__992_comb;
  wire [7:0] p7_res7__1027_comb;
  assign p7_res7__852_comb = p6_array_index_2050281 ^ p6_array_index_2050282 ^ p6_array_index_2050283 ^ p6_array_index_2050284 ^ p6_array_index_2050285 ^ p6_array_index_2050286 ^ p6_res7__838 ^ p6_array_index_2050287 ^ p6_res7__834 ^ p6_array_index_2050240 ^ p6_array_index_2050213 ^ p6_array_index_2050184 ^ p6_array_index_2050152 ^ p6_array_index_2050288 ^ p6_array_index_2050289 ^ p6_array_index_2050139;
  assign p7_array_index_2050440_comb = p6_literal_2043920[p6_res7__842];
  assign p7_res7__854_comb = p6_literal_2043910[p7_res7__852_comb] ^ p6_literal_2043912[p6_res7__850] ^ p6_literal_2043914[p6_res7__848] ^ p6_literal_2043916[p6_res7__846] ^ p6_literal_2043918[p6_res7__844] ^ p7_array_index_2050440_comb ^ p6_res7__840 ^ p6_literal_2043923[p6_res7__838] ^ p6_res7__836 ^ p6_array_index_2050252 ^ p6_array_index_2050226 ^ p6_array_index_2050198 ^ p6_array_index_2050169 ^ p6_literal_2043912[p6_array_index_2050136] ^ p6_literal_2043910[p6_array_index_2050137] ^ p6_array_index_2050138;
  assign p7_res7__856_comb = p6_literal_2043910[p7_res7__854_comb] ^ p6_literal_2043912[p7_res7__852_comb] ^ p6_literal_2043914[p6_res7__850] ^ p6_literal_2043916[p6_res7__848] ^ p6_literal_2043918[p6_res7__846] ^ p6_literal_2043920[p6_res7__844] ^ p6_res7__842 ^ p6_literal_2043923[p6_res7__840] ^ p6_res7__838 ^ p6_array_index_2050264 ^ p6_array_index_2050239 ^ p6_array_index_2050212 ^ p6_array_index_2050183 ^ p6_array_index_2050151 ^ p6_literal_2043910[p6_array_index_2050136] ^ p6_array_index_2050137;
  assign p7_res7__858_comb = p6_literal_2043910[p7_res7__856_comb] ^ p6_literal_2043912[p7_res7__854_comb] ^ p6_literal_2043914[p7_res7__852_comb] ^ p6_literal_2043916[p6_res7__850] ^ p6_literal_2043918[p6_res7__848] ^ p6_literal_2043920[p6_res7__846] ^ p6_res7__844 ^ p6_literal_2043923[p6_res7__842] ^ p6_res7__840 ^ p6_array_index_2050275 ^ p6_array_index_2050251 ^ p6_array_index_2050225 ^ p6_array_index_2050197 ^ p6_array_index_2050168 ^ p6_literal_2043910[p6_array_index_2050135] ^ p6_array_index_2050136;
  assign p7_res7__860_comb = p6_literal_2043910[p7_res7__858_comb] ^ p6_literal_2043912[p7_res7__856_comb] ^ p6_literal_2043914[p7_res7__854_comb] ^ p6_literal_2043916[p7_res7__852_comb] ^ p6_literal_2043918[p6_res7__850] ^ p6_literal_2043920[p6_res7__848] ^ p6_res7__846 ^ p6_literal_2043923[p6_res7__844] ^ p6_res7__842 ^ p6_array_index_2050286 ^ p6_array_index_2050263 ^ p6_array_index_2050238 ^ p6_array_index_2050211 ^ p6_array_index_2050182 ^ p6_array_index_2050150 ^ p6_array_index_2050135;
  assign p7_res7__862_comb = p6_literal_2043910[p7_res7__860_comb] ^ p6_literal_2043912[p7_res7__858_comb] ^ p6_literal_2043914[p7_res7__856_comb] ^ p6_literal_2043916[p7_res7__854_comb] ^ p6_literal_2043918[p7_res7__852_comb] ^ p6_literal_2043920[p6_res7__850] ^ p6_res7__848 ^ p6_literal_2043923[p6_res7__846] ^ p6_res7__844 ^ p7_array_index_2050440_comb ^ p6_array_index_2050274 ^ p6_array_index_2050250 ^ p6_array_index_2050224 ^ p6_array_index_2050196 ^ p6_array_index_2050167 ^ p6_array_index_2050134;
  assign p7_res__26_comb = {p7_res7__862_comb, p7_res7__860_comb, p7_res7__858_comb, p7_res7__856_comb, p7_res7__854_comb, p7_res7__852_comb, p6_res7__850, p6_res7__848, p6_res7__846, p6_res7__844, p6_res7__842, p6_res7__840, p6_res7__838, p6_res7__836, p6_res7__834, p6_res7__832};
  assign p7_xor_2050480_comb = p7_res__26_comb ^ p6_xor_2049900;
  assign p7_addedKey__59_comb = p7_xor_2050480_comb ^ 128'ha226_4131_9aec_d1fd_8352_9103_9b68_6b1c;
  assign p7_array_index_2050496_comb = p6_literal_2043896[p7_addedKey__59_comb[127:120]];
  assign p7_array_index_2050497_comb = p6_literal_2043896[p7_addedKey__59_comb[119:112]];
  assign p7_array_index_2050498_comb = p6_literal_2043896[p7_addedKey__59_comb[111:104]];
  assign p7_array_index_2050499_comb = p6_literal_2043896[p7_addedKey__59_comb[103:96]];
  assign p7_array_index_2050500_comb = p6_literal_2043896[p7_addedKey__59_comb[95:88]];
  assign p7_array_index_2050501_comb = p6_literal_2043896[p7_addedKey__59_comb[87:80]];
  assign p7_array_index_2050503_comb = p6_literal_2043896[p7_addedKey__59_comb[71:64]];
  assign p7_array_index_2050505_comb = p6_literal_2043896[p7_addedKey__59_comb[55:48]];
  assign p7_array_index_2050506_comb = p6_literal_2043896[p7_addedKey__59_comb[47:40]];
  assign p7_array_index_2050507_comb = p6_literal_2043896[p7_addedKey__59_comb[39:32]];
  assign p7_array_index_2050508_comb = p6_literal_2043896[p7_addedKey__59_comb[31:24]];
  assign p7_array_index_2050509_comb = p6_literal_2043896[p7_addedKey__59_comb[23:16]];
  assign p7_array_index_2050510_comb = p6_literal_2043896[p7_addedKey__59_comb[15:8]];
  assign p7_array_index_2050512_comb = p6_literal_2043910[p7_array_index_2050496_comb];
  assign p7_array_index_2050513_comb = p6_literal_2043912[p7_array_index_2050497_comb];
  assign p7_array_index_2050514_comb = p6_literal_2043914[p7_array_index_2050498_comb];
  assign p7_array_index_2050515_comb = p6_literal_2043916[p7_array_index_2050499_comb];
  assign p7_array_index_2050516_comb = p6_literal_2043918[p7_array_index_2050500_comb];
  assign p7_array_index_2050517_comb = p6_literal_2043920[p7_array_index_2050501_comb];
  assign p7_array_index_2050518_comb = p6_literal_2043896[p7_addedKey__59_comb[79:72]];
  assign p7_array_index_2050520_comb = p6_literal_2043896[p7_addedKey__59_comb[63:56]];
  assign p7_res7__864_comb = p7_array_index_2050512_comb ^ p7_array_index_2050513_comb ^ p7_array_index_2050514_comb ^ p7_array_index_2050515_comb ^ p7_array_index_2050516_comb ^ p7_array_index_2050517_comb ^ p7_array_index_2050518_comb ^ p6_literal_2043923[p7_array_index_2050503_comb] ^ p7_array_index_2050520_comb ^ p6_literal_2043920[p7_array_index_2050505_comb] ^ p6_literal_2043918[p7_array_index_2050506_comb] ^ p6_literal_2043916[p7_array_index_2050507_comb] ^ p6_literal_2043914[p7_array_index_2050508_comb] ^ p6_literal_2043912[p7_array_index_2050509_comb] ^ p6_literal_2043910[p7_array_index_2050510_comb] ^ p6_literal_2043896[p7_addedKey__59_comb[7:0]];
  assign p7_array_index_2050529_comb = p6_literal_2043910[p7_res7__864_comb];
  assign p7_array_index_2050530_comb = p6_literal_2043912[p7_array_index_2050496_comb];
  assign p7_array_index_2050531_comb = p6_literal_2043914[p7_array_index_2050497_comb];
  assign p7_array_index_2050532_comb = p6_literal_2043916[p7_array_index_2050498_comb];
  assign p7_array_index_2050533_comb = p6_literal_2043918[p7_array_index_2050499_comb];
  assign p7_array_index_2050534_comb = p6_literal_2043920[p7_array_index_2050500_comb];
  assign p7_res7__866_comb = p7_array_index_2050529_comb ^ p7_array_index_2050530_comb ^ p7_array_index_2050531_comb ^ p7_array_index_2050532_comb ^ p7_array_index_2050533_comb ^ p7_array_index_2050534_comb ^ p7_array_index_2050501_comb ^ p6_literal_2043923[p7_array_index_2050518_comb] ^ p7_array_index_2050503_comb ^ p6_literal_2043920[p7_array_index_2050520_comb] ^ p6_literal_2043918[p7_array_index_2050505_comb] ^ p6_literal_2043916[p7_array_index_2050506_comb] ^ p6_literal_2043914[p7_array_index_2050507_comb] ^ p6_literal_2043912[p7_array_index_2050508_comb] ^ p6_literal_2043910[p7_array_index_2050509_comb] ^ p7_array_index_2050510_comb;
  assign p7_array_index_2050544_comb = p6_literal_2043912[p7_res7__864_comb];
  assign p7_array_index_2050545_comb = p6_literal_2043914[p7_array_index_2050496_comb];
  assign p7_array_index_2050546_comb = p6_literal_2043916[p7_array_index_2050497_comb];
  assign p7_array_index_2050547_comb = p6_literal_2043918[p7_array_index_2050498_comb];
  assign p7_array_index_2050548_comb = p6_literal_2043920[p7_array_index_2050499_comb];
  assign p7_res7__868_comb = p6_literal_2043910[p7_res7__866_comb] ^ p7_array_index_2050544_comb ^ p7_array_index_2050545_comb ^ p7_array_index_2050546_comb ^ p7_array_index_2050547_comb ^ p7_array_index_2050548_comb ^ p7_array_index_2050500_comb ^ p6_literal_2043923[p7_array_index_2050501_comb] ^ p7_array_index_2050518_comb ^ p6_literal_2043920[p7_array_index_2050503_comb] ^ p6_literal_2043918[p7_array_index_2050520_comb] ^ p6_literal_2043916[p7_array_index_2050505_comb] ^ p6_literal_2043914[p7_array_index_2050506_comb] ^ p6_literal_2043912[p7_array_index_2050507_comb] ^ p6_literal_2043910[p7_array_index_2050508_comb] ^ p7_array_index_2050509_comb;
  assign p7_array_index_2050558_comb = p6_literal_2043912[p7_res7__866_comb];
  assign p7_array_index_2050559_comb = p6_literal_2043914[p7_res7__864_comb];
  assign p7_array_index_2050560_comb = p6_literal_2043916[p7_array_index_2050496_comb];
  assign p7_array_index_2050561_comb = p6_literal_2043918[p7_array_index_2050497_comb];
  assign p7_array_index_2050562_comb = p6_literal_2043920[p7_array_index_2050498_comb];
  assign p7_res7__870_comb = p6_literal_2043910[p7_res7__868_comb] ^ p7_array_index_2050558_comb ^ p7_array_index_2050559_comb ^ p7_array_index_2050560_comb ^ p7_array_index_2050561_comb ^ p7_array_index_2050562_comb ^ p7_array_index_2050499_comb ^ p6_literal_2043923[p7_array_index_2050500_comb] ^ p7_array_index_2050501_comb ^ p6_literal_2043920[p7_array_index_2050518_comb] ^ p6_literal_2043918[p7_array_index_2050503_comb] ^ p6_literal_2043916[p7_array_index_2050520_comb] ^ p6_literal_2043914[p7_array_index_2050505_comb] ^ p6_literal_2043912[p7_array_index_2050506_comb] ^ p6_literal_2043910[p7_array_index_2050507_comb] ^ p7_array_index_2050508_comb;
  assign p7_array_index_2050573_comb = p6_literal_2043914[p7_res7__866_comb];
  assign p7_array_index_2050574_comb = p6_literal_2043916[p7_res7__864_comb];
  assign p7_array_index_2050575_comb = p6_literal_2043918[p7_array_index_2050496_comb];
  assign p7_array_index_2050576_comb = p6_literal_2043920[p7_array_index_2050497_comb];
  assign p7_res7__872_comb = p6_literal_2043910[p7_res7__870_comb] ^ p6_literal_2043912[p7_res7__868_comb] ^ p7_array_index_2050573_comb ^ p7_array_index_2050574_comb ^ p7_array_index_2050575_comb ^ p7_array_index_2050576_comb ^ p7_array_index_2050498_comb ^ p6_literal_2043923[p7_array_index_2050499_comb] ^ p7_array_index_2050500_comb ^ p7_array_index_2050517_comb ^ p6_literal_2043918[p7_array_index_2050518_comb] ^ p6_literal_2043916[p7_array_index_2050503_comb] ^ p6_literal_2043914[p7_array_index_2050520_comb] ^ p6_literal_2043912[p7_array_index_2050505_comb] ^ p6_literal_2043910[p7_array_index_2050506_comb] ^ p7_array_index_2050507_comb;
  assign p7_array_index_2050586_comb = p6_literal_2043914[p7_res7__868_comb];
  assign p7_array_index_2050587_comb = p6_literal_2043916[p7_res7__866_comb];
  assign p7_array_index_2050588_comb = p6_literal_2043918[p7_res7__864_comb];
  assign p7_array_index_2050589_comb = p6_literal_2043920[p7_array_index_2050496_comb];
  assign p7_res7__874_comb = p6_literal_2043910[p7_res7__872_comb] ^ p6_literal_2043912[p7_res7__870_comb] ^ p7_array_index_2050586_comb ^ p7_array_index_2050587_comb ^ p7_array_index_2050588_comb ^ p7_array_index_2050589_comb ^ p7_array_index_2050497_comb ^ p6_literal_2043923[p7_array_index_2050498_comb] ^ p7_array_index_2050499_comb ^ p7_array_index_2050534_comb ^ p6_literal_2043918[p7_array_index_2050501_comb] ^ p6_literal_2043916[p7_array_index_2050518_comb] ^ p6_literal_2043914[p7_array_index_2050503_comb] ^ p6_literal_2043912[p7_array_index_2050520_comb] ^ p6_literal_2043910[p7_array_index_2050505_comb] ^ p7_array_index_2050506_comb;
  assign p7_array_index_2050600_comb = p6_literal_2043916[p7_res7__868_comb];
  assign p7_array_index_2050601_comb = p6_literal_2043918[p7_res7__866_comb];
  assign p7_array_index_2050602_comb = p6_literal_2043920[p7_res7__864_comb];
  assign p7_res7__876_comb = p6_literal_2043910[p7_res7__874_comb] ^ p6_literal_2043912[p7_res7__872_comb] ^ p6_literal_2043914[p7_res7__870_comb] ^ p7_array_index_2050600_comb ^ p7_array_index_2050601_comb ^ p7_array_index_2050602_comb ^ p7_array_index_2050496_comb ^ p6_literal_2043923[p7_array_index_2050497_comb] ^ p7_array_index_2050498_comb ^ p7_array_index_2050548_comb ^ p7_array_index_2050516_comb ^ p6_literal_2043916[p7_array_index_2050501_comb] ^ p6_literal_2043914[p7_array_index_2050518_comb] ^ p6_literal_2043912[p7_array_index_2050503_comb] ^ p6_literal_2043910[p7_array_index_2050520_comb] ^ p7_array_index_2050505_comb;
  assign p7_array_index_2050612_comb = p6_literal_2043916[p7_res7__870_comb];
  assign p7_array_index_2050613_comb = p6_literal_2043918[p7_res7__868_comb];
  assign p7_array_index_2050614_comb = p6_literal_2043920[p7_res7__866_comb];
  assign p7_res7__878_comb = p6_literal_2043910[p7_res7__876_comb] ^ p6_literal_2043912[p7_res7__874_comb] ^ p6_literal_2043914[p7_res7__872_comb] ^ p7_array_index_2050612_comb ^ p7_array_index_2050613_comb ^ p7_array_index_2050614_comb ^ p7_res7__864_comb ^ p6_literal_2043923[p7_array_index_2050496_comb] ^ p7_array_index_2050497_comb ^ p7_array_index_2050562_comb ^ p7_array_index_2050533_comb ^ p6_literal_2043916[p7_array_index_2050500_comb] ^ p6_literal_2043914[p7_array_index_2050501_comb] ^ p6_literal_2043912[p7_array_index_2050518_comb] ^ p6_literal_2043910[p7_array_index_2050503_comb] ^ p7_array_index_2050520_comb;
  assign p7_array_index_2050625_comb = p6_literal_2043918[p7_res7__870_comb];
  assign p7_array_index_2050626_comb = p6_literal_2043920[p7_res7__868_comb];
  assign p7_res7__880_comb = p6_literal_2043910[p7_res7__878_comb] ^ p6_literal_2043912[p7_res7__876_comb] ^ p6_literal_2043914[p7_res7__874_comb] ^ p6_literal_2043916[p7_res7__872_comb] ^ p7_array_index_2050625_comb ^ p7_array_index_2050626_comb ^ p7_res7__866_comb ^ p6_literal_2043923[p7_res7__864_comb] ^ p7_array_index_2050496_comb ^ p7_array_index_2050576_comb ^ p7_array_index_2050547_comb ^ p7_array_index_2050515_comb ^ p6_literal_2043914[p7_array_index_2050500_comb] ^ p6_literal_2043912[p7_array_index_2050501_comb] ^ p6_literal_2043910[p7_array_index_2050518_comb] ^ p7_array_index_2050503_comb;
  assign p7_array_index_2050636_comb = p6_literal_2043918[p7_res7__872_comb];
  assign p7_array_index_2050637_comb = p6_literal_2043920[p7_res7__870_comb];
  assign p7_res7__882_comb = p6_literal_2043910[p7_res7__880_comb] ^ p6_literal_2043912[p7_res7__878_comb] ^ p6_literal_2043914[p7_res7__876_comb] ^ p6_literal_2043916[p7_res7__874_comb] ^ p7_array_index_2050636_comb ^ p7_array_index_2050637_comb ^ p7_res7__868_comb ^ p6_literal_2043923[p7_res7__866_comb] ^ p7_res7__864_comb ^ p7_array_index_2050589_comb ^ p7_array_index_2050561_comb ^ p7_array_index_2050532_comb ^ p6_literal_2043914[p7_array_index_2050499_comb] ^ p6_literal_2043912[p7_array_index_2050500_comb] ^ p6_literal_2043910[p7_array_index_2050501_comb] ^ p7_array_index_2050518_comb;
  assign p7_array_index_2050648_comb = p6_literal_2043920[p7_res7__872_comb];
  assign p7_res7__884_comb = p6_literal_2043910[p7_res7__882_comb] ^ p6_literal_2043912[p7_res7__880_comb] ^ p6_literal_2043914[p7_res7__878_comb] ^ p6_literal_2043916[p7_res7__876_comb] ^ p6_literal_2043918[p7_res7__874_comb] ^ p7_array_index_2050648_comb ^ p7_res7__870_comb ^ p6_literal_2043923[p7_res7__868_comb] ^ p7_res7__866_comb ^ p7_array_index_2050602_comb ^ p7_array_index_2050575_comb ^ p7_array_index_2050546_comb ^ p7_array_index_2050514_comb ^ p6_literal_2043912[p7_array_index_2050499_comb] ^ p6_literal_2043910[p7_array_index_2050500_comb] ^ p7_array_index_2050501_comb;
  assign p7_array_index_2050658_comb = p6_literal_2043920[p7_res7__874_comb];
  assign p7_res7__886_comb = p6_literal_2043910[p7_res7__884_comb] ^ p6_literal_2043912[p7_res7__882_comb] ^ p6_literal_2043914[p7_res7__880_comb] ^ p6_literal_2043916[p7_res7__878_comb] ^ p6_literal_2043918[p7_res7__876_comb] ^ p7_array_index_2050658_comb ^ p7_res7__872_comb ^ p6_literal_2043923[p7_res7__870_comb] ^ p7_res7__868_comb ^ p7_array_index_2050614_comb ^ p7_array_index_2050588_comb ^ p7_array_index_2050560_comb ^ p7_array_index_2050531_comb ^ p6_literal_2043912[p7_array_index_2050498_comb] ^ p6_literal_2043910[p7_array_index_2050499_comb] ^ p7_array_index_2050500_comb;
  assign p7_res7__888_comb = p6_literal_2043910[p7_res7__886_comb] ^ p6_literal_2043912[p7_res7__884_comb] ^ p6_literal_2043914[p7_res7__882_comb] ^ p6_literal_2043916[p7_res7__880_comb] ^ p6_literal_2043918[p7_res7__878_comb] ^ p6_literal_2043920[p7_res7__876_comb] ^ p7_res7__874_comb ^ p6_literal_2043923[p7_res7__872_comb] ^ p7_res7__870_comb ^ p7_array_index_2050626_comb ^ p7_array_index_2050601_comb ^ p7_array_index_2050574_comb ^ p7_array_index_2050545_comb ^ p7_array_index_2050513_comb ^ p6_literal_2043910[p7_array_index_2050498_comb] ^ p7_array_index_2050499_comb;
  assign p7_res7__890_comb = p6_literal_2043910[p7_res7__888_comb] ^ p6_literal_2043912[p7_res7__886_comb] ^ p6_literal_2043914[p7_res7__884_comb] ^ p6_literal_2043916[p7_res7__882_comb] ^ p6_literal_2043918[p7_res7__880_comb] ^ p6_literal_2043920[p7_res7__878_comb] ^ p7_res7__876_comb ^ p6_literal_2043923[p7_res7__874_comb] ^ p7_res7__872_comb ^ p7_array_index_2050637_comb ^ p7_array_index_2050613_comb ^ p7_array_index_2050587_comb ^ p7_array_index_2050559_comb ^ p7_array_index_2050530_comb ^ p6_literal_2043910[p7_array_index_2050497_comb] ^ p7_array_index_2050498_comb;
  assign p7_res7__892_comb = p6_literal_2043910[p7_res7__890_comb] ^ p6_literal_2043912[p7_res7__888_comb] ^ p6_literal_2043914[p7_res7__886_comb] ^ p6_literal_2043916[p7_res7__884_comb] ^ p6_literal_2043918[p7_res7__882_comb] ^ p6_literal_2043920[p7_res7__880_comb] ^ p7_res7__878_comb ^ p6_literal_2043923[p7_res7__876_comb] ^ p7_res7__874_comb ^ p7_array_index_2050648_comb ^ p7_array_index_2050625_comb ^ p7_array_index_2050600_comb ^ p7_array_index_2050573_comb ^ p7_array_index_2050544_comb ^ p7_array_index_2050512_comb ^ p7_array_index_2050497_comb;
  assign p7_res7__894_comb = p6_literal_2043910[p7_res7__892_comb] ^ p6_literal_2043912[p7_res7__890_comb] ^ p6_literal_2043914[p7_res7__888_comb] ^ p6_literal_2043916[p7_res7__886_comb] ^ p6_literal_2043918[p7_res7__884_comb] ^ p6_literal_2043920[p7_res7__882_comb] ^ p7_res7__880_comb ^ p6_literal_2043923[p7_res7__878_comb] ^ p7_res7__876_comb ^ p7_array_index_2050658_comb ^ p7_array_index_2050636_comb ^ p7_array_index_2050612_comb ^ p7_array_index_2050586_comb ^ p7_array_index_2050558_comb ^ p7_array_index_2050529_comb ^ p7_array_index_2050496_comb;
  assign p7_res__27_comb = {p7_res7__894_comb, p7_res7__892_comb, p7_res7__890_comb, p7_res7__888_comb, p7_res7__886_comb, p7_res7__884_comb, p7_res7__882_comb, p7_res7__880_comb, p7_res7__878_comb, p7_res7__876_comb, p7_res7__874_comb, p7_res7__872_comb, p7_res7__870_comb, p7_res7__868_comb, p7_res7__866_comb, p7_res7__864_comb};
  assign p7_xor_2050698_comb = p7_res__27_comb ^ p6_xor_2050118;
  assign p7_addedKey__60_comb = p7_xor_2050698_comb ^ 128'hcc84_3743_f6a4_ab45_de75_2c13_46ec_ff1d;
  assign p7_array_index_2050714_comb = p6_literal_2043896[p7_addedKey__60_comb[127:120]];
  assign p7_array_index_2050715_comb = p6_literal_2043896[p7_addedKey__60_comb[119:112]];
  assign p7_array_index_2050716_comb = p6_literal_2043896[p7_addedKey__60_comb[111:104]];
  assign p7_array_index_2050717_comb = p6_literal_2043896[p7_addedKey__60_comb[103:96]];
  assign p7_array_index_2050718_comb = p6_literal_2043896[p7_addedKey__60_comb[95:88]];
  assign p7_array_index_2050719_comb = p6_literal_2043896[p7_addedKey__60_comb[87:80]];
  assign p7_array_index_2050721_comb = p6_literal_2043896[p7_addedKey__60_comb[71:64]];
  assign p7_array_index_2050723_comb = p6_literal_2043896[p7_addedKey__60_comb[55:48]];
  assign p7_array_index_2050724_comb = p6_literal_2043896[p7_addedKey__60_comb[47:40]];
  assign p7_array_index_2050725_comb = p6_literal_2043896[p7_addedKey__60_comb[39:32]];
  assign p7_array_index_2050726_comb = p6_literal_2043896[p7_addedKey__60_comb[31:24]];
  assign p7_array_index_2050727_comb = p6_literal_2043896[p7_addedKey__60_comb[23:16]];
  assign p7_array_index_2050728_comb = p6_literal_2043896[p7_addedKey__60_comb[15:8]];
  assign p7_array_index_2050730_comb = p6_literal_2043910[p7_array_index_2050714_comb];
  assign p7_array_index_2050731_comb = p6_literal_2043912[p7_array_index_2050715_comb];
  assign p7_array_index_2050732_comb = p6_literal_2043914[p7_array_index_2050716_comb];
  assign p7_array_index_2050733_comb = p6_literal_2043916[p7_array_index_2050717_comb];
  assign p7_array_index_2050734_comb = p6_literal_2043918[p7_array_index_2050718_comb];
  assign p7_array_index_2050735_comb = p6_literal_2043920[p7_array_index_2050719_comb];
  assign p7_array_index_2050736_comb = p6_literal_2043896[p7_addedKey__60_comb[79:72]];
  assign p7_array_index_2050738_comb = p6_literal_2043896[p7_addedKey__60_comb[63:56]];
  assign p7_res7__896_comb = p7_array_index_2050730_comb ^ p7_array_index_2050731_comb ^ p7_array_index_2050732_comb ^ p7_array_index_2050733_comb ^ p7_array_index_2050734_comb ^ p7_array_index_2050735_comb ^ p7_array_index_2050736_comb ^ p6_literal_2043923[p7_array_index_2050721_comb] ^ p7_array_index_2050738_comb ^ p6_literal_2043920[p7_array_index_2050723_comb] ^ p6_literal_2043918[p7_array_index_2050724_comb] ^ p6_literal_2043916[p7_array_index_2050725_comb] ^ p6_literal_2043914[p7_array_index_2050726_comb] ^ p6_literal_2043912[p7_array_index_2050727_comb] ^ p6_literal_2043910[p7_array_index_2050728_comb] ^ p6_literal_2043896[p7_addedKey__60_comb[7:0]];
  assign p7_array_index_2050747_comb = p6_literal_2043910[p7_res7__896_comb];
  assign p7_array_index_2050748_comb = p6_literal_2043912[p7_array_index_2050714_comb];
  assign p7_array_index_2050749_comb = p6_literal_2043914[p7_array_index_2050715_comb];
  assign p7_array_index_2050750_comb = p6_literal_2043916[p7_array_index_2050716_comb];
  assign p7_array_index_2050751_comb = p6_literal_2043918[p7_array_index_2050717_comb];
  assign p7_array_index_2050752_comb = p6_literal_2043920[p7_array_index_2050718_comb];
  assign p7_res7__898_comb = p7_array_index_2050747_comb ^ p7_array_index_2050748_comb ^ p7_array_index_2050749_comb ^ p7_array_index_2050750_comb ^ p7_array_index_2050751_comb ^ p7_array_index_2050752_comb ^ p7_array_index_2050719_comb ^ p6_literal_2043923[p7_array_index_2050736_comb] ^ p7_array_index_2050721_comb ^ p6_literal_2043920[p7_array_index_2050738_comb] ^ p6_literal_2043918[p7_array_index_2050723_comb] ^ p6_literal_2043916[p7_array_index_2050724_comb] ^ p6_literal_2043914[p7_array_index_2050725_comb] ^ p6_literal_2043912[p7_array_index_2050726_comb] ^ p6_literal_2043910[p7_array_index_2050727_comb] ^ p7_array_index_2050728_comb;
  assign p7_array_index_2050762_comb = p6_literal_2043912[p7_res7__896_comb];
  assign p7_array_index_2050763_comb = p6_literal_2043914[p7_array_index_2050714_comb];
  assign p7_array_index_2050764_comb = p6_literal_2043916[p7_array_index_2050715_comb];
  assign p7_array_index_2050765_comb = p6_literal_2043918[p7_array_index_2050716_comb];
  assign p7_array_index_2050766_comb = p6_literal_2043920[p7_array_index_2050717_comb];
  assign p7_res7__900_comb = p6_literal_2043910[p7_res7__898_comb] ^ p7_array_index_2050762_comb ^ p7_array_index_2050763_comb ^ p7_array_index_2050764_comb ^ p7_array_index_2050765_comb ^ p7_array_index_2050766_comb ^ p7_array_index_2050718_comb ^ p6_literal_2043923[p7_array_index_2050719_comb] ^ p7_array_index_2050736_comb ^ p6_literal_2043920[p7_array_index_2050721_comb] ^ p6_literal_2043918[p7_array_index_2050738_comb] ^ p6_literal_2043916[p7_array_index_2050723_comb] ^ p6_literal_2043914[p7_array_index_2050724_comb] ^ p6_literal_2043912[p7_array_index_2050725_comb] ^ p6_literal_2043910[p7_array_index_2050726_comb] ^ p7_array_index_2050727_comb;
  assign p7_array_index_2050776_comb = p6_literal_2043912[p7_res7__898_comb];
  assign p7_array_index_2050777_comb = p6_literal_2043914[p7_res7__896_comb];
  assign p7_array_index_2050778_comb = p6_literal_2043916[p7_array_index_2050714_comb];
  assign p7_array_index_2050779_comb = p6_literal_2043918[p7_array_index_2050715_comb];
  assign p7_array_index_2050780_comb = p6_literal_2043920[p7_array_index_2050716_comb];
  assign p7_res7__902_comb = p6_literal_2043910[p7_res7__900_comb] ^ p7_array_index_2050776_comb ^ p7_array_index_2050777_comb ^ p7_array_index_2050778_comb ^ p7_array_index_2050779_comb ^ p7_array_index_2050780_comb ^ p7_array_index_2050717_comb ^ p6_literal_2043923[p7_array_index_2050718_comb] ^ p7_array_index_2050719_comb ^ p6_literal_2043920[p7_array_index_2050736_comb] ^ p6_literal_2043918[p7_array_index_2050721_comb] ^ p6_literal_2043916[p7_array_index_2050738_comb] ^ p6_literal_2043914[p7_array_index_2050723_comb] ^ p6_literal_2043912[p7_array_index_2050724_comb] ^ p6_literal_2043910[p7_array_index_2050725_comb] ^ p7_array_index_2050726_comb;
  assign p7_array_index_2050791_comb = p6_literal_2043914[p7_res7__898_comb];
  assign p7_array_index_2050792_comb = p6_literal_2043916[p7_res7__896_comb];
  assign p7_array_index_2050793_comb = p6_literal_2043918[p7_array_index_2050714_comb];
  assign p7_array_index_2050794_comb = p6_literal_2043920[p7_array_index_2050715_comb];
  assign p7_res7__904_comb = p6_literal_2043910[p7_res7__902_comb] ^ p6_literal_2043912[p7_res7__900_comb] ^ p7_array_index_2050791_comb ^ p7_array_index_2050792_comb ^ p7_array_index_2050793_comb ^ p7_array_index_2050794_comb ^ p7_array_index_2050716_comb ^ p6_literal_2043923[p7_array_index_2050717_comb] ^ p7_array_index_2050718_comb ^ p7_array_index_2050735_comb ^ p6_literal_2043918[p7_array_index_2050736_comb] ^ p6_literal_2043916[p7_array_index_2050721_comb] ^ p6_literal_2043914[p7_array_index_2050738_comb] ^ p6_literal_2043912[p7_array_index_2050723_comb] ^ p6_literal_2043910[p7_array_index_2050724_comb] ^ p7_array_index_2050725_comb;
  assign p7_array_index_2050804_comb = p6_literal_2043914[p7_res7__900_comb];
  assign p7_array_index_2050805_comb = p6_literal_2043916[p7_res7__898_comb];
  assign p7_array_index_2050806_comb = p6_literal_2043918[p7_res7__896_comb];
  assign p7_array_index_2050807_comb = p6_literal_2043920[p7_array_index_2050714_comb];
  assign p7_res7__906_comb = p6_literal_2043910[p7_res7__904_comb] ^ p6_literal_2043912[p7_res7__902_comb] ^ p7_array_index_2050804_comb ^ p7_array_index_2050805_comb ^ p7_array_index_2050806_comb ^ p7_array_index_2050807_comb ^ p7_array_index_2050715_comb ^ p6_literal_2043923[p7_array_index_2050716_comb] ^ p7_array_index_2050717_comb ^ p7_array_index_2050752_comb ^ p6_literal_2043918[p7_array_index_2050719_comb] ^ p6_literal_2043916[p7_array_index_2050736_comb] ^ p6_literal_2043914[p7_array_index_2050721_comb] ^ p6_literal_2043912[p7_array_index_2050738_comb] ^ p6_literal_2043910[p7_array_index_2050723_comb] ^ p7_array_index_2050724_comb;
  assign p7_array_index_2050818_comb = p6_literal_2043916[p7_res7__900_comb];
  assign p7_array_index_2050819_comb = p6_literal_2043918[p7_res7__898_comb];
  assign p7_array_index_2050820_comb = p6_literal_2043920[p7_res7__896_comb];
  assign p7_res7__908_comb = p6_literal_2043910[p7_res7__906_comb] ^ p6_literal_2043912[p7_res7__904_comb] ^ p6_literal_2043914[p7_res7__902_comb] ^ p7_array_index_2050818_comb ^ p7_array_index_2050819_comb ^ p7_array_index_2050820_comb ^ p7_array_index_2050714_comb ^ p6_literal_2043923[p7_array_index_2050715_comb] ^ p7_array_index_2050716_comb ^ p7_array_index_2050766_comb ^ p7_array_index_2050734_comb ^ p6_literal_2043916[p7_array_index_2050719_comb] ^ p6_literal_2043914[p7_array_index_2050736_comb] ^ p6_literal_2043912[p7_array_index_2050721_comb] ^ p6_literal_2043910[p7_array_index_2050738_comb] ^ p7_array_index_2050723_comb;
  assign p7_array_index_2050830_comb = p6_literal_2043916[p7_res7__902_comb];
  assign p7_array_index_2050831_comb = p6_literal_2043918[p7_res7__900_comb];
  assign p7_array_index_2050832_comb = p6_literal_2043920[p7_res7__898_comb];
  assign p7_res7__910_comb = p6_literal_2043910[p7_res7__908_comb] ^ p6_literal_2043912[p7_res7__906_comb] ^ p6_literal_2043914[p7_res7__904_comb] ^ p7_array_index_2050830_comb ^ p7_array_index_2050831_comb ^ p7_array_index_2050832_comb ^ p7_res7__896_comb ^ p6_literal_2043923[p7_array_index_2050714_comb] ^ p7_array_index_2050715_comb ^ p7_array_index_2050780_comb ^ p7_array_index_2050751_comb ^ p6_literal_2043916[p7_array_index_2050718_comb] ^ p6_literal_2043914[p7_array_index_2050719_comb] ^ p6_literal_2043912[p7_array_index_2050736_comb] ^ p6_literal_2043910[p7_array_index_2050721_comb] ^ p7_array_index_2050738_comb;
  assign p7_array_index_2050843_comb = p6_literal_2043918[p7_res7__902_comb];
  assign p7_array_index_2050844_comb = p6_literal_2043920[p7_res7__900_comb];
  assign p7_res7__912_comb = p6_literal_2043910[p7_res7__910_comb] ^ p6_literal_2043912[p7_res7__908_comb] ^ p6_literal_2043914[p7_res7__906_comb] ^ p6_literal_2043916[p7_res7__904_comb] ^ p7_array_index_2050843_comb ^ p7_array_index_2050844_comb ^ p7_res7__898_comb ^ p6_literal_2043923[p7_res7__896_comb] ^ p7_array_index_2050714_comb ^ p7_array_index_2050794_comb ^ p7_array_index_2050765_comb ^ p7_array_index_2050733_comb ^ p6_literal_2043914[p7_array_index_2050718_comb] ^ p6_literal_2043912[p7_array_index_2050719_comb] ^ p6_literal_2043910[p7_array_index_2050736_comb] ^ p7_array_index_2050721_comb;
  assign p7_array_index_2050854_comb = p6_literal_2043918[p7_res7__904_comb];
  assign p7_array_index_2050855_comb = p6_literal_2043920[p7_res7__902_comb];
  assign p7_res7__914_comb = p6_literal_2043910[p7_res7__912_comb] ^ p6_literal_2043912[p7_res7__910_comb] ^ p6_literal_2043914[p7_res7__908_comb] ^ p6_literal_2043916[p7_res7__906_comb] ^ p7_array_index_2050854_comb ^ p7_array_index_2050855_comb ^ p7_res7__900_comb ^ p6_literal_2043923[p7_res7__898_comb] ^ p7_res7__896_comb ^ p7_array_index_2050807_comb ^ p7_array_index_2050779_comb ^ p7_array_index_2050750_comb ^ p6_literal_2043914[p7_array_index_2050717_comb] ^ p6_literal_2043912[p7_array_index_2050718_comb] ^ p6_literal_2043910[p7_array_index_2050719_comb] ^ p7_array_index_2050736_comb;
  assign p7_array_index_2050866_comb = p6_literal_2043920[p7_res7__904_comb];
  assign p7_res7__916_comb = p6_literal_2043910[p7_res7__914_comb] ^ p6_literal_2043912[p7_res7__912_comb] ^ p6_literal_2043914[p7_res7__910_comb] ^ p6_literal_2043916[p7_res7__908_comb] ^ p6_literal_2043918[p7_res7__906_comb] ^ p7_array_index_2050866_comb ^ p7_res7__902_comb ^ p6_literal_2043923[p7_res7__900_comb] ^ p7_res7__898_comb ^ p7_array_index_2050820_comb ^ p7_array_index_2050793_comb ^ p7_array_index_2050764_comb ^ p7_array_index_2050732_comb ^ p6_literal_2043912[p7_array_index_2050717_comb] ^ p6_literal_2043910[p7_array_index_2050718_comb] ^ p7_array_index_2050719_comb;
  assign p7_array_index_2050876_comb = p6_literal_2043920[p7_res7__906_comb];
  assign p7_res7__918_comb = p6_literal_2043910[p7_res7__916_comb] ^ p6_literal_2043912[p7_res7__914_comb] ^ p6_literal_2043914[p7_res7__912_comb] ^ p6_literal_2043916[p7_res7__910_comb] ^ p6_literal_2043918[p7_res7__908_comb] ^ p7_array_index_2050876_comb ^ p7_res7__904_comb ^ p6_literal_2043923[p7_res7__902_comb] ^ p7_res7__900_comb ^ p7_array_index_2050832_comb ^ p7_array_index_2050806_comb ^ p7_array_index_2050778_comb ^ p7_array_index_2050749_comb ^ p6_literal_2043912[p7_array_index_2050716_comb] ^ p6_literal_2043910[p7_array_index_2050717_comb] ^ p7_array_index_2050718_comb;
  assign p7_res7__920_comb = p6_literal_2043910[p7_res7__918_comb] ^ p6_literal_2043912[p7_res7__916_comb] ^ p6_literal_2043914[p7_res7__914_comb] ^ p6_literal_2043916[p7_res7__912_comb] ^ p6_literal_2043918[p7_res7__910_comb] ^ p6_literal_2043920[p7_res7__908_comb] ^ p7_res7__906_comb ^ p6_literal_2043923[p7_res7__904_comb] ^ p7_res7__902_comb ^ p7_array_index_2050844_comb ^ p7_array_index_2050819_comb ^ p7_array_index_2050792_comb ^ p7_array_index_2050763_comb ^ p7_array_index_2050731_comb ^ p6_literal_2043910[p7_array_index_2050716_comb] ^ p7_array_index_2050717_comb;
  assign p7_res7__922_comb = p6_literal_2043910[p7_res7__920_comb] ^ p6_literal_2043912[p7_res7__918_comb] ^ p6_literal_2043914[p7_res7__916_comb] ^ p6_literal_2043916[p7_res7__914_comb] ^ p6_literal_2043918[p7_res7__912_comb] ^ p6_literal_2043920[p7_res7__910_comb] ^ p7_res7__908_comb ^ p6_literal_2043923[p7_res7__906_comb] ^ p7_res7__904_comb ^ p7_array_index_2050855_comb ^ p7_array_index_2050831_comb ^ p7_array_index_2050805_comb ^ p7_array_index_2050777_comb ^ p7_array_index_2050748_comb ^ p6_literal_2043910[p7_array_index_2050715_comb] ^ p7_array_index_2050716_comb;
  assign p7_res7__924_comb = p6_literal_2043910[p7_res7__922_comb] ^ p6_literal_2043912[p7_res7__920_comb] ^ p6_literal_2043914[p7_res7__918_comb] ^ p6_literal_2043916[p7_res7__916_comb] ^ p6_literal_2043918[p7_res7__914_comb] ^ p6_literal_2043920[p7_res7__912_comb] ^ p7_res7__910_comb ^ p6_literal_2043923[p7_res7__908_comb] ^ p7_res7__906_comb ^ p7_array_index_2050866_comb ^ p7_array_index_2050843_comb ^ p7_array_index_2050818_comb ^ p7_array_index_2050791_comb ^ p7_array_index_2050762_comb ^ p7_array_index_2050730_comb ^ p7_array_index_2050715_comb;
  assign p7_res7__926_comb = p6_literal_2043910[p7_res7__924_comb] ^ p6_literal_2043912[p7_res7__922_comb] ^ p6_literal_2043914[p7_res7__920_comb] ^ p6_literal_2043916[p7_res7__918_comb] ^ p6_literal_2043918[p7_res7__916_comb] ^ p6_literal_2043920[p7_res7__914_comb] ^ p7_res7__912_comb ^ p6_literal_2043923[p7_res7__910_comb] ^ p7_res7__908_comb ^ p7_array_index_2050876_comb ^ p7_array_index_2050854_comb ^ p7_array_index_2050830_comb ^ p7_array_index_2050804_comb ^ p7_array_index_2050776_comb ^ p7_array_index_2050747_comb ^ p7_array_index_2050714_comb;
  assign p7_res__28_comb = {p7_res7__926_comb, p7_res7__924_comb, p7_res7__922_comb, p7_res7__920_comb, p7_res7__918_comb, p7_res7__916_comb, p7_res7__914_comb, p7_res7__912_comb, p7_res7__910_comb, p7_res7__908_comb, p7_res7__906_comb, p7_res7__904_comb, p7_res7__902_comb, p7_res7__900_comb, p7_res7__898_comb, p7_res7__896_comb};
  assign p7_xor_2050916_comb = p7_res__28_comb ^ p7_xor_2050480_comb;
  assign p7_addedKey__61_comb = p7_xor_2050916_comb ^ 128'h7ea1_add5_427c_254e_391c_2823_e2a3_801e;
  assign p7_array_index_2050932_comb = p6_literal_2043896[p7_addedKey__61_comb[127:120]];
  assign p7_array_index_2050933_comb = p6_literal_2043896[p7_addedKey__61_comb[119:112]];
  assign p7_array_index_2050934_comb = p6_literal_2043896[p7_addedKey__61_comb[111:104]];
  assign p7_array_index_2050935_comb = p6_literal_2043896[p7_addedKey__61_comb[103:96]];
  assign p7_array_index_2050936_comb = p6_literal_2043896[p7_addedKey__61_comb[95:88]];
  assign p7_array_index_2050937_comb = p6_literal_2043896[p7_addedKey__61_comb[87:80]];
  assign p7_array_index_2050939_comb = p6_literal_2043896[p7_addedKey__61_comb[71:64]];
  assign p7_array_index_2050941_comb = p6_literal_2043896[p7_addedKey__61_comb[55:48]];
  assign p7_array_index_2050942_comb = p6_literal_2043896[p7_addedKey__61_comb[47:40]];
  assign p7_array_index_2050943_comb = p6_literal_2043896[p7_addedKey__61_comb[39:32]];
  assign p7_array_index_2050944_comb = p6_literal_2043896[p7_addedKey__61_comb[31:24]];
  assign p7_array_index_2050945_comb = p6_literal_2043896[p7_addedKey__61_comb[23:16]];
  assign p7_array_index_2050946_comb = p6_literal_2043896[p7_addedKey__61_comb[15:8]];
  assign p7_array_index_2050948_comb = p6_literal_2043910[p7_array_index_2050932_comb];
  assign p7_array_index_2050949_comb = p6_literal_2043912[p7_array_index_2050933_comb];
  assign p7_array_index_2050950_comb = p6_literal_2043914[p7_array_index_2050934_comb];
  assign p7_array_index_2050951_comb = p6_literal_2043916[p7_array_index_2050935_comb];
  assign p7_array_index_2050952_comb = p6_literal_2043918[p7_array_index_2050936_comb];
  assign p7_array_index_2050953_comb = p6_literal_2043920[p7_array_index_2050937_comb];
  assign p7_array_index_2050954_comb = p6_literal_2043896[p7_addedKey__61_comb[79:72]];
  assign p7_array_index_2050956_comb = p6_literal_2043896[p7_addedKey__61_comb[63:56]];
  assign p7_res7__928_comb = p7_array_index_2050948_comb ^ p7_array_index_2050949_comb ^ p7_array_index_2050950_comb ^ p7_array_index_2050951_comb ^ p7_array_index_2050952_comb ^ p7_array_index_2050953_comb ^ p7_array_index_2050954_comb ^ p6_literal_2043923[p7_array_index_2050939_comb] ^ p7_array_index_2050956_comb ^ p6_literal_2043920[p7_array_index_2050941_comb] ^ p6_literal_2043918[p7_array_index_2050942_comb] ^ p6_literal_2043916[p7_array_index_2050943_comb] ^ p6_literal_2043914[p7_array_index_2050944_comb] ^ p6_literal_2043912[p7_array_index_2050945_comb] ^ p6_literal_2043910[p7_array_index_2050946_comb] ^ p6_literal_2043896[p7_addedKey__61_comb[7:0]];
  assign p7_array_index_2050965_comb = p6_literal_2043910[p7_res7__928_comb];
  assign p7_array_index_2050966_comb = p6_literal_2043912[p7_array_index_2050932_comb];
  assign p7_array_index_2050967_comb = p6_literal_2043914[p7_array_index_2050933_comb];
  assign p7_array_index_2050968_comb = p6_literal_2043916[p7_array_index_2050934_comb];
  assign p7_array_index_2050969_comb = p6_literal_2043918[p7_array_index_2050935_comb];
  assign p7_array_index_2050970_comb = p6_literal_2043920[p7_array_index_2050936_comb];
  assign p7_res7__930_comb = p7_array_index_2050965_comb ^ p7_array_index_2050966_comb ^ p7_array_index_2050967_comb ^ p7_array_index_2050968_comb ^ p7_array_index_2050969_comb ^ p7_array_index_2050970_comb ^ p7_array_index_2050937_comb ^ p6_literal_2043923[p7_array_index_2050954_comb] ^ p7_array_index_2050939_comb ^ p6_literal_2043920[p7_array_index_2050956_comb] ^ p6_literal_2043918[p7_array_index_2050941_comb] ^ p6_literal_2043916[p7_array_index_2050942_comb] ^ p6_literal_2043914[p7_array_index_2050943_comb] ^ p6_literal_2043912[p7_array_index_2050944_comb] ^ p6_literal_2043910[p7_array_index_2050945_comb] ^ p7_array_index_2050946_comb;
  assign p7_array_index_2050980_comb = p6_literal_2043912[p7_res7__928_comb];
  assign p7_array_index_2050981_comb = p6_literal_2043914[p7_array_index_2050932_comb];
  assign p7_array_index_2050982_comb = p6_literal_2043916[p7_array_index_2050933_comb];
  assign p7_array_index_2050983_comb = p6_literal_2043918[p7_array_index_2050934_comb];
  assign p7_array_index_2050984_comb = p6_literal_2043920[p7_array_index_2050935_comb];
  assign p7_res7__932_comb = p6_literal_2043910[p7_res7__930_comb] ^ p7_array_index_2050980_comb ^ p7_array_index_2050981_comb ^ p7_array_index_2050982_comb ^ p7_array_index_2050983_comb ^ p7_array_index_2050984_comb ^ p7_array_index_2050936_comb ^ p6_literal_2043923[p7_array_index_2050937_comb] ^ p7_array_index_2050954_comb ^ p6_literal_2043920[p7_array_index_2050939_comb] ^ p6_literal_2043918[p7_array_index_2050956_comb] ^ p6_literal_2043916[p7_array_index_2050941_comb] ^ p6_literal_2043914[p7_array_index_2050942_comb] ^ p6_literal_2043912[p7_array_index_2050943_comb] ^ p6_literal_2043910[p7_array_index_2050944_comb] ^ p7_array_index_2050945_comb;
  assign p7_array_index_2050994_comb = p6_literal_2043912[p7_res7__930_comb];
  assign p7_array_index_2050995_comb = p6_literal_2043914[p7_res7__928_comb];
  assign p7_array_index_2050996_comb = p6_literal_2043916[p7_array_index_2050932_comb];
  assign p7_array_index_2050997_comb = p6_literal_2043918[p7_array_index_2050933_comb];
  assign p7_array_index_2050998_comb = p6_literal_2043920[p7_array_index_2050934_comb];
  assign p7_res7__934_comb = p6_literal_2043910[p7_res7__932_comb] ^ p7_array_index_2050994_comb ^ p7_array_index_2050995_comb ^ p7_array_index_2050996_comb ^ p7_array_index_2050997_comb ^ p7_array_index_2050998_comb ^ p7_array_index_2050935_comb ^ p6_literal_2043923[p7_array_index_2050936_comb] ^ p7_array_index_2050937_comb ^ p6_literal_2043920[p7_array_index_2050954_comb] ^ p6_literal_2043918[p7_array_index_2050939_comb] ^ p6_literal_2043916[p7_array_index_2050956_comb] ^ p6_literal_2043914[p7_array_index_2050941_comb] ^ p6_literal_2043912[p7_array_index_2050942_comb] ^ p6_literal_2043910[p7_array_index_2050943_comb] ^ p7_array_index_2050944_comb;
  assign p7_array_index_2051009_comb = p6_literal_2043914[p7_res7__930_comb];
  assign p7_array_index_2051010_comb = p6_literal_2043916[p7_res7__928_comb];
  assign p7_array_index_2051011_comb = p6_literal_2043918[p7_array_index_2050932_comb];
  assign p7_array_index_2051012_comb = p6_literal_2043920[p7_array_index_2050933_comb];
  assign p7_res7__936_comb = p6_literal_2043910[p7_res7__934_comb] ^ p6_literal_2043912[p7_res7__932_comb] ^ p7_array_index_2051009_comb ^ p7_array_index_2051010_comb ^ p7_array_index_2051011_comb ^ p7_array_index_2051012_comb ^ p7_array_index_2050934_comb ^ p6_literal_2043923[p7_array_index_2050935_comb] ^ p7_array_index_2050936_comb ^ p7_array_index_2050953_comb ^ p6_literal_2043918[p7_array_index_2050954_comb] ^ p6_literal_2043916[p7_array_index_2050939_comb] ^ p6_literal_2043914[p7_array_index_2050956_comb] ^ p6_literal_2043912[p7_array_index_2050941_comb] ^ p6_literal_2043910[p7_array_index_2050942_comb] ^ p7_array_index_2050943_comb;
  assign p7_array_index_2051022_comb = p6_literal_2043914[p7_res7__932_comb];
  assign p7_array_index_2051023_comb = p6_literal_2043916[p7_res7__930_comb];
  assign p7_array_index_2051024_comb = p6_literal_2043918[p7_res7__928_comb];
  assign p7_array_index_2051025_comb = p6_literal_2043920[p7_array_index_2050932_comb];
  assign p7_res7__938_comb = p6_literal_2043910[p7_res7__936_comb] ^ p6_literal_2043912[p7_res7__934_comb] ^ p7_array_index_2051022_comb ^ p7_array_index_2051023_comb ^ p7_array_index_2051024_comb ^ p7_array_index_2051025_comb ^ p7_array_index_2050933_comb ^ p6_literal_2043923[p7_array_index_2050934_comb] ^ p7_array_index_2050935_comb ^ p7_array_index_2050970_comb ^ p6_literal_2043918[p7_array_index_2050937_comb] ^ p6_literal_2043916[p7_array_index_2050954_comb] ^ p6_literal_2043914[p7_array_index_2050939_comb] ^ p6_literal_2043912[p7_array_index_2050956_comb] ^ p6_literal_2043910[p7_array_index_2050941_comb] ^ p7_array_index_2050942_comb;
  assign p7_array_index_2051036_comb = p6_literal_2043916[p7_res7__932_comb];
  assign p7_array_index_2051037_comb = p6_literal_2043918[p7_res7__930_comb];
  assign p7_array_index_2051038_comb = p6_literal_2043920[p7_res7__928_comb];
  assign p7_res7__940_comb = p6_literal_2043910[p7_res7__938_comb] ^ p6_literal_2043912[p7_res7__936_comb] ^ p6_literal_2043914[p7_res7__934_comb] ^ p7_array_index_2051036_comb ^ p7_array_index_2051037_comb ^ p7_array_index_2051038_comb ^ p7_array_index_2050932_comb ^ p6_literal_2043923[p7_array_index_2050933_comb] ^ p7_array_index_2050934_comb ^ p7_array_index_2050984_comb ^ p7_array_index_2050952_comb ^ p6_literal_2043916[p7_array_index_2050937_comb] ^ p6_literal_2043914[p7_array_index_2050954_comb] ^ p6_literal_2043912[p7_array_index_2050939_comb] ^ p6_literal_2043910[p7_array_index_2050956_comb] ^ p7_array_index_2050941_comb;
  assign p7_array_index_2051048_comb = p6_literal_2043916[p7_res7__934_comb];
  assign p7_array_index_2051049_comb = p6_literal_2043918[p7_res7__932_comb];
  assign p7_array_index_2051050_comb = p6_literal_2043920[p7_res7__930_comb];
  assign p7_res7__942_comb = p6_literal_2043910[p7_res7__940_comb] ^ p6_literal_2043912[p7_res7__938_comb] ^ p6_literal_2043914[p7_res7__936_comb] ^ p7_array_index_2051048_comb ^ p7_array_index_2051049_comb ^ p7_array_index_2051050_comb ^ p7_res7__928_comb ^ p6_literal_2043923[p7_array_index_2050932_comb] ^ p7_array_index_2050933_comb ^ p7_array_index_2050998_comb ^ p7_array_index_2050969_comb ^ p6_literal_2043916[p7_array_index_2050936_comb] ^ p6_literal_2043914[p7_array_index_2050937_comb] ^ p6_literal_2043912[p7_array_index_2050954_comb] ^ p6_literal_2043910[p7_array_index_2050939_comb] ^ p7_array_index_2050956_comb;
  assign p7_array_index_2051061_comb = p6_literal_2043918[p7_res7__934_comb];
  assign p7_array_index_2051062_comb = p6_literal_2043920[p7_res7__932_comb];
  assign p7_res7__944_comb = p6_literal_2043910[p7_res7__942_comb] ^ p6_literal_2043912[p7_res7__940_comb] ^ p6_literal_2043914[p7_res7__938_comb] ^ p6_literal_2043916[p7_res7__936_comb] ^ p7_array_index_2051061_comb ^ p7_array_index_2051062_comb ^ p7_res7__930_comb ^ p6_literal_2043923[p7_res7__928_comb] ^ p7_array_index_2050932_comb ^ p7_array_index_2051012_comb ^ p7_array_index_2050983_comb ^ p7_array_index_2050951_comb ^ p6_literal_2043914[p7_array_index_2050936_comb] ^ p6_literal_2043912[p7_array_index_2050937_comb] ^ p6_literal_2043910[p7_array_index_2050954_comb] ^ p7_array_index_2050939_comb;
  assign p7_array_index_2051072_comb = p6_literal_2043918[p7_res7__936_comb];
  assign p7_array_index_2051073_comb = p6_literal_2043920[p7_res7__934_comb];
  assign p7_res7__946_comb = p6_literal_2043910[p7_res7__944_comb] ^ p6_literal_2043912[p7_res7__942_comb] ^ p6_literal_2043914[p7_res7__940_comb] ^ p6_literal_2043916[p7_res7__938_comb] ^ p7_array_index_2051072_comb ^ p7_array_index_2051073_comb ^ p7_res7__932_comb ^ p6_literal_2043923[p7_res7__930_comb] ^ p7_res7__928_comb ^ p7_array_index_2051025_comb ^ p7_array_index_2050997_comb ^ p7_array_index_2050968_comb ^ p6_literal_2043914[p7_array_index_2050935_comb] ^ p6_literal_2043912[p7_array_index_2050936_comb] ^ p6_literal_2043910[p7_array_index_2050937_comb] ^ p7_array_index_2050954_comb;
  assign p7_array_index_2051084_comb = p6_literal_2043920[p7_res7__936_comb];
  assign p7_res7__948_comb = p6_literal_2043910[p7_res7__946_comb] ^ p6_literal_2043912[p7_res7__944_comb] ^ p6_literal_2043914[p7_res7__942_comb] ^ p6_literal_2043916[p7_res7__940_comb] ^ p6_literal_2043918[p7_res7__938_comb] ^ p7_array_index_2051084_comb ^ p7_res7__934_comb ^ p6_literal_2043923[p7_res7__932_comb] ^ p7_res7__930_comb ^ p7_array_index_2051038_comb ^ p7_array_index_2051011_comb ^ p7_array_index_2050982_comb ^ p7_array_index_2050950_comb ^ p6_literal_2043912[p7_array_index_2050935_comb] ^ p6_literal_2043910[p7_array_index_2050936_comb] ^ p7_array_index_2050937_comb;
  assign p7_array_index_2051094_comb = p6_literal_2043920[p7_res7__938_comb];
  assign p7_res7__950_comb = p6_literal_2043910[p7_res7__948_comb] ^ p6_literal_2043912[p7_res7__946_comb] ^ p6_literal_2043914[p7_res7__944_comb] ^ p6_literal_2043916[p7_res7__942_comb] ^ p6_literal_2043918[p7_res7__940_comb] ^ p7_array_index_2051094_comb ^ p7_res7__936_comb ^ p6_literal_2043923[p7_res7__934_comb] ^ p7_res7__932_comb ^ p7_array_index_2051050_comb ^ p7_array_index_2051024_comb ^ p7_array_index_2050996_comb ^ p7_array_index_2050967_comb ^ p6_literal_2043912[p7_array_index_2050934_comb] ^ p6_literal_2043910[p7_array_index_2050935_comb] ^ p7_array_index_2050936_comb;
  assign p7_res7__952_comb = p6_literal_2043910[p7_res7__950_comb] ^ p6_literal_2043912[p7_res7__948_comb] ^ p6_literal_2043914[p7_res7__946_comb] ^ p6_literal_2043916[p7_res7__944_comb] ^ p6_literal_2043918[p7_res7__942_comb] ^ p6_literal_2043920[p7_res7__940_comb] ^ p7_res7__938_comb ^ p6_literal_2043923[p7_res7__936_comb] ^ p7_res7__934_comb ^ p7_array_index_2051062_comb ^ p7_array_index_2051037_comb ^ p7_array_index_2051010_comb ^ p7_array_index_2050981_comb ^ p7_array_index_2050949_comb ^ p6_literal_2043910[p7_array_index_2050934_comb] ^ p7_array_index_2050935_comb;
  assign p7_res7__954_comb = p6_literal_2043910[p7_res7__952_comb] ^ p6_literal_2043912[p7_res7__950_comb] ^ p6_literal_2043914[p7_res7__948_comb] ^ p6_literal_2043916[p7_res7__946_comb] ^ p6_literal_2043918[p7_res7__944_comb] ^ p6_literal_2043920[p7_res7__942_comb] ^ p7_res7__940_comb ^ p6_literal_2043923[p7_res7__938_comb] ^ p7_res7__936_comb ^ p7_array_index_2051073_comb ^ p7_array_index_2051049_comb ^ p7_array_index_2051023_comb ^ p7_array_index_2050995_comb ^ p7_array_index_2050966_comb ^ p6_literal_2043910[p7_array_index_2050933_comb] ^ p7_array_index_2050934_comb;
  assign p7_res7__956_comb = p6_literal_2043910[p7_res7__954_comb] ^ p6_literal_2043912[p7_res7__952_comb] ^ p6_literal_2043914[p7_res7__950_comb] ^ p6_literal_2043916[p7_res7__948_comb] ^ p6_literal_2043918[p7_res7__946_comb] ^ p6_literal_2043920[p7_res7__944_comb] ^ p7_res7__942_comb ^ p6_literal_2043923[p7_res7__940_comb] ^ p7_res7__938_comb ^ p7_array_index_2051084_comb ^ p7_array_index_2051061_comb ^ p7_array_index_2051036_comb ^ p7_array_index_2051009_comb ^ p7_array_index_2050980_comb ^ p7_array_index_2050948_comb ^ p7_array_index_2050933_comb;
  assign p7_res7__958_comb = p6_literal_2043910[p7_res7__956_comb] ^ p6_literal_2043912[p7_res7__954_comb] ^ p6_literal_2043914[p7_res7__952_comb] ^ p6_literal_2043916[p7_res7__950_comb] ^ p6_literal_2043918[p7_res7__948_comb] ^ p6_literal_2043920[p7_res7__946_comb] ^ p7_res7__944_comb ^ p6_literal_2043923[p7_res7__942_comb] ^ p7_res7__940_comb ^ p7_array_index_2051094_comb ^ p7_array_index_2051072_comb ^ p7_array_index_2051048_comb ^ p7_array_index_2051022_comb ^ p7_array_index_2050994_comb ^ p7_array_index_2050965_comb ^ p7_array_index_2050932_comb;
  assign p7_res__29_comb = {p7_res7__958_comb, p7_res7__956_comb, p7_res7__954_comb, p7_res7__952_comb, p7_res7__950_comb, p7_res7__948_comb, p7_res7__946_comb, p7_res7__944_comb, p7_res7__942_comb, p7_res7__940_comb, p7_res7__938_comb, p7_res7__936_comb, p7_res7__934_comb, p7_res7__932_comb, p7_res7__930_comb, p7_res7__928_comb};
  assign p7_xor_2051134_comb = p7_res__29_comb ^ p7_xor_2050698_comb;
  assign p7_addedKey__62_comb = p7_xor_2051134_comb ^ 128'h1003_dba7_2e34_5ff6_643b_9533_3f27_141f;
  assign p7_array_index_2051150_comb = p6_literal_2043896[p7_addedKey__62_comb[127:120]];
  assign p7_array_index_2051151_comb = p6_literal_2043896[p7_addedKey__62_comb[119:112]];
  assign p7_array_index_2051152_comb = p6_literal_2043896[p7_addedKey__62_comb[111:104]];
  assign p7_array_index_2051153_comb = p6_literal_2043896[p7_addedKey__62_comb[103:96]];
  assign p7_array_index_2051154_comb = p6_literal_2043896[p7_addedKey__62_comb[95:88]];
  assign p7_array_index_2051155_comb = p6_literal_2043896[p7_addedKey__62_comb[87:80]];
  assign p7_array_index_2051157_comb = p6_literal_2043896[p7_addedKey__62_comb[71:64]];
  assign p7_array_index_2051159_comb = p6_literal_2043896[p7_addedKey__62_comb[55:48]];
  assign p7_array_index_2051160_comb = p6_literal_2043896[p7_addedKey__62_comb[47:40]];
  assign p7_array_index_2051161_comb = p6_literal_2043896[p7_addedKey__62_comb[39:32]];
  assign p7_array_index_2051162_comb = p6_literal_2043896[p7_addedKey__62_comb[31:24]];
  assign p7_array_index_2051163_comb = p6_literal_2043896[p7_addedKey__62_comb[23:16]];
  assign p7_array_index_2051164_comb = p6_literal_2043896[p7_addedKey__62_comb[15:8]];
  assign p7_array_index_2051166_comb = p6_literal_2043910[p7_array_index_2051150_comb];
  assign p7_array_index_2051167_comb = p6_literal_2043912[p7_array_index_2051151_comb];
  assign p7_array_index_2051168_comb = p6_literal_2043914[p7_array_index_2051152_comb];
  assign p7_array_index_2051169_comb = p6_literal_2043916[p7_array_index_2051153_comb];
  assign p7_array_index_2051170_comb = p6_literal_2043918[p7_array_index_2051154_comb];
  assign p7_array_index_2051171_comb = p6_literal_2043920[p7_array_index_2051155_comb];
  assign p7_array_index_2051172_comb = p6_literal_2043896[p7_addedKey__62_comb[79:72]];
  assign p7_array_index_2051174_comb = p6_literal_2043896[p7_addedKey__62_comb[63:56]];
  assign p7_res7__960_comb = p7_array_index_2051166_comb ^ p7_array_index_2051167_comb ^ p7_array_index_2051168_comb ^ p7_array_index_2051169_comb ^ p7_array_index_2051170_comb ^ p7_array_index_2051171_comb ^ p7_array_index_2051172_comb ^ p6_literal_2043923[p7_array_index_2051157_comb] ^ p7_array_index_2051174_comb ^ p6_literal_2043920[p7_array_index_2051159_comb] ^ p6_literal_2043918[p7_array_index_2051160_comb] ^ p6_literal_2043916[p7_array_index_2051161_comb] ^ p6_literal_2043914[p7_array_index_2051162_comb] ^ p6_literal_2043912[p7_array_index_2051163_comb] ^ p6_literal_2043910[p7_array_index_2051164_comb] ^ p6_literal_2043896[p7_addedKey__62_comb[7:0]];
  assign p7_array_index_2051183_comb = p6_literal_2043910[p7_res7__960_comb];
  assign p7_array_index_2051184_comb = p6_literal_2043912[p7_array_index_2051150_comb];
  assign p7_array_index_2051185_comb = p6_literal_2043914[p7_array_index_2051151_comb];
  assign p7_array_index_2051186_comb = p6_literal_2043916[p7_array_index_2051152_comb];
  assign p7_array_index_2051187_comb = p6_literal_2043918[p7_array_index_2051153_comb];
  assign p7_array_index_2051188_comb = p6_literal_2043920[p7_array_index_2051154_comb];
  assign p7_res7__962_comb = p7_array_index_2051183_comb ^ p7_array_index_2051184_comb ^ p7_array_index_2051185_comb ^ p7_array_index_2051186_comb ^ p7_array_index_2051187_comb ^ p7_array_index_2051188_comb ^ p7_array_index_2051155_comb ^ p6_literal_2043923[p7_array_index_2051172_comb] ^ p7_array_index_2051157_comb ^ p6_literal_2043920[p7_array_index_2051174_comb] ^ p6_literal_2043918[p7_array_index_2051159_comb] ^ p6_literal_2043916[p7_array_index_2051160_comb] ^ p6_literal_2043914[p7_array_index_2051161_comb] ^ p6_literal_2043912[p7_array_index_2051162_comb] ^ p6_literal_2043910[p7_array_index_2051163_comb] ^ p7_array_index_2051164_comb;
  assign p7_array_index_2051198_comb = p6_literal_2043912[p7_res7__960_comb];
  assign p7_array_index_2051199_comb = p6_literal_2043914[p7_array_index_2051150_comb];
  assign p7_array_index_2051200_comb = p6_literal_2043916[p7_array_index_2051151_comb];
  assign p7_array_index_2051201_comb = p6_literal_2043918[p7_array_index_2051152_comb];
  assign p7_array_index_2051202_comb = p6_literal_2043920[p7_array_index_2051153_comb];
  assign p7_res7__964_comb = p6_literal_2043910[p7_res7__962_comb] ^ p7_array_index_2051198_comb ^ p7_array_index_2051199_comb ^ p7_array_index_2051200_comb ^ p7_array_index_2051201_comb ^ p7_array_index_2051202_comb ^ p7_array_index_2051154_comb ^ p6_literal_2043923[p7_array_index_2051155_comb] ^ p7_array_index_2051172_comb ^ p6_literal_2043920[p7_array_index_2051157_comb] ^ p6_literal_2043918[p7_array_index_2051174_comb] ^ p6_literal_2043916[p7_array_index_2051159_comb] ^ p6_literal_2043914[p7_array_index_2051160_comb] ^ p6_literal_2043912[p7_array_index_2051161_comb] ^ p6_literal_2043910[p7_array_index_2051162_comb] ^ p7_array_index_2051163_comb;
  assign p7_array_index_2051212_comb = p6_literal_2043912[p7_res7__962_comb];
  assign p7_array_index_2051213_comb = p6_literal_2043914[p7_res7__960_comb];
  assign p7_array_index_2051214_comb = p6_literal_2043916[p7_array_index_2051150_comb];
  assign p7_array_index_2051215_comb = p6_literal_2043918[p7_array_index_2051151_comb];
  assign p7_array_index_2051216_comb = p6_literal_2043920[p7_array_index_2051152_comb];
  assign p7_res7__966_comb = p6_literal_2043910[p7_res7__964_comb] ^ p7_array_index_2051212_comb ^ p7_array_index_2051213_comb ^ p7_array_index_2051214_comb ^ p7_array_index_2051215_comb ^ p7_array_index_2051216_comb ^ p7_array_index_2051153_comb ^ p6_literal_2043923[p7_array_index_2051154_comb] ^ p7_array_index_2051155_comb ^ p6_literal_2043920[p7_array_index_2051172_comb] ^ p6_literal_2043918[p7_array_index_2051157_comb] ^ p6_literal_2043916[p7_array_index_2051174_comb] ^ p6_literal_2043914[p7_array_index_2051159_comb] ^ p6_literal_2043912[p7_array_index_2051160_comb] ^ p6_literal_2043910[p7_array_index_2051161_comb] ^ p7_array_index_2051162_comb;
  assign p7_array_index_2051227_comb = p6_literal_2043914[p7_res7__962_comb];
  assign p7_array_index_2051228_comb = p6_literal_2043916[p7_res7__960_comb];
  assign p7_array_index_2051229_comb = p6_literal_2043918[p7_array_index_2051150_comb];
  assign p7_array_index_2051230_comb = p6_literal_2043920[p7_array_index_2051151_comb];
  assign p7_res7__968_comb = p6_literal_2043910[p7_res7__966_comb] ^ p6_literal_2043912[p7_res7__964_comb] ^ p7_array_index_2051227_comb ^ p7_array_index_2051228_comb ^ p7_array_index_2051229_comb ^ p7_array_index_2051230_comb ^ p7_array_index_2051152_comb ^ p6_literal_2043923[p7_array_index_2051153_comb] ^ p7_array_index_2051154_comb ^ p7_array_index_2051171_comb ^ p6_literal_2043918[p7_array_index_2051172_comb] ^ p6_literal_2043916[p7_array_index_2051157_comb] ^ p6_literal_2043914[p7_array_index_2051174_comb] ^ p6_literal_2043912[p7_array_index_2051159_comb] ^ p6_literal_2043910[p7_array_index_2051160_comb] ^ p7_array_index_2051161_comb;
  assign p7_array_index_2051240_comb = p6_literal_2043914[p7_res7__964_comb];
  assign p7_array_index_2051241_comb = p6_literal_2043916[p7_res7__962_comb];
  assign p7_array_index_2051242_comb = p6_literal_2043918[p7_res7__960_comb];
  assign p7_array_index_2051243_comb = p6_literal_2043920[p7_array_index_2051150_comb];
  assign p7_res7__970_comb = p6_literal_2043910[p7_res7__968_comb] ^ p6_literal_2043912[p7_res7__966_comb] ^ p7_array_index_2051240_comb ^ p7_array_index_2051241_comb ^ p7_array_index_2051242_comb ^ p7_array_index_2051243_comb ^ p7_array_index_2051151_comb ^ p6_literal_2043923[p7_array_index_2051152_comb] ^ p7_array_index_2051153_comb ^ p7_array_index_2051188_comb ^ p6_literal_2043918[p7_array_index_2051155_comb] ^ p6_literal_2043916[p7_array_index_2051172_comb] ^ p6_literal_2043914[p7_array_index_2051157_comb] ^ p6_literal_2043912[p7_array_index_2051174_comb] ^ p6_literal_2043910[p7_array_index_2051159_comb] ^ p7_array_index_2051160_comb;
  assign p7_array_index_2051254_comb = p6_literal_2043916[p7_res7__964_comb];
  assign p7_array_index_2051255_comb = p6_literal_2043918[p7_res7__962_comb];
  assign p7_array_index_2051256_comb = p6_literal_2043920[p7_res7__960_comb];
  assign p7_res7__972_comb = p6_literal_2043910[p7_res7__970_comb] ^ p6_literal_2043912[p7_res7__968_comb] ^ p6_literal_2043914[p7_res7__966_comb] ^ p7_array_index_2051254_comb ^ p7_array_index_2051255_comb ^ p7_array_index_2051256_comb ^ p7_array_index_2051150_comb ^ p6_literal_2043923[p7_array_index_2051151_comb] ^ p7_array_index_2051152_comb ^ p7_array_index_2051202_comb ^ p7_array_index_2051170_comb ^ p6_literal_2043916[p7_array_index_2051155_comb] ^ p6_literal_2043914[p7_array_index_2051172_comb] ^ p6_literal_2043912[p7_array_index_2051157_comb] ^ p6_literal_2043910[p7_array_index_2051174_comb] ^ p7_array_index_2051159_comb;
  assign p7_array_index_2051266_comb = p6_literal_2043916[p7_res7__966_comb];
  assign p7_array_index_2051267_comb = p6_literal_2043918[p7_res7__964_comb];
  assign p7_array_index_2051268_comb = p6_literal_2043920[p7_res7__962_comb];
  assign p7_res7__974_comb = p6_literal_2043910[p7_res7__972_comb] ^ p6_literal_2043912[p7_res7__970_comb] ^ p6_literal_2043914[p7_res7__968_comb] ^ p7_array_index_2051266_comb ^ p7_array_index_2051267_comb ^ p7_array_index_2051268_comb ^ p7_res7__960_comb ^ p6_literal_2043923[p7_array_index_2051150_comb] ^ p7_array_index_2051151_comb ^ p7_array_index_2051216_comb ^ p7_array_index_2051187_comb ^ p6_literal_2043916[p7_array_index_2051154_comb] ^ p6_literal_2043914[p7_array_index_2051155_comb] ^ p6_literal_2043912[p7_array_index_2051172_comb] ^ p6_literal_2043910[p7_array_index_2051157_comb] ^ p7_array_index_2051174_comb;
  assign p7_array_index_2051279_comb = p6_literal_2043918[p7_res7__966_comb];
  assign p7_array_index_2051280_comb = p6_literal_2043920[p7_res7__964_comb];
  assign p7_res7__976_comb = p6_literal_2043910[p7_res7__974_comb] ^ p6_literal_2043912[p7_res7__972_comb] ^ p6_literal_2043914[p7_res7__970_comb] ^ p6_literal_2043916[p7_res7__968_comb] ^ p7_array_index_2051279_comb ^ p7_array_index_2051280_comb ^ p7_res7__962_comb ^ p6_literal_2043923[p7_res7__960_comb] ^ p7_array_index_2051150_comb ^ p7_array_index_2051230_comb ^ p7_array_index_2051201_comb ^ p7_array_index_2051169_comb ^ p6_literal_2043914[p7_array_index_2051154_comb] ^ p6_literal_2043912[p7_array_index_2051155_comb] ^ p6_literal_2043910[p7_array_index_2051172_comb] ^ p7_array_index_2051157_comb;
  assign p7_array_index_2051290_comb = p6_literal_2043918[p7_res7__968_comb];
  assign p7_array_index_2051291_comb = p6_literal_2043920[p7_res7__966_comb];
  assign p7_res7__978_comb = p6_literal_2043910[p7_res7__976_comb] ^ p6_literal_2043912[p7_res7__974_comb] ^ p6_literal_2043914[p7_res7__972_comb] ^ p6_literal_2043916[p7_res7__970_comb] ^ p7_array_index_2051290_comb ^ p7_array_index_2051291_comb ^ p7_res7__964_comb ^ p6_literal_2043923[p7_res7__962_comb] ^ p7_res7__960_comb ^ p7_array_index_2051243_comb ^ p7_array_index_2051215_comb ^ p7_array_index_2051186_comb ^ p6_literal_2043914[p7_array_index_2051153_comb] ^ p6_literal_2043912[p7_array_index_2051154_comb] ^ p6_literal_2043910[p7_array_index_2051155_comb] ^ p7_array_index_2051172_comb;
  assign p7_array_index_2051302_comb = p6_literal_2043920[p7_res7__968_comb];
  assign p7_res7__980_comb = p6_literal_2043910[p7_res7__978_comb] ^ p6_literal_2043912[p7_res7__976_comb] ^ p6_literal_2043914[p7_res7__974_comb] ^ p6_literal_2043916[p7_res7__972_comb] ^ p6_literal_2043918[p7_res7__970_comb] ^ p7_array_index_2051302_comb ^ p7_res7__966_comb ^ p6_literal_2043923[p7_res7__964_comb] ^ p7_res7__962_comb ^ p7_array_index_2051256_comb ^ p7_array_index_2051229_comb ^ p7_array_index_2051200_comb ^ p7_array_index_2051168_comb ^ p6_literal_2043912[p7_array_index_2051153_comb] ^ p6_literal_2043910[p7_array_index_2051154_comb] ^ p7_array_index_2051155_comb;
  assign p7_array_index_2051312_comb = p6_literal_2043920[p7_res7__970_comb];
  assign p7_res7__982_comb = p6_literal_2043910[p7_res7__980_comb] ^ p6_literal_2043912[p7_res7__978_comb] ^ p6_literal_2043914[p7_res7__976_comb] ^ p6_literal_2043916[p7_res7__974_comb] ^ p6_literal_2043918[p7_res7__972_comb] ^ p7_array_index_2051312_comb ^ p7_res7__968_comb ^ p6_literal_2043923[p7_res7__966_comb] ^ p7_res7__964_comb ^ p7_array_index_2051268_comb ^ p7_array_index_2051242_comb ^ p7_array_index_2051214_comb ^ p7_array_index_2051185_comb ^ p6_literal_2043912[p7_array_index_2051152_comb] ^ p6_literal_2043910[p7_array_index_2051153_comb] ^ p7_array_index_2051154_comb;
  assign p7_res7__984_comb = p6_literal_2043910[p7_res7__982_comb] ^ p6_literal_2043912[p7_res7__980_comb] ^ p6_literal_2043914[p7_res7__978_comb] ^ p6_literal_2043916[p7_res7__976_comb] ^ p6_literal_2043918[p7_res7__974_comb] ^ p6_literal_2043920[p7_res7__972_comb] ^ p7_res7__970_comb ^ p6_literal_2043923[p7_res7__968_comb] ^ p7_res7__966_comb ^ p7_array_index_2051280_comb ^ p7_array_index_2051255_comb ^ p7_array_index_2051228_comb ^ p7_array_index_2051199_comb ^ p7_array_index_2051167_comb ^ p6_literal_2043910[p7_array_index_2051152_comb] ^ p7_array_index_2051153_comb;
  assign p7_res7__986_comb = p6_literal_2043910[p7_res7__984_comb] ^ p6_literal_2043912[p7_res7__982_comb] ^ p6_literal_2043914[p7_res7__980_comb] ^ p6_literal_2043916[p7_res7__978_comb] ^ p6_literal_2043918[p7_res7__976_comb] ^ p6_literal_2043920[p7_res7__974_comb] ^ p7_res7__972_comb ^ p6_literal_2043923[p7_res7__970_comb] ^ p7_res7__968_comb ^ p7_array_index_2051291_comb ^ p7_array_index_2051267_comb ^ p7_array_index_2051241_comb ^ p7_array_index_2051213_comb ^ p7_array_index_2051184_comb ^ p6_literal_2043910[p7_array_index_2051151_comb] ^ p7_array_index_2051152_comb;
  assign p7_res7__988_comb = p6_literal_2043910[p7_res7__986_comb] ^ p6_literal_2043912[p7_res7__984_comb] ^ p6_literal_2043914[p7_res7__982_comb] ^ p6_literal_2043916[p7_res7__980_comb] ^ p6_literal_2043918[p7_res7__978_comb] ^ p6_literal_2043920[p7_res7__976_comb] ^ p7_res7__974_comb ^ p6_literal_2043923[p7_res7__972_comb] ^ p7_res7__970_comb ^ p7_array_index_2051302_comb ^ p7_array_index_2051279_comb ^ p7_array_index_2051254_comb ^ p7_array_index_2051227_comb ^ p7_array_index_2051198_comb ^ p7_array_index_2051166_comb ^ p7_array_index_2051151_comb;
  assign p7_res7__990_comb = p6_literal_2043910[p7_res7__988_comb] ^ p6_literal_2043912[p7_res7__986_comb] ^ p6_literal_2043914[p7_res7__984_comb] ^ p6_literal_2043916[p7_res7__982_comb] ^ p6_literal_2043918[p7_res7__980_comb] ^ p6_literal_2043920[p7_res7__978_comb] ^ p7_res7__976_comb ^ p6_literal_2043923[p7_res7__974_comb] ^ p7_res7__972_comb ^ p7_array_index_2051312_comb ^ p7_array_index_2051290_comb ^ p7_array_index_2051266_comb ^ p7_array_index_2051240_comb ^ p7_array_index_2051212_comb ^ p7_array_index_2051183_comb ^ p7_array_index_2051150_comb;
  assign p7_res__30_comb = {p7_res7__990_comb, p7_res7__988_comb, p7_res7__986_comb, p7_res7__984_comb, p7_res7__982_comb, p7_res7__980_comb, p7_res7__978_comb, p7_res7__976_comb, p7_res7__974_comb, p7_res7__972_comb, p7_res7__970_comb, p7_res7__968_comb, p7_res7__966_comb, p7_res7__964_comb, p7_res7__962_comb, p7_res7__960_comb};
  assign p7_k9_comb = p7_res__30_comb ^ p7_xor_2050916_comb;
  assign p7_xor_2051355_comb = p6_encoded ^ p7_k9_comb;
  assign p7_addedKey__63_comb = p7_k9_comb ^ 128'h5ea7_d858_1e14_9b61_f16a_c145_9ced_a820;
  assign p7_bit_slice_2051370_comb = p7_xor_2051355_comb[111:104];
  assign p7_bit_slice_2051371_comb = p7_xor_2051355_comb[103:96];
  assign p7_bit_slice_2051372_comb = p7_xor_2051355_comb[95:88];
  assign p7_bit_slice_2051373_comb = p7_xor_2051355_comb[87:80];
  assign p7_bit_slice_2051374_comb = p7_xor_2051355_comb[79:72];
  assign p7_bit_slice_2051375_comb = p7_xor_2051355_comb[63:56];
  assign p7_bit_slice_2051376_comb = p7_xor_2051355_comb[47:40];
  assign p7_bit_slice_2051377_comb = p7_xor_2051355_comb[39:32];
  assign p7_bit_slice_2051378_comb = p7_xor_2051355_comb[31:24];
  assign p7_bit_slice_2051379_comb = p7_xor_2051355_comb[23:16];
  assign p7_bit_slice_2051380_comb = p7_xor_2051355_comb[15:8];
  assign p7_bit_slice_2051381_comb = p7_xor_2051355_comb[7:0];
  assign p7_bit_slice_2051404_comb = p7_xor_2051355_comb[71:64];
  assign p7_bit_slice_2051406_comb = p7_xor_2051355_comb[55:48];
  assign p7_array_index_2051407_comb = p6_literal_2043920[p7_bit_slice_2051376_comb];
  assign p7_array_index_2051408_comb = p6_literal_2043918[p7_bit_slice_2051377_comb];
  assign p7_array_index_2051409_comb = p6_literal_2043916[p7_bit_slice_2051378_comb];
  assign p7_array_index_2051410_comb = p6_literal_2043914[p7_bit_slice_2051379_comb];
  assign p7_array_index_2051411_comb = p6_literal_2043912[p7_bit_slice_2051380_comb];
  assign p7_array_index_2051412_comb = p6_literal_2043910[p7_bit_slice_2051381_comb];
  assign p7_array_index_2051382_comb = p6_literal_2043896[p7_addedKey__63_comb[127:120]];
  assign p7_array_index_2051383_comb = p6_literal_2043896[p7_addedKey__63_comb[119:112]];
  assign p7_array_index_2051384_comb = p6_literal_2043896[p7_addedKey__63_comb[111:104]];
  assign p7_array_index_2051385_comb = p6_literal_2043896[p7_addedKey__63_comb[103:96]];
  assign p7_array_index_2051386_comb = p6_literal_2043896[p7_addedKey__63_comb[95:88]];
  assign p7_array_index_2051387_comb = p6_literal_2043896[p7_addedKey__63_comb[87:80]];
  assign p7_array_index_2051389_comb = p6_literal_2043896[p7_addedKey__63_comb[71:64]];
  assign p7_array_index_2051391_comb = p6_literal_2043896[p7_addedKey__63_comb[55:48]];
  assign p7_array_index_2051392_comb = p6_literal_2043896[p7_addedKey__63_comb[47:40]];
  assign p7_array_index_2051393_comb = p6_literal_2043896[p7_addedKey__63_comb[39:32]];
  assign p7_array_index_2051394_comb = p6_literal_2043896[p7_addedKey__63_comb[31:24]];
  assign p7_array_index_2051395_comb = p6_literal_2043896[p7_addedKey__63_comb[23:16]];
  assign p7_array_index_2051396_comb = p6_literal_2043896[p7_addedKey__63_comb[15:8]];
  assign p7_res7__1025_comb = p6_literal_2043910[p7_xor_2051355_comb[119:112]] ^ p6_literal_2043912[p7_bit_slice_2051370_comb] ^ p6_literal_2043914[p7_bit_slice_2051371_comb] ^ p6_literal_2043916[p7_bit_slice_2051372_comb] ^ p6_literal_2043918[p7_bit_slice_2051373_comb] ^ p6_literal_2043920[p7_bit_slice_2051374_comb] ^ p7_bit_slice_2051404_comb ^ p6_literal_2043923[p7_bit_slice_2051375_comb] ^ p7_bit_slice_2051406_comb ^ p7_array_index_2051407_comb ^ p7_array_index_2051408_comb ^ p7_array_index_2051409_comb ^ p7_array_index_2051410_comb ^ p7_array_index_2051411_comb ^ p7_array_index_2051412_comb ^ p7_xor_2051355_comb[127:120];
  assign p7_array_index_2051414_comb = p6_literal_2043910[p7_array_index_2051382_comb];
  assign p7_array_index_2051415_comb = p6_literal_2043912[p7_array_index_2051383_comb];
  assign p7_array_index_2051416_comb = p6_literal_2043914[p7_array_index_2051384_comb];
  assign p7_array_index_2051417_comb = p6_literal_2043916[p7_array_index_2051385_comb];
  assign p7_array_index_2051418_comb = p6_literal_2043918[p7_array_index_2051386_comb];
  assign p7_array_index_2051419_comb = p6_literal_2043920[p7_array_index_2051387_comb];
  assign p7_array_index_2051420_comb = p6_literal_2043896[p7_addedKey__63_comb[79:72]];
  assign p7_array_index_2051422_comb = p6_literal_2043896[p7_addedKey__63_comb[63:56]];
  assign p7_array_index_2051439_comb = p6_literal_2043920[p7_bit_slice_2051377_comb];
  assign p7_array_index_2051440_comb = p6_literal_2043918[p7_bit_slice_2051378_comb];
  assign p7_array_index_2051441_comb = p6_literal_2043916[p7_bit_slice_2051379_comb];
  assign p7_array_index_2051442_comb = p6_literal_2043914[p7_bit_slice_2051380_comb];
  assign p7_array_index_2051443_comb = p6_literal_2043912[p7_bit_slice_2051381_comb];
  assign p7_array_index_2051444_comb = p6_literal_2043910[p7_res7__1025_comb];
  assign p7_res7__992_comb = p7_array_index_2051414_comb ^ p7_array_index_2051415_comb ^ p7_array_index_2051416_comb ^ p7_array_index_2051417_comb ^ p7_array_index_2051418_comb ^ p7_array_index_2051419_comb ^ p7_array_index_2051420_comb ^ p6_literal_2043923[p7_array_index_2051389_comb] ^ p7_array_index_2051422_comb ^ p6_literal_2043920[p7_array_index_2051391_comb] ^ p6_literal_2043918[p7_array_index_2051392_comb] ^ p6_literal_2043916[p7_array_index_2051393_comb] ^ p6_literal_2043914[p7_array_index_2051394_comb] ^ p6_literal_2043912[p7_array_index_2051395_comb] ^ p6_literal_2043910[p7_array_index_2051396_comb] ^ p6_literal_2043896[p7_addedKey__63_comb[7:0]];
  assign p7_res7__1027_comb = p6_literal_2043910[p7_bit_slice_2051370_comb] ^ p6_literal_2043912[p7_bit_slice_2051371_comb] ^ p6_literal_2043914[p7_bit_slice_2051372_comb] ^ p6_literal_2043916[p7_bit_slice_2051373_comb] ^ p6_literal_2043918[p7_bit_slice_2051374_comb] ^ p6_literal_2043920[p7_bit_slice_2051404_comb] ^ p7_bit_slice_2051375_comb ^ p6_literal_2043923[p7_bit_slice_2051406_comb] ^ p7_bit_slice_2051376_comb ^ p7_array_index_2051439_comb ^ p7_array_index_2051440_comb ^ p7_array_index_2051441_comb ^ p7_array_index_2051442_comb ^ p7_array_index_2051443_comb ^ p7_array_index_2051444_comb ^ p7_xor_2051355_comb[119:112];

  // Registers for pipe stage 7:
  reg [127:0] p7_bit_slice_2043893;
  reg [127:0] p7_bit_slice_2044119;
  reg [127:0] p7_k3;
  reg [127:0] p7_k2;
  reg [127:0] p7_k5;
  reg [127:0] p7_k4;
  reg [127:0] p7_k7;
  reg [127:0] p7_k6;
  reg [127:0] p7_xor_2051134;
  reg [7:0] p7_bit_slice_2051370;
  reg [7:0] p7_bit_slice_2051371;
  reg [7:0] p7_bit_slice_2051372;
  reg [7:0] p7_bit_slice_2051373;
  reg [7:0] p7_bit_slice_2051374;
  reg [7:0] p7_bit_slice_2051375;
  reg [7:0] p7_bit_slice_2051376;
  reg [7:0] p7_bit_slice_2051377;
  reg [7:0] p7_bit_slice_2051378;
  reg [7:0] p7_bit_slice_2051379;
  reg [7:0] p7_bit_slice_2051380;
  reg [7:0] p7_bit_slice_2051381;
  reg [7:0] p7_array_index_2051382;
  reg [7:0] p7_array_index_2051383;
  reg [7:0] p7_array_index_2051384;
  reg [7:0] p7_array_index_2051385;
  reg [7:0] p7_array_index_2051386;
  reg [7:0] p7_array_index_2051387;
  reg [7:0] p7_array_index_2051389;
  reg [7:0] p7_array_index_2051391;
  reg [7:0] p7_array_index_2051392;
  reg [7:0] p7_array_index_2051393;
  reg [7:0] p7_array_index_2051394;
  reg [7:0] p7_array_index_2051395;
  reg [7:0] p7_array_index_2051396;
  reg [7:0] p7_bit_slice_2051404;
  reg [7:0] p7_bit_slice_2051406;
  reg [7:0] p7_array_index_2051407;
  reg [7:0] p7_array_index_2051408;
  reg [7:0] p7_array_index_2051409;
  reg [7:0] p7_array_index_2051410;
  reg [7:0] p7_array_index_2051411;
  reg [7:0] p7_array_index_2051412;
  reg [7:0] p7_array_index_2051414;
  reg [7:0] p7_array_index_2051415;
  reg [7:0] p7_array_index_2051416;
  reg [7:0] p7_array_index_2051417;
  reg [7:0] p7_array_index_2051418;
  reg [7:0] p7_array_index_2051419;
  reg [7:0] p7_array_index_2051420;
  reg [7:0] p7_array_index_2051422;
  reg [7:0] p7_res7__1025;
  reg [7:0] p7_res7__992;
  reg [7:0] p7_array_index_2051439;
  reg [7:0] p7_array_index_2051440;
  reg [7:0] p7_array_index_2051441;
  reg [7:0] p7_array_index_2051442;
  reg [7:0] p7_array_index_2051443;
  reg [7:0] p7_array_index_2051444;
  reg [7:0] p7_res7__1027;
  reg [7:0] p8_literal_2043910[256];
  reg [7:0] p8_literal_2043912[256];
  reg [7:0] p8_literal_2043914[256];
  reg [7:0] p8_literal_2043916[256];
  reg [7:0] p8_literal_2043918[256];
  reg [7:0] p8_literal_2043920[256];
  reg [7:0] p8_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p7_bit_slice_2043893 <= p6_bit_slice_2043893;
    p7_bit_slice_2044119 <= p6_bit_slice_2044119;
    p7_k3 <= p6_k3;
    p7_k2 <= p6_k2;
    p7_k5 <= p6_k5;
    p7_k4 <= p6_k4;
    p7_k7 <= p6_k7;
    p7_k6 <= p6_k6;
    p7_xor_2051134 <= p7_xor_2051134_comb;
    p7_bit_slice_2051370 <= p7_bit_slice_2051370_comb;
    p7_bit_slice_2051371 <= p7_bit_slice_2051371_comb;
    p7_bit_slice_2051372 <= p7_bit_slice_2051372_comb;
    p7_bit_slice_2051373 <= p7_bit_slice_2051373_comb;
    p7_bit_slice_2051374 <= p7_bit_slice_2051374_comb;
    p7_bit_slice_2051375 <= p7_bit_slice_2051375_comb;
    p7_bit_slice_2051376 <= p7_bit_slice_2051376_comb;
    p7_bit_slice_2051377 <= p7_bit_slice_2051377_comb;
    p7_bit_slice_2051378 <= p7_bit_slice_2051378_comb;
    p7_bit_slice_2051379 <= p7_bit_slice_2051379_comb;
    p7_bit_slice_2051380 <= p7_bit_slice_2051380_comb;
    p7_bit_slice_2051381 <= p7_bit_slice_2051381_comb;
    p7_array_index_2051382 <= p7_array_index_2051382_comb;
    p7_array_index_2051383 <= p7_array_index_2051383_comb;
    p7_array_index_2051384 <= p7_array_index_2051384_comb;
    p7_array_index_2051385 <= p7_array_index_2051385_comb;
    p7_array_index_2051386 <= p7_array_index_2051386_comb;
    p7_array_index_2051387 <= p7_array_index_2051387_comb;
    p7_array_index_2051389 <= p7_array_index_2051389_comb;
    p7_array_index_2051391 <= p7_array_index_2051391_comb;
    p7_array_index_2051392 <= p7_array_index_2051392_comb;
    p7_array_index_2051393 <= p7_array_index_2051393_comb;
    p7_array_index_2051394 <= p7_array_index_2051394_comb;
    p7_array_index_2051395 <= p7_array_index_2051395_comb;
    p7_array_index_2051396 <= p7_array_index_2051396_comb;
    p7_bit_slice_2051404 <= p7_bit_slice_2051404_comb;
    p7_bit_slice_2051406 <= p7_bit_slice_2051406_comb;
    p7_array_index_2051407 <= p7_array_index_2051407_comb;
    p7_array_index_2051408 <= p7_array_index_2051408_comb;
    p7_array_index_2051409 <= p7_array_index_2051409_comb;
    p7_array_index_2051410 <= p7_array_index_2051410_comb;
    p7_array_index_2051411 <= p7_array_index_2051411_comb;
    p7_array_index_2051412 <= p7_array_index_2051412_comb;
    p7_array_index_2051414 <= p7_array_index_2051414_comb;
    p7_array_index_2051415 <= p7_array_index_2051415_comb;
    p7_array_index_2051416 <= p7_array_index_2051416_comb;
    p7_array_index_2051417 <= p7_array_index_2051417_comb;
    p7_array_index_2051418 <= p7_array_index_2051418_comb;
    p7_array_index_2051419 <= p7_array_index_2051419_comb;
    p7_array_index_2051420 <= p7_array_index_2051420_comb;
    p7_array_index_2051422 <= p7_array_index_2051422_comb;
    p7_res7__1025 <= p7_res7__1025_comb;
    p7_res7__992 <= p7_res7__992_comb;
    p7_array_index_2051439 <= p7_array_index_2051439_comb;
    p7_array_index_2051440 <= p7_array_index_2051440_comb;
    p7_array_index_2051441 <= p7_array_index_2051441_comb;
    p7_array_index_2051442 <= p7_array_index_2051442_comb;
    p7_array_index_2051443 <= p7_array_index_2051443_comb;
    p7_array_index_2051444 <= p7_array_index_2051444_comb;
    p7_res7__1027 <= p7_res7__1027_comb;
    p8_literal_2043910 <= p7_literal_2043910;
    p8_literal_2043912 <= p7_literal_2043912;
    p8_literal_2043914 <= p7_literal_2043914;
    p8_literal_2043916 <= p7_literal_2043916;
    p8_literal_2043918 <= p7_literal_2043918;
    p8_literal_2043920 <= p7_literal_2043920;
    p8_literal_2043923 <= p7_literal_2043923;
  end

  // ===== Pipe stage 8:
  wire [7:0] p8_array_index_2051578_comb;
  wire [7:0] p8_array_index_2051579_comb;
  wire [7:0] p8_array_index_2051580_comb;
  wire [7:0] p8_array_index_2051581_comb;
  wire [7:0] p8_array_index_2051582_comb;
  wire [7:0] p8_array_index_2051583_comb;
  wire [7:0] p8_res7__994_comb;
  wire [7:0] p8_array_index_2051599_comb;
  wire [7:0] p8_array_index_2051600_comb;
  wire [7:0] p8_array_index_2051601_comb;
  wire [7:0] p8_array_index_2051602_comb;
  wire [7:0] p8_array_index_2051603_comb;
  wire [7:0] p8_array_index_2051606_comb;
  wire [7:0] p8_array_index_2051607_comb;
  wire [7:0] p8_array_index_2051608_comb;
  wire [7:0] p8_array_index_2051609_comb;
  wire [7:0] p8_array_index_2051610_comb;
  wire [7:0] p8_res7__1029_comb;
  wire [7:0] p8_res7__996_comb;
  wire [7:0] p8_array_index_2051627_comb;
  wire [7:0] p8_array_index_2051628_comb;
  wire [7:0] p8_array_index_2051629_comb;
  wire [7:0] p8_array_index_2051630_comb;
  wire [7:0] p8_array_index_2051631_comb;
  wire [7:0] p8_array_index_2051634_comb;
  wire [7:0] p8_array_index_2051635_comb;
  wire [7:0] p8_array_index_2051636_comb;
  wire [7:0] p8_array_index_2051637_comb;
  wire [7:0] p8_array_index_2051638_comb;
  wire [7:0] p8_res7__1031_comb;
  wire [7:0] p8_res7__998_comb;
  wire [7:0] p8_array_index_2051654_comb;
  wire [7:0] p8_array_index_2051655_comb;
  wire [7:0] p8_array_index_2051656_comb;
  wire [7:0] p8_array_index_2051657_comb;
  wire [7:0] p8_array_index_2051662_comb;
  wire [7:0] p8_array_index_2051663_comb;
  wire [7:0] p8_array_index_2051664_comb;
  wire [7:0] p8_array_index_2051665_comb;
  wire [7:0] p8_res7__1033_comb;
  wire [7:0] p8_res7__1000_comb;
  wire [7:0] p8_array_index_2051680_comb;
  wire [7:0] p8_array_index_2051681_comb;
  wire [7:0] p8_array_index_2051682_comb;
  wire [7:0] p8_array_index_2051683_comb;
  wire [7:0] p8_array_index_2051688_comb;
  wire [7:0] p8_array_index_2051689_comb;
  wire [7:0] p8_array_index_2051690_comb;
  wire [7:0] p8_array_index_2051691_comb;
  wire [7:0] p8_res7__1035_comb;
  wire [7:0] p8_res7__1002_comb;
  wire [7:0] p8_array_index_2051705_comb;
  wire [7:0] p8_array_index_2051706_comb;
  wire [7:0] p8_array_index_2051707_comb;
  wire [7:0] p8_array_index_2051714_comb;
  wire [7:0] p8_array_index_2051715_comb;
  wire [7:0] p8_array_index_2051716_comb;
  wire [7:0] p8_res7__1037_comb;
  wire [7:0] p8_res7__1004_comb;
  wire [7:0] p8_array_index_2051729_comb;
  wire [7:0] p8_array_index_2051730_comb;
  wire [7:0] p8_array_index_2051731_comb;
  wire [7:0] p8_array_index_2051738_comb;
  wire [7:0] p8_array_index_2051739_comb;
  wire [7:0] p8_array_index_2051740_comb;
  wire [7:0] p8_res7__1039_comb;
  wire [7:0] p8_res7__1006_comb;
  wire [7:0] p8_array_index_2051752_comb;
  wire [7:0] p8_array_index_2051753_comb;
  wire [7:0] p8_array_index_2051762_comb;
  wire [7:0] p8_array_index_2051763_comb;
  wire [7:0] p8_res7__1041_comb;
  wire [7:0] p8_res7__1008_comb;
  wire [7:0] p8_array_index_2051774_comb;
  wire [7:0] p8_array_index_2051775_comb;
  wire [7:0] p8_array_index_2051784_comb;
  wire [7:0] p8_array_index_2051785_comb;
  wire [7:0] p8_res7__1043_comb;
  wire [7:0] p8_res7__1010_comb;
  wire [7:0] p8_array_index_2051795_comb;
  wire [7:0] p8_array_index_2051806_comb;
  wire [7:0] p8_res7__1045_comb;
  wire [7:0] p8_res7__1012_comb;
  wire [7:0] p8_array_index_2051815_comb;
  wire [7:0] p8_array_index_2051826_comb;
  wire [7:0] p8_res7__1047_comb;
  wire [7:0] p8_res7__1014_comb;
  wire [7:0] p8_res7__1049_comb;
  wire [7:0] p8_res7__1016_comb;
  wire [7:0] p8_res7__1051_comb;
  wire [7:0] p8_res7__1018_comb;
  wire [7:0] p8_res7__1053_comb;
  wire [7:0] p8_res7__1020_comb;
  wire [7:0] p8_res7__1055_comb;
  wire [7:0] p8_res7__1022_comb;
  wire [127:0] p8_res__31_comb;
  wire [127:0] p8_permut__32_comb;
  wire [127:0] p8_xor_2051919_comb;
  wire [7:0] p8_array_index_2051942_comb;
  wire [7:0] p8_array_index_2051943_comb;
  wire [7:0] p8_array_index_2051944_comb;
  wire [7:0] p8_array_index_2051945_comb;
  wire [7:0] p8_array_index_2051946_comb;
  wire [7:0] p8_array_index_2051947_comb;
  wire [7:0] p8_res7__1057_comb;
  wire [7:0] p8_array_index_2051957_comb;
  wire [7:0] p8_array_index_2051958_comb;
  wire [7:0] p8_array_index_2051959_comb;
  wire [7:0] p8_array_index_2051960_comb;
  wire [7:0] p8_array_index_2051961_comb;
  wire [7:0] p8_array_index_2051962_comb;
  wire [7:0] p8_res7__1059_comb;
  wire [7:0] p8_array_index_2051971_comb;
  wire [7:0] p8_array_index_2051972_comb;
  wire [7:0] p8_array_index_2051973_comb;
  wire [7:0] p8_array_index_2051974_comb;
  wire [7:0] p8_array_index_2051975_comb;
  wire [7:0] p8_res7__1061_comb;
  wire [7:0] p8_array_index_2051985_comb;
  wire [7:0] p8_array_index_2051986_comb;
  wire [7:0] p8_array_index_2051987_comb;
  wire [7:0] p8_array_index_2051988_comb;
  wire [7:0] p8_array_index_2051989_comb;
  wire [7:0] p8_res7__1063_comb;
  wire [7:0] p8_array_index_2051998_comb;
  wire [7:0] p8_array_index_2051999_comb;
  wire [7:0] p8_array_index_2052000_comb;
  wire [7:0] p8_array_index_2052001_comb;
  wire [7:0] p8_res7__1065_comb;
  wire [7:0] p8_array_index_2052011_comb;
  wire [7:0] p8_array_index_2052012_comb;
  wire [7:0] p8_array_index_2052013_comb;
  wire [7:0] p8_array_index_2052014_comb;
  wire [7:0] p8_res7__1067_comb;
  wire [7:0] p8_array_index_2052023_comb;
  wire [7:0] p8_array_index_2052024_comb;
  wire [7:0] p8_array_index_2052025_comb;
  wire [7:0] p8_res7__1069_comb;
  wire [7:0] p8_array_index_2052035_comb;
  wire [7:0] p8_array_index_2052036_comb;
  wire [7:0] p8_array_index_2052037_comb;
  wire [7:0] p8_res7__1071_comb;
  wire [7:0] p8_array_index_2052046_comb;
  wire [7:0] p8_array_index_2052047_comb;
  wire [7:0] p8_res7__1073_comb;
  wire [7:0] p8_array_index_2052057_comb;
  wire [7:0] p8_array_index_2052058_comb;
  wire [7:0] p8_res7__1075_comb;
  wire [7:0] p8_array_index_2052067_comb;
  wire [7:0] p8_res7__1077_comb;
  wire [7:0] p8_array_index_2052077_comb;
  wire [7:0] p8_res7__1079_comb;
  wire [7:0] p8_res7__1081_comb;
  wire [7:0] p8_res7__1083_comb;
  wire [7:0] p8_res7__1085_comb;
  wire [7:0] p8_res7__1087_comb;
  wire [127:0] p8_permut__33_comb;
  wire [127:0] p8_xor_2052135_comb;
  wire [7:0] p8_array_index_2052158_comb;
  wire [7:0] p8_array_index_2052159_comb;
  wire [7:0] p8_array_index_2052160_comb;
  wire [7:0] p8_array_index_2052161_comb;
  wire [7:0] p8_array_index_2052162_comb;
  wire [7:0] p8_array_index_2052163_comb;
  wire [7:0] p8_res7__1089_comb;
  wire [7:0] p8_array_index_2052173_comb;
  wire [7:0] p8_array_index_2052174_comb;
  wire [7:0] p8_array_index_2052175_comb;
  wire [7:0] p8_array_index_2052176_comb;
  wire [7:0] p8_array_index_2052177_comb;
  wire [7:0] p8_array_index_2052178_comb;
  wire [7:0] p8_res7__1091_comb;
  wire [7:0] p8_array_index_2052187_comb;
  wire [7:0] p8_array_index_2052188_comb;
  wire [7:0] p8_array_index_2052189_comb;
  wire [7:0] p8_array_index_2052190_comb;
  wire [7:0] p8_array_index_2052191_comb;
  wire [7:0] p8_res7__1093_comb;
  wire [7:0] p8_array_index_2052201_comb;
  wire [7:0] p8_array_index_2052202_comb;
  wire [7:0] p8_array_index_2052203_comb;
  wire [7:0] p8_array_index_2052204_comb;
  wire [7:0] p8_array_index_2052205_comb;
  wire [7:0] p8_res7__1095_comb;
  wire [7:0] p8_array_index_2052214_comb;
  wire [7:0] p8_array_index_2052215_comb;
  wire [7:0] p8_array_index_2052216_comb;
  wire [7:0] p8_array_index_2052217_comb;
  wire [7:0] p8_res7__1097_comb;
  wire [7:0] p8_array_index_2052227_comb;
  wire [7:0] p8_array_index_2052228_comb;
  wire [7:0] p8_array_index_2052229_comb;
  wire [7:0] p8_array_index_2052230_comb;
  wire [7:0] p8_res7__1099_comb;
  wire [7:0] p8_array_index_2052239_comb;
  wire [7:0] p8_array_index_2052240_comb;
  wire [7:0] p8_array_index_2052241_comb;
  wire [7:0] p8_res7__1101_comb;
  wire [7:0] p8_array_index_2052251_comb;
  wire [7:0] p8_array_index_2052252_comb;
  wire [7:0] p8_array_index_2052253_comb;
  wire [7:0] p8_res7__1103_comb;
  wire [7:0] p8_array_index_2052262_comb;
  wire [7:0] p8_array_index_2052263_comb;
  wire [7:0] p8_res7__1105_comb;
  wire [7:0] p8_array_index_2052273_comb;
  wire [7:0] p8_array_index_2052274_comb;
  wire [7:0] p8_res7__1107_comb;
  wire [7:0] p8_array_index_2052283_comb;
  wire [7:0] p8_res7__1109_comb;
  wire [7:0] p8_array_index_2052293_comb;
  wire [7:0] p8_res7__1111_comb;
  wire [7:0] p8_res7__1113_comb;
  wire [7:0] p8_res7__1115_comb;
  wire [7:0] p8_res7__1117_comb;
  wire [7:0] p8_res7__1119_comb;
  wire [127:0] p8_permut__34_comb;
  wire [127:0] p8_xor_2052351_comb;
  wire [7:0] p8_array_index_2052374_comb;
  wire [7:0] p8_array_index_2052375_comb;
  wire [7:0] p8_array_index_2052376_comb;
  wire [7:0] p8_array_index_2052377_comb;
  wire [7:0] p8_array_index_2052378_comb;
  wire [7:0] p8_array_index_2052379_comb;
  wire [7:0] p8_res7__1121_comb;
  wire [7:0] p8_array_index_2052389_comb;
  wire [7:0] p8_array_index_2052390_comb;
  wire [7:0] p8_array_index_2052391_comb;
  wire [7:0] p8_array_index_2052392_comb;
  wire [7:0] p8_array_index_2052393_comb;
  wire [7:0] p8_array_index_2052394_comb;
  wire [7:0] p8_res7__1123_comb;
  wire [7:0] p8_array_index_2052403_comb;
  wire [7:0] p8_array_index_2052404_comb;
  wire [7:0] p8_array_index_2052405_comb;
  wire [7:0] p8_array_index_2052406_comb;
  wire [7:0] p8_array_index_2052407_comb;
  wire [7:0] p8_res7__1125_comb;
  wire [7:0] p8_array_index_2052417_comb;
  wire [7:0] p8_array_index_2052418_comb;
  wire [7:0] p8_array_index_2052419_comb;
  wire [7:0] p8_array_index_2052420_comb;
  wire [7:0] p8_array_index_2052421_comb;
  wire [7:0] p8_res7__1127_comb;
  wire [7:0] p8_array_index_2052430_comb;
  wire [7:0] p8_array_index_2052431_comb;
  wire [7:0] p8_array_index_2052432_comb;
  wire [7:0] p8_array_index_2052433_comb;
  wire [7:0] p8_res7__1129_comb;
  wire [7:0] p8_array_index_2052443_comb;
  wire [7:0] p8_array_index_2052444_comb;
  wire [7:0] p8_array_index_2052445_comb;
  wire [7:0] p8_array_index_2052446_comb;
  wire [7:0] p8_res7__1131_comb;
  wire [7:0] p8_array_index_2052455_comb;
  wire [7:0] p8_array_index_2052456_comb;
  wire [7:0] p8_array_index_2052457_comb;
  wire [7:0] p8_res7__1133_comb;
  wire [7:0] p8_array_index_2052467_comb;
  wire [7:0] p8_array_index_2052468_comb;
  wire [7:0] p8_array_index_2052469_comb;
  wire [7:0] p8_res7__1135_comb;
  wire [7:0] p8_array_index_2052478_comb;
  wire [7:0] p8_array_index_2052479_comb;
  wire [7:0] p8_res7__1137_comb;
  wire [7:0] p8_array_index_2052489_comb;
  wire [7:0] p8_array_index_2052490_comb;
  wire [7:0] p8_res7__1139_comb;
  wire [7:0] p8_array_index_2052499_comb;
  wire [7:0] p8_res7__1141_comb;
  wire [7:0] p8_array_index_2052509_comb;
  wire [7:0] p8_res7__1143_comb;
  wire [7:0] p8_res7__1145_comb;
  wire [7:0] p8_res7__1147_comb;
  wire [7:0] p8_res7__1149_comb;
  wire [7:0] p8_res7__1151_comb;
  wire [127:0] p8_permut__35_comb;
  wire [127:0] p8_xor_2052567_comb;
  wire [7:0] p8_bit_slice_2052575_comb;
  wire [7:0] p8_bit_slice_2052576_comb;
  wire [7:0] p8_bit_slice_2052577_comb;
  wire [7:0] p8_bit_slice_2052578_comb;
  wire [7:0] p8_bit_slice_2052579_comb;
  wire [7:0] p8_bit_slice_2052580_comb;
  wire [7:0] p8_bit_slice_2052589_comb;
  wire [7:0] p8_array_index_2052590_comb;
  wire [7:0] p8_array_index_2052591_comb;
  wire [7:0] p8_array_index_2052592_comb;
  wire [7:0] p8_array_index_2052593_comb;
  wire [7:0] p8_array_index_2052594_comb;
  wire [7:0] p8_array_index_2052595_comb;
  wire [7:0] p8_res7__1153_comb;
  wire [7:0] p8_array_index_2052605_comb;
  wire [7:0] p8_array_index_2052606_comb;
  wire [7:0] p8_array_index_2052607_comb;
  wire [7:0] p8_array_index_2052608_comb;
  wire [7:0] p8_array_index_2052609_comb;
  wire [7:0] p8_array_index_2052610_comb;
  wire [7:0] p8_res7__1155_comb;
  wire [7:0] p8_array_index_2052619_comb;
  wire [7:0] p8_array_index_2052620_comb;
  wire [7:0] p8_array_index_2052621_comb;
  wire [7:0] p8_array_index_2052622_comb;
  wire [7:0] p8_array_index_2052623_comb;
  wire [7:0] p8_res7__1157_comb;
  wire [7:0] p8_array_index_2052633_comb;
  wire [7:0] p8_array_index_2052634_comb;
  wire [7:0] p8_array_index_2052635_comb;
  wire [7:0] p8_array_index_2052636_comb;
  wire [7:0] p8_array_index_2052637_comb;
  wire [7:0] p8_res7__1159_comb;
  wire [7:0] p8_array_index_2052646_comb;
  wire [7:0] p8_array_index_2052647_comb;
  wire [7:0] p8_array_index_2052648_comb;
  wire [7:0] p8_array_index_2052649_comb;
  wire [7:0] p8_res7__1161_comb;
  wire [7:0] p8_array_index_2052659_comb;
  wire [7:0] p8_array_index_2052660_comb;
  wire [7:0] p8_array_index_2052661_comb;
  wire [7:0] p8_array_index_2052662_comb;
  wire [7:0] p8_res7__1163_comb;
  wire [7:0] p8_array_index_2052671_comb;
  wire [7:0] p8_array_index_2052672_comb;
  wire [7:0] p8_array_index_2052673_comb;
  wire [7:0] p8_res7__1165_comb;
  wire [7:0] p8_array_index_2052683_comb;
  wire [7:0] p8_array_index_2052684_comb;
  wire [7:0] p8_array_index_2052685_comb;
  wire [7:0] p8_res7__1167_comb;
  wire [7:0] p8_array_index_2052694_comb;
  wire [7:0] p8_array_index_2052695_comb;
  wire [7:0] p8_res7__1169_comb;
  assign p8_array_index_2051578_comb = p7_literal_2043910[p7_res7__992];
  assign p8_array_index_2051579_comb = p7_literal_2043912[p7_array_index_2051382];
  assign p8_array_index_2051580_comb = p7_literal_2043914[p7_array_index_2051383];
  assign p8_array_index_2051581_comb = p7_literal_2043916[p7_array_index_2051384];
  assign p8_array_index_2051582_comb = p7_literal_2043918[p7_array_index_2051385];
  assign p8_array_index_2051583_comb = p7_literal_2043920[p7_array_index_2051386];
  assign p8_res7__994_comb = p8_array_index_2051578_comb ^ p8_array_index_2051579_comb ^ p8_array_index_2051580_comb ^ p8_array_index_2051581_comb ^ p8_array_index_2051582_comb ^ p8_array_index_2051583_comb ^ p7_array_index_2051387 ^ p7_literal_2043923[p7_array_index_2051420] ^ p7_array_index_2051389 ^ p7_literal_2043920[p7_array_index_2051422] ^ p7_literal_2043918[p7_array_index_2051391] ^ p7_literal_2043916[p7_array_index_2051392] ^ p7_literal_2043914[p7_array_index_2051393] ^ p7_literal_2043912[p7_array_index_2051394] ^ p7_literal_2043910[p7_array_index_2051395] ^ p7_array_index_2051396;
  assign p8_array_index_2051599_comb = p7_literal_2043920[p7_bit_slice_2051378];
  assign p8_array_index_2051600_comb = p7_literal_2043918[p7_bit_slice_2051379];
  assign p8_array_index_2051601_comb = p7_literal_2043916[p7_bit_slice_2051380];
  assign p8_array_index_2051602_comb = p7_literal_2043914[p7_bit_slice_2051381];
  assign p8_array_index_2051603_comb = p7_literal_2043912[p7_res7__1025];
  assign p8_array_index_2051606_comb = p7_literal_2043912[p7_res7__992];
  assign p8_array_index_2051607_comb = p7_literal_2043914[p7_array_index_2051382];
  assign p8_array_index_2051608_comb = p7_literal_2043916[p7_array_index_2051383];
  assign p8_array_index_2051609_comb = p7_literal_2043918[p7_array_index_2051384];
  assign p8_array_index_2051610_comb = p7_literal_2043920[p7_array_index_2051385];
  assign p8_res7__1029_comb = p7_literal_2043910[p7_bit_slice_2051371] ^ p7_literal_2043912[p7_bit_slice_2051372] ^ p7_literal_2043914[p7_bit_slice_2051373] ^ p7_literal_2043916[p7_bit_slice_2051374] ^ p7_literal_2043918[p7_bit_slice_2051404] ^ p7_literal_2043920[p7_bit_slice_2051375] ^ p7_bit_slice_2051406 ^ p7_literal_2043923[p7_bit_slice_2051376] ^ p7_bit_slice_2051377 ^ p8_array_index_2051599_comb ^ p8_array_index_2051600_comb ^ p8_array_index_2051601_comb ^ p8_array_index_2051602_comb ^ p8_array_index_2051603_comb ^ p7_literal_2043910[p7_res7__1027] ^ p7_bit_slice_2051370;
  assign p8_res7__996_comb = p7_literal_2043910[p8_res7__994_comb] ^ p8_array_index_2051606_comb ^ p8_array_index_2051607_comb ^ p8_array_index_2051608_comb ^ p8_array_index_2051609_comb ^ p8_array_index_2051610_comb ^ p7_array_index_2051386 ^ p7_literal_2043923[p7_array_index_2051387] ^ p7_array_index_2051420 ^ p7_literal_2043920[p7_array_index_2051389] ^ p7_literal_2043918[p7_array_index_2051422] ^ p7_literal_2043916[p7_array_index_2051391] ^ p7_literal_2043914[p7_array_index_2051392] ^ p7_literal_2043912[p7_array_index_2051393] ^ p7_literal_2043910[p7_array_index_2051394] ^ p7_array_index_2051395;
  assign p8_array_index_2051627_comb = p7_literal_2043920[p7_bit_slice_2051379];
  assign p8_array_index_2051628_comb = p7_literal_2043918[p7_bit_slice_2051380];
  assign p8_array_index_2051629_comb = p7_literal_2043916[p7_bit_slice_2051381];
  assign p8_array_index_2051630_comb = p7_literal_2043914[p7_res7__1025];
  assign p8_array_index_2051631_comb = p7_literal_2043912[p7_res7__1027];
  assign p8_array_index_2051634_comb = p7_literal_2043912[p8_res7__994_comb];
  assign p8_array_index_2051635_comb = p7_literal_2043914[p7_res7__992];
  assign p8_array_index_2051636_comb = p7_literal_2043916[p7_array_index_2051382];
  assign p8_array_index_2051637_comb = p7_literal_2043918[p7_array_index_2051383];
  assign p8_array_index_2051638_comb = p7_literal_2043920[p7_array_index_2051384];
  assign p8_res7__1031_comb = p7_literal_2043910[p7_bit_slice_2051372] ^ p7_literal_2043912[p7_bit_slice_2051373] ^ p7_literal_2043914[p7_bit_slice_2051374] ^ p7_literal_2043916[p7_bit_slice_2051404] ^ p7_literal_2043918[p7_bit_slice_2051375] ^ p7_literal_2043920[p7_bit_slice_2051406] ^ p7_bit_slice_2051376 ^ p7_literal_2043923[p7_bit_slice_2051377] ^ p7_bit_slice_2051378 ^ p8_array_index_2051627_comb ^ p8_array_index_2051628_comb ^ p8_array_index_2051629_comb ^ p8_array_index_2051630_comb ^ p8_array_index_2051631_comb ^ p7_literal_2043910[p8_res7__1029_comb] ^ p7_bit_slice_2051371;
  assign p8_res7__998_comb = p7_literal_2043910[p8_res7__996_comb] ^ p8_array_index_2051634_comb ^ p8_array_index_2051635_comb ^ p8_array_index_2051636_comb ^ p8_array_index_2051637_comb ^ p8_array_index_2051638_comb ^ p7_array_index_2051385 ^ p7_literal_2043923[p7_array_index_2051386] ^ p7_array_index_2051387 ^ p7_literal_2043920[p7_array_index_2051420] ^ p7_literal_2043918[p7_array_index_2051389] ^ p7_literal_2043916[p7_array_index_2051422] ^ p7_literal_2043914[p7_array_index_2051391] ^ p7_literal_2043912[p7_array_index_2051392] ^ p7_literal_2043910[p7_array_index_2051393] ^ p7_array_index_2051394;
  assign p8_array_index_2051654_comb = p7_literal_2043920[p7_bit_slice_2051380];
  assign p8_array_index_2051655_comb = p7_literal_2043918[p7_bit_slice_2051381];
  assign p8_array_index_2051656_comb = p7_literal_2043916[p7_res7__1025];
  assign p8_array_index_2051657_comb = p7_literal_2043914[p7_res7__1027];
  assign p8_array_index_2051662_comb = p7_literal_2043914[p8_res7__994_comb];
  assign p8_array_index_2051663_comb = p7_literal_2043916[p7_res7__992];
  assign p8_array_index_2051664_comb = p7_literal_2043918[p7_array_index_2051382];
  assign p8_array_index_2051665_comb = p7_literal_2043920[p7_array_index_2051383];
  assign p8_res7__1033_comb = p7_literal_2043910[p7_bit_slice_2051373] ^ p7_literal_2043912[p7_bit_slice_2051374] ^ p7_literal_2043914[p7_bit_slice_2051404] ^ p7_literal_2043916[p7_bit_slice_2051375] ^ p7_literal_2043918[p7_bit_slice_2051406] ^ p7_array_index_2051407 ^ p7_bit_slice_2051377 ^ p7_literal_2043923[p7_bit_slice_2051378] ^ p7_bit_slice_2051379 ^ p8_array_index_2051654_comb ^ p8_array_index_2051655_comb ^ p8_array_index_2051656_comb ^ p8_array_index_2051657_comb ^ p7_literal_2043912[p8_res7__1029_comb] ^ p7_literal_2043910[p8_res7__1031_comb] ^ p7_bit_slice_2051372;
  assign p8_res7__1000_comb = p7_literal_2043910[p8_res7__998_comb] ^ p7_literal_2043912[p8_res7__996_comb] ^ p8_array_index_2051662_comb ^ p8_array_index_2051663_comb ^ p8_array_index_2051664_comb ^ p8_array_index_2051665_comb ^ p7_array_index_2051384 ^ p7_literal_2043923[p7_array_index_2051385] ^ p7_array_index_2051386 ^ p7_array_index_2051419 ^ p7_literal_2043918[p7_array_index_2051420] ^ p7_literal_2043916[p7_array_index_2051389] ^ p7_literal_2043914[p7_array_index_2051422] ^ p7_literal_2043912[p7_array_index_2051391] ^ p7_literal_2043910[p7_array_index_2051392] ^ p7_array_index_2051393;
  assign p8_array_index_2051680_comb = p7_literal_2043920[p7_bit_slice_2051381];
  assign p8_array_index_2051681_comb = p7_literal_2043918[p7_res7__1025];
  assign p8_array_index_2051682_comb = p7_literal_2043916[p7_res7__1027];
  assign p8_array_index_2051683_comb = p7_literal_2043914[p8_res7__1029_comb];
  assign p8_array_index_2051688_comb = p7_literal_2043914[p8_res7__996_comb];
  assign p8_array_index_2051689_comb = p7_literal_2043916[p8_res7__994_comb];
  assign p8_array_index_2051690_comb = p7_literal_2043918[p7_res7__992];
  assign p8_array_index_2051691_comb = p7_literal_2043920[p7_array_index_2051382];
  assign p8_res7__1035_comb = p7_literal_2043910[p7_bit_slice_2051374] ^ p7_literal_2043912[p7_bit_slice_2051404] ^ p7_literal_2043914[p7_bit_slice_2051375] ^ p7_literal_2043916[p7_bit_slice_2051406] ^ p7_literal_2043918[p7_bit_slice_2051376] ^ p7_array_index_2051439 ^ p7_bit_slice_2051378 ^ p7_literal_2043923[p7_bit_slice_2051379] ^ p7_bit_slice_2051380 ^ p8_array_index_2051680_comb ^ p8_array_index_2051681_comb ^ p8_array_index_2051682_comb ^ p8_array_index_2051683_comb ^ p7_literal_2043912[p8_res7__1031_comb] ^ p7_literal_2043910[p8_res7__1033_comb] ^ p7_bit_slice_2051373;
  assign p8_res7__1002_comb = p7_literal_2043910[p8_res7__1000_comb] ^ p7_literal_2043912[p8_res7__998_comb] ^ p8_array_index_2051688_comb ^ p8_array_index_2051689_comb ^ p8_array_index_2051690_comb ^ p8_array_index_2051691_comb ^ p7_array_index_2051383 ^ p7_literal_2043923[p7_array_index_2051384] ^ p7_array_index_2051385 ^ p8_array_index_2051583_comb ^ p7_literal_2043918[p7_array_index_2051387] ^ p7_literal_2043916[p7_array_index_2051420] ^ p7_literal_2043914[p7_array_index_2051389] ^ p7_literal_2043912[p7_array_index_2051422] ^ p7_literal_2043910[p7_array_index_2051391] ^ p7_array_index_2051392;
  assign p8_array_index_2051705_comb = p7_literal_2043920[p7_res7__1025];
  assign p8_array_index_2051706_comb = p7_literal_2043918[p7_res7__1027];
  assign p8_array_index_2051707_comb = p7_literal_2043916[p8_res7__1029_comb];
  assign p8_array_index_2051714_comb = p7_literal_2043916[p8_res7__996_comb];
  assign p8_array_index_2051715_comb = p7_literal_2043918[p8_res7__994_comb];
  assign p8_array_index_2051716_comb = p7_literal_2043920[p7_res7__992];
  assign p8_res7__1037_comb = p7_literal_2043910[p7_bit_slice_2051404] ^ p7_literal_2043912[p7_bit_slice_2051375] ^ p7_literal_2043914[p7_bit_slice_2051406] ^ p7_literal_2043916[p7_bit_slice_2051376] ^ p7_array_index_2051408 ^ p8_array_index_2051599_comb ^ p7_bit_slice_2051379 ^ p7_literal_2043923[p7_bit_slice_2051380] ^ p7_bit_slice_2051381 ^ p8_array_index_2051705_comb ^ p8_array_index_2051706_comb ^ p8_array_index_2051707_comb ^ p7_literal_2043914[p8_res7__1031_comb] ^ p7_literal_2043912[p8_res7__1033_comb] ^ p7_literal_2043910[p8_res7__1035_comb] ^ p7_bit_slice_2051374;
  assign p8_res7__1004_comb = p7_literal_2043910[p8_res7__1002_comb] ^ p7_literal_2043912[p8_res7__1000_comb] ^ p7_literal_2043914[p8_res7__998_comb] ^ p8_array_index_2051714_comb ^ p8_array_index_2051715_comb ^ p8_array_index_2051716_comb ^ p7_array_index_2051382 ^ p7_literal_2043923[p7_array_index_2051383] ^ p7_array_index_2051384 ^ p8_array_index_2051610_comb ^ p7_array_index_2051418 ^ p7_literal_2043916[p7_array_index_2051387] ^ p7_literal_2043914[p7_array_index_2051420] ^ p7_literal_2043912[p7_array_index_2051389] ^ p7_literal_2043910[p7_array_index_2051422] ^ p7_array_index_2051391;
  assign p8_array_index_2051729_comb = p7_literal_2043920[p7_res7__1027];
  assign p8_array_index_2051730_comb = p7_literal_2043918[p8_res7__1029_comb];
  assign p8_array_index_2051731_comb = p7_literal_2043916[p8_res7__1031_comb];
  assign p8_array_index_2051738_comb = p7_literal_2043916[p8_res7__998_comb];
  assign p8_array_index_2051739_comb = p7_literal_2043918[p8_res7__996_comb];
  assign p8_array_index_2051740_comb = p7_literal_2043920[p8_res7__994_comb];
  assign p8_res7__1039_comb = p7_literal_2043910[p7_bit_slice_2051375] ^ p7_literal_2043912[p7_bit_slice_2051406] ^ p7_literal_2043914[p7_bit_slice_2051376] ^ p7_literal_2043916[p7_bit_slice_2051377] ^ p7_array_index_2051440 ^ p8_array_index_2051627_comb ^ p7_bit_slice_2051380 ^ p7_literal_2043923[p7_bit_slice_2051381] ^ p7_res7__1025 ^ p8_array_index_2051729_comb ^ p8_array_index_2051730_comb ^ p8_array_index_2051731_comb ^ p7_literal_2043914[p8_res7__1033_comb] ^ p7_literal_2043912[p8_res7__1035_comb] ^ p7_literal_2043910[p8_res7__1037_comb] ^ p7_bit_slice_2051404;
  assign p8_res7__1006_comb = p7_literal_2043910[p8_res7__1004_comb] ^ p7_literal_2043912[p8_res7__1002_comb] ^ p7_literal_2043914[p8_res7__1000_comb] ^ p8_array_index_2051738_comb ^ p8_array_index_2051739_comb ^ p8_array_index_2051740_comb ^ p7_res7__992 ^ p7_literal_2043923[p7_array_index_2051382] ^ p7_array_index_2051383 ^ p8_array_index_2051638_comb ^ p8_array_index_2051582_comb ^ p7_literal_2043916[p7_array_index_2051386] ^ p7_literal_2043914[p7_array_index_2051387] ^ p7_literal_2043912[p7_array_index_2051420] ^ p7_literal_2043910[p7_array_index_2051389] ^ p7_array_index_2051422;
  assign p8_array_index_2051752_comb = p7_literal_2043920[p8_res7__1029_comb];
  assign p8_array_index_2051753_comb = p7_literal_2043918[p8_res7__1031_comb];
  assign p8_array_index_2051762_comb = p7_literal_2043918[p8_res7__998_comb];
  assign p8_array_index_2051763_comb = p7_literal_2043920[p8_res7__996_comb];
  assign p8_res7__1041_comb = p7_literal_2043910[p7_bit_slice_2051406] ^ p7_literal_2043912[p7_bit_slice_2051376] ^ p7_literal_2043914[p7_bit_slice_2051377] ^ p7_array_index_2051409 ^ p8_array_index_2051600_comb ^ p8_array_index_2051654_comb ^ p7_bit_slice_2051381 ^ p7_literal_2043923[p7_res7__1025] ^ p7_res7__1027 ^ p8_array_index_2051752_comb ^ p8_array_index_2051753_comb ^ p7_literal_2043916[p8_res7__1033_comb] ^ p7_literal_2043914[p8_res7__1035_comb] ^ p7_literal_2043912[p8_res7__1037_comb] ^ p7_literal_2043910[p8_res7__1039_comb] ^ p7_bit_slice_2051375;
  assign p8_res7__1008_comb = p7_literal_2043910[p8_res7__1006_comb] ^ p7_literal_2043912[p8_res7__1004_comb] ^ p7_literal_2043914[p8_res7__1002_comb] ^ p7_literal_2043916[p8_res7__1000_comb] ^ p8_array_index_2051762_comb ^ p8_array_index_2051763_comb ^ p8_res7__994_comb ^ p7_literal_2043923[p7_res7__992] ^ p7_array_index_2051382 ^ p8_array_index_2051665_comb ^ p8_array_index_2051609_comb ^ p7_array_index_2051417 ^ p7_literal_2043914[p7_array_index_2051386] ^ p7_literal_2043912[p7_array_index_2051387] ^ p7_literal_2043910[p7_array_index_2051420] ^ p7_array_index_2051389;
  assign p8_array_index_2051774_comb = p7_literal_2043920[p8_res7__1031_comb];
  assign p8_array_index_2051775_comb = p7_literal_2043918[p8_res7__1033_comb];
  assign p8_array_index_2051784_comb = p7_literal_2043918[p8_res7__1000_comb];
  assign p8_array_index_2051785_comb = p7_literal_2043920[p8_res7__998_comb];
  assign p8_res7__1043_comb = p7_literal_2043910[p7_bit_slice_2051376] ^ p7_literal_2043912[p7_bit_slice_2051377] ^ p7_literal_2043914[p7_bit_slice_2051378] ^ p7_array_index_2051441 ^ p8_array_index_2051628_comb ^ p8_array_index_2051680_comb ^ p7_res7__1025 ^ p7_literal_2043923[p7_res7__1027] ^ p8_res7__1029_comb ^ p8_array_index_2051774_comb ^ p8_array_index_2051775_comb ^ p7_literal_2043916[p8_res7__1035_comb] ^ p7_literal_2043914[p8_res7__1037_comb] ^ p7_literal_2043912[p8_res7__1039_comb] ^ p7_literal_2043910[p8_res7__1041_comb] ^ p7_bit_slice_2051406;
  assign p8_res7__1010_comb = p7_literal_2043910[p8_res7__1008_comb] ^ p7_literal_2043912[p8_res7__1006_comb] ^ p7_literal_2043914[p8_res7__1004_comb] ^ p7_literal_2043916[p8_res7__1002_comb] ^ p8_array_index_2051784_comb ^ p8_array_index_2051785_comb ^ p8_res7__996_comb ^ p7_literal_2043923[p8_res7__994_comb] ^ p7_res7__992 ^ p8_array_index_2051691_comb ^ p8_array_index_2051637_comb ^ p8_array_index_2051581_comb ^ p7_literal_2043914[p7_array_index_2051385] ^ p7_literal_2043912[p7_array_index_2051386] ^ p7_literal_2043910[p7_array_index_2051387] ^ p7_array_index_2051420;
  assign p8_array_index_2051795_comb = p7_literal_2043920[p8_res7__1033_comb];
  assign p8_array_index_2051806_comb = p7_literal_2043920[p8_res7__1000_comb];
  assign p8_res7__1045_comb = p7_literal_2043910[p7_bit_slice_2051377] ^ p7_literal_2043912[p7_bit_slice_2051378] ^ p7_array_index_2051410 ^ p8_array_index_2051601_comb ^ p8_array_index_2051655_comb ^ p8_array_index_2051705_comb ^ p7_res7__1027 ^ p7_literal_2043923[p8_res7__1029_comb] ^ p8_res7__1031_comb ^ p8_array_index_2051795_comb ^ p7_literal_2043918[p8_res7__1035_comb] ^ p7_literal_2043916[p8_res7__1037_comb] ^ p7_literal_2043914[p8_res7__1039_comb] ^ p7_literal_2043912[p8_res7__1041_comb] ^ p7_literal_2043910[p8_res7__1043_comb] ^ p7_bit_slice_2051376;
  assign p8_res7__1012_comb = p7_literal_2043910[p8_res7__1010_comb] ^ p7_literal_2043912[p8_res7__1008_comb] ^ p7_literal_2043914[p8_res7__1006_comb] ^ p7_literal_2043916[p8_res7__1004_comb] ^ p7_literal_2043918[p8_res7__1002_comb] ^ p8_array_index_2051806_comb ^ p8_res7__998_comb ^ p7_literal_2043923[p8_res7__996_comb] ^ p8_res7__994_comb ^ p8_array_index_2051716_comb ^ p8_array_index_2051664_comb ^ p8_array_index_2051608_comb ^ p7_array_index_2051416 ^ p7_literal_2043912[p7_array_index_2051385] ^ p7_literal_2043910[p7_array_index_2051386] ^ p7_array_index_2051387;
  assign p8_array_index_2051815_comb = p7_literal_2043920[p8_res7__1035_comb];
  assign p8_array_index_2051826_comb = p7_literal_2043920[p8_res7__1002_comb];
  assign p8_res7__1047_comb = p7_literal_2043910[p7_bit_slice_2051378] ^ p7_literal_2043912[p7_bit_slice_2051379] ^ p7_array_index_2051442 ^ p8_array_index_2051629_comb ^ p8_array_index_2051681_comb ^ p8_array_index_2051729_comb ^ p8_res7__1029_comb ^ p7_literal_2043923[p8_res7__1031_comb] ^ p8_res7__1033_comb ^ p8_array_index_2051815_comb ^ p7_literal_2043918[p8_res7__1037_comb] ^ p7_literal_2043916[p8_res7__1039_comb] ^ p7_literal_2043914[p8_res7__1041_comb] ^ p7_literal_2043912[p8_res7__1043_comb] ^ p7_literal_2043910[p8_res7__1045_comb] ^ p7_bit_slice_2051377;
  assign p8_res7__1014_comb = p7_literal_2043910[p8_res7__1012_comb] ^ p7_literal_2043912[p8_res7__1010_comb] ^ p7_literal_2043914[p8_res7__1008_comb] ^ p7_literal_2043916[p8_res7__1006_comb] ^ p7_literal_2043918[p8_res7__1004_comb] ^ p8_array_index_2051826_comb ^ p8_res7__1000_comb ^ p7_literal_2043923[p8_res7__998_comb] ^ p8_res7__996_comb ^ p8_array_index_2051740_comb ^ p8_array_index_2051690_comb ^ p8_array_index_2051636_comb ^ p8_array_index_2051580_comb ^ p7_literal_2043912[p7_array_index_2051384] ^ p7_literal_2043910[p7_array_index_2051385] ^ p7_array_index_2051386;
  assign p8_res7__1049_comb = p7_literal_2043910[p7_bit_slice_2051379] ^ p7_array_index_2051411 ^ p8_array_index_2051602_comb ^ p8_array_index_2051656_comb ^ p8_array_index_2051706_comb ^ p8_array_index_2051752_comb ^ p8_res7__1031_comb ^ p7_literal_2043923[p8_res7__1033_comb] ^ p8_res7__1035_comb ^ p7_literal_2043920[p8_res7__1037_comb] ^ p7_literal_2043918[p8_res7__1039_comb] ^ p7_literal_2043916[p8_res7__1041_comb] ^ p7_literal_2043914[p8_res7__1043_comb] ^ p7_literal_2043912[p8_res7__1045_comb] ^ p7_literal_2043910[p8_res7__1047_comb] ^ p7_bit_slice_2051378;
  assign p8_res7__1016_comb = p7_literal_2043910[p8_res7__1014_comb] ^ p7_literal_2043912[p8_res7__1012_comb] ^ p7_literal_2043914[p8_res7__1010_comb] ^ p7_literal_2043916[p8_res7__1008_comb] ^ p7_literal_2043918[p8_res7__1006_comb] ^ p7_literal_2043920[p8_res7__1004_comb] ^ p8_res7__1002_comb ^ p7_literal_2043923[p8_res7__1000_comb] ^ p8_res7__998_comb ^ p8_array_index_2051763_comb ^ p8_array_index_2051715_comb ^ p8_array_index_2051663_comb ^ p8_array_index_2051607_comb ^ p7_array_index_2051415 ^ p7_literal_2043910[p7_array_index_2051384] ^ p7_array_index_2051385;
  assign p8_res7__1051_comb = p7_literal_2043910[p7_bit_slice_2051380] ^ p7_array_index_2051443 ^ p8_array_index_2051630_comb ^ p8_array_index_2051682_comb ^ p8_array_index_2051730_comb ^ p8_array_index_2051774_comb ^ p8_res7__1033_comb ^ p7_literal_2043923[p8_res7__1035_comb] ^ p8_res7__1037_comb ^ p7_literal_2043920[p8_res7__1039_comb] ^ p7_literal_2043918[p8_res7__1041_comb] ^ p7_literal_2043916[p8_res7__1043_comb] ^ p7_literal_2043914[p8_res7__1045_comb] ^ p7_literal_2043912[p8_res7__1047_comb] ^ p7_literal_2043910[p8_res7__1049_comb] ^ p7_bit_slice_2051379;
  assign p8_res7__1018_comb = p7_literal_2043910[p8_res7__1016_comb] ^ p7_literal_2043912[p8_res7__1014_comb] ^ p7_literal_2043914[p8_res7__1012_comb] ^ p7_literal_2043916[p8_res7__1010_comb] ^ p7_literal_2043918[p8_res7__1008_comb] ^ p7_literal_2043920[p8_res7__1006_comb] ^ p8_res7__1004_comb ^ p7_literal_2043923[p8_res7__1002_comb] ^ p8_res7__1000_comb ^ p8_array_index_2051785_comb ^ p8_array_index_2051739_comb ^ p8_array_index_2051689_comb ^ p8_array_index_2051635_comb ^ p8_array_index_2051579_comb ^ p7_literal_2043910[p7_array_index_2051383] ^ p7_array_index_2051384;
  assign p8_res7__1053_comb = p7_array_index_2051412 ^ p8_array_index_2051603_comb ^ p8_array_index_2051657_comb ^ p8_array_index_2051707_comb ^ p8_array_index_2051753_comb ^ p8_array_index_2051795_comb ^ p8_res7__1035_comb ^ p7_literal_2043923[p8_res7__1037_comb] ^ p8_res7__1039_comb ^ p7_literal_2043920[p8_res7__1041_comb] ^ p7_literal_2043918[p8_res7__1043_comb] ^ p7_literal_2043916[p8_res7__1045_comb] ^ p7_literal_2043914[p8_res7__1047_comb] ^ p7_literal_2043912[p8_res7__1049_comb] ^ p7_literal_2043910[p8_res7__1051_comb] ^ p7_bit_slice_2051380;
  assign p8_res7__1020_comb = p7_literal_2043910[p8_res7__1018_comb] ^ p7_literal_2043912[p8_res7__1016_comb] ^ p7_literal_2043914[p8_res7__1014_comb] ^ p7_literal_2043916[p8_res7__1012_comb] ^ p7_literal_2043918[p8_res7__1010_comb] ^ p7_literal_2043920[p8_res7__1008_comb] ^ p8_res7__1006_comb ^ p7_literal_2043923[p8_res7__1004_comb] ^ p8_res7__1002_comb ^ p8_array_index_2051806_comb ^ p8_array_index_2051762_comb ^ p8_array_index_2051714_comb ^ p8_array_index_2051662_comb ^ p8_array_index_2051606_comb ^ p7_array_index_2051414 ^ p7_array_index_2051383;
  assign p8_res7__1055_comb = p7_array_index_2051444 ^ p8_array_index_2051631_comb ^ p8_array_index_2051683_comb ^ p8_array_index_2051731_comb ^ p8_array_index_2051775_comb ^ p8_array_index_2051815_comb ^ p8_res7__1037_comb ^ p7_literal_2043923[p8_res7__1039_comb] ^ p8_res7__1041_comb ^ p7_literal_2043920[p8_res7__1043_comb] ^ p7_literal_2043918[p8_res7__1045_comb] ^ p7_literal_2043916[p8_res7__1047_comb] ^ p7_literal_2043914[p8_res7__1049_comb] ^ p7_literal_2043912[p8_res7__1051_comb] ^ p7_literal_2043910[p8_res7__1053_comb] ^ p7_bit_slice_2051381;
  assign p8_res7__1022_comb = p7_literal_2043910[p8_res7__1020_comb] ^ p7_literal_2043912[p8_res7__1018_comb] ^ p7_literal_2043914[p8_res7__1016_comb] ^ p7_literal_2043916[p8_res7__1014_comb] ^ p7_literal_2043918[p8_res7__1012_comb] ^ p7_literal_2043920[p8_res7__1010_comb] ^ p8_res7__1008_comb ^ p7_literal_2043923[p8_res7__1006_comb] ^ p8_res7__1004_comb ^ p8_array_index_2051826_comb ^ p8_array_index_2051784_comb ^ p8_array_index_2051738_comb ^ p8_array_index_2051688_comb ^ p8_array_index_2051634_comb ^ p8_array_index_2051578_comb ^ p7_array_index_2051382;
  assign p8_res__31_comb = {p8_res7__1022_comb, p8_res7__1020_comb, p8_res7__1018_comb, p8_res7__1016_comb, p8_res7__1014_comb, p8_res7__1012_comb, p8_res7__1010_comb, p8_res7__1008_comb, p8_res7__1006_comb, p8_res7__1004_comb, p8_res7__1002_comb, p8_res7__1000_comb, p8_res7__998_comb, p8_res7__996_comb, p8_res7__994_comb, p7_res7__992};
  assign p8_permut__32_comb = {literal_2051898[p7_res7__1025], literal_2051898[p7_res7__1027], literal_2051898[p8_res7__1029_comb], literal_2051898[p8_res7__1031_comb], literal_2051898[p8_res7__1033_comb], literal_2051898[p8_res7__1035_comb], literal_2051898[p8_res7__1037_comb], literal_2051898[p8_res7__1039_comb], literal_2051898[p8_res7__1041_comb], literal_2051898[p8_res7__1043_comb], literal_2051898[p8_res7__1045_comb], literal_2051898[p8_res7__1047_comb], literal_2051898[p8_res7__1049_comb], literal_2051898[p8_res7__1051_comb], literal_2051898[p8_res7__1053_comb], literal_2051898[p8_res7__1055_comb]};
  assign p8_xor_2051919_comb = p8_res__31_comb ^ p7_xor_2051134 ^ p8_permut__32_comb;
  assign p8_array_index_2051942_comb = p7_literal_2043920[p8_xor_2051919_comb[47:40]];
  assign p8_array_index_2051943_comb = p7_literal_2043918[p8_xor_2051919_comb[39:32]];
  assign p8_array_index_2051944_comb = p7_literal_2043916[p8_xor_2051919_comb[31:24]];
  assign p8_array_index_2051945_comb = p7_literal_2043914[p8_xor_2051919_comb[23:16]];
  assign p8_array_index_2051946_comb = p7_literal_2043912[p8_xor_2051919_comb[15:8]];
  assign p8_array_index_2051947_comb = p7_literal_2043910[p8_xor_2051919_comb[7:0]];
  assign p8_res7__1057_comb = p7_literal_2043910[p8_xor_2051919_comb[119:112]] ^ p7_literal_2043912[p8_xor_2051919_comb[111:104]] ^ p7_literal_2043914[p8_xor_2051919_comb[103:96]] ^ p7_literal_2043916[p8_xor_2051919_comb[95:88]] ^ p7_literal_2043918[p8_xor_2051919_comb[87:80]] ^ p7_literal_2043920[p8_xor_2051919_comb[79:72]] ^ p8_xor_2051919_comb[71:64] ^ p7_literal_2043923[p8_xor_2051919_comb[63:56]] ^ p8_xor_2051919_comb[55:48] ^ p8_array_index_2051942_comb ^ p8_array_index_2051943_comb ^ p8_array_index_2051944_comb ^ p8_array_index_2051945_comb ^ p8_array_index_2051946_comb ^ p8_array_index_2051947_comb ^ p8_xor_2051919_comb[127:120];
  assign p8_array_index_2051957_comb = p7_literal_2043920[p8_xor_2051919_comb[39:32]];
  assign p8_array_index_2051958_comb = p7_literal_2043918[p8_xor_2051919_comb[31:24]];
  assign p8_array_index_2051959_comb = p7_literal_2043916[p8_xor_2051919_comb[23:16]];
  assign p8_array_index_2051960_comb = p7_literal_2043914[p8_xor_2051919_comb[15:8]];
  assign p8_array_index_2051961_comb = p7_literal_2043912[p8_xor_2051919_comb[7:0]];
  assign p8_array_index_2051962_comb = p7_literal_2043910[p8_res7__1057_comb];
  assign p8_res7__1059_comb = p7_literal_2043910[p8_xor_2051919_comb[111:104]] ^ p7_literal_2043912[p8_xor_2051919_comb[103:96]] ^ p7_literal_2043914[p8_xor_2051919_comb[95:88]] ^ p7_literal_2043916[p8_xor_2051919_comb[87:80]] ^ p7_literal_2043918[p8_xor_2051919_comb[79:72]] ^ p7_literal_2043920[p8_xor_2051919_comb[71:64]] ^ p8_xor_2051919_comb[63:56] ^ p7_literal_2043923[p8_xor_2051919_comb[55:48]] ^ p8_xor_2051919_comb[47:40] ^ p8_array_index_2051957_comb ^ p8_array_index_2051958_comb ^ p8_array_index_2051959_comb ^ p8_array_index_2051960_comb ^ p8_array_index_2051961_comb ^ p8_array_index_2051962_comb ^ p8_xor_2051919_comb[119:112];
  assign p8_array_index_2051971_comb = p7_literal_2043920[p8_xor_2051919_comb[31:24]];
  assign p8_array_index_2051972_comb = p7_literal_2043918[p8_xor_2051919_comb[23:16]];
  assign p8_array_index_2051973_comb = p7_literal_2043916[p8_xor_2051919_comb[15:8]];
  assign p8_array_index_2051974_comb = p7_literal_2043914[p8_xor_2051919_comb[7:0]];
  assign p8_array_index_2051975_comb = p7_literal_2043912[p8_res7__1057_comb];
  assign p8_res7__1061_comb = p7_literal_2043910[p8_xor_2051919_comb[103:96]] ^ p7_literal_2043912[p8_xor_2051919_comb[95:88]] ^ p7_literal_2043914[p8_xor_2051919_comb[87:80]] ^ p7_literal_2043916[p8_xor_2051919_comb[79:72]] ^ p7_literal_2043918[p8_xor_2051919_comb[71:64]] ^ p7_literal_2043920[p8_xor_2051919_comb[63:56]] ^ p8_xor_2051919_comb[55:48] ^ p7_literal_2043923[p8_xor_2051919_comb[47:40]] ^ p8_xor_2051919_comb[39:32] ^ p8_array_index_2051971_comb ^ p8_array_index_2051972_comb ^ p8_array_index_2051973_comb ^ p8_array_index_2051974_comb ^ p8_array_index_2051975_comb ^ p7_literal_2043910[p8_res7__1059_comb] ^ p8_xor_2051919_comb[111:104];
  assign p8_array_index_2051985_comb = p7_literal_2043920[p8_xor_2051919_comb[23:16]];
  assign p8_array_index_2051986_comb = p7_literal_2043918[p8_xor_2051919_comb[15:8]];
  assign p8_array_index_2051987_comb = p7_literal_2043916[p8_xor_2051919_comb[7:0]];
  assign p8_array_index_2051988_comb = p7_literal_2043914[p8_res7__1057_comb];
  assign p8_array_index_2051989_comb = p7_literal_2043912[p8_res7__1059_comb];
  assign p8_res7__1063_comb = p7_literal_2043910[p8_xor_2051919_comb[95:88]] ^ p7_literal_2043912[p8_xor_2051919_comb[87:80]] ^ p7_literal_2043914[p8_xor_2051919_comb[79:72]] ^ p7_literal_2043916[p8_xor_2051919_comb[71:64]] ^ p7_literal_2043918[p8_xor_2051919_comb[63:56]] ^ p7_literal_2043920[p8_xor_2051919_comb[55:48]] ^ p8_xor_2051919_comb[47:40] ^ p7_literal_2043923[p8_xor_2051919_comb[39:32]] ^ p8_xor_2051919_comb[31:24] ^ p8_array_index_2051985_comb ^ p8_array_index_2051986_comb ^ p8_array_index_2051987_comb ^ p8_array_index_2051988_comb ^ p8_array_index_2051989_comb ^ p7_literal_2043910[p8_res7__1061_comb] ^ p8_xor_2051919_comb[103:96];
  assign p8_array_index_2051998_comb = p7_literal_2043920[p8_xor_2051919_comb[15:8]];
  assign p8_array_index_2051999_comb = p7_literal_2043918[p8_xor_2051919_comb[7:0]];
  assign p8_array_index_2052000_comb = p7_literal_2043916[p8_res7__1057_comb];
  assign p8_array_index_2052001_comb = p7_literal_2043914[p8_res7__1059_comb];
  assign p8_res7__1065_comb = p7_literal_2043910[p8_xor_2051919_comb[87:80]] ^ p7_literal_2043912[p8_xor_2051919_comb[79:72]] ^ p7_literal_2043914[p8_xor_2051919_comb[71:64]] ^ p7_literal_2043916[p8_xor_2051919_comb[63:56]] ^ p7_literal_2043918[p8_xor_2051919_comb[55:48]] ^ p8_array_index_2051942_comb ^ p8_xor_2051919_comb[39:32] ^ p7_literal_2043923[p8_xor_2051919_comb[31:24]] ^ p8_xor_2051919_comb[23:16] ^ p8_array_index_2051998_comb ^ p8_array_index_2051999_comb ^ p8_array_index_2052000_comb ^ p8_array_index_2052001_comb ^ p7_literal_2043912[p8_res7__1061_comb] ^ p7_literal_2043910[p8_res7__1063_comb] ^ p8_xor_2051919_comb[95:88];
  assign p8_array_index_2052011_comb = p7_literal_2043920[p8_xor_2051919_comb[7:0]];
  assign p8_array_index_2052012_comb = p7_literal_2043918[p8_res7__1057_comb];
  assign p8_array_index_2052013_comb = p7_literal_2043916[p8_res7__1059_comb];
  assign p8_array_index_2052014_comb = p7_literal_2043914[p8_res7__1061_comb];
  assign p8_res7__1067_comb = p7_literal_2043910[p8_xor_2051919_comb[79:72]] ^ p7_literal_2043912[p8_xor_2051919_comb[71:64]] ^ p7_literal_2043914[p8_xor_2051919_comb[63:56]] ^ p7_literal_2043916[p8_xor_2051919_comb[55:48]] ^ p7_literal_2043918[p8_xor_2051919_comb[47:40]] ^ p8_array_index_2051957_comb ^ p8_xor_2051919_comb[31:24] ^ p7_literal_2043923[p8_xor_2051919_comb[23:16]] ^ p8_xor_2051919_comb[15:8] ^ p8_array_index_2052011_comb ^ p8_array_index_2052012_comb ^ p8_array_index_2052013_comb ^ p8_array_index_2052014_comb ^ p7_literal_2043912[p8_res7__1063_comb] ^ p7_literal_2043910[p8_res7__1065_comb] ^ p8_xor_2051919_comb[87:80];
  assign p8_array_index_2052023_comb = p7_literal_2043920[p8_res7__1057_comb];
  assign p8_array_index_2052024_comb = p7_literal_2043918[p8_res7__1059_comb];
  assign p8_array_index_2052025_comb = p7_literal_2043916[p8_res7__1061_comb];
  assign p8_res7__1069_comb = p7_literal_2043910[p8_xor_2051919_comb[71:64]] ^ p7_literal_2043912[p8_xor_2051919_comb[63:56]] ^ p7_literal_2043914[p8_xor_2051919_comb[55:48]] ^ p7_literal_2043916[p8_xor_2051919_comb[47:40]] ^ p8_array_index_2051943_comb ^ p8_array_index_2051971_comb ^ p8_xor_2051919_comb[23:16] ^ p7_literal_2043923[p8_xor_2051919_comb[15:8]] ^ p8_xor_2051919_comb[7:0] ^ p8_array_index_2052023_comb ^ p8_array_index_2052024_comb ^ p8_array_index_2052025_comb ^ p7_literal_2043914[p8_res7__1063_comb] ^ p7_literal_2043912[p8_res7__1065_comb] ^ p7_literal_2043910[p8_res7__1067_comb] ^ p8_xor_2051919_comb[79:72];
  assign p8_array_index_2052035_comb = p7_literal_2043920[p8_res7__1059_comb];
  assign p8_array_index_2052036_comb = p7_literal_2043918[p8_res7__1061_comb];
  assign p8_array_index_2052037_comb = p7_literal_2043916[p8_res7__1063_comb];
  assign p8_res7__1071_comb = p7_literal_2043910[p8_xor_2051919_comb[63:56]] ^ p7_literal_2043912[p8_xor_2051919_comb[55:48]] ^ p7_literal_2043914[p8_xor_2051919_comb[47:40]] ^ p7_literal_2043916[p8_xor_2051919_comb[39:32]] ^ p8_array_index_2051958_comb ^ p8_array_index_2051985_comb ^ p8_xor_2051919_comb[15:8] ^ p7_literal_2043923[p8_xor_2051919_comb[7:0]] ^ p8_res7__1057_comb ^ p8_array_index_2052035_comb ^ p8_array_index_2052036_comb ^ p8_array_index_2052037_comb ^ p7_literal_2043914[p8_res7__1065_comb] ^ p7_literal_2043912[p8_res7__1067_comb] ^ p7_literal_2043910[p8_res7__1069_comb] ^ p8_xor_2051919_comb[71:64];
  assign p8_array_index_2052046_comb = p7_literal_2043920[p8_res7__1061_comb];
  assign p8_array_index_2052047_comb = p7_literal_2043918[p8_res7__1063_comb];
  assign p8_res7__1073_comb = p7_literal_2043910[p8_xor_2051919_comb[55:48]] ^ p7_literal_2043912[p8_xor_2051919_comb[47:40]] ^ p7_literal_2043914[p8_xor_2051919_comb[39:32]] ^ p8_array_index_2051944_comb ^ p8_array_index_2051972_comb ^ p8_array_index_2051998_comb ^ p8_xor_2051919_comb[7:0] ^ p7_literal_2043923[p8_res7__1057_comb] ^ p8_res7__1059_comb ^ p8_array_index_2052046_comb ^ p8_array_index_2052047_comb ^ p7_literal_2043916[p8_res7__1065_comb] ^ p7_literal_2043914[p8_res7__1067_comb] ^ p7_literal_2043912[p8_res7__1069_comb] ^ p7_literal_2043910[p8_res7__1071_comb] ^ p8_xor_2051919_comb[63:56];
  assign p8_array_index_2052057_comb = p7_literal_2043920[p8_res7__1063_comb];
  assign p8_array_index_2052058_comb = p7_literal_2043918[p8_res7__1065_comb];
  assign p8_res7__1075_comb = p7_literal_2043910[p8_xor_2051919_comb[47:40]] ^ p7_literal_2043912[p8_xor_2051919_comb[39:32]] ^ p7_literal_2043914[p8_xor_2051919_comb[31:24]] ^ p8_array_index_2051959_comb ^ p8_array_index_2051986_comb ^ p8_array_index_2052011_comb ^ p8_res7__1057_comb ^ p7_literal_2043923[p8_res7__1059_comb] ^ p8_res7__1061_comb ^ p8_array_index_2052057_comb ^ p8_array_index_2052058_comb ^ p7_literal_2043916[p8_res7__1067_comb] ^ p7_literal_2043914[p8_res7__1069_comb] ^ p7_literal_2043912[p8_res7__1071_comb] ^ p7_literal_2043910[p8_res7__1073_comb] ^ p8_xor_2051919_comb[55:48];
  assign p8_array_index_2052067_comb = p7_literal_2043920[p8_res7__1065_comb];
  assign p8_res7__1077_comb = p7_literal_2043910[p8_xor_2051919_comb[39:32]] ^ p7_literal_2043912[p8_xor_2051919_comb[31:24]] ^ p8_array_index_2051945_comb ^ p8_array_index_2051973_comb ^ p8_array_index_2051999_comb ^ p8_array_index_2052023_comb ^ p8_res7__1059_comb ^ p7_literal_2043923[p8_res7__1061_comb] ^ p8_res7__1063_comb ^ p8_array_index_2052067_comb ^ p7_literal_2043918[p8_res7__1067_comb] ^ p7_literal_2043916[p8_res7__1069_comb] ^ p7_literal_2043914[p8_res7__1071_comb] ^ p7_literal_2043912[p8_res7__1073_comb] ^ p7_literal_2043910[p8_res7__1075_comb] ^ p8_xor_2051919_comb[47:40];
  assign p8_array_index_2052077_comb = p7_literal_2043920[p8_res7__1067_comb];
  assign p8_res7__1079_comb = p7_literal_2043910[p8_xor_2051919_comb[31:24]] ^ p7_literal_2043912[p8_xor_2051919_comb[23:16]] ^ p8_array_index_2051960_comb ^ p8_array_index_2051987_comb ^ p8_array_index_2052012_comb ^ p8_array_index_2052035_comb ^ p8_res7__1061_comb ^ p7_literal_2043923[p8_res7__1063_comb] ^ p8_res7__1065_comb ^ p8_array_index_2052077_comb ^ p7_literal_2043918[p8_res7__1069_comb] ^ p7_literal_2043916[p8_res7__1071_comb] ^ p7_literal_2043914[p8_res7__1073_comb] ^ p7_literal_2043912[p8_res7__1075_comb] ^ p7_literal_2043910[p8_res7__1077_comb] ^ p8_xor_2051919_comb[39:32];
  assign p8_res7__1081_comb = p7_literal_2043910[p8_xor_2051919_comb[23:16]] ^ p8_array_index_2051946_comb ^ p8_array_index_2051974_comb ^ p8_array_index_2052000_comb ^ p8_array_index_2052024_comb ^ p8_array_index_2052046_comb ^ p8_res7__1063_comb ^ p7_literal_2043923[p8_res7__1065_comb] ^ p8_res7__1067_comb ^ p7_literal_2043920[p8_res7__1069_comb] ^ p7_literal_2043918[p8_res7__1071_comb] ^ p7_literal_2043916[p8_res7__1073_comb] ^ p7_literal_2043914[p8_res7__1075_comb] ^ p7_literal_2043912[p8_res7__1077_comb] ^ p7_literal_2043910[p8_res7__1079_comb] ^ p8_xor_2051919_comb[31:24];
  assign p8_res7__1083_comb = p7_literal_2043910[p8_xor_2051919_comb[15:8]] ^ p8_array_index_2051961_comb ^ p8_array_index_2051988_comb ^ p8_array_index_2052013_comb ^ p8_array_index_2052036_comb ^ p8_array_index_2052057_comb ^ p8_res7__1065_comb ^ p7_literal_2043923[p8_res7__1067_comb] ^ p8_res7__1069_comb ^ p7_literal_2043920[p8_res7__1071_comb] ^ p7_literal_2043918[p8_res7__1073_comb] ^ p7_literal_2043916[p8_res7__1075_comb] ^ p7_literal_2043914[p8_res7__1077_comb] ^ p7_literal_2043912[p8_res7__1079_comb] ^ p7_literal_2043910[p8_res7__1081_comb] ^ p8_xor_2051919_comb[23:16];
  assign p8_res7__1085_comb = p8_array_index_2051947_comb ^ p8_array_index_2051975_comb ^ p8_array_index_2052001_comb ^ p8_array_index_2052025_comb ^ p8_array_index_2052047_comb ^ p8_array_index_2052067_comb ^ p8_res7__1067_comb ^ p7_literal_2043923[p8_res7__1069_comb] ^ p8_res7__1071_comb ^ p7_literal_2043920[p8_res7__1073_comb] ^ p7_literal_2043918[p8_res7__1075_comb] ^ p7_literal_2043916[p8_res7__1077_comb] ^ p7_literal_2043914[p8_res7__1079_comb] ^ p7_literal_2043912[p8_res7__1081_comb] ^ p7_literal_2043910[p8_res7__1083_comb] ^ p8_xor_2051919_comb[15:8];
  assign p8_res7__1087_comb = p8_array_index_2051962_comb ^ p8_array_index_2051989_comb ^ p8_array_index_2052014_comb ^ p8_array_index_2052037_comb ^ p8_array_index_2052058_comb ^ p8_array_index_2052077_comb ^ p8_res7__1069_comb ^ p7_literal_2043923[p8_res7__1071_comb] ^ p8_res7__1073_comb ^ p7_literal_2043920[p8_res7__1075_comb] ^ p7_literal_2043918[p8_res7__1077_comb] ^ p7_literal_2043916[p8_res7__1079_comb] ^ p7_literal_2043914[p8_res7__1081_comb] ^ p7_literal_2043912[p8_res7__1083_comb] ^ p7_literal_2043910[p8_res7__1085_comb] ^ p8_xor_2051919_comb[7:0];
  assign p8_permut__33_comb = {literal_2051898[p8_res7__1057_comb], literal_2051898[p8_res7__1059_comb], literal_2051898[p8_res7__1061_comb], literal_2051898[p8_res7__1063_comb], literal_2051898[p8_res7__1065_comb], literal_2051898[p8_res7__1067_comb], literal_2051898[p8_res7__1069_comb], literal_2051898[p8_res7__1071_comb], literal_2051898[p8_res7__1073_comb], literal_2051898[p8_res7__1075_comb], literal_2051898[p8_res7__1077_comb], literal_2051898[p8_res7__1079_comb], literal_2051898[p8_res7__1081_comb], literal_2051898[p8_res7__1083_comb], literal_2051898[p8_res7__1085_comb], literal_2051898[p8_res7__1087_comb]};
  assign p8_xor_2052135_comb = p7_k7 ^ p8_permut__33_comb;
  assign p8_array_index_2052158_comb = p7_literal_2043920[p8_xor_2052135_comb[47:40]];
  assign p8_array_index_2052159_comb = p7_literal_2043918[p8_xor_2052135_comb[39:32]];
  assign p8_array_index_2052160_comb = p7_literal_2043916[p8_xor_2052135_comb[31:24]];
  assign p8_array_index_2052161_comb = p7_literal_2043914[p8_xor_2052135_comb[23:16]];
  assign p8_array_index_2052162_comb = p7_literal_2043912[p8_xor_2052135_comb[15:8]];
  assign p8_array_index_2052163_comb = p7_literal_2043910[p8_xor_2052135_comb[7:0]];
  assign p8_res7__1089_comb = p7_literal_2043910[p8_xor_2052135_comb[119:112]] ^ p7_literal_2043912[p8_xor_2052135_comb[111:104]] ^ p7_literal_2043914[p8_xor_2052135_comb[103:96]] ^ p7_literal_2043916[p8_xor_2052135_comb[95:88]] ^ p7_literal_2043918[p8_xor_2052135_comb[87:80]] ^ p7_literal_2043920[p8_xor_2052135_comb[79:72]] ^ p8_xor_2052135_comb[71:64] ^ p7_literal_2043923[p8_xor_2052135_comb[63:56]] ^ p8_xor_2052135_comb[55:48] ^ p8_array_index_2052158_comb ^ p8_array_index_2052159_comb ^ p8_array_index_2052160_comb ^ p8_array_index_2052161_comb ^ p8_array_index_2052162_comb ^ p8_array_index_2052163_comb ^ p8_xor_2052135_comb[127:120];
  assign p8_array_index_2052173_comb = p7_literal_2043920[p8_xor_2052135_comb[39:32]];
  assign p8_array_index_2052174_comb = p7_literal_2043918[p8_xor_2052135_comb[31:24]];
  assign p8_array_index_2052175_comb = p7_literal_2043916[p8_xor_2052135_comb[23:16]];
  assign p8_array_index_2052176_comb = p7_literal_2043914[p8_xor_2052135_comb[15:8]];
  assign p8_array_index_2052177_comb = p7_literal_2043912[p8_xor_2052135_comb[7:0]];
  assign p8_array_index_2052178_comb = p7_literal_2043910[p8_res7__1089_comb];
  assign p8_res7__1091_comb = p7_literal_2043910[p8_xor_2052135_comb[111:104]] ^ p7_literal_2043912[p8_xor_2052135_comb[103:96]] ^ p7_literal_2043914[p8_xor_2052135_comb[95:88]] ^ p7_literal_2043916[p8_xor_2052135_comb[87:80]] ^ p7_literal_2043918[p8_xor_2052135_comb[79:72]] ^ p7_literal_2043920[p8_xor_2052135_comb[71:64]] ^ p8_xor_2052135_comb[63:56] ^ p7_literal_2043923[p8_xor_2052135_comb[55:48]] ^ p8_xor_2052135_comb[47:40] ^ p8_array_index_2052173_comb ^ p8_array_index_2052174_comb ^ p8_array_index_2052175_comb ^ p8_array_index_2052176_comb ^ p8_array_index_2052177_comb ^ p8_array_index_2052178_comb ^ p8_xor_2052135_comb[119:112];
  assign p8_array_index_2052187_comb = p7_literal_2043920[p8_xor_2052135_comb[31:24]];
  assign p8_array_index_2052188_comb = p7_literal_2043918[p8_xor_2052135_comb[23:16]];
  assign p8_array_index_2052189_comb = p7_literal_2043916[p8_xor_2052135_comb[15:8]];
  assign p8_array_index_2052190_comb = p7_literal_2043914[p8_xor_2052135_comb[7:0]];
  assign p8_array_index_2052191_comb = p7_literal_2043912[p8_res7__1089_comb];
  assign p8_res7__1093_comb = p7_literal_2043910[p8_xor_2052135_comb[103:96]] ^ p7_literal_2043912[p8_xor_2052135_comb[95:88]] ^ p7_literal_2043914[p8_xor_2052135_comb[87:80]] ^ p7_literal_2043916[p8_xor_2052135_comb[79:72]] ^ p7_literal_2043918[p8_xor_2052135_comb[71:64]] ^ p7_literal_2043920[p8_xor_2052135_comb[63:56]] ^ p8_xor_2052135_comb[55:48] ^ p7_literal_2043923[p8_xor_2052135_comb[47:40]] ^ p8_xor_2052135_comb[39:32] ^ p8_array_index_2052187_comb ^ p8_array_index_2052188_comb ^ p8_array_index_2052189_comb ^ p8_array_index_2052190_comb ^ p8_array_index_2052191_comb ^ p7_literal_2043910[p8_res7__1091_comb] ^ p8_xor_2052135_comb[111:104];
  assign p8_array_index_2052201_comb = p7_literal_2043920[p8_xor_2052135_comb[23:16]];
  assign p8_array_index_2052202_comb = p7_literal_2043918[p8_xor_2052135_comb[15:8]];
  assign p8_array_index_2052203_comb = p7_literal_2043916[p8_xor_2052135_comb[7:0]];
  assign p8_array_index_2052204_comb = p7_literal_2043914[p8_res7__1089_comb];
  assign p8_array_index_2052205_comb = p7_literal_2043912[p8_res7__1091_comb];
  assign p8_res7__1095_comb = p7_literal_2043910[p8_xor_2052135_comb[95:88]] ^ p7_literal_2043912[p8_xor_2052135_comb[87:80]] ^ p7_literal_2043914[p8_xor_2052135_comb[79:72]] ^ p7_literal_2043916[p8_xor_2052135_comb[71:64]] ^ p7_literal_2043918[p8_xor_2052135_comb[63:56]] ^ p7_literal_2043920[p8_xor_2052135_comb[55:48]] ^ p8_xor_2052135_comb[47:40] ^ p7_literal_2043923[p8_xor_2052135_comb[39:32]] ^ p8_xor_2052135_comb[31:24] ^ p8_array_index_2052201_comb ^ p8_array_index_2052202_comb ^ p8_array_index_2052203_comb ^ p8_array_index_2052204_comb ^ p8_array_index_2052205_comb ^ p7_literal_2043910[p8_res7__1093_comb] ^ p8_xor_2052135_comb[103:96];
  assign p8_array_index_2052214_comb = p7_literal_2043920[p8_xor_2052135_comb[15:8]];
  assign p8_array_index_2052215_comb = p7_literal_2043918[p8_xor_2052135_comb[7:0]];
  assign p8_array_index_2052216_comb = p7_literal_2043916[p8_res7__1089_comb];
  assign p8_array_index_2052217_comb = p7_literal_2043914[p8_res7__1091_comb];
  assign p8_res7__1097_comb = p7_literal_2043910[p8_xor_2052135_comb[87:80]] ^ p7_literal_2043912[p8_xor_2052135_comb[79:72]] ^ p7_literal_2043914[p8_xor_2052135_comb[71:64]] ^ p7_literal_2043916[p8_xor_2052135_comb[63:56]] ^ p7_literal_2043918[p8_xor_2052135_comb[55:48]] ^ p8_array_index_2052158_comb ^ p8_xor_2052135_comb[39:32] ^ p7_literal_2043923[p8_xor_2052135_comb[31:24]] ^ p8_xor_2052135_comb[23:16] ^ p8_array_index_2052214_comb ^ p8_array_index_2052215_comb ^ p8_array_index_2052216_comb ^ p8_array_index_2052217_comb ^ p7_literal_2043912[p8_res7__1093_comb] ^ p7_literal_2043910[p8_res7__1095_comb] ^ p8_xor_2052135_comb[95:88];
  assign p8_array_index_2052227_comb = p7_literal_2043920[p8_xor_2052135_comb[7:0]];
  assign p8_array_index_2052228_comb = p7_literal_2043918[p8_res7__1089_comb];
  assign p8_array_index_2052229_comb = p7_literal_2043916[p8_res7__1091_comb];
  assign p8_array_index_2052230_comb = p7_literal_2043914[p8_res7__1093_comb];
  assign p8_res7__1099_comb = p7_literal_2043910[p8_xor_2052135_comb[79:72]] ^ p7_literal_2043912[p8_xor_2052135_comb[71:64]] ^ p7_literal_2043914[p8_xor_2052135_comb[63:56]] ^ p7_literal_2043916[p8_xor_2052135_comb[55:48]] ^ p7_literal_2043918[p8_xor_2052135_comb[47:40]] ^ p8_array_index_2052173_comb ^ p8_xor_2052135_comb[31:24] ^ p7_literal_2043923[p8_xor_2052135_comb[23:16]] ^ p8_xor_2052135_comb[15:8] ^ p8_array_index_2052227_comb ^ p8_array_index_2052228_comb ^ p8_array_index_2052229_comb ^ p8_array_index_2052230_comb ^ p7_literal_2043912[p8_res7__1095_comb] ^ p7_literal_2043910[p8_res7__1097_comb] ^ p8_xor_2052135_comb[87:80];
  assign p8_array_index_2052239_comb = p7_literal_2043920[p8_res7__1089_comb];
  assign p8_array_index_2052240_comb = p7_literal_2043918[p8_res7__1091_comb];
  assign p8_array_index_2052241_comb = p7_literal_2043916[p8_res7__1093_comb];
  assign p8_res7__1101_comb = p7_literal_2043910[p8_xor_2052135_comb[71:64]] ^ p7_literal_2043912[p8_xor_2052135_comb[63:56]] ^ p7_literal_2043914[p8_xor_2052135_comb[55:48]] ^ p7_literal_2043916[p8_xor_2052135_comb[47:40]] ^ p8_array_index_2052159_comb ^ p8_array_index_2052187_comb ^ p8_xor_2052135_comb[23:16] ^ p7_literal_2043923[p8_xor_2052135_comb[15:8]] ^ p8_xor_2052135_comb[7:0] ^ p8_array_index_2052239_comb ^ p8_array_index_2052240_comb ^ p8_array_index_2052241_comb ^ p7_literal_2043914[p8_res7__1095_comb] ^ p7_literal_2043912[p8_res7__1097_comb] ^ p7_literal_2043910[p8_res7__1099_comb] ^ p8_xor_2052135_comb[79:72];
  assign p8_array_index_2052251_comb = p7_literal_2043920[p8_res7__1091_comb];
  assign p8_array_index_2052252_comb = p7_literal_2043918[p8_res7__1093_comb];
  assign p8_array_index_2052253_comb = p7_literal_2043916[p8_res7__1095_comb];
  assign p8_res7__1103_comb = p7_literal_2043910[p8_xor_2052135_comb[63:56]] ^ p7_literal_2043912[p8_xor_2052135_comb[55:48]] ^ p7_literal_2043914[p8_xor_2052135_comb[47:40]] ^ p7_literal_2043916[p8_xor_2052135_comb[39:32]] ^ p8_array_index_2052174_comb ^ p8_array_index_2052201_comb ^ p8_xor_2052135_comb[15:8] ^ p7_literal_2043923[p8_xor_2052135_comb[7:0]] ^ p8_res7__1089_comb ^ p8_array_index_2052251_comb ^ p8_array_index_2052252_comb ^ p8_array_index_2052253_comb ^ p7_literal_2043914[p8_res7__1097_comb] ^ p7_literal_2043912[p8_res7__1099_comb] ^ p7_literal_2043910[p8_res7__1101_comb] ^ p8_xor_2052135_comb[71:64];
  assign p8_array_index_2052262_comb = p7_literal_2043920[p8_res7__1093_comb];
  assign p8_array_index_2052263_comb = p7_literal_2043918[p8_res7__1095_comb];
  assign p8_res7__1105_comb = p7_literal_2043910[p8_xor_2052135_comb[55:48]] ^ p7_literal_2043912[p8_xor_2052135_comb[47:40]] ^ p7_literal_2043914[p8_xor_2052135_comb[39:32]] ^ p8_array_index_2052160_comb ^ p8_array_index_2052188_comb ^ p8_array_index_2052214_comb ^ p8_xor_2052135_comb[7:0] ^ p7_literal_2043923[p8_res7__1089_comb] ^ p8_res7__1091_comb ^ p8_array_index_2052262_comb ^ p8_array_index_2052263_comb ^ p7_literal_2043916[p8_res7__1097_comb] ^ p7_literal_2043914[p8_res7__1099_comb] ^ p7_literal_2043912[p8_res7__1101_comb] ^ p7_literal_2043910[p8_res7__1103_comb] ^ p8_xor_2052135_comb[63:56];
  assign p8_array_index_2052273_comb = p7_literal_2043920[p8_res7__1095_comb];
  assign p8_array_index_2052274_comb = p7_literal_2043918[p8_res7__1097_comb];
  assign p8_res7__1107_comb = p7_literal_2043910[p8_xor_2052135_comb[47:40]] ^ p7_literal_2043912[p8_xor_2052135_comb[39:32]] ^ p7_literal_2043914[p8_xor_2052135_comb[31:24]] ^ p8_array_index_2052175_comb ^ p8_array_index_2052202_comb ^ p8_array_index_2052227_comb ^ p8_res7__1089_comb ^ p7_literal_2043923[p8_res7__1091_comb] ^ p8_res7__1093_comb ^ p8_array_index_2052273_comb ^ p8_array_index_2052274_comb ^ p7_literal_2043916[p8_res7__1099_comb] ^ p7_literal_2043914[p8_res7__1101_comb] ^ p7_literal_2043912[p8_res7__1103_comb] ^ p7_literal_2043910[p8_res7__1105_comb] ^ p8_xor_2052135_comb[55:48];
  assign p8_array_index_2052283_comb = p7_literal_2043920[p8_res7__1097_comb];
  assign p8_res7__1109_comb = p7_literal_2043910[p8_xor_2052135_comb[39:32]] ^ p7_literal_2043912[p8_xor_2052135_comb[31:24]] ^ p8_array_index_2052161_comb ^ p8_array_index_2052189_comb ^ p8_array_index_2052215_comb ^ p8_array_index_2052239_comb ^ p8_res7__1091_comb ^ p7_literal_2043923[p8_res7__1093_comb] ^ p8_res7__1095_comb ^ p8_array_index_2052283_comb ^ p7_literal_2043918[p8_res7__1099_comb] ^ p7_literal_2043916[p8_res7__1101_comb] ^ p7_literal_2043914[p8_res7__1103_comb] ^ p7_literal_2043912[p8_res7__1105_comb] ^ p7_literal_2043910[p8_res7__1107_comb] ^ p8_xor_2052135_comb[47:40];
  assign p8_array_index_2052293_comb = p7_literal_2043920[p8_res7__1099_comb];
  assign p8_res7__1111_comb = p7_literal_2043910[p8_xor_2052135_comb[31:24]] ^ p7_literal_2043912[p8_xor_2052135_comb[23:16]] ^ p8_array_index_2052176_comb ^ p8_array_index_2052203_comb ^ p8_array_index_2052228_comb ^ p8_array_index_2052251_comb ^ p8_res7__1093_comb ^ p7_literal_2043923[p8_res7__1095_comb] ^ p8_res7__1097_comb ^ p8_array_index_2052293_comb ^ p7_literal_2043918[p8_res7__1101_comb] ^ p7_literal_2043916[p8_res7__1103_comb] ^ p7_literal_2043914[p8_res7__1105_comb] ^ p7_literal_2043912[p8_res7__1107_comb] ^ p7_literal_2043910[p8_res7__1109_comb] ^ p8_xor_2052135_comb[39:32];
  assign p8_res7__1113_comb = p7_literal_2043910[p8_xor_2052135_comb[23:16]] ^ p8_array_index_2052162_comb ^ p8_array_index_2052190_comb ^ p8_array_index_2052216_comb ^ p8_array_index_2052240_comb ^ p8_array_index_2052262_comb ^ p8_res7__1095_comb ^ p7_literal_2043923[p8_res7__1097_comb] ^ p8_res7__1099_comb ^ p7_literal_2043920[p8_res7__1101_comb] ^ p7_literal_2043918[p8_res7__1103_comb] ^ p7_literal_2043916[p8_res7__1105_comb] ^ p7_literal_2043914[p8_res7__1107_comb] ^ p7_literal_2043912[p8_res7__1109_comb] ^ p7_literal_2043910[p8_res7__1111_comb] ^ p8_xor_2052135_comb[31:24];
  assign p8_res7__1115_comb = p7_literal_2043910[p8_xor_2052135_comb[15:8]] ^ p8_array_index_2052177_comb ^ p8_array_index_2052204_comb ^ p8_array_index_2052229_comb ^ p8_array_index_2052252_comb ^ p8_array_index_2052273_comb ^ p8_res7__1097_comb ^ p7_literal_2043923[p8_res7__1099_comb] ^ p8_res7__1101_comb ^ p7_literal_2043920[p8_res7__1103_comb] ^ p7_literal_2043918[p8_res7__1105_comb] ^ p7_literal_2043916[p8_res7__1107_comb] ^ p7_literal_2043914[p8_res7__1109_comb] ^ p7_literal_2043912[p8_res7__1111_comb] ^ p7_literal_2043910[p8_res7__1113_comb] ^ p8_xor_2052135_comb[23:16];
  assign p8_res7__1117_comb = p8_array_index_2052163_comb ^ p8_array_index_2052191_comb ^ p8_array_index_2052217_comb ^ p8_array_index_2052241_comb ^ p8_array_index_2052263_comb ^ p8_array_index_2052283_comb ^ p8_res7__1099_comb ^ p7_literal_2043923[p8_res7__1101_comb] ^ p8_res7__1103_comb ^ p7_literal_2043920[p8_res7__1105_comb] ^ p7_literal_2043918[p8_res7__1107_comb] ^ p7_literal_2043916[p8_res7__1109_comb] ^ p7_literal_2043914[p8_res7__1111_comb] ^ p7_literal_2043912[p8_res7__1113_comb] ^ p7_literal_2043910[p8_res7__1115_comb] ^ p8_xor_2052135_comb[15:8];
  assign p8_res7__1119_comb = p8_array_index_2052178_comb ^ p8_array_index_2052205_comb ^ p8_array_index_2052230_comb ^ p8_array_index_2052253_comb ^ p8_array_index_2052274_comb ^ p8_array_index_2052293_comb ^ p8_res7__1101_comb ^ p7_literal_2043923[p8_res7__1103_comb] ^ p8_res7__1105_comb ^ p7_literal_2043920[p8_res7__1107_comb] ^ p7_literal_2043918[p8_res7__1109_comb] ^ p7_literal_2043916[p8_res7__1111_comb] ^ p7_literal_2043914[p8_res7__1113_comb] ^ p7_literal_2043912[p8_res7__1115_comb] ^ p7_literal_2043910[p8_res7__1117_comb] ^ p8_xor_2052135_comb[7:0];
  assign p8_permut__34_comb = {literal_2051898[p8_res7__1089_comb], literal_2051898[p8_res7__1091_comb], literal_2051898[p8_res7__1093_comb], literal_2051898[p8_res7__1095_comb], literal_2051898[p8_res7__1097_comb], literal_2051898[p8_res7__1099_comb], literal_2051898[p8_res7__1101_comb], literal_2051898[p8_res7__1103_comb], literal_2051898[p8_res7__1105_comb], literal_2051898[p8_res7__1107_comb], literal_2051898[p8_res7__1109_comb], literal_2051898[p8_res7__1111_comb], literal_2051898[p8_res7__1113_comb], literal_2051898[p8_res7__1115_comb], literal_2051898[p8_res7__1117_comb], literal_2051898[p8_res7__1119_comb]};
  assign p8_xor_2052351_comb = p7_k6 ^ p8_permut__34_comb;
  assign p8_array_index_2052374_comb = p7_literal_2043920[p8_xor_2052351_comb[47:40]];
  assign p8_array_index_2052375_comb = p7_literal_2043918[p8_xor_2052351_comb[39:32]];
  assign p8_array_index_2052376_comb = p7_literal_2043916[p8_xor_2052351_comb[31:24]];
  assign p8_array_index_2052377_comb = p7_literal_2043914[p8_xor_2052351_comb[23:16]];
  assign p8_array_index_2052378_comb = p7_literal_2043912[p8_xor_2052351_comb[15:8]];
  assign p8_array_index_2052379_comb = p7_literal_2043910[p8_xor_2052351_comb[7:0]];
  assign p8_res7__1121_comb = p7_literal_2043910[p8_xor_2052351_comb[119:112]] ^ p7_literal_2043912[p8_xor_2052351_comb[111:104]] ^ p7_literal_2043914[p8_xor_2052351_comb[103:96]] ^ p7_literal_2043916[p8_xor_2052351_comb[95:88]] ^ p7_literal_2043918[p8_xor_2052351_comb[87:80]] ^ p7_literal_2043920[p8_xor_2052351_comb[79:72]] ^ p8_xor_2052351_comb[71:64] ^ p7_literal_2043923[p8_xor_2052351_comb[63:56]] ^ p8_xor_2052351_comb[55:48] ^ p8_array_index_2052374_comb ^ p8_array_index_2052375_comb ^ p8_array_index_2052376_comb ^ p8_array_index_2052377_comb ^ p8_array_index_2052378_comb ^ p8_array_index_2052379_comb ^ p8_xor_2052351_comb[127:120];
  assign p8_array_index_2052389_comb = p7_literal_2043920[p8_xor_2052351_comb[39:32]];
  assign p8_array_index_2052390_comb = p7_literal_2043918[p8_xor_2052351_comb[31:24]];
  assign p8_array_index_2052391_comb = p7_literal_2043916[p8_xor_2052351_comb[23:16]];
  assign p8_array_index_2052392_comb = p7_literal_2043914[p8_xor_2052351_comb[15:8]];
  assign p8_array_index_2052393_comb = p7_literal_2043912[p8_xor_2052351_comb[7:0]];
  assign p8_array_index_2052394_comb = p7_literal_2043910[p8_res7__1121_comb];
  assign p8_res7__1123_comb = p7_literal_2043910[p8_xor_2052351_comb[111:104]] ^ p7_literal_2043912[p8_xor_2052351_comb[103:96]] ^ p7_literal_2043914[p8_xor_2052351_comb[95:88]] ^ p7_literal_2043916[p8_xor_2052351_comb[87:80]] ^ p7_literal_2043918[p8_xor_2052351_comb[79:72]] ^ p7_literal_2043920[p8_xor_2052351_comb[71:64]] ^ p8_xor_2052351_comb[63:56] ^ p7_literal_2043923[p8_xor_2052351_comb[55:48]] ^ p8_xor_2052351_comb[47:40] ^ p8_array_index_2052389_comb ^ p8_array_index_2052390_comb ^ p8_array_index_2052391_comb ^ p8_array_index_2052392_comb ^ p8_array_index_2052393_comb ^ p8_array_index_2052394_comb ^ p8_xor_2052351_comb[119:112];
  assign p8_array_index_2052403_comb = p7_literal_2043920[p8_xor_2052351_comb[31:24]];
  assign p8_array_index_2052404_comb = p7_literal_2043918[p8_xor_2052351_comb[23:16]];
  assign p8_array_index_2052405_comb = p7_literal_2043916[p8_xor_2052351_comb[15:8]];
  assign p8_array_index_2052406_comb = p7_literal_2043914[p8_xor_2052351_comb[7:0]];
  assign p8_array_index_2052407_comb = p7_literal_2043912[p8_res7__1121_comb];
  assign p8_res7__1125_comb = p7_literal_2043910[p8_xor_2052351_comb[103:96]] ^ p7_literal_2043912[p8_xor_2052351_comb[95:88]] ^ p7_literal_2043914[p8_xor_2052351_comb[87:80]] ^ p7_literal_2043916[p8_xor_2052351_comb[79:72]] ^ p7_literal_2043918[p8_xor_2052351_comb[71:64]] ^ p7_literal_2043920[p8_xor_2052351_comb[63:56]] ^ p8_xor_2052351_comb[55:48] ^ p7_literal_2043923[p8_xor_2052351_comb[47:40]] ^ p8_xor_2052351_comb[39:32] ^ p8_array_index_2052403_comb ^ p8_array_index_2052404_comb ^ p8_array_index_2052405_comb ^ p8_array_index_2052406_comb ^ p8_array_index_2052407_comb ^ p7_literal_2043910[p8_res7__1123_comb] ^ p8_xor_2052351_comb[111:104];
  assign p8_array_index_2052417_comb = p7_literal_2043920[p8_xor_2052351_comb[23:16]];
  assign p8_array_index_2052418_comb = p7_literal_2043918[p8_xor_2052351_comb[15:8]];
  assign p8_array_index_2052419_comb = p7_literal_2043916[p8_xor_2052351_comb[7:0]];
  assign p8_array_index_2052420_comb = p7_literal_2043914[p8_res7__1121_comb];
  assign p8_array_index_2052421_comb = p7_literal_2043912[p8_res7__1123_comb];
  assign p8_res7__1127_comb = p7_literal_2043910[p8_xor_2052351_comb[95:88]] ^ p7_literal_2043912[p8_xor_2052351_comb[87:80]] ^ p7_literal_2043914[p8_xor_2052351_comb[79:72]] ^ p7_literal_2043916[p8_xor_2052351_comb[71:64]] ^ p7_literal_2043918[p8_xor_2052351_comb[63:56]] ^ p7_literal_2043920[p8_xor_2052351_comb[55:48]] ^ p8_xor_2052351_comb[47:40] ^ p7_literal_2043923[p8_xor_2052351_comb[39:32]] ^ p8_xor_2052351_comb[31:24] ^ p8_array_index_2052417_comb ^ p8_array_index_2052418_comb ^ p8_array_index_2052419_comb ^ p8_array_index_2052420_comb ^ p8_array_index_2052421_comb ^ p7_literal_2043910[p8_res7__1125_comb] ^ p8_xor_2052351_comb[103:96];
  assign p8_array_index_2052430_comb = p7_literal_2043920[p8_xor_2052351_comb[15:8]];
  assign p8_array_index_2052431_comb = p7_literal_2043918[p8_xor_2052351_comb[7:0]];
  assign p8_array_index_2052432_comb = p7_literal_2043916[p8_res7__1121_comb];
  assign p8_array_index_2052433_comb = p7_literal_2043914[p8_res7__1123_comb];
  assign p8_res7__1129_comb = p7_literal_2043910[p8_xor_2052351_comb[87:80]] ^ p7_literal_2043912[p8_xor_2052351_comb[79:72]] ^ p7_literal_2043914[p8_xor_2052351_comb[71:64]] ^ p7_literal_2043916[p8_xor_2052351_comb[63:56]] ^ p7_literal_2043918[p8_xor_2052351_comb[55:48]] ^ p8_array_index_2052374_comb ^ p8_xor_2052351_comb[39:32] ^ p7_literal_2043923[p8_xor_2052351_comb[31:24]] ^ p8_xor_2052351_comb[23:16] ^ p8_array_index_2052430_comb ^ p8_array_index_2052431_comb ^ p8_array_index_2052432_comb ^ p8_array_index_2052433_comb ^ p7_literal_2043912[p8_res7__1125_comb] ^ p7_literal_2043910[p8_res7__1127_comb] ^ p8_xor_2052351_comb[95:88];
  assign p8_array_index_2052443_comb = p7_literal_2043920[p8_xor_2052351_comb[7:0]];
  assign p8_array_index_2052444_comb = p7_literal_2043918[p8_res7__1121_comb];
  assign p8_array_index_2052445_comb = p7_literal_2043916[p8_res7__1123_comb];
  assign p8_array_index_2052446_comb = p7_literal_2043914[p8_res7__1125_comb];
  assign p8_res7__1131_comb = p7_literal_2043910[p8_xor_2052351_comb[79:72]] ^ p7_literal_2043912[p8_xor_2052351_comb[71:64]] ^ p7_literal_2043914[p8_xor_2052351_comb[63:56]] ^ p7_literal_2043916[p8_xor_2052351_comb[55:48]] ^ p7_literal_2043918[p8_xor_2052351_comb[47:40]] ^ p8_array_index_2052389_comb ^ p8_xor_2052351_comb[31:24] ^ p7_literal_2043923[p8_xor_2052351_comb[23:16]] ^ p8_xor_2052351_comb[15:8] ^ p8_array_index_2052443_comb ^ p8_array_index_2052444_comb ^ p8_array_index_2052445_comb ^ p8_array_index_2052446_comb ^ p7_literal_2043912[p8_res7__1127_comb] ^ p7_literal_2043910[p8_res7__1129_comb] ^ p8_xor_2052351_comb[87:80];
  assign p8_array_index_2052455_comb = p7_literal_2043920[p8_res7__1121_comb];
  assign p8_array_index_2052456_comb = p7_literal_2043918[p8_res7__1123_comb];
  assign p8_array_index_2052457_comb = p7_literal_2043916[p8_res7__1125_comb];
  assign p8_res7__1133_comb = p7_literal_2043910[p8_xor_2052351_comb[71:64]] ^ p7_literal_2043912[p8_xor_2052351_comb[63:56]] ^ p7_literal_2043914[p8_xor_2052351_comb[55:48]] ^ p7_literal_2043916[p8_xor_2052351_comb[47:40]] ^ p8_array_index_2052375_comb ^ p8_array_index_2052403_comb ^ p8_xor_2052351_comb[23:16] ^ p7_literal_2043923[p8_xor_2052351_comb[15:8]] ^ p8_xor_2052351_comb[7:0] ^ p8_array_index_2052455_comb ^ p8_array_index_2052456_comb ^ p8_array_index_2052457_comb ^ p7_literal_2043914[p8_res7__1127_comb] ^ p7_literal_2043912[p8_res7__1129_comb] ^ p7_literal_2043910[p8_res7__1131_comb] ^ p8_xor_2052351_comb[79:72];
  assign p8_array_index_2052467_comb = p7_literal_2043920[p8_res7__1123_comb];
  assign p8_array_index_2052468_comb = p7_literal_2043918[p8_res7__1125_comb];
  assign p8_array_index_2052469_comb = p7_literal_2043916[p8_res7__1127_comb];
  assign p8_res7__1135_comb = p7_literal_2043910[p8_xor_2052351_comb[63:56]] ^ p7_literal_2043912[p8_xor_2052351_comb[55:48]] ^ p7_literal_2043914[p8_xor_2052351_comb[47:40]] ^ p7_literal_2043916[p8_xor_2052351_comb[39:32]] ^ p8_array_index_2052390_comb ^ p8_array_index_2052417_comb ^ p8_xor_2052351_comb[15:8] ^ p7_literal_2043923[p8_xor_2052351_comb[7:0]] ^ p8_res7__1121_comb ^ p8_array_index_2052467_comb ^ p8_array_index_2052468_comb ^ p8_array_index_2052469_comb ^ p7_literal_2043914[p8_res7__1129_comb] ^ p7_literal_2043912[p8_res7__1131_comb] ^ p7_literal_2043910[p8_res7__1133_comb] ^ p8_xor_2052351_comb[71:64];
  assign p8_array_index_2052478_comb = p7_literal_2043920[p8_res7__1125_comb];
  assign p8_array_index_2052479_comb = p7_literal_2043918[p8_res7__1127_comb];
  assign p8_res7__1137_comb = p7_literal_2043910[p8_xor_2052351_comb[55:48]] ^ p7_literal_2043912[p8_xor_2052351_comb[47:40]] ^ p7_literal_2043914[p8_xor_2052351_comb[39:32]] ^ p8_array_index_2052376_comb ^ p8_array_index_2052404_comb ^ p8_array_index_2052430_comb ^ p8_xor_2052351_comb[7:0] ^ p7_literal_2043923[p8_res7__1121_comb] ^ p8_res7__1123_comb ^ p8_array_index_2052478_comb ^ p8_array_index_2052479_comb ^ p7_literal_2043916[p8_res7__1129_comb] ^ p7_literal_2043914[p8_res7__1131_comb] ^ p7_literal_2043912[p8_res7__1133_comb] ^ p7_literal_2043910[p8_res7__1135_comb] ^ p8_xor_2052351_comb[63:56];
  assign p8_array_index_2052489_comb = p7_literal_2043920[p8_res7__1127_comb];
  assign p8_array_index_2052490_comb = p7_literal_2043918[p8_res7__1129_comb];
  assign p8_res7__1139_comb = p7_literal_2043910[p8_xor_2052351_comb[47:40]] ^ p7_literal_2043912[p8_xor_2052351_comb[39:32]] ^ p7_literal_2043914[p8_xor_2052351_comb[31:24]] ^ p8_array_index_2052391_comb ^ p8_array_index_2052418_comb ^ p8_array_index_2052443_comb ^ p8_res7__1121_comb ^ p7_literal_2043923[p8_res7__1123_comb] ^ p8_res7__1125_comb ^ p8_array_index_2052489_comb ^ p8_array_index_2052490_comb ^ p7_literal_2043916[p8_res7__1131_comb] ^ p7_literal_2043914[p8_res7__1133_comb] ^ p7_literal_2043912[p8_res7__1135_comb] ^ p7_literal_2043910[p8_res7__1137_comb] ^ p8_xor_2052351_comb[55:48];
  assign p8_array_index_2052499_comb = p7_literal_2043920[p8_res7__1129_comb];
  assign p8_res7__1141_comb = p7_literal_2043910[p8_xor_2052351_comb[39:32]] ^ p7_literal_2043912[p8_xor_2052351_comb[31:24]] ^ p8_array_index_2052377_comb ^ p8_array_index_2052405_comb ^ p8_array_index_2052431_comb ^ p8_array_index_2052455_comb ^ p8_res7__1123_comb ^ p7_literal_2043923[p8_res7__1125_comb] ^ p8_res7__1127_comb ^ p8_array_index_2052499_comb ^ p7_literal_2043918[p8_res7__1131_comb] ^ p7_literal_2043916[p8_res7__1133_comb] ^ p7_literal_2043914[p8_res7__1135_comb] ^ p7_literal_2043912[p8_res7__1137_comb] ^ p7_literal_2043910[p8_res7__1139_comb] ^ p8_xor_2052351_comb[47:40];
  assign p8_array_index_2052509_comb = p7_literal_2043920[p8_res7__1131_comb];
  assign p8_res7__1143_comb = p7_literal_2043910[p8_xor_2052351_comb[31:24]] ^ p7_literal_2043912[p8_xor_2052351_comb[23:16]] ^ p8_array_index_2052392_comb ^ p8_array_index_2052419_comb ^ p8_array_index_2052444_comb ^ p8_array_index_2052467_comb ^ p8_res7__1125_comb ^ p7_literal_2043923[p8_res7__1127_comb] ^ p8_res7__1129_comb ^ p8_array_index_2052509_comb ^ p7_literal_2043918[p8_res7__1133_comb] ^ p7_literal_2043916[p8_res7__1135_comb] ^ p7_literal_2043914[p8_res7__1137_comb] ^ p7_literal_2043912[p8_res7__1139_comb] ^ p7_literal_2043910[p8_res7__1141_comb] ^ p8_xor_2052351_comb[39:32];
  assign p8_res7__1145_comb = p7_literal_2043910[p8_xor_2052351_comb[23:16]] ^ p8_array_index_2052378_comb ^ p8_array_index_2052406_comb ^ p8_array_index_2052432_comb ^ p8_array_index_2052456_comb ^ p8_array_index_2052478_comb ^ p8_res7__1127_comb ^ p7_literal_2043923[p8_res7__1129_comb] ^ p8_res7__1131_comb ^ p7_literal_2043920[p8_res7__1133_comb] ^ p7_literal_2043918[p8_res7__1135_comb] ^ p7_literal_2043916[p8_res7__1137_comb] ^ p7_literal_2043914[p8_res7__1139_comb] ^ p7_literal_2043912[p8_res7__1141_comb] ^ p7_literal_2043910[p8_res7__1143_comb] ^ p8_xor_2052351_comb[31:24];
  assign p8_res7__1147_comb = p7_literal_2043910[p8_xor_2052351_comb[15:8]] ^ p8_array_index_2052393_comb ^ p8_array_index_2052420_comb ^ p8_array_index_2052445_comb ^ p8_array_index_2052468_comb ^ p8_array_index_2052489_comb ^ p8_res7__1129_comb ^ p7_literal_2043923[p8_res7__1131_comb] ^ p8_res7__1133_comb ^ p7_literal_2043920[p8_res7__1135_comb] ^ p7_literal_2043918[p8_res7__1137_comb] ^ p7_literal_2043916[p8_res7__1139_comb] ^ p7_literal_2043914[p8_res7__1141_comb] ^ p7_literal_2043912[p8_res7__1143_comb] ^ p7_literal_2043910[p8_res7__1145_comb] ^ p8_xor_2052351_comb[23:16];
  assign p8_res7__1149_comb = p8_array_index_2052379_comb ^ p8_array_index_2052407_comb ^ p8_array_index_2052433_comb ^ p8_array_index_2052457_comb ^ p8_array_index_2052479_comb ^ p8_array_index_2052499_comb ^ p8_res7__1131_comb ^ p7_literal_2043923[p8_res7__1133_comb] ^ p8_res7__1135_comb ^ p7_literal_2043920[p8_res7__1137_comb] ^ p7_literal_2043918[p8_res7__1139_comb] ^ p7_literal_2043916[p8_res7__1141_comb] ^ p7_literal_2043914[p8_res7__1143_comb] ^ p7_literal_2043912[p8_res7__1145_comb] ^ p7_literal_2043910[p8_res7__1147_comb] ^ p8_xor_2052351_comb[15:8];
  assign p8_res7__1151_comb = p8_array_index_2052394_comb ^ p8_array_index_2052421_comb ^ p8_array_index_2052446_comb ^ p8_array_index_2052469_comb ^ p8_array_index_2052490_comb ^ p8_array_index_2052509_comb ^ p8_res7__1133_comb ^ p7_literal_2043923[p8_res7__1135_comb] ^ p8_res7__1137_comb ^ p7_literal_2043920[p8_res7__1139_comb] ^ p7_literal_2043918[p8_res7__1141_comb] ^ p7_literal_2043916[p8_res7__1143_comb] ^ p7_literal_2043914[p8_res7__1145_comb] ^ p7_literal_2043912[p8_res7__1147_comb] ^ p7_literal_2043910[p8_res7__1149_comb] ^ p8_xor_2052351_comb[7:0];
  assign p8_permut__35_comb = {literal_2051898[p8_res7__1121_comb], literal_2051898[p8_res7__1123_comb], literal_2051898[p8_res7__1125_comb], literal_2051898[p8_res7__1127_comb], literal_2051898[p8_res7__1129_comb], literal_2051898[p8_res7__1131_comb], literal_2051898[p8_res7__1133_comb], literal_2051898[p8_res7__1135_comb], literal_2051898[p8_res7__1137_comb], literal_2051898[p8_res7__1139_comb], literal_2051898[p8_res7__1141_comb], literal_2051898[p8_res7__1143_comb], literal_2051898[p8_res7__1145_comb], literal_2051898[p8_res7__1147_comb], literal_2051898[p8_res7__1149_comb], literal_2051898[p8_res7__1151_comb]};
  assign p8_xor_2052567_comb = p7_k5 ^ p8_permut__35_comb;
  assign p8_bit_slice_2052575_comb = p8_xor_2052567_comb[47:40];
  assign p8_bit_slice_2052576_comb = p8_xor_2052567_comb[39:32];
  assign p8_bit_slice_2052577_comb = p8_xor_2052567_comb[31:24];
  assign p8_bit_slice_2052578_comb = p8_xor_2052567_comb[23:16];
  assign p8_bit_slice_2052579_comb = p8_xor_2052567_comb[15:8];
  assign p8_bit_slice_2052580_comb = p8_xor_2052567_comb[7:0];
  assign p8_bit_slice_2052589_comb = p8_xor_2052567_comb[55:48];
  assign p8_array_index_2052590_comb = p7_literal_2043920[p8_bit_slice_2052575_comb];
  assign p8_array_index_2052591_comb = p7_literal_2043918[p8_bit_slice_2052576_comb];
  assign p8_array_index_2052592_comb = p7_literal_2043916[p8_bit_slice_2052577_comb];
  assign p8_array_index_2052593_comb = p7_literal_2043914[p8_bit_slice_2052578_comb];
  assign p8_array_index_2052594_comb = p7_literal_2043912[p8_bit_slice_2052579_comb];
  assign p8_array_index_2052595_comb = p7_literal_2043910[p8_bit_slice_2052580_comb];
  assign p8_res7__1153_comb = p7_literal_2043910[p8_xor_2052567_comb[119:112]] ^ p7_literal_2043912[p8_xor_2052567_comb[111:104]] ^ p7_literal_2043914[p8_xor_2052567_comb[103:96]] ^ p7_literal_2043916[p8_xor_2052567_comb[95:88]] ^ p7_literal_2043918[p8_xor_2052567_comb[87:80]] ^ p7_literal_2043920[p8_xor_2052567_comb[79:72]] ^ p8_xor_2052567_comb[71:64] ^ p7_literal_2043923[p8_xor_2052567_comb[63:56]] ^ p8_bit_slice_2052589_comb ^ p8_array_index_2052590_comb ^ p8_array_index_2052591_comb ^ p8_array_index_2052592_comb ^ p8_array_index_2052593_comb ^ p8_array_index_2052594_comb ^ p8_array_index_2052595_comb ^ p8_xor_2052567_comb[127:120];
  assign p8_array_index_2052605_comb = p7_literal_2043920[p8_bit_slice_2052576_comb];
  assign p8_array_index_2052606_comb = p7_literal_2043918[p8_bit_slice_2052577_comb];
  assign p8_array_index_2052607_comb = p7_literal_2043916[p8_bit_slice_2052578_comb];
  assign p8_array_index_2052608_comb = p7_literal_2043914[p8_bit_slice_2052579_comb];
  assign p8_array_index_2052609_comb = p7_literal_2043912[p8_bit_slice_2052580_comb];
  assign p8_array_index_2052610_comb = p7_literal_2043910[p8_res7__1153_comb];
  assign p8_res7__1155_comb = p7_literal_2043910[p8_xor_2052567_comb[111:104]] ^ p7_literal_2043912[p8_xor_2052567_comb[103:96]] ^ p7_literal_2043914[p8_xor_2052567_comb[95:88]] ^ p7_literal_2043916[p8_xor_2052567_comb[87:80]] ^ p7_literal_2043918[p8_xor_2052567_comb[79:72]] ^ p7_literal_2043920[p8_xor_2052567_comb[71:64]] ^ p8_xor_2052567_comb[63:56] ^ p7_literal_2043923[p8_bit_slice_2052589_comb] ^ p8_bit_slice_2052575_comb ^ p8_array_index_2052605_comb ^ p8_array_index_2052606_comb ^ p8_array_index_2052607_comb ^ p8_array_index_2052608_comb ^ p8_array_index_2052609_comb ^ p8_array_index_2052610_comb ^ p8_xor_2052567_comb[119:112];
  assign p8_array_index_2052619_comb = p7_literal_2043920[p8_bit_slice_2052577_comb];
  assign p8_array_index_2052620_comb = p7_literal_2043918[p8_bit_slice_2052578_comb];
  assign p8_array_index_2052621_comb = p7_literal_2043916[p8_bit_slice_2052579_comb];
  assign p8_array_index_2052622_comb = p7_literal_2043914[p8_bit_slice_2052580_comb];
  assign p8_array_index_2052623_comb = p7_literal_2043912[p8_res7__1153_comb];
  assign p8_res7__1157_comb = p7_literal_2043910[p8_xor_2052567_comb[103:96]] ^ p7_literal_2043912[p8_xor_2052567_comb[95:88]] ^ p7_literal_2043914[p8_xor_2052567_comb[87:80]] ^ p7_literal_2043916[p8_xor_2052567_comb[79:72]] ^ p7_literal_2043918[p8_xor_2052567_comb[71:64]] ^ p7_literal_2043920[p8_xor_2052567_comb[63:56]] ^ p8_bit_slice_2052589_comb ^ p7_literal_2043923[p8_bit_slice_2052575_comb] ^ p8_bit_slice_2052576_comb ^ p8_array_index_2052619_comb ^ p8_array_index_2052620_comb ^ p8_array_index_2052621_comb ^ p8_array_index_2052622_comb ^ p8_array_index_2052623_comb ^ p7_literal_2043910[p8_res7__1155_comb] ^ p8_xor_2052567_comb[111:104];
  assign p8_array_index_2052633_comb = p7_literal_2043920[p8_bit_slice_2052578_comb];
  assign p8_array_index_2052634_comb = p7_literal_2043918[p8_bit_slice_2052579_comb];
  assign p8_array_index_2052635_comb = p7_literal_2043916[p8_bit_slice_2052580_comb];
  assign p8_array_index_2052636_comb = p7_literal_2043914[p8_res7__1153_comb];
  assign p8_array_index_2052637_comb = p7_literal_2043912[p8_res7__1155_comb];
  assign p8_res7__1159_comb = p7_literal_2043910[p8_xor_2052567_comb[95:88]] ^ p7_literal_2043912[p8_xor_2052567_comb[87:80]] ^ p7_literal_2043914[p8_xor_2052567_comb[79:72]] ^ p7_literal_2043916[p8_xor_2052567_comb[71:64]] ^ p7_literal_2043918[p8_xor_2052567_comb[63:56]] ^ p7_literal_2043920[p8_bit_slice_2052589_comb] ^ p8_bit_slice_2052575_comb ^ p7_literal_2043923[p8_bit_slice_2052576_comb] ^ p8_bit_slice_2052577_comb ^ p8_array_index_2052633_comb ^ p8_array_index_2052634_comb ^ p8_array_index_2052635_comb ^ p8_array_index_2052636_comb ^ p8_array_index_2052637_comb ^ p7_literal_2043910[p8_res7__1157_comb] ^ p8_xor_2052567_comb[103:96];
  assign p8_array_index_2052646_comb = p7_literal_2043920[p8_bit_slice_2052579_comb];
  assign p8_array_index_2052647_comb = p7_literal_2043918[p8_bit_slice_2052580_comb];
  assign p8_array_index_2052648_comb = p7_literal_2043916[p8_res7__1153_comb];
  assign p8_array_index_2052649_comb = p7_literal_2043914[p8_res7__1155_comb];
  assign p8_res7__1161_comb = p7_literal_2043910[p8_xor_2052567_comb[87:80]] ^ p7_literal_2043912[p8_xor_2052567_comb[79:72]] ^ p7_literal_2043914[p8_xor_2052567_comb[71:64]] ^ p7_literal_2043916[p8_xor_2052567_comb[63:56]] ^ p7_literal_2043918[p8_bit_slice_2052589_comb] ^ p8_array_index_2052590_comb ^ p8_bit_slice_2052576_comb ^ p7_literal_2043923[p8_bit_slice_2052577_comb] ^ p8_bit_slice_2052578_comb ^ p8_array_index_2052646_comb ^ p8_array_index_2052647_comb ^ p8_array_index_2052648_comb ^ p8_array_index_2052649_comb ^ p7_literal_2043912[p8_res7__1157_comb] ^ p7_literal_2043910[p8_res7__1159_comb] ^ p8_xor_2052567_comb[95:88];
  assign p8_array_index_2052659_comb = p7_literal_2043920[p8_bit_slice_2052580_comb];
  assign p8_array_index_2052660_comb = p7_literal_2043918[p8_res7__1153_comb];
  assign p8_array_index_2052661_comb = p7_literal_2043916[p8_res7__1155_comb];
  assign p8_array_index_2052662_comb = p7_literal_2043914[p8_res7__1157_comb];
  assign p8_res7__1163_comb = p7_literal_2043910[p8_xor_2052567_comb[79:72]] ^ p7_literal_2043912[p8_xor_2052567_comb[71:64]] ^ p7_literal_2043914[p8_xor_2052567_comb[63:56]] ^ p7_literal_2043916[p8_bit_slice_2052589_comb] ^ p7_literal_2043918[p8_bit_slice_2052575_comb] ^ p8_array_index_2052605_comb ^ p8_bit_slice_2052577_comb ^ p7_literal_2043923[p8_bit_slice_2052578_comb] ^ p8_bit_slice_2052579_comb ^ p8_array_index_2052659_comb ^ p8_array_index_2052660_comb ^ p8_array_index_2052661_comb ^ p8_array_index_2052662_comb ^ p7_literal_2043912[p8_res7__1159_comb] ^ p7_literal_2043910[p8_res7__1161_comb] ^ p8_xor_2052567_comb[87:80];
  assign p8_array_index_2052671_comb = p7_literal_2043920[p8_res7__1153_comb];
  assign p8_array_index_2052672_comb = p7_literal_2043918[p8_res7__1155_comb];
  assign p8_array_index_2052673_comb = p7_literal_2043916[p8_res7__1157_comb];
  assign p8_res7__1165_comb = p7_literal_2043910[p8_xor_2052567_comb[71:64]] ^ p7_literal_2043912[p8_xor_2052567_comb[63:56]] ^ p7_literal_2043914[p8_bit_slice_2052589_comb] ^ p7_literal_2043916[p8_bit_slice_2052575_comb] ^ p8_array_index_2052591_comb ^ p8_array_index_2052619_comb ^ p8_bit_slice_2052578_comb ^ p7_literal_2043923[p8_bit_slice_2052579_comb] ^ p8_bit_slice_2052580_comb ^ p8_array_index_2052671_comb ^ p8_array_index_2052672_comb ^ p8_array_index_2052673_comb ^ p7_literal_2043914[p8_res7__1159_comb] ^ p7_literal_2043912[p8_res7__1161_comb] ^ p7_literal_2043910[p8_res7__1163_comb] ^ p8_xor_2052567_comb[79:72];
  assign p8_array_index_2052683_comb = p7_literal_2043920[p8_res7__1155_comb];
  assign p8_array_index_2052684_comb = p7_literal_2043918[p8_res7__1157_comb];
  assign p8_array_index_2052685_comb = p7_literal_2043916[p8_res7__1159_comb];
  assign p8_res7__1167_comb = p7_literal_2043910[p8_xor_2052567_comb[63:56]] ^ p7_literal_2043912[p8_bit_slice_2052589_comb] ^ p7_literal_2043914[p8_bit_slice_2052575_comb] ^ p7_literal_2043916[p8_bit_slice_2052576_comb] ^ p8_array_index_2052606_comb ^ p8_array_index_2052633_comb ^ p8_bit_slice_2052579_comb ^ p7_literal_2043923[p8_bit_slice_2052580_comb] ^ p8_res7__1153_comb ^ p8_array_index_2052683_comb ^ p8_array_index_2052684_comb ^ p8_array_index_2052685_comb ^ p7_literal_2043914[p8_res7__1161_comb] ^ p7_literal_2043912[p8_res7__1163_comb] ^ p7_literal_2043910[p8_res7__1165_comb] ^ p8_xor_2052567_comb[71:64];
  assign p8_array_index_2052694_comb = p7_literal_2043920[p8_res7__1157_comb];
  assign p8_array_index_2052695_comb = p7_literal_2043918[p8_res7__1159_comb];
  assign p8_res7__1169_comb = p7_literal_2043910[p8_bit_slice_2052589_comb] ^ p7_literal_2043912[p8_bit_slice_2052575_comb] ^ p7_literal_2043914[p8_bit_slice_2052576_comb] ^ p8_array_index_2052592_comb ^ p8_array_index_2052620_comb ^ p8_array_index_2052646_comb ^ p8_bit_slice_2052580_comb ^ p7_literal_2043923[p8_res7__1153_comb] ^ p8_res7__1155_comb ^ p8_array_index_2052694_comb ^ p8_array_index_2052695_comb ^ p7_literal_2043916[p8_res7__1161_comb] ^ p7_literal_2043914[p8_res7__1163_comb] ^ p7_literal_2043912[p8_res7__1165_comb] ^ p7_literal_2043910[p8_res7__1167_comb] ^ p8_xor_2052567_comb[63:56];

  // Registers for pipe stage 8:
  reg [127:0] p8_bit_slice_2043893;
  reg [127:0] p8_bit_slice_2044119;
  reg [127:0] p8_k3;
  reg [127:0] p8_k2;
  reg [127:0] p8_k4;
  reg [7:0] p8_bit_slice_2052575;
  reg [7:0] p8_bit_slice_2052576;
  reg [7:0] p8_bit_slice_2052577;
  reg [7:0] p8_bit_slice_2052578;
  reg [7:0] p8_bit_slice_2052579;
  reg [7:0] p8_bit_slice_2052580;
  reg [7:0] p8_bit_slice_2052589;
  reg [7:0] p8_array_index_2052593;
  reg [7:0] p8_array_index_2052594;
  reg [7:0] p8_array_index_2052595;
  reg [7:0] p8_res7__1153;
  reg [7:0] p8_array_index_2052607;
  reg [7:0] p8_array_index_2052608;
  reg [7:0] p8_array_index_2052609;
  reg [7:0] p8_array_index_2052610;
  reg [7:0] p8_res7__1155;
  reg [7:0] p8_array_index_2052621;
  reg [7:0] p8_array_index_2052622;
  reg [7:0] p8_array_index_2052623;
  reg [7:0] p8_res7__1157;
  reg [7:0] p8_array_index_2052634;
  reg [7:0] p8_array_index_2052635;
  reg [7:0] p8_array_index_2052636;
  reg [7:0] p8_array_index_2052637;
  reg [7:0] p8_res7__1159;
  reg [7:0] p8_array_index_2052647;
  reg [7:0] p8_array_index_2052648;
  reg [7:0] p8_array_index_2052649;
  reg [7:0] p8_res7__1161;
  reg [7:0] p8_array_index_2052659;
  reg [7:0] p8_array_index_2052660;
  reg [7:0] p8_array_index_2052661;
  reg [7:0] p8_array_index_2052662;
  reg [7:0] p8_res7__1163;
  reg [7:0] p8_array_index_2052671;
  reg [7:0] p8_array_index_2052672;
  reg [7:0] p8_array_index_2052673;
  reg [7:0] p8_res7__1165;
  reg [7:0] p8_array_index_2052683;
  reg [7:0] p8_array_index_2052684;
  reg [7:0] p8_array_index_2052685;
  reg [7:0] p8_res7__1167;
  reg [7:0] p8_array_index_2052694;
  reg [7:0] p8_array_index_2052695;
  reg [7:0] p8_res7__1169;
  always_ff @ (posedge clk) begin
    p8_bit_slice_2043893 <= p7_bit_slice_2043893;
    p8_bit_slice_2044119 <= p7_bit_slice_2044119;
    p8_k3 <= p7_k3;
    p8_k2 <= p7_k2;
    p8_k4 <= p7_k4;
    p8_bit_slice_2052575 <= p8_bit_slice_2052575_comb;
    p8_bit_slice_2052576 <= p8_bit_slice_2052576_comb;
    p8_bit_slice_2052577 <= p8_bit_slice_2052577_comb;
    p8_bit_slice_2052578 <= p8_bit_slice_2052578_comb;
    p8_bit_slice_2052579 <= p8_bit_slice_2052579_comb;
    p8_bit_slice_2052580 <= p8_bit_slice_2052580_comb;
    p8_bit_slice_2052589 <= p8_bit_slice_2052589_comb;
    p8_array_index_2052593 <= p8_array_index_2052593_comb;
    p8_array_index_2052594 <= p8_array_index_2052594_comb;
    p8_array_index_2052595 <= p8_array_index_2052595_comb;
    p8_res7__1153 <= p8_res7__1153_comb;
    p8_array_index_2052607 <= p8_array_index_2052607_comb;
    p8_array_index_2052608 <= p8_array_index_2052608_comb;
    p8_array_index_2052609 <= p8_array_index_2052609_comb;
    p8_array_index_2052610 <= p8_array_index_2052610_comb;
    p8_res7__1155 <= p8_res7__1155_comb;
    p8_array_index_2052621 <= p8_array_index_2052621_comb;
    p8_array_index_2052622 <= p8_array_index_2052622_comb;
    p8_array_index_2052623 <= p8_array_index_2052623_comb;
    p8_res7__1157 <= p8_res7__1157_comb;
    p8_array_index_2052634 <= p8_array_index_2052634_comb;
    p8_array_index_2052635 <= p8_array_index_2052635_comb;
    p8_array_index_2052636 <= p8_array_index_2052636_comb;
    p8_array_index_2052637 <= p8_array_index_2052637_comb;
    p8_res7__1159 <= p8_res7__1159_comb;
    p8_array_index_2052647 <= p8_array_index_2052647_comb;
    p8_array_index_2052648 <= p8_array_index_2052648_comb;
    p8_array_index_2052649 <= p8_array_index_2052649_comb;
    p8_res7__1161 <= p8_res7__1161_comb;
    p8_array_index_2052659 <= p8_array_index_2052659_comb;
    p8_array_index_2052660 <= p8_array_index_2052660_comb;
    p8_array_index_2052661 <= p8_array_index_2052661_comb;
    p8_array_index_2052662 <= p8_array_index_2052662_comb;
    p8_res7__1163 <= p8_res7__1163_comb;
    p8_array_index_2052671 <= p8_array_index_2052671_comb;
    p8_array_index_2052672 <= p8_array_index_2052672_comb;
    p8_array_index_2052673 <= p8_array_index_2052673_comb;
    p8_res7__1165 <= p8_res7__1165_comb;
    p8_array_index_2052683 <= p8_array_index_2052683_comb;
    p8_array_index_2052684 <= p8_array_index_2052684_comb;
    p8_array_index_2052685 <= p8_array_index_2052685_comb;
    p8_res7__1167 <= p8_res7__1167_comb;
    p8_array_index_2052694 <= p8_array_index_2052694_comb;
    p8_array_index_2052695 <= p8_array_index_2052695_comb;
    p8_res7__1169 <= p8_res7__1169_comb;
  end

  // ===== Pipe stage 9:
  wire [7:0] p9_array_index_2052821_comb;
  wire [7:0] p9_array_index_2052822_comb;
  wire [7:0] p9_res7__1171_comb;
  wire [7:0] p9_array_index_2052831_comb;
  wire [7:0] p9_res7__1173_comb;
  wire [7:0] p9_array_index_2052841_comb;
  wire [7:0] p9_res7__1175_comb;
  wire [7:0] p9_res7__1177_comb;
  wire [7:0] p9_res7__1179_comb;
  wire [7:0] p9_res7__1181_comb;
  wire [7:0] p9_res7__1183_comb;
  wire [127:0] p9_permut__36_comb;
  wire [127:0] p9_xor_2052899_comb;
  wire [7:0] p9_array_index_2052922_comb;
  wire [7:0] p9_array_index_2052923_comb;
  wire [7:0] p9_array_index_2052924_comb;
  wire [7:0] p9_array_index_2052925_comb;
  wire [7:0] p9_array_index_2052926_comb;
  wire [7:0] p9_array_index_2052927_comb;
  wire [7:0] p9_res7__1185_comb;
  wire [7:0] p9_array_index_2052937_comb;
  wire [7:0] p9_array_index_2052938_comb;
  wire [7:0] p9_array_index_2052939_comb;
  wire [7:0] p9_array_index_2052940_comb;
  wire [7:0] p9_array_index_2052941_comb;
  wire [7:0] p9_array_index_2052942_comb;
  wire [7:0] p9_res7__1187_comb;
  wire [7:0] p9_array_index_2052951_comb;
  wire [7:0] p9_array_index_2052952_comb;
  wire [7:0] p9_array_index_2052953_comb;
  wire [7:0] p9_array_index_2052954_comb;
  wire [7:0] p9_array_index_2052955_comb;
  wire [7:0] p9_res7__1189_comb;
  wire [7:0] p9_array_index_2052965_comb;
  wire [7:0] p9_array_index_2052966_comb;
  wire [7:0] p9_array_index_2052967_comb;
  wire [7:0] p9_array_index_2052968_comb;
  wire [7:0] p9_array_index_2052969_comb;
  wire [7:0] p9_res7__1191_comb;
  wire [7:0] p9_array_index_2052978_comb;
  wire [7:0] p9_array_index_2052979_comb;
  wire [7:0] p9_array_index_2052980_comb;
  wire [7:0] p9_array_index_2052981_comb;
  wire [7:0] p9_res7__1193_comb;
  wire [7:0] p9_array_index_2052991_comb;
  wire [7:0] p9_array_index_2052992_comb;
  wire [7:0] p9_array_index_2052993_comb;
  wire [7:0] p9_array_index_2052994_comb;
  wire [7:0] p9_res7__1195_comb;
  wire [7:0] p9_array_index_2053003_comb;
  wire [7:0] p9_array_index_2053004_comb;
  wire [7:0] p9_array_index_2053005_comb;
  wire [7:0] p9_res7__1197_comb;
  wire [7:0] p9_array_index_2053015_comb;
  wire [7:0] p9_array_index_2053016_comb;
  wire [7:0] p9_array_index_2053017_comb;
  wire [7:0] p9_res7__1199_comb;
  wire [7:0] p9_array_index_2053026_comb;
  wire [7:0] p9_array_index_2053027_comb;
  wire [7:0] p9_res7__1201_comb;
  wire [7:0] p9_array_index_2053037_comb;
  wire [7:0] p9_array_index_2053038_comb;
  wire [7:0] p9_res7__1203_comb;
  wire [7:0] p9_array_index_2053047_comb;
  wire [7:0] p9_res7__1205_comb;
  wire [7:0] p9_array_index_2053057_comb;
  wire [7:0] p9_res7__1207_comb;
  wire [7:0] p9_res7__1209_comb;
  wire [7:0] p9_res7__1211_comb;
  wire [7:0] p9_res7__1213_comb;
  wire [7:0] p9_res7__1215_comb;
  wire [127:0] p9_permut__37_comb;
  wire [127:0] p9_xor_2053115_comb;
  wire [7:0] p9_array_index_2053138_comb;
  wire [7:0] p9_array_index_2053139_comb;
  wire [7:0] p9_array_index_2053140_comb;
  wire [7:0] p9_array_index_2053141_comb;
  wire [7:0] p9_array_index_2053142_comb;
  wire [7:0] p9_array_index_2053143_comb;
  wire [7:0] p9_res7__1217_comb;
  wire [7:0] p9_array_index_2053153_comb;
  wire [7:0] p9_array_index_2053154_comb;
  wire [7:0] p9_array_index_2053155_comb;
  wire [7:0] p9_array_index_2053156_comb;
  wire [7:0] p9_array_index_2053157_comb;
  wire [7:0] p9_array_index_2053158_comb;
  wire [7:0] p9_res7__1219_comb;
  wire [7:0] p9_array_index_2053167_comb;
  wire [7:0] p9_array_index_2053168_comb;
  wire [7:0] p9_array_index_2053169_comb;
  wire [7:0] p9_array_index_2053170_comb;
  wire [7:0] p9_array_index_2053171_comb;
  wire [7:0] p9_res7__1221_comb;
  wire [7:0] p9_array_index_2053181_comb;
  wire [7:0] p9_array_index_2053182_comb;
  wire [7:0] p9_array_index_2053183_comb;
  wire [7:0] p9_array_index_2053184_comb;
  wire [7:0] p9_array_index_2053185_comb;
  wire [7:0] p9_res7__1223_comb;
  wire [7:0] p9_array_index_2053194_comb;
  wire [7:0] p9_array_index_2053195_comb;
  wire [7:0] p9_array_index_2053196_comb;
  wire [7:0] p9_array_index_2053197_comb;
  wire [7:0] p9_res7__1225_comb;
  wire [7:0] p9_array_index_2053207_comb;
  wire [7:0] p9_array_index_2053208_comb;
  wire [7:0] p9_array_index_2053209_comb;
  wire [7:0] p9_array_index_2053210_comb;
  wire [7:0] p9_res7__1227_comb;
  wire [7:0] p9_array_index_2053219_comb;
  wire [7:0] p9_array_index_2053220_comb;
  wire [7:0] p9_array_index_2053221_comb;
  wire [7:0] p9_res7__1229_comb;
  wire [7:0] p9_array_index_2053231_comb;
  wire [7:0] p9_array_index_2053232_comb;
  wire [7:0] p9_array_index_2053233_comb;
  wire [7:0] p9_res7__1231_comb;
  wire [7:0] p9_array_index_2053242_comb;
  wire [7:0] p9_array_index_2053243_comb;
  wire [7:0] p9_res7__1233_comb;
  wire [7:0] p9_array_index_2053253_comb;
  wire [7:0] p9_array_index_2053254_comb;
  wire [7:0] p9_res7__1235_comb;
  wire [7:0] p9_array_index_2053263_comb;
  wire [7:0] p9_res7__1237_comb;
  wire [7:0] p9_array_index_2053273_comb;
  wire [7:0] p9_res7__1239_comb;
  wire [7:0] p9_res7__1241_comb;
  wire [7:0] p9_res7__1243_comb;
  wire [7:0] p9_res7__1245_comb;
  wire [7:0] p9_res7__1247_comb;
  wire [127:0] p9_permut__38_comb;
  wire [127:0] p9_xor_2053331_comb;
  wire [7:0] p9_array_index_2053354_comb;
  wire [7:0] p9_array_index_2053355_comb;
  wire [7:0] p9_array_index_2053356_comb;
  wire [7:0] p9_array_index_2053357_comb;
  wire [7:0] p9_array_index_2053358_comb;
  wire [7:0] p9_array_index_2053359_comb;
  wire [7:0] p9_res7__1249_comb;
  wire [7:0] p9_array_index_2053369_comb;
  wire [7:0] p9_array_index_2053370_comb;
  wire [7:0] p9_array_index_2053371_comb;
  wire [7:0] p9_array_index_2053372_comb;
  wire [7:0] p9_array_index_2053373_comb;
  wire [7:0] p9_array_index_2053374_comb;
  wire [7:0] p9_res7__1251_comb;
  wire [7:0] p9_array_index_2053383_comb;
  wire [7:0] p9_array_index_2053384_comb;
  wire [7:0] p9_array_index_2053385_comb;
  wire [7:0] p9_array_index_2053386_comb;
  wire [7:0] p9_array_index_2053387_comb;
  wire [7:0] p9_res7__1253_comb;
  wire [7:0] p9_array_index_2053397_comb;
  wire [7:0] p9_array_index_2053398_comb;
  wire [7:0] p9_array_index_2053399_comb;
  wire [7:0] p9_array_index_2053400_comb;
  wire [7:0] p9_array_index_2053401_comb;
  wire [7:0] p9_res7__1255_comb;
  wire [7:0] p9_array_index_2053410_comb;
  wire [7:0] p9_array_index_2053411_comb;
  wire [7:0] p9_array_index_2053412_comb;
  wire [7:0] p9_array_index_2053413_comb;
  wire [7:0] p9_res7__1257_comb;
  wire [7:0] p9_array_index_2053423_comb;
  wire [7:0] p9_array_index_2053424_comb;
  wire [7:0] p9_array_index_2053425_comb;
  wire [7:0] p9_array_index_2053426_comb;
  wire [7:0] p9_res7__1259_comb;
  wire [7:0] p9_array_index_2053435_comb;
  wire [7:0] p9_array_index_2053436_comb;
  wire [7:0] p9_array_index_2053437_comb;
  wire [7:0] p9_res7__1261_comb;
  wire [7:0] p9_array_index_2053447_comb;
  wire [7:0] p9_array_index_2053448_comb;
  wire [7:0] p9_array_index_2053449_comb;
  wire [7:0] p9_res7__1263_comb;
  wire [7:0] p9_array_index_2053458_comb;
  wire [7:0] p9_array_index_2053459_comb;
  wire [7:0] p9_res7__1265_comb;
  wire [7:0] p9_array_index_2053469_comb;
  wire [7:0] p9_array_index_2053470_comb;
  wire [7:0] p9_res7__1267_comb;
  wire [7:0] p9_array_index_2053479_comb;
  wire [7:0] p9_res7__1269_comb;
  wire [7:0] p9_array_index_2053489_comb;
  wire [7:0] p9_res7__1271_comb;
  wire [7:0] p9_res7__1273_comb;
  wire [7:0] p9_res7__1275_comb;
  wire [7:0] p9_res7__1277_comb;
  wire [7:0] p9_res7__1279_comb;
  wire [127:0] p9_permut__39_comb;
  wire [127:0] p9_xor_2053547_comb;
  wire [7:0] p9_array_index_2053570_comb;
  wire [7:0] p9_array_index_2053571_comb;
  wire [7:0] p9_array_index_2053572_comb;
  wire [7:0] p9_array_index_2053573_comb;
  wire [7:0] p9_array_index_2053574_comb;
  wire [7:0] p9_array_index_2053575_comb;
  wire [7:0] p9_res7__1281_comb;
  wire [7:0] p9_array_index_2053585_comb;
  wire [7:0] p9_array_index_2053586_comb;
  wire [7:0] p9_array_index_2053587_comb;
  wire [7:0] p9_array_index_2053588_comb;
  wire [7:0] p9_array_index_2053589_comb;
  wire [7:0] p9_array_index_2053590_comb;
  wire [7:0] p9_res7__1283_comb;
  wire [7:0] p9_array_index_2053599_comb;
  wire [7:0] p9_array_index_2053600_comb;
  wire [7:0] p9_array_index_2053601_comb;
  wire [7:0] p9_array_index_2053602_comb;
  wire [7:0] p9_array_index_2053603_comb;
  wire [7:0] p9_res7__1285_comb;
  wire [7:0] p9_array_index_2053613_comb;
  wire [7:0] p9_array_index_2053614_comb;
  wire [7:0] p9_array_index_2053615_comb;
  wire [7:0] p9_array_index_2053616_comb;
  wire [7:0] p9_array_index_2053617_comb;
  wire [7:0] p9_res7__1287_comb;
  wire [7:0] p9_array_index_2053626_comb;
  wire [7:0] p9_array_index_2053627_comb;
  wire [7:0] p9_array_index_2053628_comb;
  wire [7:0] p9_array_index_2053629_comb;
  wire [7:0] p9_res7__1289_comb;
  wire [7:0] p9_array_index_2053639_comb;
  wire [7:0] p9_array_index_2053640_comb;
  wire [7:0] p9_array_index_2053641_comb;
  wire [7:0] p9_array_index_2053642_comb;
  wire [7:0] p9_res7__1291_comb;
  wire [7:0] p9_array_index_2053651_comb;
  wire [7:0] p9_array_index_2053652_comb;
  wire [7:0] p9_array_index_2053653_comb;
  wire [7:0] p9_res7__1293_comb;
  wire [7:0] p9_array_index_2053663_comb;
  wire [7:0] p9_array_index_2053664_comb;
  wire [7:0] p9_array_index_2053665_comb;
  wire [7:0] p9_res7__1295_comb;
  wire [7:0] p9_array_index_2053674_comb;
  wire [7:0] p9_array_index_2053675_comb;
  wire [7:0] p9_res7__1297_comb;
  wire [7:0] p9_array_index_2053685_comb;
  wire [7:0] p9_array_index_2053686_comb;
  wire [7:0] p9_res7__1299_comb;
  wire [7:0] p9_array_index_2053695_comb;
  wire [7:0] p9_res7__1301_comb;
  wire [7:0] p9_array_index_2053705_comb;
  wire [7:0] p9_res7__1303_comb;
  wire [7:0] p9_res7__1305_comb;
  wire [7:0] p9_res7__1307_comb;
  wire [7:0] p9_res7__1309_comb;
  wire [7:0] p9_res7__1311_comb;
  wire [127:0] p9_permut__40_comb;
  wire [127:0] p9_newValue_comb;
  assign p9_array_index_2052821_comb = p8_literal_2043920[p8_res7__1159];
  assign p9_array_index_2052822_comb = p8_literal_2043918[p8_res7__1161];
  assign p9_res7__1171_comb = p8_literal_2043910[p8_bit_slice_2052575] ^ p8_literal_2043912[p8_bit_slice_2052576] ^ p8_literal_2043914[p8_bit_slice_2052577] ^ p8_array_index_2052607 ^ p8_array_index_2052634 ^ p8_array_index_2052659 ^ p8_res7__1153 ^ p8_literal_2043923[p8_res7__1155] ^ p8_res7__1157 ^ p9_array_index_2052821_comb ^ p9_array_index_2052822_comb ^ p8_literal_2043916[p8_res7__1163] ^ p8_literal_2043914[p8_res7__1165] ^ p8_literal_2043912[p8_res7__1167] ^ p8_literal_2043910[p8_res7__1169] ^ p8_bit_slice_2052589;
  assign p9_array_index_2052831_comb = p8_literal_2043920[p8_res7__1161];
  assign p9_res7__1173_comb = p8_literal_2043910[p8_bit_slice_2052576] ^ p8_literal_2043912[p8_bit_slice_2052577] ^ p8_array_index_2052593 ^ p8_array_index_2052621 ^ p8_array_index_2052647 ^ p8_array_index_2052671 ^ p8_res7__1155 ^ p8_literal_2043923[p8_res7__1157] ^ p8_res7__1159 ^ p9_array_index_2052831_comb ^ p8_literal_2043918[p8_res7__1163] ^ p8_literal_2043916[p8_res7__1165] ^ p8_literal_2043914[p8_res7__1167] ^ p8_literal_2043912[p8_res7__1169] ^ p8_literal_2043910[p9_res7__1171_comb] ^ p8_bit_slice_2052575;
  assign p9_array_index_2052841_comb = p8_literal_2043920[p8_res7__1163];
  assign p9_res7__1175_comb = p8_literal_2043910[p8_bit_slice_2052577] ^ p8_literal_2043912[p8_bit_slice_2052578] ^ p8_array_index_2052608 ^ p8_array_index_2052635 ^ p8_array_index_2052660 ^ p8_array_index_2052683 ^ p8_res7__1157 ^ p8_literal_2043923[p8_res7__1159] ^ p8_res7__1161 ^ p9_array_index_2052841_comb ^ p8_literal_2043918[p8_res7__1165] ^ p8_literal_2043916[p8_res7__1167] ^ p8_literal_2043914[p8_res7__1169] ^ p8_literal_2043912[p9_res7__1171_comb] ^ p8_literal_2043910[p9_res7__1173_comb] ^ p8_bit_slice_2052576;
  assign p9_res7__1177_comb = p8_literal_2043910[p8_bit_slice_2052578] ^ p8_array_index_2052594 ^ p8_array_index_2052622 ^ p8_array_index_2052648 ^ p8_array_index_2052672 ^ p8_array_index_2052694 ^ p8_res7__1159 ^ p8_literal_2043923[p8_res7__1161] ^ p8_res7__1163 ^ p8_literal_2043920[p8_res7__1165] ^ p8_literal_2043918[p8_res7__1167] ^ p8_literal_2043916[p8_res7__1169] ^ p8_literal_2043914[p9_res7__1171_comb] ^ p8_literal_2043912[p9_res7__1173_comb] ^ p8_literal_2043910[p9_res7__1175_comb] ^ p8_bit_slice_2052577;
  assign p9_res7__1179_comb = p8_literal_2043910[p8_bit_slice_2052579] ^ p8_array_index_2052609 ^ p8_array_index_2052636 ^ p8_array_index_2052661 ^ p8_array_index_2052684 ^ p9_array_index_2052821_comb ^ p8_res7__1161 ^ p8_literal_2043923[p8_res7__1163] ^ p8_res7__1165 ^ p8_literal_2043920[p8_res7__1167] ^ p8_literal_2043918[p8_res7__1169] ^ p8_literal_2043916[p9_res7__1171_comb] ^ p8_literal_2043914[p9_res7__1173_comb] ^ p8_literal_2043912[p9_res7__1175_comb] ^ p8_literal_2043910[p9_res7__1177_comb] ^ p8_bit_slice_2052578;
  assign p9_res7__1181_comb = p8_array_index_2052595 ^ p8_array_index_2052623 ^ p8_array_index_2052649 ^ p8_array_index_2052673 ^ p8_array_index_2052695 ^ p9_array_index_2052831_comb ^ p8_res7__1163 ^ p8_literal_2043923[p8_res7__1165] ^ p8_res7__1167 ^ p8_literal_2043920[p8_res7__1169] ^ p8_literal_2043918[p9_res7__1171_comb] ^ p8_literal_2043916[p9_res7__1173_comb] ^ p8_literal_2043914[p9_res7__1175_comb] ^ p8_literal_2043912[p9_res7__1177_comb] ^ p8_literal_2043910[p9_res7__1179_comb] ^ p8_bit_slice_2052579;
  assign p9_res7__1183_comb = p8_array_index_2052610 ^ p8_array_index_2052637 ^ p8_array_index_2052662 ^ p8_array_index_2052685 ^ p9_array_index_2052822_comb ^ p9_array_index_2052841_comb ^ p8_res7__1165 ^ p8_literal_2043923[p8_res7__1167] ^ p8_res7__1169 ^ p8_literal_2043920[p9_res7__1171_comb] ^ p8_literal_2043918[p9_res7__1173_comb] ^ p8_literal_2043916[p9_res7__1175_comb] ^ p8_literal_2043914[p9_res7__1177_comb] ^ p8_literal_2043912[p9_res7__1179_comb] ^ p8_literal_2043910[p9_res7__1181_comb] ^ p8_bit_slice_2052580;
  assign p9_permut__36_comb = {p8_literal_2051898[p8_res7__1153], p8_literal_2051898[p8_res7__1155], p8_literal_2051898[p8_res7__1157], p8_literal_2051898[p8_res7__1159], p8_literal_2051898[p8_res7__1161], p8_literal_2051898[p8_res7__1163], p8_literal_2051898[p8_res7__1165], p8_literal_2051898[p8_res7__1167], p8_literal_2051898[p8_res7__1169], p8_literal_2051898[p9_res7__1171_comb], p8_literal_2051898[p9_res7__1173_comb], p8_literal_2051898[p9_res7__1175_comb], p8_literal_2051898[p9_res7__1177_comb], p8_literal_2051898[p9_res7__1179_comb], p8_literal_2051898[p9_res7__1181_comb], p8_literal_2051898[p9_res7__1183_comb]};
  assign p9_xor_2052899_comb = p8_k4 ^ p9_permut__36_comb;
  assign p9_array_index_2052922_comb = p8_literal_2043920[p9_xor_2052899_comb[47:40]];
  assign p9_array_index_2052923_comb = p8_literal_2043918[p9_xor_2052899_comb[39:32]];
  assign p9_array_index_2052924_comb = p8_literal_2043916[p9_xor_2052899_comb[31:24]];
  assign p9_array_index_2052925_comb = p8_literal_2043914[p9_xor_2052899_comb[23:16]];
  assign p9_array_index_2052926_comb = p8_literal_2043912[p9_xor_2052899_comb[15:8]];
  assign p9_array_index_2052927_comb = p8_literal_2043910[p9_xor_2052899_comb[7:0]];
  assign p9_res7__1185_comb = p8_literal_2043910[p9_xor_2052899_comb[119:112]] ^ p8_literal_2043912[p9_xor_2052899_comb[111:104]] ^ p8_literal_2043914[p9_xor_2052899_comb[103:96]] ^ p8_literal_2043916[p9_xor_2052899_comb[95:88]] ^ p8_literal_2043918[p9_xor_2052899_comb[87:80]] ^ p8_literal_2043920[p9_xor_2052899_comb[79:72]] ^ p9_xor_2052899_comb[71:64] ^ p8_literal_2043923[p9_xor_2052899_comb[63:56]] ^ p9_xor_2052899_comb[55:48] ^ p9_array_index_2052922_comb ^ p9_array_index_2052923_comb ^ p9_array_index_2052924_comb ^ p9_array_index_2052925_comb ^ p9_array_index_2052926_comb ^ p9_array_index_2052927_comb ^ p9_xor_2052899_comb[127:120];
  assign p9_array_index_2052937_comb = p8_literal_2043920[p9_xor_2052899_comb[39:32]];
  assign p9_array_index_2052938_comb = p8_literal_2043918[p9_xor_2052899_comb[31:24]];
  assign p9_array_index_2052939_comb = p8_literal_2043916[p9_xor_2052899_comb[23:16]];
  assign p9_array_index_2052940_comb = p8_literal_2043914[p9_xor_2052899_comb[15:8]];
  assign p9_array_index_2052941_comb = p8_literal_2043912[p9_xor_2052899_comb[7:0]];
  assign p9_array_index_2052942_comb = p8_literal_2043910[p9_res7__1185_comb];
  assign p9_res7__1187_comb = p8_literal_2043910[p9_xor_2052899_comb[111:104]] ^ p8_literal_2043912[p9_xor_2052899_comb[103:96]] ^ p8_literal_2043914[p9_xor_2052899_comb[95:88]] ^ p8_literal_2043916[p9_xor_2052899_comb[87:80]] ^ p8_literal_2043918[p9_xor_2052899_comb[79:72]] ^ p8_literal_2043920[p9_xor_2052899_comb[71:64]] ^ p9_xor_2052899_comb[63:56] ^ p8_literal_2043923[p9_xor_2052899_comb[55:48]] ^ p9_xor_2052899_comb[47:40] ^ p9_array_index_2052937_comb ^ p9_array_index_2052938_comb ^ p9_array_index_2052939_comb ^ p9_array_index_2052940_comb ^ p9_array_index_2052941_comb ^ p9_array_index_2052942_comb ^ p9_xor_2052899_comb[119:112];
  assign p9_array_index_2052951_comb = p8_literal_2043920[p9_xor_2052899_comb[31:24]];
  assign p9_array_index_2052952_comb = p8_literal_2043918[p9_xor_2052899_comb[23:16]];
  assign p9_array_index_2052953_comb = p8_literal_2043916[p9_xor_2052899_comb[15:8]];
  assign p9_array_index_2052954_comb = p8_literal_2043914[p9_xor_2052899_comb[7:0]];
  assign p9_array_index_2052955_comb = p8_literal_2043912[p9_res7__1185_comb];
  assign p9_res7__1189_comb = p8_literal_2043910[p9_xor_2052899_comb[103:96]] ^ p8_literal_2043912[p9_xor_2052899_comb[95:88]] ^ p8_literal_2043914[p9_xor_2052899_comb[87:80]] ^ p8_literal_2043916[p9_xor_2052899_comb[79:72]] ^ p8_literal_2043918[p9_xor_2052899_comb[71:64]] ^ p8_literal_2043920[p9_xor_2052899_comb[63:56]] ^ p9_xor_2052899_comb[55:48] ^ p8_literal_2043923[p9_xor_2052899_comb[47:40]] ^ p9_xor_2052899_comb[39:32] ^ p9_array_index_2052951_comb ^ p9_array_index_2052952_comb ^ p9_array_index_2052953_comb ^ p9_array_index_2052954_comb ^ p9_array_index_2052955_comb ^ p8_literal_2043910[p9_res7__1187_comb] ^ p9_xor_2052899_comb[111:104];
  assign p9_array_index_2052965_comb = p8_literal_2043920[p9_xor_2052899_comb[23:16]];
  assign p9_array_index_2052966_comb = p8_literal_2043918[p9_xor_2052899_comb[15:8]];
  assign p9_array_index_2052967_comb = p8_literal_2043916[p9_xor_2052899_comb[7:0]];
  assign p9_array_index_2052968_comb = p8_literal_2043914[p9_res7__1185_comb];
  assign p9_array_index_2052969_comb = p8_literal_2043912[p9_res7__1187_comb];
  assign p9_res7__1191_comb = p8_literal_2043910[p9_xor_2052899_comb[95:88]] ^ p8_literal_2043912[p9_xor_2052899_comb[87:80]] ^ p8_literal_2043914[p9_xor_2052899_comb[79:72]] ^ p8_literal_2043916[p9_xor_2052899_comb[71:64]] ^ p8_literal_2043918[p9_xor_2052899_comb[63:56]] ^ p8_literal_2043920[p9_xor_2052899_comb[55:48]] ^ p9_xor_2052899_comb[47:40] ^ p8_literal_2043923[p9_xor_2052899_comb[39:32]] ^ p9_xor_2052899_comb[31:24] ^ p9_array_index_2052965_comb ^ p9_array_index_2052966_comb ^ p9_array_index_2052967_comb ^ p9_array_index_2052968_comb ^ p9_array_index_2052969_comb ^ p8_literal_2043910[p9_res7__1189_comb] ^ p9_xor_2052899_comb[103:96];
  assign p9_array_index_2052978_comb = p8_literal_2043920[p9_xor_2052899_comb[15:8]];
  assign p9_array_index_2052979_comb = p8_literal_2043918[p9_xor_2052899_comb[7:0]];
  assign p9_array_index_2052980_comb = p8_literal_2043916[p9_res7__1185_comb];
  assign p9_array_index_2052981_comb = p8_literal_2043914[p9_res7__1187_comb];
  assign p9_res7__1193_comb = p8_literal_2043910[p9_xor_2052899_comb[87:80]] ^ p8_literal_2043912[p9_xor_2052899_comb[79:72]] ^ p8_literal_2043914[p9_xor_2052899_comb[71:64]] ^ p8_literal_2043916[p9_xor_2052899_comb[63:56]] ^ p8_literal_2043918[p9_xor_2052899_comb[55:48]] ^ p9_array_index_2052922_comb ^ p9_xor_2052899_comb[39:32] ^ p8_literal_2043923[p9_xor_2052899_comb[31:24]] ^ p9_xor_2052899_comb[23:16] ^ p9_array_index_2052978_comb ^ p9_array_index_2052979_comb ^ p9_array_index_2052980_comb ^ p9_array_index_2052981_comb ^ p8_literal_2043912[p9_res7__1189_comb] ^ p8_literal_2043910[p9_res7__1191_comb] ^ p9_xor_2052899_comb[95:88];
  assign p9_array_index_2052991_comb = p8_literal_2043920[p9_xor_2052899_comb[7:0]];
  assign p9_array_index_2052992_comb = p8_literal_2043918[p9_res7__1185_comb];
  assign p9_array_index_2052993_comb = p8_literal_2043916[p9_res7__1187_comb];
  assign p9_array_index_2052994_comb = p8_literal_2043914[p9_res7__1189_comb];
  assign p9_res7__1195_comb = p8_literal_2043910[p9_xor_2052899_comb[79:72]] ^ p8_literal_2043912[p9_xor_2052899_comb[71:64]] ^ p8_literal_2043914[p9_xor_2052899_comb[63:56]] ^ p8_literal_2043916[p9_xor_2052899_comb[55:48]] ^ p8_literal_2043918[p9_xor_2052899_comb[47:40]] ^ p9_array_index_2052937_comb ^ p9_xor_2052899_comb[31:24] ^ p8_literal_2043923[p9_xor_2052899_comb[23:16]] ^ p9_xor_2052899_comb[15:8] ^ p9_array_index_2052991_comb ^ p9_array_index_2052992_comb ^ p9_array_index_2052993_comb ^ p9_array_index_2052994_comb ^ p8_literal_2043912[p9_res7__1191_comb] ^ p8_literal_2043910[p9_res7__1193_comb] ^ p9_xor_2052899_comb[87:80];
  assign p9_array_index_2053003_comb = p8_literal_2043920[p9_res7__1185_comb];
  assign p9_array_index_2053004_comb = p8_literal_2043918[p9_res7__1187_comb];
  assign p9_array_index_2053005_comb = p8_literal_2043916[p9_res7__1189_comb];
  assign p9_res7__1197_comb = p8_literal_2043910[p9_xor_2052899_comb[71:64]] ^ p8_literal_2043912[p9_xor_2052899_comb[63:56]] ^ p8_literal_2043914[p9_xor_2052899_comb[55:48]] ^ p8_literal_2043916[p9_xor_2052899_comb[47:40]] ^ p9_array_index_2052923_comb ^ p9_array_index_2052951_comb ^ p9_xor_2052899_comb[23:16] ^ p8_literal_2043923[p9_xor_2052899_comb[15:8]] ^ p9_xor_2052899_comb[7:0] ^ p9_array_index_2053003_comb ^ p9_array_index_2053004_comb ^ p9_array_index_2053005_comb ^ p8_literal_2043914[p9_res7__1191_comb] ^ p8_literal_2043912[p9_res7__1193_comb] ^ p8_literal_2043910[p9_res7__1195_comb] ^ p9_xor_2052899_comb[79:72];
  assign p9_array_index_2053015_comb = p8_literal_2043920[p9_res7__1187_comb];
  assign p9_array_index_2053016_comb = p8_literal_2043918[p9_res7__1189_comb];
  assign p9_array_index_2053017_comb = p8_literal_2043916[p9_res7__1191_comb];
  assign p9_res7__1199_comb = p8_literal_2043910[p9_xor_2052899_comb[63:56]] ^ p8_literal_2043912[p9_xor_2052899_comb[55:48]] ^ p8_literal_2043914[p9_xor_2052899_comb[47:40]] ^ p8_literal_2043916[p9_xor_2052899_comb[39:32]] ^ p9_array_index_2052938_comb ^ p9_array_index_2052965_comb ^ p9_xor_2052899_comb[15:8] ^ p8_literal_2043923[p9_xor_2052899_comb[7:0]] ^ p9_res7__1185_comb ^ p9_array_index_2053015_comb ^ p9_array_index_2053016_comb ^ p9_array_index_2053017_comb ^ p8_literal_2043914[p9_res7__1193_comb] ^ p8_literal_2043912[p9_res7__1195_comb] ^ p8_literal_2043910[p9_res7__1197_comb] ^ p9_xor_2052899_comb[71:64];
  assign p9_array_index_2053026_comb = p8_literal_2043920[p9_res7__1189_comb];
  assign p9_array_index_2053027_comb = p8_literal_2043918[p9_res7__1191_comb];
  assign p9_res7__1201_comb = p8_literal_2043910[p9_xor_2052899_comb[55:48]] ^ p8_literal_2043912[p9_xor_2052899_comb[47:40]] ^ p8_literal_2043914[p9_xor_2052899_comb[39:32]] ^ p9_array_index_2052924_comb ^ p9_array_index_2052952_comb ^ p9_array_index_2052978_comb ^ p9_xor_2052899_comb[7:0] ^ p8_literal_2043923[p9_res7__1185_comb] ^ p9_res7__1187_comb ^ p9_array_index_2053026_comb ^ p9_array_index_2053027_comb ^ p8_literal_2043916[p9_res7__1193_comb] ^ p8_literal_2043914[p9_res7__1195_comb] ^ p8_literal_2043912[p9_res7__1197_comb] ^ p8_literal_2043910[p9_res7__1199_comb] ^ p9_xor_2052899_comb[63:56];
  assign p9_array_index_2053037_comb = p8_literal_2043920[p9_res7__1191_comb];
  assign p9_array_index_2053038_comb = p8_literal_2043918[p9_res7__1193_comb];
  assign p9_res7__1203_comb = p8_literal_2043910[p9_xor_2052899_comb[47:40]] ^ p8_literal_2043912[p9_xor_2052899_comb[39:32]] ^ p8_literal_2043914[p9_xor_2052899_comb[31:24]] ^ p9_array_index_2052939_comb ^ p9_array_index_2052966_comb ^ p9_array_index_2052991_comb ^ p9_res7__1185_comb ^ p8_literal_2043923[p9_res7__1187_comb] ^ p9_res7__1189_comb ^ p9_array_index_2053037_comb ^ p9_array_index_2053038_comb ^ p8_literal_2043916[p9_res7__1195_comb] ^ p8_literal_2043914[p9_res7__1197_comb] ^ p8_literal_2043912[p9_res7__1199_comb] ^ p8_literal_2043910[p9_res7__1201_comb] ^ p9_xor_2052899_comb[55:48];
  assign p9_array_index_2053047_comb = p8_literal_2043920[p9_res7__1193_comb];
  assign p9_res7__1205_comb = p8_literal_2043910[p9_xor_2052899_comb[39:32]] ^ p8_literal_2043912[p9_xor_2052899_comb[31:24]] ^ p9_array_index_2052925_comb ^ p9_array_index_2052953_comb ^ p9_array_index_2052979_comb ^ p9_array_index_2053003_comb ^ p9_res7__1187_comb ^ p8_literal_2043923[p9_res7__1189_comb] ^ p9_res7__1191_comb ^ p9_array_index_2053047_comb ^ p8_literal_2043918[p9_res7__1195_comb] ^ p8_literal_2043916[p9_res7__1197_comb] ^ p8_literal_2043914[p9_res7__1199_comb] ^ p8_literal_2043912[p9_res7__1201_comb] ^ p8_literal_2043910[p9_res7__1203_comb] ^ p9_xor_2052899_comb[47:40];
  assign p9_array_index_2053057_comb = p8_literal_2043920[p9_res7__1195_comb];
  assign p9_res7__1207_comb = p8_literal_2043910[p9_xor_2052899_comb[31:24]] ^ p8_literal_2043912[p9_xor_2052899_comb[23:16]] ^ p9_array_index_2052940_comb ^ p9_array_index_2052967_comb ^ p9_array_index_2052992_comb ^ p9_array_index_2053015_comb ^ p9_res7__1189_comb ^ p8_literal_2043923[p9_res7__1191_comb] ^ p9_res7__1193_comb ^ p9_array_index_2053057_comb ^ p8_literal_2043918[p9_res7__1197_comb] ^ p8_literal_2043916[p9_res7__1199_comb] ^ p8_literal_2043914[p9_res7__1201_comb] ^ p8_literal_2043912[p9_res7__1203_comb] ^ p8_literal_2043910[p9_res7__1205_comb] ^ p9_xor_2052899_comb[39:32];
  assign p9_res7__1209_comb = p8_literal_2043910[p9_xor_2052899_comb[23:16]] ^ p9_array_index_2052926_comb ^ p9_array_index_2052954_comb ^ p9_array_index_2052980_comb ^ p9_array_index_2053004_comb ^ p9_array_index_2053026_comb ^ p9_res7__1191_comb ^ p8_literal_2043923[p9_res7__1193_comb] ^ p9_res7__1195_comb ^ p8_literal_2043920[p9_res7__1197_comb] ^ p8_literal_2043918[p9_res7__1199_comb] ^ p8_literal_2043916[p9_res7__1201_comb] ^ p8_literal_2043914[p9_res7__1203_comb] ^ p8_literal_2043912[p9_res7__1205_comb] ^ p8_literal_2043910[p9_res7__1207_comb] ^ p9_xor_2052899_comb[31:24];
  assign p9_res7__1211_comb = p8_literal_2043910[p9_xor_2052899_comb[15:8]] ^ p9_array_index_2052941_comb ^ p9_array_index_2052968_comb ^ p9_array_index_2052993_comb ^ p9_array_index_2053016_comb ^ p9_array_index_2053037_comb ^ p9_res7__1193_comb ^ p8_literal_2043923[p9_res7__1195_comb] ^ p9_res7__1197_comb ^ p8_literal_2043920[p9_res7__1199_comb] ^ p8_literal_2043918[p9_res7__1201_comb] ^ p8_literal_2043916[p9_res7__1203_comb] ^ p8_literal_2043914[p9_res7__1205_comb] ^ p8_literal_2043912[p9_res7__1207_comb] ^ p8_literal_2043910[p9_res7__1209_comb] ^ p9_xor_2052899_comb[23:16];
  assign p9_res7__1213_comb = p9_array_index_2052927_comb ^ p9_array_index_2052955_comb ^ p9_array_index_2052981_comb ^ p9_array_index_2053005_comb ^ p9_array_index_2053027_comb ^ p9_array_index_2053047_comb ^ p9_res7__1195_comb ^ p8_literal_2043923[p9_res7__1197_comb] ^ p9_res7__1199_comb ^ p8_literal_2043920[p9_res7__1201_comb] ^ p8_literal_2043918[p9_res7__1203_comb] ^ p8_literal_2043916[p9_res7__1205_comb] ^ p8_literal_2043914[p9_res7__1207_comb] ^ p8_literal_2043912[p9_res7__1209_comb] ^ p8_literal_2043910[p9_res7__1211_comb] ^ p9_xor_2052899_comb[15:8];
  assign p9_res7__1215_comb = p9_array_index_2052942_comb ^ p9_array_index_2052969_comb ^ p9_array_index_2052994_comb ^ p9_array_index_2053017_comb ^ p9_array_index_2053038_comb ^ p9_array_index_2053057_comb ^ p9_res7__1197_comb ^ p8_literal_2043923[p9_res7__1199_comb] ^ p9_res7__1201_comb ^ p8_literal_2043920[p9_res7__1203_comb] ^ p8_literal_2043918[p9_res7__1205_comb] ^ p8_literal_2043916[p9_res7__1207_comb] ^ p8_literal_2043914[p9_res7__1209_comb] ^ p8_literal_2043912[p9_res7__1211_comb] ^ p8_literal_2043910[p9_res7__1213_comb] ^ p9_xor_2052899_comb[7:0];
  assign p9_permut__37_comb = {p8_literal_2051898[p9_res7__1185_comb], p8_literal_2051898[p9_res7__1187_comb], p8_literal_2051898[p9_res7__1189_comb], p8_literal_2051898[p9_res7__1191_comb], p8_literal_2051898[p9_res7__1193_comb], p8_literal_2051898[p9_res7__1195_comb], p8_literal_2051898[p9_res7__1197_comb], p8_literal_2051898[p9_res7__1199_comb], p8_literal_2051898[p9_res7__1201_comb], p8_literal_2051898[p9_res7__1203_comb], p8_literal_2051898[p9_res7__1205_comb], p8_literal_2051898[p9_res7__1207_comb], p8_literal_2051898[p9_res7__1209_comb], p8_literal_2051898[p9_res7__1211_comb], p8_literal_2051898[p9_res7__1213_comb], p8_literal_2051898[p9_res7__1215_comb]};
  assign p9_xor_2053115_comb = p8_k3 ^ p9_permut__37_comb;
  assign p9_array_index_2053138_comb = p8_literal_2043920[p9_xor_2053115_comb[47:40]];
  assign p9_array_index_2053139_comb = p8_literal_2043918[p9_xor_2053115_comb[39:32]];
  assign p9_array_index_2053140_comb = p8_literal_2043916[p9_xor_2053115_comb[31:24]];
  assign p9_array_index_2053141_comb = p8_literal_2043914[p9_xor_2053115_comb[23:16]];
  assign p9_array_index_2053142_comb = p8_literal_2043912[p9_xor_2053115_comb[15:8]];
  assign p9_array_index_2053143_comb = p8_literal_2043910[p9_xor_2053115_comb[7:0]];
  assign p9_res7__1217_comb = p8_literal_2043910[p9_xor_2053115_comb[119:112]] ^ p8_literal_2043912[p9_xor_2053115_comb[111:104]] ^ p8_literal_2043914[p9_xor_2053115_comb[103:96]] ^ p8_literal_2043916[p9_xor_2053115_comb[95:88]] ^ p8_literal_2043918[p9_xor_2053115_comb[87:80]] ^ p8_literal_2043920[p9_xor_2053115_comb[79:72]] ^ p9_xor_2053115_comb[71:64] ^ p8_literal_2043923[p9_xor_2053115_comb[63:56]] ^ p9_xor_2053115_comb[55:48] ^ p9_array_index_2053138_comb ^ p9_array_index_2053139_comb ^ p9_array_index_2053140_comb ^ p9_array_index_2053141_comb ^ p9_array_index_2053142_comb ^ p9_array_index_2053143_comb ^ p9_xor_2053115_comb[127:120];
  assign p9_array_index_2053153_comb = p8_literal_2043920[p9_xor_2053115_comb[39:32]];
  assign p9_array_index_2053154_comb = p8_literal_2043918[p9_xor_2053115_comb[31:24]];
  assign p9_array_index_2053155_comb = p8_literal_2043916[p9_xor_2053115_comb[23:16]];
  assign p9_array_index_2053156_comb = p8_literal_2043914[p9_xor_2053115_comb[15:8]];
  assign p9_array_index_2053157_comb = p8_literal_2043912[p9_xor_2053115_comb[7:0]];
  assign p9_array_index_2053158_comb = p8_literal_2043910[p9_res7__1217_comb];
  assign p9_res7__1219_comb = p8_literal_2043910[p9_xor_2053115_comb[111:104]] ^ p8_literal_2043912[p9_xor_2053115_comb[103:96]] ^ p8_literal_2043914[p9_xor_2053115_comb[95:88]] ^ p8_literal_2043916[p9_xor_2053115_comb[87:80]] ^ p8_literal_2043918[p9_xor_2053115_comb[79:72]] ^ p8_literal_2043920[p9_xor_2053115_comb[71:64]] ^ p9_xor_2053115_comb[63:56] ^ p8_literal_2043923[p9_xor_2053115_comb[55:48]] ^ p9_xor_2053115_comb[47:40] ^ p9_array_index_2053153_comb ^ p9_array_index_2053154_comb ^ p9_array_index_2053155_comb ^ p9_array_index_2053156_comb ^ p9_array_index_2053157_comb ^ p9_array_index_2053158_comb ^ p9_xor_2053115_comb[119:112];
  assign p9_array_index_2053167_comb = p8_literal_2043920[p9_xor_2053115_comb[31:24]];
  assign p9_array_index_2053168_comb = p8_literal_2043918[p9_xor_2053115_comb[23:16]];
  assign p9_array_index_2053169_comb = p8_literal_2043916[p9_xor_2053115_comb[15:8]];
  assign p9_array_index_2053170_comb = p8_literal_2043914[p9_xor_2053115_comb[7:0]];
  assign p9_array_index_2053171_comb = p8_literal_2043912[p9_res7__1217_comb];
  assign p9_res7__1221_comb = p8_literal_2043910[p9_xor_2053115_comb[103:96]] ^ p8_literal_2043912[p9_xor_2053115_comb[95:88]] ^ p8_literal_2043914[p9_xor_2053115_comb[87:80]] ^ p8_literal_2043916[p9_xor_2053115_comb[79:72]] ^ p8_literal_2043918[p9_xor_2053115_comb[71:64]] ^ p8_literal_2043920[p9_xor_2053115_comb[63:56]] ^ p9_xor_2053115_comb[55:48] ^ p8_literal_2043923[p9_xor_2053115_comb[47:40]] ^ p9_xor_2053115_comb[39:32] ^ p9_array_index_2053167_comb ^ p9_array_index_2053168_comb ^ p9_array_index_2053169_comb ^ p9_array_index_2053170_comb ^ p9_array_index_2053171_comb ^ p8_literal_2043910[p9_res7__1219_comb] ^ p9_xor_2053115_comb[111:104];
  assign p9_array_index_2053181_comb = p8_literal_2043920[p9_xor_2053115_comb[23:16]];
  assign p9_array_index_2053182_comb = p8_literal_2043918[p9_xor_2053115_comb[15:8]];
  assign p9_array_index_2053183_comb = p8_literal_2043916[p9_xor_2053115_comb[7:0]];
  assign p9_array_index_2053184_comb = p8_literal_2043914[p9_res7__1217_comb];
  assign p9_array_index_2053185_comb = p8_literal_2043912[p9_res7__1219_comb];
  assign p9_res7__1223_comb = p8_literal_2043910[p9_xor_2053115_comb[95:88]] ^ p8_literal_2043912[p9_xor_2053115_comb[87:80]] ^ p8_literal_2043914[p9_xor_2053115_comb[79:72]] ^ p8_literal_2043916[p9_xor_2053115_comb[71:64]] ^ p8_literal_2043918[p9_xor_2053115_comb[63:56]] ^ p8_literal_2043920[p9_xor_2053115_comb[55:48]] ^ p9_xor_2053115_comb[47:40] ^ p8_literal_2043923[p9_xor_2053115_comb[39:32]] ^ p9_xor_2053115_comb[31:24] ^ p9_array_index_2053181_comb ^ p9_array_index_2053182_comb ^ p9_array_index_2053183_comb ^ p9_array_index_2053184_comb ^ p9_array_index_2053185_comb ^ p8_literal_2043910[p9_res7__1221_comb] ^ p9_xor_2053115_comb[103:96];
  assign p9_array_index_2053194_comb = p8_literal_2043920[p9_xor_2053115_comb[15:8]];
  assign p9_array_index_2053195_comb = p8_literal_2043918[p9_xor_2053115_comb[7:0]];
  assign p9_array_index_2053196_comb = p8_literal_2043916[p9_res7__1217_comb];
  assign p9_array_index_2053197_comb = p8_literal_2043914[p9_res7__1219_comb];
  assign p9_res7__1225_comb = p8_literal_2043910[p9_xor_2053115_comb[87:80]] ^ p8_literal_2043912[p9_xor_2053115_comb[79:72]] ^ p8_literal_2043914[p9_xor_2053115_comb[71:64]] ^ p8_literal_2043916[p9_xor_2053115_comb[63:56]] ^ p8_literal_2043918[p9_xor_2053115_comb[55:48]] ^ p9_array_index_2053138_comb ^ p9_xor_2053115_comb[39:32] ^ p8_literal_2043923[p9_xor_2053115_comb[31:24]] ^ p9_xor_2053115_comb[23:16] ^ p9_array_index_2053194_comb ^ p9_array_index_2053195_comb ^ p9_array_index_2053196_comb ^ p9_array_index_2053197_comb ^ p8_literal_2043912[p9_res7__1221_comb] ^ p8_literal_2043910[p9_res7__1223_comb] ^ p9_xor_2053115_comb[95:88];
  assign p9_array_index_2053207_comb = p8_literal_2043920[p9_xor_2053115_comb[7:0]];
  assign p9_array_index_2053208_comb = p8_literal_2043918[p9_res7__1217_comb];
  assign p9_array_index_2053209_comb = p8_literal_2043916[p9_res7__1219_comb];
  assign p9_array_index_2053210_comb = p8_literal_2043914[p9_res7__1221_comb];
  assign p9_res7__1227_comb = p8_literal_2043910[p9_xor_2053115_comb[79:72]] ^ p8_literal_2043912[p9_xor_2053115_comb[71:64]] ^ p8_literal_2043914[p9_xor_2053115_comb[63:56]] ^ p8_literal_2043916[p9_xor_2053115_comb[55:48]] ^ p8_literal_2043918[p9_xor_2053115_comb[47:40]] ^ p9_array_index_2053153_comb ^ p9_xor_2053115_comb[31:24] ^ p8_literal_2043923[p9_xor_2053115_comb[23:16]] ^ p9_xor_2053115_comb[15:8] ^ p9_array_index_2053207_comb ^ p9_array_index_2053208_comb ^ p9_array_index_2053209_comb ^ p9_array_index_2053210_comb ^ p8_literal_2043912[p9_res7__1223_comb] ^ p8_literal_2043910[p9_res7__1225_comb] ^ p9_xor_2053115_comb[87:80];
  assign p9_array_index_2053219_comb = p8_literal_2043920[p9_res7__1217_comb];
  assign p9_array_index_2053220_comb = p8_literal_2043918[p9_res7__1219_comb];
  assign p9_array_index_2053221_comb = p8_literal_2043916[p9_res7__1221_comb];
  assign p9_res7__1229_comb = p8_literal_2043910[p9_xor_2053115_comb[71:64]] ^ p8_literal_2043912[p9_xor_2053115_comb[63:56]] ^ p8_literal_2043914[p9_xor_2053115_comb[55:48]] ^ p8_literal_2043916[p9_xor_2053115_comb[47:40]] ^ p9_array_index_2053139_comb ^ p9_array_index_2053167_comb ^ p9_xor_2053115_comb[23:16] ^ p8_literal_2043923[p9_xor_2053115_comb[15:8]] ^ p9_xor_2053115_comb[7:0] ^ p9_array_index_2053219_comb ^ p9_array_index_2053220_comb ^ p9_array_index_2053221_comb ^ p8_literal_2043914[p9_res7__1223_comb] ^ p8_literal_2043912[p9_res7__1225_comb] ^ p8_literal_2043910[p9_res7__1227_comb] ^ p9_xor_2053115_comb[79:72];
  assign p9_array_index_2053231_comb = p8_literal_2043920[p9_res7__1219_comb];
  assign p9_array_index_2053232_comb = p8_literal_2043918[p9_res7__1221_comb];
  assign p9_array_index_2053233_comb = p8_literal_2043916[p9_res7__1223_comb];
  assign p9_res7__1231_comb = p8_literal_2043910[p9_xor_2053115_comb[63:56]] ^ p8_literal_2043912[p9_xor_2053115_comb[55:48]] ^ p8_literal_2043914[p9_xor_2053115_comb[47:40]] ^ p8_literal_2043916[p9_xor_2053115_comb[39:32]] ^ p9_array_index_2053154_comb ^ p9_array_index_2053181_comb ^ p9_xor_2053115_comb[15:8] ^ p8_literal_2043923[p9_xor_2053115_comb[7:0]] ^ p9_res7__1217_comb ^ p9_array_index_2053231_comb ^ p9_array_index_2053232_comb ^ p9_array_index_2053233_comb ^ p8_literal_2043914[p9_res7__1225_comb] ^ p8_literal_2043912[p9_res7__1227_comb] ^ p8_literal_2043910[p9_res7__1229_comb] ^ p9_xor_2053115_comb[71:64];
  assign p9_array_index_2053242_comb = p8_literal_2043920[p9_res7__1221_comb];
  assign p9_array_index_2053243_comb = p8_literal_2043918[p9_res7__1223_comb];
  assign p9_res7__1233_comb = p8_literal_2043910[p9_xor_2053115_comb[55:48]] ^ p8_literal_2043912[p9_xor_2053115_comb[47:40]] ^ p8_literal_2043914[p9_xor_2053115_comb[39:32]] ^ p9_array_index_2053140_comb ^ p9_array_index_2053168_comb ^ p9_array_index_2053194_comb ^ p9_xor_2053115_comb[7:0] ^ p8_literal_2043923[p9_res7__1217_comb] ^ p9_res7__1219_comb ^ p9_array_index_2053242_comb ^ p9_array_index_2053243_comb ^ p8_literal_2043916[p9_res7__1225_comb] ^ p8_literal_2043914[p9_res7__1227_comb] ^ p8_literal_2043912[p9_res7__1229_comb] ^ p8_literal_2043910[p9_res7__1231_comb] ^ p9_xor_2053115_comb[63:56];
  assign p9_array_index_2053253_comb = p8_literal_2043920[p9_res7__1223_comb];
  assign p9_array_index_2053254_comb = p8_literal_2043918[p9_res7__1225_comb];
  assign p9_res7__1235_comb = p8_literal_2043910[p9_xor_2053115_comb[47:40]] ^ p8_literal_2043912[p9_xor_2053115_comb[39:32]] ^ p8_literal_2043914[p9_xor_2053115_comb[31:24]] ^ p9_array_index_2053155_comb ^ p9_array_index_2053182_comb ^ p9_array_index_2053207_comb ^ p9_res7__1217_comb ^ p8_literal_2043923[p9_res7__1219_comb] ^ p9_res7__1221_comb ^ p9_array_index_2053253_comb ^ p9_array_index_2053254_comb ^ p8_literal_2043916[p9_res7__1227_comb] ^ p8_literal_2043914[p9_res7__1229_comb] ^ p8_literal_2043912[p9_res7__1231_comb] ^ p8_literal_2043910[p9_res7__1233_comb] ^ p9_xor_2053115_comb[55:48];
  assign p9_array_index_2053263_comb = p8_literal_2043920[p9_res7__1225_comb];
  assign p9_res7__1237_comb = p8_literal_2043910[p9_xor_2053115_comb[39:32]] ^ p8_literal_2043912[p9_xor_2053115_comb[31:24]] ^ p9_array_index_2053141_comb ^ p9_array_index_2053169_comb ^ p9_array_index_2053195_comb ^ p9_array_index_2053219_comb ^ p9_res7__1219_comb ^ p8_literal_2043923[p9_res7__1221_comb] ^ p9_res7__1223_comb ^ p9_array_index_2053263_comb ^ p8_literal_2043918[p9_res7__1227_comb] ^ p8_literal_2043916[p9_res7__1229_comb] ^ p8_literal_2043914[p9_res7__1231_comb] ^ p8_literal_2043912[p9_res7__1233_comb] ^ p8_literal_2043910[p9_res7__1235_comb] ^ p9_xor_2053115_comb[47:40];
  assign p9_array_index_2053273_comb = p8_literal_2043920[p9_res7__1227_comb];
  assign p9_res7__1239_comb = p8_literal_2043910[p9_xor_2053115_comb[31:24]] ^ p8_literal_2043912[p9_xor_2053115_comb[23:16]] ^ p9_array_index_2053156_comb ^ p9_array_index_2053183_comb ^ p9_array_index_2053208_comb ^ p9_array_index_2053231_comb ^ p9_res7__1221_comb ^ p8_literal_2043923[p9_res7__1223_comb] ^ p9_res7__1225_comb ^ p9_array_index_2053273_comb ^ p8_literal_2043918[p9_res7__1229_comb] ^ p8_literal_2043916[p9_res7__1231_comb] ^ p8_literal_2043914[p9_res7__1233_comb] ^ p8_literal_2043912[p9_res7__1235_comb] ^ p8_literal_2043910[p9_res7__1237_comb] ^ p9_xor_2053115_comb[39:32];
  assign p9_res7__1241_comb = p8_literal_2043910[p9_xor_2053115_comb[23:16]] ^ p9_array_index_2053142_comb ^ p9_array_index_2053170_comb ^ p9_array_index_2053196_comb ^ p9_array_index_2053220_comb ^ p9_array_index_2053242_comb ^ p9_res7__1223_comb ^ p8_literal_2043923[p9_res7__1225_comb] ^ p9_res7__1227_comb ^ p8_literal_2043920[p9_res7__1229_comb] ^ p8_literal_2043918[p9_res7__1231_comb] ^ p8_literal_2043916[p9_res7__1233_comb] ^ p8_literal_2043914[p9_res7__1235_comb] ^ p8_literal_2043912[p9_res7__1237_comb] ^ p8_literal_2043910[p9_res7__1239_comb] ^ p9_xor_2053115_comb[31:24];
  assign p9_res7__1243_comb = p8_literal_2043910[p9_xor_2053115_comb[15:8]] ^ p9_array_index_2053157_comb ^ p9_array_index_2053184_comb ^ p9_array_index_2053209_comb ^ p9_array_index_2053232_comb ^ p9_array_index_2053253_comb ^ p9_res7__1225_comb ^ p8_literal_2043923[p9_res7__1227_comb] ^ p9_res7__1229_comb ^ p8_literal_2043920[p9_res7__1231_comb] ^ p8_literal_2043918[p9_res7__1233_comb] ^ p8_literal_2043916[p9_res7__1235_comb] ^ p8_literal_2043914[p9_res7__1237_comb] ^ p8_literal_2043912[p9_res7__1239_comb] ^ p8_literal_2043910[p9_res7__1241_comb] ^ p9_xor_2053115_comb[23:16];
  assign p9_res7__1245_comb = p9_array_index_2053143_comb ^ p9_array_index_2053171_comb ^ p9_array_index_2053197_comb ^ p9_array_index_2053221_comb ^ p9_array_index_2053243_comb ^ p9_array_index_2053263_comb ^ p9_res7__1227_comb ^ p8_literal_2043923[p9_res7__1229_comb] ^ p9_res7__1231_comb ^ p8_literal_2043920[p9_res7__1233_comb] ^ p8_literal_2043918[p9_res7__1235_comb] ^ p8_literal_2043916[p9_res7__1237_comb] ^ p8_literal_2043914[p9_res7__1239_comb] ^ p8_literal_2043912[p9_res7__1241_comb] ^ p8_literal_2043910[p9_res7__1243_comb] ^ p9_xor_2053115_comb[15:8];
  assign p9_res7__1247_comb = p9_array_index_2053158_comb ^ p9_array_index_2053185_comb ^ p9_array_index_2053210_comb ^ p9_array_index_2053233_comb ^ p9_array_index_2053254_comb ^ p9_array_index_2053273_comb ^ p9_res7__1229_comb ^ p8_literal_2043923[p9_res7__1231_comb] ^ p9_res7__1233_comb ^ p8_literal_2043920[p9_res7__1235_comb] ^ p8_literal_2043918[p9_res7__1237_comb] ^ p8_literal_2043916[p9_res7__1239_comb] ^ p8_literal_2043914[p9_res7__1241_comb] ^ p8_literal_2043912[p9_res7__1243_comb] ^ p8_literal_2043910[p9_res7__1245_comb] ^ p9_xor_2053115_comb[7:0];
  assign p9_permut__38_comb = {p8_literal_2051898[p9_res7__1217_comb], p8_literal_2051898[p9_res7__1219_comb], p8_literal_2051898[p9_res7__1221_comb], p8_literal_2051898[p9_res7__1223_comb], p8_literal_2051898[p9_res7__1225_comb], p8_literal_2051898[p9_res7__1227_comb], p8_literal_2051898[p9_res7__1229_comb], p8_literal_2051898[p9_res7__1231_comb], p8_literal_2051898[p9_res7__1233_comb], p8_literal_2051898[p9_res7__1235_comb], p8_literal_2051898[p9_res7__1237_comb], p8_literal_2051898[p9_res7__1239_comb], p8_literal_2051898[p9_res7__1241_comb], p8_literal_2051898[p9_res7__1243_comb], p8_literal_2051898[p9_res7__1245_comb], p8_literal_2051898[p9_res7__1247_comb]};
  assign p9_xor_2053331_comb = p8_k2 ^ p9_permut__38_comb;
  assign p9_array_index_2053354_comb = p8_literal_2043920[p9_xor_2053331_comb[47:40]];
  assign p9_array_index_2053355_comb = p8_literal_2043918[p9_xor_2053331_comb[39:32]];
  assign p9_array_index_2053356_comb = p8_literal_2043916[p9_xor_2053331_comb[31:24]];
  assign p9_array_index_2053357_comb = p8_literal_2043914[p9_xor_2053331_comb[23:16]];
  assign p9_array_index_2053358_comb = p8_literal_2043912[p9_xor_2053331_comb[15:8]];
  assign p9_array_index_2053359_comb = p8_literal_2043910[p9_xor_2053331_comb[7:0]];
  assign p9_res7__1249_comb = p8_literal_2043910[p9_xor_2053331_comb[119:112]] ^ p8_literal_2043912[p9_xor_2053331_comb[111:104]] ^ p8_literal_2043914[p9_xor_2053331_comb[103:96]] ^ p8_literal_2043916[p9_xor_2053331_comb[95:88]] ^ p8_literal_2043918[p9_xor_2053331_comb[87:80]] ^ p8_literal_2043920[p9_xor_2053331_comb[79:72]] ^ p9_xor_2053331_comb[71:64] ^ p8_literal_2043923[p9_xor_2053331_comb[63:56]] ^ p9_xor_2053331_comb[55:48] ^ p9_array_index_2053354_comb ^ p9_array_index_2053355_comb ^ p9_array_index_2053356_comb ^ p9_array_index_2053357_comb ^ p9_array_index_2053358_comb ^ p9_array_index_2053359_comb ^ p9_xor_2053331_comb[127:120];
  assign p9_array_index_2053369_comb = p8_literal_2043920[p9_xor_2053331_comb[39:32]];
  assign p9_array_index_2053370_comb = p8_literal_2043918[p9_xor_2053331_comb[31:24]];
  assign p9_array_index_2053371_comb = p8_literal_2043916[p9_xor_2053331_comb[23:16]];
  assign p9_array_index_2053372_comb = p8_literal_2043914[p9_xor_2053331_comb[15:8]];
  assign p9_array_index_2053373_comb = p8_literal_2043912[p9_xor_2053331_comb[7:0]];
  assign p9_array_index_2053374_comb = p8_literal_2043910[p9_res7__1249_comb];
  assign p9_res7__1251_comb = p8_literal_2043910[p9_xor_2053331_comb[111:104]] ^ p8_literal_2043912[p9_xor_2053331_comb[103:96]] ^ p8_literal_2043914[p9_xor_2053331_comb[95:88]] ^ p8_literal_2043916[p9_xor_2053331_comb[87:80]] ^ p8_literal_2043918[p9_xor_2053331_comb[79:72]] ^ p8_literal_2043920[p9_xor_2053331_comb[71:64]] ^ p9_xor_2053331_comb[63:56] ^ p8_literal_2043923[p9_xor_2053331_comb[55:48]] ^ p9_xor_2053331_comb[47:40] ^ p9_array_index_2053369_comb ^ p9_array_index_2053370_comb ^ p9_array_index_2053371_comb ^ p9_array_index_2053372_comb ^ p9_array_index_2053373_comb ^ p9_array_index_2053374_comb ^ p9_xor_2053331_comb[119:112];
  assign p9_array_index_2053383_comb = p8_literal_2043920[p9_xor_2053331_comb[31:24]];
  assign p9_array_index_2053384_comb = p8_literal_2043918[p9_xor_2053331_comb[23:16]];
  assign p9_array_index_2053385_comb = p8_literal_2043916[p9_xor_2053331_comb[15:8]];
  assign p9_array_index_2053386_comb = p8_literal_2043914[p9_xor_2053331_comb[7:0]];
  assign p9_array_index_2053387_comb = p8_literal_2043912[p9_res7__1249_comb];
  assign p9_res7__1253_comb = p8_literal_2043910[p9_xor_2053331_comb[103:96]] ^ p8_literal_2043912[p9_xor_2053331_comb[95:88]] ^ p8_literal_2043914[p9_xor_2053331_comb[87:80]] ^ p8_literal_2043916[p9_xor_2053331_comb[79:72]] ^ p8_literal_2043918[p9_xor_2053331_comb[71:64]] ^ p8_literal_2043920[p9_xor_2053331_comb[63:56]] ^ p9_xor_2053331_comb[55:48] ^ p8_literal_2043923[p9_xor_2053331_comb[47:40]] ^ p9_xor_2053331_comb[39:32] ^ p9_array_index_2053383_comb ^ p9_array_index_2053384_comb ^ p9_array_index_2053385_comb ^ p9_array_index_2053386_comb ^ p9_array_index_2053387_comb ^ p8_literal_2043910[p9_res7__1251_comb] ^ p9_xor_2053331_comb[111:104];
  assign p9_array_index_2053397_comb = p8_literal_2043920[p9_xor_2053331_comb[23:16]];
  assign p9_array_index_2053398_comb = p8_literal_2043918[p9_xor_2053331_comb[15:8]];
  assign p9_array_index_2053399_comb = p8_literal_2043916[p9_xor_2053331_comb[7:0]];
  assign p9_array_index_2053400_comb = p8_literal_2043914[p9_res7__1249_comb];
  assign p9_array_index_2053401_comb = p8_literal_2043912[p9_res7__1251_comb];
  assign p9_res7__1255_comb = p8_literal_2043910[p9_xor_2053331_comb[95:88]] ^ p8_literal_2043912[p9_xor_2053331_comb[87:80]] ^ p8_literal_2043914[p9_xor_2053331_comb[79:72]] ^ p8_literal_2043916[p9_xor_2053331_comb[71:64]] ^ p8_literal_2043918[p9_xor_2053331_comb[63:56]] ^ p8_literal_2043920[p9_xor_2053331_comb[55:48]] ^ p9_xor_2053331_comb[47:40] ^ p8_literal_2043923[p9_xor_2053331_comb[39:32]] ^ p9_xor_2053331_comb[31:24] ^ p9_array_index_2053397_comb ^ p9_array_index_2053398_comb ^ p9_array_index_2053399_comb ^ p9_array_index_2053400_comb ^ p9_array_index_2053401_comb ^ p8_literal_2043910[p9_res7__1253_comb] ^ p9_xor_2053331_comb[103:96];
  assign p9_array_index_2053410_comb = p8_literal_2043920[p9_xor_2053331_comb[15:8]];
  assign p9_array_index_2053411_comb = p8_literal_2043918[p9_xor_2053331_comb[7:0]];
  assign p9_array_index_2053412_comb = p8_literal_2043916[p9_res7__1249_comb];
  assign p9_array_index_2053413_comb = p8_literal_2043914[p9_res7__1251_comb];
  assign p9_res7__1257_comb = p8_literal_2043910[p9_xor_2053331_comb[87:80]] ^ p8_literal_2043912[p9_xor_2053331_comb[79:72]] ^ p8_literal_2043914[p9_xor_2053331_comb[71:64]] ^ p8_literal_2043916[p9_xor_2053331_comb[63:56]] ^ p8_literal_2043918[p9_xor_2053331_comb[55:48]] ^ p9_array_index_2053354_comb ^ p9_xor_2053331_comb[39:32] ^ p8_literal_2043923[p9_xor_2053331_comb[31:24]] ^ p9_xor_2053331_comb[23:16] ^ p9_array_index_2053410_comb ^ p9_array_index_2053411_comb ^ p9_array_index_2053412_comb ^ p9_array_index_2053413_comb ^ p8_literal_2043912[p9_res7__1253_comb] ^ p8_literal_2043910[p9_res7__1255_comb] ^ p9_xor_2053331_comb[95:88];
  assign p9_array_index_2053423_comb = p8_literal_2043920[p9_xor_2053331_comb[7:0]];
  assign p9_array_index_2053424_comb = p8_literal_2043918[p9_res7__1249_comb];
  assign p9_array_index_2053425_comb = p8_literal_2043916[p9_res7__1251_comb];
  assign p9_array_index_2053426_comb = p8_literal_2043914[p9_res7__1253_comb];
  assign p9_res7__1259_comb = p8_literal_2043910[p9_xor_2053331_comb[79:72]] ^ p8_literal_2043912[p9_xor_2053331_comb[71:64]] ^ p8_literal_2043914[p9_xor_2053331_comb[63:56]] ^ p8_literal_2043916[p9_xor_2053331_comb[55:48]] ^ p8_literal_2043918[p9_xor_2053331_comb[47:40]] ^ p9_array_index_2053369_comb ^ p9_xor_2053331_comb[31:24] ^ p8_literal_2043923[p9_xor_2053331_comb[23:16]] ^ p9_xor_2053331_comb[15:8] ^ p9_array_index_2053423_comb ^ p9_array_index_2053424_comb ^ p9_array_index_2053425_comb ^ p9_array_index_2053426_comb ^ p8_literal_2043912[p9_res7__1255_comb] ^ p8_literal_2043910[p9_res7__1257_comb] ^ p9_xor_2053331_comb[87:80];
  assign p9_array_index_2053435_comb = p8_literal_2043920[p9_res7__1249_comb];
  assign p9_array_index_2053436_comb = p8_literal_2043918[p9_res7__1251_comb];
  assign p9_array_index_2053437_comb = p8_literal_2043916[p9_res7__1253_comb];
  assign p9_res7__1261_comb = p8_literal_2043910[p9_xor_2053331_comb[71:64]] ^ p8_literal_2043912[p9_xor_2053331_comb[63:56]] ^ p8_literal_2043914[p9_xor_2053331_comb[55:48]] ^ p8_literal_2043916[p9_xor_2053331_comb[47:40]] ^ p9_array_index_2053355_comb ^ p9_array_index_2053383_comb ^ p9_xor_2053331_comb[23:16] ^ p8_literal_2043923[p9_xor_2053331_comb[15:8]] ^ p9_xor_2053331_comb[7:0] ^ p9_array_index_2053435_comb ^ p9_array_index_2053436_comb ^ p9_array_index_2053437_comb ^ p8_literal_2043914[p9_res7__1255_comb] ^ p8_literal_2043912[p9_res7__1257_comb] ^ p8_literal_2043910[p9_res7__1259_comb] ^ p9_xor_2053331_comb[79:72];
  assign p9_array_index_2053447_comb = p8_literal_2043920[p9_res7__1251_comb];
  assign p9_array_index_2053448_comb = p8_literal_2043918[p9_res7__1253_comb];
  assign p9_array_index_2053449_comb = p8_literal_2043916[p9_res7__1255_comb];
  assign p9_res7__1263_comb = p8_literal_2043910[p9_xor_2053331_comb[63:56]] ^ p8_literal_2043912[p9_xor_2053331_comb[55:48]] ^ p8_literal_2043914[p9_xor_2053331_comb[47:40]] ^ p8_literal_2043916[p9_xor_2053331_comb[39:32]] ^ p9_array_index_2053370_comb ^ p9_array_index_2053397_comb ^ p9_xor_2053331_comb[15:8] ^ p8_literal_2043923[p9_xor_2053331_comb[7:0]] ^ p9_res7__1249_comb ^ p9_array_index_2053447_comb ^ p9_array_index_2053448_comb ^ p9_array_index_2053449_comb ^ p8_literal_2043914[p9_res7__1257_comb] ^ p8_literal_2043912[p9_res7__1259_comb] ^ p8_literal_2043910[p9_res7__1261_comb] ^ p9_xor_2053331_comb[71:64];
  assign p9_array_index_2053458_comb = p8_literal_2043920[p9_res7__1253_comb];
  assign p9_array_index_2053459_comb = p8_literal_2043918[p9_res7__1255_comb];
  assign p9_res7__1265_comb = p8_literal_2043910[p9_xor_2053331_comb[55:48]] ^ p8_literal_2043912[p9_xor_2053331_comb[47:40]] ^ p8_literal_2043914[p9_xor_2053331_comb[39:32]] ^ p9_array_index_2053356_comb ^ p9_array_index_2053384_comb ^ p9_array_index_2053410_comb ^ p9_xor_2053331_comb[7:0] ^ p8_literal_2043923[p9_res7__1249_comb] ^ p9_res7__1251_comb ^ p9_array_index_2053458_comb ^ p9_array_index_2053459_comb ^ p8_literal_2043916[p9_res7__1257_comb] ^ p8_literal_2043914[p9_res7__1259_comb] ^ p8_literal_2043912[p9_res7__1261_comb] ^ p8_literal_2043910[p9_res7__1263_comb] ^ p9_xor_2053331_comb[63:56];
  assign p9_array_index_2053469_comb = p8_literal_2043920[p9_res7__1255_comb];
  assign p9_array_index_2053470_comb = p8_literal_2043918[p9_res7__1257_comb];
  assign p9_res7__1267_comb = p8_literal_2043910[p9_xor_2053331_comb[47:40]] ^ p8_literal_2043912[p9_xor_2053331_comb[39:32]] ^ p8_literal_2043914[p9_xor_2053331_comb[31:24]] ^ p9_array_index_2053371_comb ^ p9_array_index_2053398_comb ^ p9_array_index_2053423_comb ^ p9_res7__1249_comb ^ p8_literal_2043923[p9_res7__1251_comb] ^ p9_res7__1253_comb ^ p9_array_index_2053469_comb ^ p9_array_index_2053470_comb ^ p8_literal_2043916[p9_res7__1259_comb] ^ p8_literal_2043914[p9_res7__1261_comb] ^ p8_literal_2043912[p9_res7__1263_comb] ^ p8_literal_2043910[p9_res7__1265_comb] ^ p9_xor_2053331_comb[55:48];
  assign p9_array_index_2053479_comb = p8_literal_2043920[p9_res7__1257_comb];
  assign p9_res7__1269_comb = p8_literal_2043910[p9_xor_2053331_comb[39:32]] ^ p8_literal_2043912[p9_xor_2053331_comb[31:24]] ^ p9_array_index_2053357_comb ^ p9_array_index_2053385_comb ^ p9_array_index_2053411_comb ^ p9_array_index_2053435_comb ^ p9_res7__1251_comb ^ p8_literal_2043923[p9_res7__1253_comb] ^ p9_res7__1255_comb ^ p9_array_index_2053479_comb ^ p8_literal_2043918[p9_res7__1259_comb] ^ p8_literal_2043916[p9_res7__1261_comb] ^ p8_literal_2043914[p9_res7__1263_comb] ^ p8_literal_2043912[p9_res7__1265_comb] ^ p8_literal_2043910[p9_res7__1267_comb] ^ p9_xor_2053331_comb[47:40];
  assign p9_array_index_2053489_comb = p8_literal_2043920[p9_res7__1259_comb];
  assign p9_res7__1271_comb = p8_literal_2043910[p9_xor_2053331_comb[31:24]] ^ p8_literal_2043912[p9_xor_2053331_comb[23:16]] ^ p9_array_index_2053372_comb ^ p9_array_index_2053399_comb ^ p9_array_index_2053424_comb ^ p9_array_index_2053447_comb ^ p9_res7__1253_comb ^ p8_literal_2043923[p9_res7__1255_comb] ^ p9_res7__1257_comb ^ p9_array_index_2053489_comb ^ p8_literal_2043918[p9_res7__1261_comb] ^ p8_literal_2043916[p9_res7__1263_comb] ^ p8_literal_2043914[p9_res7__1265_comb] ^ p8_literal_2043912[p9_res7__1267_comb] ^ p8_literal_2043910[p9_res7__1269_comb] ^ p9_xor_2053331_comb[39:32];
  assign p9_res7__1273_comb = p8_literal_2043910[p9_xor_2053331_comb[23:16]] ^ p9_array_index_2053358_comb ^ p9_array_index_2053386_comb ^ p9_array_index_2053412_comb ^ p9_array_index_2053436_comb ^ p9_array_index_2053458_comb ^ p9_res7__1255_comb ^ p8_literal_2043923[p9_res7__1257_comb] ^ p9_res7__1259_comb ^ p8_literal_2043920[p9_res7__1261_comb] ^ p8_literal_2043918[p9_res7__1263_comb] ^ p8_literal_2043916[p9_res7__1265_comb] ^ p8_literal_2043914[p9_res7__1267_comb] ^ p8_literal_2043912[p9_res7__1269_comb] ^ p8_literal_2043910[p9_res7__1271_comb] ^ p9_xor_2053331_comb[31:24];
  assign p9_res7__1275_comb = p8_literal_2043910[p9_xor_2053331_comb[15:8]] ^ p9_array_index_2053373_comb ^ p9_array_index_2053400_comb ^ p9_array_index_2053425_comb ^ p9_array_index_2053448_comb ^ p9_array_index_2053469_comb ^ p9_res7__1257_comb ^ p8_literal_2043923[p9_res7__1259_comb] ^ p9_res7__1261_comb ^ p8_literal_2043920[p9_res7__1263_comb] ^ p8_literal_2043918[p9_res7__1265_comb] ^ p8_literal_2043916[p9_res7__1267_comb] ^ p8_literal_2043914[p9_res7__1269_comb] ^ p8_literal_2043912[p9_res7__1271_comb] ^ p8_literal_2043910[p9_res7__1273_comb] ^ p9_xor_2053331_comb[23:16];
  assign p9_res7__1277_comb = p9_array_index_2053359_comb ^ p9_array_index_2053387_comb ^ p9_array_index_2053413_comb ^ p9_array_index_2053437_comb ^ p9_array_index_2053459_comb ^ p9_array_index_2053479_comb ^ p9_res7__1259_comb ^ p8_literal_2043923[p9_res7__1261_comb] ^ p9_res7__1263_comb ^ p8_literal_2043920[p9_res7__1265_comb] ^ p8_literal_2043918[p9_res7__1267_comb] ^ p8_literal_2043916[p9_res7__1269_comb] ^ p8_literal_2043914[p9_res7__1271_comb] ^ p8_literal_2043912[p9_res7__1273_comb] ^ p8_literal_2043910[p9_res7__1275_comb] ^ p9_xor_2053331_comb[15:8];
  assign p9_res7__1279_comb = p9_array_index_2053374_comb ^ p9_array_index_2053401_comb ^ p9_array_index_2053426_comb ^ p9_array_index_2053449_comb ^ p9_array_index_2053470_comb ^ p9_array_index_2053489_comb ^ p9_res7__1261_comb ^ p8_literal_2043923[p9_res7__1263_comb] ^ p9_res7__1265_comb ^ p8_literal_2043920[p9_res7__1267_comb] ^ p8_literal_2043918[p9_res7__1269_comb] ^ p8_literal_2043916[p9_res7__1271_comb] ^ p8_literal_2043914[p9_res7__1273_comb] ^ p8_literal_2043912[p9_res7__1275_comb] ^ p8_literal_2043910[p9_res7__1277_comb] ^ p9_xor_2053331_comb[7:0];
  assign p9_permut__39_comb = {p8_literal_2051898[p9_res7__1249_comb], p8_literal_2051898[p9_res7__1251_comb], p8_literal_2051898[p9_res7__1253_comb], p8_literal_2051898[p9_res7__1255_comb], p8_literal_2051898[p9_res7__1257_comb], p8_literal_2051898[p9_res7__1259_comb], p8_literal_2051898[p9_res7__1261_comb], p8_literal_2051898[p9_res7__1263_comb], p8_literal_2051898[p9_res7__1265_comb], p8_literal_2051898[p9_res7__1267_comb], p8_literal_2051898[p9_res7__1269_comb], p8_literal_2051898[p9_res7__1271_comb], p8_literal_2051898[p9_res7__1273_comb], p8_literal_2051898[p9_res7__1275_comb], p8_literal_2051898[p9_res7__1277_comb], p8_literal_2051898[p9_res7__1279_comb]};
  assign p9_xor_2053547_comb = p8_bit_slice_2044119 ^ p9_permut__39_comb;
  assign p9_array_index_2053570_comb = p8_literal_2043920[p9_xor_2053547_comb[47:40]];
  assign p9_array_index_2053571_comb = p8_literal_2043918[p9_xor_2053547_comb[39:32]];
  assign p9_array_index_2053572_comb = p8_literal_2043916[p9_xor_2053547_comb[31:24]];
  assign p9_array_index_2053573_comb = p8_literal_2043914[p9_xor_2053547_comb[23:16]];
  assign p9_array_index_2053574_comb = p8_literal_2043912[p9_xor_2053547_comb[15:8]];
  assign p9_array_index_2053575_comb = p8_literal_2043910[p9_xor_2053547_comb[7:0]];
  assign p9_res7__1281_comb = p8_literal_2043910[p9_xor_2053547_comb[119:112]] ^ p8_literal_2043912[p9_xor_2053547_comb[111:104]] ^ p8_literal_2043914[p9_xor_2053547_comb[103:96]] ^ p8_literal_2043916[p9_xor_2053547_comb[95:88]] ^ p8_literal_2043918[p9_xor_2053547_comb[87:80]] ^ p8_literal_2043920[p9_xor_2053547_comb[79:72]] ^ p9_xor_2053547_comb[71:64] ^ p8_literal_2043923[p9_xor_2053547_comb[63:56]] ^ p9_xor_2053547_comb[55:48] ^ p9_array_index_2053570_comb ^ p9_array_index_2053571_comb ^ p9_array_index_2053572_comb ^ p9_array_index_2053573_comb ^ p9_array_index_2053574_comb ^ p9_array_index_2053575_comb ^ p9_xor_2053547_comb[127:120];
  assign p9_array_index_2053585_comb = p8_literal_2043920[p9_xor_2053547_comb[39:32]];
  assign p9_array_index_2053586_comb = p8_literal_2043918[p9_xor_2053547_comb[31:24]];
  assign p9_array_index_2053587_comb = p8_literal_2043916[p9_xor_2053547_comb[23:16]];
  assign p9_array_index_2053588_comb = p8_literal_2043914[p9_xor_2053547_comb[15:8]];
  assign p9_array_index_2053589_comb = p8_literal_2043912[p9_xor_2053547_comb[7:0]];
  assign p9_array_index_2053590_comb = p8_literal_2043910[p9_res7__1281_comb];
  assign p9_res7__1283_comb = p8_literal_2043910[p9_xor_2053547_comb[111:104]] ^ p8_literal_2043912[p9_xor_2053547_comb[103:96]] ^ p8_literal_2043914[p9_xor_2053547_comb[95:88]] ^ p8_literal_2043916[p9_xor_2053547_comb[87:80]] ^ p8_literal_2043918[p9_xor_2053547_comb[79:72]] ^ p8_literal_2043920[p9_xor_2053547_comb[71:64]] ^ p9_xor_2053547_comb[63:56] ^ p8_literal_2043923[p9_xor_2053547_comb[55:48]] ^ p9_xor_2053547_comb[47:40] ^ p9_array_index_2053585_comb ^ p9_array_index_2053586_comb ^ p9_array_index_2053587_comb ^ p9_array_index_2053588_comb ^ p9_array_index_2053589_comb ^ p9_array_index_2053590_comb ^ p9_xor_2053547_comb[119:112];
  assign p9_array_index_2053599_comb = p8_literal_2043920[p9_xor_2053547_comb[31:24]];
  assign p9_array_index_2053600_comb = p8_literal_2043918[p9_xor_2053547_comb[23:16]];
  assign p9_array_index_2053601_comb = p8_literal_2043916[p9_xor_2053547_comb[15:8]];
  assign p9_array_index_2053602_comb = p8_literal_2043914[p9_xor_2053547_comb[7:0]];
  assign p9_array_index_2053603_comb = p8_literal_2043912[p9_res7__1281_comb];
  assign p9_res7__1285_comb = p8_literal_2043910[p9_xor_2053547_comb[103:96]] ^ p8_literal_2043912[p9_xor_2053547_comb[95:88]] ^ p8_literal_2043914[p9_xor_2053547_comb[87:80]] ^ p8_literal_2043916[p9_xor_2053547_comb[79:72]] ^ p8_literal_2043918[p9_xor_2053547_comb[71:64]] ^ p8_literal_2043920[p9_xor_2053547_comb[63:56]] ^ p9_xor_2053547_comb[55:48] ^ p8_literal_2043923[p9_xor_2053547_comb[47:40]] ^ p9_xor_2053547_comb[39:32] ^ p9_array_index_2053599_comb ^ p9_array_index_2053600_comb ^ p9_array_index_2053601_comb ^ p9_array_index_2053602_comb ^ p9_array_index_2053603_comb ^ p8_literal_2043910[p9_res7__1283_comb] ^ p9_xor_2053547_comb[111:104];
  assign p9_array_index_2053613_comb = p8_literal_2043920[p9_xor_2053547_comb[23:16]];
  assign p9_array_index_2053614_comb = p8_literal_2043918[p9_xor_2053547_comb[15:8]];
  assign p9_array_index_2053615_comb = p8_literal_2043916[p9_xor_2053547_comb[7:0]];
  assign p9_array_index_2053616_comb = p8_literal_2043914[p9_res7__1281_comb];
  assign p9_array_index_2053617_comb = p8_literal_2043912[p9_res7__1283_comb];
  assign p9_res7__1287_comb = p8_literal_2043910[p9_xor_2053547_comb[95:88]] ^ p8_literal_2043912[p9_xor_2053547_comb[87:80]] ^ p8_literal_2043914[p9_xor_2053547_comb[79:72]] ^ p8_literal_2043916[p9_xor_2053547_comb[71:64]] ^ p8_literal_2043918[p9_xor_2053547_comb[63:56]] ^ p8_literal_2043920[p9_xor_2053547_comb[55:48]] ^ p9_xor_2053547_comb[47:40] ^ p8_literal_2043923[p9_xor_2053547_comb[39:32]] ^ p9_xor_2053547_comb[31:24] ^ p9_array_index_2053613_comb ^ p9_array_index_2053614_comb ^ p9_array_index_2053615_comb ^ p9_array_index_2053616_comb ^ p9_array_index_2053617_comb ^ p8_literal_2043910[p9_res7__1285_comb] ^ p9_xor_2053547_comb[103:96];
  assign p9_array_index_2053626_comb = p8_literal_2043920[p9_xor_2053547_comb[15:8]];
  assign p9_array_index_2053627_comb = p8_literal_2043918[p9_xor_2053547_comb[7:0]];
  assign p9_array_index_2053628_comb = p8_literal_2043916[p9_res7__1281_comb];
  assign p9_array_index_2053629_comb = p8_literal_2043914[p9_res7__1283_comb];
  assign p9_res7__1289_comb = p8_literal_2043910[p9_xor_2053547_comb[87:80]] ^ p8_literal_2043912[p9_xor_2053547_comb[79:72]] ^ p8_literal_2043914[p9_xor_2053547_comb[71:64]] ^ p8_literal_2043916[p9_xor_2053547_comb[63:56]] ^ p8_literal_2043918[p9_xor_2053547_comb[55:48]] ^ p9_array_index_2053570_comb ^ p9_xor_2053547_comb[39:32] ^ p8_literal_2043923[p9_xor_2053547_comb[31:24]] ^ p9_xor_2053547_comb[23:16] ^ p9_array_index_2053626_comb ^ p9_array_index_2053627_comb ^ p9_array_index_2053628_comb ^ p9_array_index_2053629_comb ^ p8_literal_2043912[p9_res7__1285_comb] ^ p8_literal_2043910[p9_res7__1287_comb] ^ p9_xor_2053547_comb[95:88];
  assign p9_array_index_2053639_comb = p8_literal_2043920[p9_xor_2053547_comb[7:0]];
  assign p9_array_index_2053640_comb = p8_literal_2043918[p9_res7__1281_comb];
  assign p9_array_index_2053641_comb = p8_literal_2043916[p9_res7__1283_comb];
  assign p9_array_index_2053642_comb = p8_literal_2043914[p9_res7__1285_comb];
  assign p9_res7__1291_comb = p8_literal_2043910[p9_xor_2053547_comb[79:72]] ^ p8_literal_2043912[p9_xor_2053547_comb[71:64]] ^ p8_literal_2043914[p9_xor_2053547_comb[63:56]] ^ p8_literal_2043916[p9_xor_2053547_comb[55:48]] ^ p8_literal_2043918[p9_xor_2053547_comb[47:40]] ^ p9_array_index_2053585_comb ^ p9_xor_2053547_comb[31:24] ^ p8_literal_2043923[p9_xor_2053547_comb[23:16]] ^ p9_xor_2053547_comb[15:8] ^ p9_array_index_2053639_comb ^ p9_array_index_2053640_comb ^ p9_array_index_2053641_comb ^ p9_array_index_2053642_comb ^ p8_literal_2043912[p9_res7__1287_comb] ^ p8_literal_2043910[p9_res7__1289_comb] ^ p9_xor_2053547_comb[87:80];
  assign p9_array_index_2053651_comb = p8_literal_2043920[p9_res7__1281_comb];
  assign p9_array_index_2053652_comb = p8_literal_2043918[p9_res7__1283_comb];
  assign p9_array_index_2053653_comb = p8_literal_2043916[p9_res7__1285_comb];
  assign p9_res7__1293_comb = p8_literal_2043910[p9_xor_2053547_comb[71:64]] ^ p8_literal_2043912[p9_xor_2053547_comb[63:56]] ^ p8_literal_2043914[p9_xor_2053547_comb[55:48]] ^ p8_literal_2043916[p9_xor_2053547_comb[47:40]] ^ p9_array_index_2053571_comb ^ p9_array_index_2053599_comb ^ p9_xor_2053547_comb[23:16] ^ p8_literal_2043923[p9_xor_2053547_comb[15:8]] ^ p9_xor_2053547_comb[7:0] ^ p9_array_index_2053651_comb ^ p9_array_index_2053652_comb ^ p9_array_index_2053653_comb ^ p8_literal_2043914[p9_res7__1287_comb] ^ p8_literal_2043912[p9_res7__1289_comb] ^ p8_literal_2043910[p9_res7__1291_comb] ^ p9_xor_2053547_comb[79:72];
  assign p9_array_index_2053663_comb = p8_literal_2043920[p9_res7__1283_comb];
  assign p9_array_index_2053664_comb = p8_literal_2043918[p9_res7__1285_comb];
  assign p9_array_index_2053665_comb = p8_literal_2043916[p9_res7__1287_comb];
  assign p9_res7__1295_comb = p8_literal_2043910[p9_xor_2053547_comb[63:56]] ^ p8_literal_2043912[p9_xor_2053547_comb[55:48]] ^ p8_literal_2043914[p9_xor_2053547_comb[47:40]] ^ p8_literal_2043916[p9_xor_2053547_comb[39:32]] ^ p9_array_index_2053586_comb ^ p9_array_index_2053613_comb ^ p9_xor_2053547_comb[15:8] ^ p8_literal_2043923[p9_xor_2053547_comb[7:0]] ^ p9_res7__1281_comb ^ p9_array_index_2053663_comb ^ p9_array_index_2053664_comb ^ p9_array_index_2053665_comb ^ p8_literal_2043914[p9_res7__1289_comb] ^ p8_literal_2043912[p9_res7__1291_comb] ^ p8_literal_2043910[p9_res7__1293_comb] ^ p9_xor_2053547_comb[71:64];
  assign p9_array_index_2053674_comb = p8_literal_2043920[p9_res7__1285_comb];
  assign p9_array_index_2053675_comb = p8_literal_2043918[p9_res7__1287_comb];
  assign p9_res7__1297_comb = p8_literal_2043910[p9_xor_2053547_comb[55:48]] ^ p8_literal_2043912[p9_xor_2053547_comb[47:40]] ^ p8_literal_2043914[p9_xor_2053547_comb[39:32]] ^ p9_array_index_2053572_comb ^ p9_array_index_2053600_comb ^ p9_array_index_2053626_comb ^ p9_xor_2053547_comb[7:0] ^ p8_literal_2043923[p9_res7__1281_comb] ^ p9_res7__1283_comb ^ p9_array_index_2053674_comb ^ p9_array_index_2053675_comb ^ p8_literal_2043916[p9_res7__1289_comb] ^ p8_literal_2043914[p9_res7__1291_comb] ^ p8_literal_2043912[p9_res7__1293_comb] ^ p8_literal_2043910[p9_res7__1295_comb] ^ p9_xor_2053547_comb[63:56];
  assign p9_array_index_2053685_comb = p8_literal_2043920[p9_res7__1287_comb];
  assign p9_array_index_2053686_comb = p8_literal_2043918[p9_res7__1289_comb];
  assign p9_res7__1299_comb = p8_literal_2043910[p9_xor_2053547_comb[47:40]] ^ p8_literal_2043912[p9_xor_2053547_comb[39:32]] ^ p8_literal_2043914[p9_xor_2053547_comb[31:24]] ^ p9_array_index_2053587_comb ^ p9_array_index_2053614_comb ^ p9_array_index_2053639_comb ^ p9_res7__1281_comb ^ p8_literal_2043923[p9_res7__1283_comb] ^ p9_res7__1285_comb ^ p9_array_index_2053685_comb ^ p9_array_index_2053686_comb ^ p8_literal_2043916[p9_res7__1291_comb] ^ p8_literal_2043914[p9_res7__1293_comb] ^ p8_literal_2043912[p9_res7__1295_comb] ^ p8_literal_2043910[p9_res7__1297_comb] ^ p9_xor_2053547_comb[55:48];
  assign p9_array_index_2053695_comb = p8_literal_2043920[p9_res7__1289_comb];
  assign p9_res7__1301_comb = p8_literal_2043910[p9_xor_2053547_comb[39:32]] ^ p8_literal_2043912[p9_xor_2053547_comb[31:24]] ^ p9_array_index_2053573_comb ^ p9_array_index_2053601_comb ^ p9_array_index_2053627_comb ^ p9_array_index_2053651_comb ^ p9_res7__1283_comb ^ p8_literal_2043923[p9_res7__1285_comb] ^ p9_res7__1287_comb ^ p9_array_index_2053695_comb ^ p8_literal_2043918[p9_res7__1291_comb] ^ p8_literal_2043916[p9_res7__1293_comb] ^ p8_literal_2043914[p9_res7__1295_comb] ^ p8_literal_2043912[p9_res7__1297_comb] ^ p8_literal_2043910[p9_res7__1299_comb] ^ p9_xor_2053547_comb[47:40];
  assign p9_array_index_2053705_comb = p8_literal_2043920[p9_res7__1291_comb];
  assign p9_res7__1303_comb = p8_literal_2043910[p9_xor_2053547_comb[31:24]] ^ p8_literal_2043912[p9_xor_2053547_comb[23:16]] ^ p9_array_index_2053588_comb ^ p9_array_index_2053615_comb ^ p9_array_index_2053640_comb ^ p9_array_index_2053663_comb ^ p9_res7__1285_comb ^ p8_literal_2043923[p9_res7__1287_comb] ^ p9_res7__1289_comb ^ p9_array_index_2053705_comb ^ p8_literal_2043918[p9_res7__1293_comb] ^ p8_literal_2043916[p9_res7__1295_comb] ^ p8_literal_2043914[p9_res7__1297_comb] ^ p8_literal_2043912[p9_res7__1299_comb] ^ p8_literal_2043910[p9_res7__1301_comb] ^ p9_xor_2053547_comb[39:32];
  assign p9_res7__1305_comb = p8_literal_2043910[p9_xor_2053547_comb[23:16]] ^ p9_array_index_2053574_comb ^ p9_array_index_2053602_comb ^ p9_array_index_2053628_comb ^ p9_array_index_2053652_comb ^ p9_array_index_2053674_comb ^ p9_res7__1287_comb ^ p8_literal_2043923[p9_res7__1289_comb] ^ p9_res7__1291_comb ^ p8_literal_2043920[p9_res7__1293_comb] ^ p8_literal_2043918[p9_res7__1295_comb] ^ p8_literal_2043916[p9_res7__1297_comb] ^ p8_literal_2043914[p9_res7__1299_comb] ^ p8_literal_2043912[p9_res7__1301_comb] ^ p8_literal_2043910[p9_res7__1303_comb] ^ p9_xor_2053547_comb[31:24];
  assign p9_res7__1307_comb = p8_literal_2043910[p9_xor_2053547_comb[15:8]] ^ p9_array_index_2053589_comb ^ p9_array_index_2053616_comb ^ p9_array_index_2053641_comb ^ p9_array_index_2053664_comb ^ p9_array_index_2053685_comb ^ p9_res7__1289_comb ^ p8_literal_2043923[p9_res7__1291_comb] ^ p9_res7__1293_comb ^ p8_literal_2043920[p9_res7__1295_comb] ^ p8_literal_2043918[p9_res7__1297_comb] ^ p8_literal_2043916[p9_res7__1299_comb] ^ p8_literal_2043914[p9_res7__1301_comb] ^ p8_literal_2043912[p9_res7__1303_comb] ^ p8_literal_2043910[p9_res7__1305_comb] ^ p9_xor_2053547_comb[23:16];
  assign p9_res7__1309_comb = p9_array_index_2053575_comb ^ p9_array_index_2053603_comb ^ p9_array_index_2053629_comb ^ p9_array_index_2053653_comb ^ p9_array_index_2053675_comb ^ p9_array_index_2053695_comb ^ p9_res7__1291_comb ^ p8_literal_2043923[p9_res7__1293_comb] ^ p9_res7__1295_comb ^ p8_literal_2043920[p9_res7__1297_comb] ^ p8_literal_2043918[p9_res7__1299_comb] ^ p8_literal_2043916[p9_res7__1301_comb] ^ p8_literal_2043914[p9_res7__1303_comb] ^ p8_literal_2043912[p9_res7__1305_comb] ^ p8_literal_2043910[p9_res7__1307_comb] ^ p9_xor_2053547_comb[15:8];
  assign p9_res7__1311_comb = p9_array_index_2053590_comb ^ p9_array_index_2053617_comb ^ p9_array_index_2053642_comb ^ p9_array_index_2053665_comb ^ p9_array_index_2053686_comb ^ p9_array_index_2053705_comb ^ p9_res7__1293_comb ^ p8_literal_2043923[p9_res7__1295_comb] ^ p9_res7__1297_comb ^ p8_literal_2043920[p9_res7__1299_comb] ^ p8_literal_2043918[p9_res7__1301_comb] ^ p8_literal_2043916[p9_res7__1303_comb] ^ p8_literal_2043914[p9_res7__1305_comb] ^ p8_literal_2043912[p9_res7__1307_comb] ^ p8_literal_2043910[p9_res7__1309_comb] ^ p9_xor_2053547_comb[7:0];
  assign p9_permut__40_comb = {p8_literal_2051898[p9_res7__1281_comb], p8_literal_2051898[p9_res7__1283_comb], p8_literal_2051898[p9_res7__1285_comb], p8_literal_2051898[p9_res7__1287_comb], p8_literal_2051898[p9_res7__1289_comb], p8_literal_2051898[p9_res7__1291_comb], p8_literal_2051898[p9_res7__1293_comb], p8_literal_2051898[p9_res7__1295_comb], p8_literal_2051898[p9_res7__1297_comb], p8_literal_2051898[p9_res7__1299_comb], p8_literal_2051898[p9_res7__1301_comb], p8_literal_2051898[p9_res7__1303_comb], p8_literal_2051898[p9_res7__1305_comb], p8_literal_2051898[p9_res7__1307_comb], p8_literal_2051898[p9_res7__1309_comb], p8_literal_2051898[p9_res7__1311_comb]};
  assign p9_newValue_comb = p8_bit_slice_2043893 ^ p9_permut__40_comb;

  // Registers for pipe stage 9:
  reg [127:0] p9_newValue;
  always_ff @ (posedge clk) begin
    p9_newValue <= p9_newValue_comb;
  end
  assign out = p9_newValue;
endmodule
