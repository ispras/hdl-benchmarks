// IWLS benchmark module "t481" printed on Wed May 29 17:28:14 2002
module t481(v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, \v16.0 );
input
  v10,
  v11,
  v12,
  v13,
  v14,
  v15,
  v0,
  v1,
  v2,
  v3,
  v4,
  v5,
  v6,
  v7,
  v8,
  v9;
output
  \v16.0 ;
wire
  \[8612] ,
  \[12396] ,
  \[11535] ,
  \[10348] ,
  \[14053] ,
  \[4566] ,
  \[14056] ,
  \[6956] ,
  \[13200] ,
  \[4900] ,
  \[12737] ,
  \[13597] ,
  \[10344] ,
  \[9477] ,
  \[3375] ,
  \[8281] ,
  \[4905] ,
  \[5765] ,
  \[12005] ,
  \[1322] ,
  \[5037] ,
  \[12740] ,
  \[10352] ,
  \[12012] ,
  \[7427] ,
  \[13937] ,
  \[7090] ,
  \[6231] ,
  \[8620] ,
  \[8289] ,
  \[3715] ,
  \[584] ,
  \[4575] ,
  \[11545] ,
  \[6964] ,
  \[13206] ,
  \[1329] ,
  \[14065] ,
  \[9484] ,
  \[4910] ,
  \[11552] ,
  \[7098] ,
  \[6239] ,
  \[12749] ,
  \[14072] ,
  \[14071] ,
  \[5773] ,
  \[3385] ,
  \[2526] ,
  \[8629] ,
  \[21807] ,
  \[12745] ,
  \[21471] ,
  \[926] ,
  \[21809] ,
  \[12020] ,
  \[13948] ,
  \[2193] ,
  \[21803] ,
  \[12752] ,
  \[13219] ,
  \[21805] ,
  \[8299] ,
  \[3725] ,
  \[21477] ,
  \[4585] ,
  \[13216] ,
  \[21479] ,
  \[21811] ,
  \[12028] ,
  \[2531] ,
  \[597] ,
  \[10702] ,
  \[14075] ,
  \[21473] ,
  \[11561] ,
  \[4922] ,
  \[6249] ,
  \[14082] ,
  \[21475] ,
  \[3394] ,
  \[14081] ,
  \[5783] ,
  \[933] ,
  \[8639] ,
  \[204] ,
  \[21817] ,
  \[5055] ,
  \[205] ,
  \[11568] ,
  \[206] ,
  \[3000] ,
  \[21481] ,
  \[21819] ,
  \[4927] ,
  \[12760] ,
  \[207] ,
  \[13958] ,
  \[13227] ,
  \[21813] ,
  \[1344] ,
  \[3733] ,
  \[9107] ,
  \[4593] ,
  \[21815] ,
  \[6982] ,
  \[21487] ,
  \[10378] ,
  \[3008] ,
  \[21489] ,
  \[21821] ,
  \[14085] ,
  \[12037] ,
  \[6257] ,
  \[10711] ,
  \[21483] ,
  \[940] ,
  \[4931] ,
  \[2543] ,
  \[11571] ,
  \[211] ,
  \[5791] ,
  \[8647] ,
  \[12769] ,
  \[212] ,
  \[11904] ,
  \[21485] ,
  \[213] ,
  \[10376] ,
  \[214] ,
  \[21827] ,
  \[9841] ,
  \[215] ,
  \[216] ,
  \[21491] ,
  \[21829] ,
  \[7455] ,
  \[217] ,
  \[9844] ,
  \[13968] ,
  \[218] ,
  \[4209] ,
  \[21823] ,
  \[11579] ,
  \[12041] ,
  \[3743] ,
  \[21825] ,
  \[13969] ,
  \[11576] ,
  \[21497] ,
  \[13963] ,
  \[5405] ,
  \[14093] ,
  \[10387] ,
  \[3018] ,
  \[6995] ,
  \[14096] ,
  \[21499] ,
  \[13235] ,
  \[21831] ,
  \[2551] ,
  \[6267] ,
  \[21493] ,
  \[11581] ,
  \[8657] ,
  \[13972] ,
  \[12779] ,
  \[10383] ,
  \[11914] ,
  \[21495] ,
  \[223] ,
  \[4944] ,
  \[224] ,
  \[954] ,
  \[12776] ,
  \[225] ,
  \[10728] ,
  \[1361] ,
  \[4217] ,
  \[12050] ,
  \[11587] ,
  \[13248] ,
  \[3751] ,
  \[13978] ,
  \[6607] ,
  \[4949] ,
  \[11921] ,
  \[10724] ,
  \[6272] ,
  \[13979] ,
  \[13244] ,
  \[3026] ,
  \[7803] ,
  \[22307] ,
  \[13245] ,
  \[2561] ,
  \[6276] ,
  \[22309] ,
  \[11591] ,
  \[13982] ,
  \[12789] ,
  \[11924] ,
  \[12784] ,
  \[9130] ,
  \[4954] ,
  \[12056] ,
  \[9861] ,
  \[10738] ,
  \[7474] ,
  \[10007] ,
  \[6615] ,
  \[11930] ,
  \[21849] ,
  \[2569] ,
  \[22311] ,
  \[3761] ,
  \[11202] ,
  \[2902] ,
  \[13988] ,
  \[1374] ,
  \[12792] ,
  \[10733] ,
  \[13989] ,
  \[11593] ,
  \[13254] ,
  \[3036] ,
  \[10735] ,
  \[9869] ,
  \[1710] ,
  \[22317] ,
  \[13256] ,
  \[11208] ,
  \[11938] ,
  \[21851] ,
  \[12068] ,
  \[8674] ,
  \[12400] ,
  \[22319] ,
  \[5427] ,
  \[10741] ,
  \[22313] ,
  \[971] ,
  \[13262] ,
  \[6289] ,
  \[13992] ,
  \[22315] ,
  \[5094] ,
  \[7483] ,
  \[12796] ,
  \[12065] ,
  \[1381] ,
  \[11210] ,
  \[6625] ,
  \[4237] ,
  \[10747] ,
  \[9143] ,
  \[3770] ,
  \[2579] ,
  \[12408] ,
  \[22321] ,
  \[11212] ,
  \[13998] ,
  \[10749] ,
  \[21853] ,
  \[12071] ,
  \[12409] ,
  \[3044] ,
  \[21855] ,
  \[13264] ,
  \[1388] ,
  \[6294] ,
  \[7823] ,
  \[22327] ,
  \[11218] ,
  \[2918] ,
  \[1721] ,
  \[11948] ,
  \[3778] ,
  \[22329] ,
  \[10752] ,
  \[13270] ,
  \[12077] ,
  \[8685] ,
  \[10021] ,
  \[4971] ,
  \[12412] ,
  \[6298] ,
  \[22323] ,
  \[12079] ,
  \[22325] ,
  \[6633] ,
  \[21867] ,
  \[2587] ,
  \[7493] ,
  \[10028] ,
  \[10758] ,
  \[985] ,
  \[256] ,
  \[21869] ,
  \[13605] ,
  \[12418] ,
  \[257] ,
  \[22331] ,
  \[13610] ,
  \[258] ,
  \[21863] ,
  \[259] ,
  \[12419] ,
  \[3054] ,
  \[21865] ,
  \[7833] ,
  \[22337] ,
  \[3787] ,
  \[11958] ,
  \[21871] ,
  \[12088] ,
  \[1732] ,
  \[22339] ,
  \[10762] ,
  \[260] ,
  \[12422] ,
  \[261] ,
  \[22333] ,
  \[5449] ,
  \[7108] ,
  \[11224] ,
  \[262] ,
  \[992] ,
  \[263] ,
  \[22335] ,
  \[1737] ,
  \[9161] ,
  \[21877] ,
  \[2597] ,
  \[12085] ,
  \[2931] ,
  \[22341] ,
  \[268] ,
  \[4259] ,
  \[3062] ,
  \[21873] ,
  \[269] ,
  \[10764] ,
  \[999] ,
  \[13622] ,
  \[12429] ,
  \[21875] ,
  \[7841] ,
  \[604] ,
  \[13283] ,
  \[12098] ,
  \[12430] ,
  \[1742] ,
  \[11967] ,
  \[7116] ,
  \[270] ,
  \[3402] ,
  \[13627] ,
  \[13291] ,
  \[4993] ,
  \[8310] ,
  \[12094] ,
  \[11233] ,
  \[6653] ,
  \[11966] ,
  \[21887] ,
  \[10777] ,
  \[21889] ,
  \[8314] ,
  \[3071] ,
  \[10049] ,
  \[11241] ,
  \[279] ,
  \[611] ,
  \[10774] ,
  \[9176] ,
  \[13632] ,
  \[12439] ,
  \[4603] ,
  \[2215] ,
  \[7851] ,
  \[13294] ,
  \[12433] ,
  \[2946] ,
  \[21891] ,
  \[12440] ,
  \[22359] ,
  \[3411] ,
  \[7126] ,
  \[280] ,
  \[1754] ,
  \[281] ,
  \[282] ,
  \[8320] ,
  \[7859] ,
  \[13634] ,
  \[11976] ,
  \[11250] ,
  \[10057] ,
  \[1759] ,
  \[286] ,
  \[10787] ,
  \[21501] ,
  \[287] ,
  \[22361] ,
  \[3081] ,
  \[9184] ,
  \[288] ,
  \[289] ,
  \[5471] ,
  \[5809] ,
  \[12449] ,
  \[2954] ,
  \[13641] ,
  \[4614] ,
  \[12443] ,
  \[1030] ,
  \[14103] ,
  \[7134] ,
  \[14106] ,
  \[11257] ,
  \[4280] ,
  \[627] ,
  \[3421] ,
  \[1033] ,
  \[13648] ,
  \[1763] ,
  \[290] ,
  \[11259] ,
  \[291] ,
  \[22363] ,
  \[292] ,
  \[7869] ,
  \[293] ,
  \[22365] ,
  \[8331] ,
  \[11986] ,
  \[13646] ,
  \[6675] ,
  \[10797] ,
  \[4288] ,
  \[9194] ,
  \[298] ,
  \[2963] ,
  \[299] ,
  \[3093] ,
  \[14117] ,
  \[13651] ,
  \[12454] ,
  \[634] ,
  \[10795] ,
  \[14114] ,
  \[4625] ,
  \[2237] ,
  \[7143] ,
  \[11600] ,
  \[21519] ,
  \[3430] ,
  \[11602] ,
  \[5488] ,
  \[13657] ,
  \[7877] ,
  \[1776] ,
  \[11993] ,
  \[11266] ,
  \[11608] ,
  \[21521] ,
  \[3438] ,
  \[4298] ,
  \[5827] ,
  \[10079] ,
  \[2973] ,
  \[641] ,
  \[14127] ,
  \[13661] ,
  \[5493] ,
  \[14124] ,
  \[7153] ,
  \[12466] ,
  \[4636] ,
  \[1781] ,
  \[11610] ,
  \[22389] ,
  \[5100] ,
  \[5498] ,
  \[21523] ,
  \[7887] ,
  \[14132] ,
  \[21525] ,
  \[8350] ,
  \[1786] ,
  \[10416] ,
  \[13663] ,
  \[11275] ,
  \[12806] ,
  \[3447] ,
  \[6695] ,
  \[22391] ,
  \[2982] ,
  \[14138] ,
  \[11619] ,
  \[14137] ,
  \[13672] ,
  \[12479] ,
  \[7162] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[4647] ,
  \[2259] ,
  \[22001] ,
  \[7895] ,
  \[19] ,
  \[1063] ,
  \[12817] ,
  \[22393] ,
  \[7501] ,
  \[10426] ,
  \[22395] ,
  \[14141] ,
  \[11285] ,
  \[1798] ,
  \[5845] ,
  \[3457] ,
  \[2990] ,
  \[20] ,
  \[11627] ,
  \[21] ,
  \[13680] ,
  \[11292] ,
  \[22] ,
  \[14148] ,
  \[1404] ,
  \[22003] ,
  \[12822] ,
  \[23] ,
  \[7170] ,
  \[12489] ,
  \[6311] ,
  \[8368] ,
  \[22005] ,
  \[10095] ,
  \[4656] ,
  \[28] ,
  \[21549] ,
  \[29] ,
  \[7176] ,
  \[8707] ,
  \[11294] ,
  \[6319] ,
  \[14152] ,
  \[1076] ,
  \[2605] ,
  \[7511] ,
  \[12824] ,
  \[14151] ,
  \[3465] ,
  \[10435] ,
  \[9569] ,
  \[22017] ,
  \[5855] ,
  \[13686] ,
  \[30] ,
  \[21551] ,
  \[12100] ,
  \[22019] ,
  \[31] ,
  \[10441] ,
  \[32] ,
  \[14158] ,
  \[22013] ,
  \[12832] ,
  \[33] ,
  \[14157] ,
  \[7180] ,
  \[12499] ,
  \[34] ,
  \[672] ,
  \[12494] ,
  \[7519] ,
  \[22015] ,
  \[35] ,
  \[4664] ,
  \[2276] ,
  \[3805] ,
  \[36] ,
  \[11635] ,
  \[37] ,
  \[38] ,
  \[12108] ,
  \[22021] ,
  \[1083] ,
  \[10449] ,
  \[21553] ,
  \[11641] ,
  \[10444] ,
  \[6329] ,
  \[21555] ,
  \[2615] ,
  \[5863] ,
  \[3475] ,
  \[13694] ,
  \[9579] ,
  \[22027] ,
  \[13696] ,
  \[1421] ,
  \[2281] ,
  \[12110] ,
  \[11647] ,
  \[10452] ,
  \[13308] ,
  \[5138] ,
  \[22023] ,
  \[11649] ,
  \[43] ,
  \[8387] ,
  \[44] ,
  \[7529] ,
  \[22025] ,
  \[11643] ,
  \[45] ,
  \[4674] ,
  \[2286] ,
  \[21567] ,
  \[1090] ,
  \[7193] ,
  \[10457] ,
  \[686] ,
  \[14166] ,
  \[21569] ,
  \[3480] ,
  \[12118] ,
  \[12848] ,
  \[6337] ,
  \[10459] ,
  \[21563] ,
  \[2623] ,
  \[10454] ,
  \[21565] ,
  \[3484] ,
  \[13311] ,
  \[5873] ,
  \[12843] ,
  \[9589] ,
  \[12116] ,
  \[22037] ,
  \[21571] ,
  \[21909] ,
  \[22039] ,
  \[11657] ,
  \[13318] ,
  \[1434] ,
  \[7537] ,
  \[14177] ,
  \[4682] ,
  \[8397] ,
  \[3823] ,
  \[12851] ,
  \[54] ,
  \[55] ,
  \[8731] ,
  \[56] ,
  \[21577] ,
  \[11655] ,
  \[57] ,
  \[2298] ,
  \[21911] ,
  \[22041] ,
  \[12127] ,
  \[6347] ,
  \[300] ,
  \[21573] ,
  \[2633] ,
  \[301] ,
  \[10464] ,
  \[5881] ,
  \[12859] ,
  \[302] ,
  \[21575] ,
  \[303] ,
  \[10466] ,
  \[12853] ,
  \[304] ,
  \[305] ,
  \[9202] ,
  \[3497] ,
  \[12125] ,
  \[1441] ,
  \[306] ,
  \[12130] ,
  \[307] ,
  \[61] ,
  \[308] ,
  \[62] ,
  \[10809] ,
  \[21913] ,
  \[7547] ,
  \[63] ,
  \[14187] ,
  \[12861] ,
  \[11664] ,
  \[64] ,
  \[3104] ,
  \[10803] ,
  \[21915] ,
  \[65] ,
  \[4694] ,
  \[8011] ,
  \[11666] ,
  \[66] ,
  \[10805] ,
  \[21587] ,
  \[1448] ,
  \[67] ,
  \[13326] ,
  \[6355] ,
  \[68] ,
  \[21589] ,
  \[2641] ,
  \[5160] ,
  \[12867] ,
  \[11672] ,
  \[8746] ,
  \[5891] ,
  \[12139] ,
  \[10473] ,
  \[313] ,
  \[12133] ,
  \[7552] ,
  \[314] ,
  \[10475] ,
  \[21927] ,
  \[315] ,
  \[4306] ,
  \[9212] ,
  \[10817] ,
  \[5896] ,
  \[21591] ,
  \[21929] ,
  \[22059] ,
  \[3841] ,
  \[10481] ,
  \[14198] ,
  \[21923] ,
  \[7557] ,
  \[12872] ,
  \[73] ,
  \[11674] ,
  \[74] ,
  \[21925] ,
  \[75] ,
  \[10815] ,
  \[10820] ,
  \[6365] ,
  \[13335] ,
  \[21931] ,
  \[2651] ,
  \[8754] ,
  \[22061] ,
  \[12878] ,
  \[13340] ,
  \[10483] ,
  \[12874] ,
  \[9220] ,
  \[8029] ,
  \[21937] ,
  \[12146] ,
  \[4316] ,
  \[10828] ,
  \[11688] ,
  \[6705] ,
  \[21939] ,
  \[2659] ,
  \[13348] ,
  \[21933] ,
  \[9955] ,
  \[1464] ,
  \[22063] ,
  \[11689] ,
  \[5512] ,
  \[84] ,
  \[21935] ,
  \[7569] ,
  \[22065] ,
  \[11683] ,
  \[85] ,
  \[10826] ,
  \[9958] ,
  \[6373] ,
  \[86] ,
  \[3126] ,
  \[22407] ,
  \[87] ,
  \[10830] ,
  \[8763] ,
  \[21941] ,
  \[22409] ,
  \[5517] ,
  \[1803] ,
  \[11692] ,
  \[331] ,
  \[22403] ,
  \[5182] ,
  \[332] ,
  \[10493] ,
  \[12884] ,
  \[333] ,
  \[22405] ,
  \[4324] ,
  \[12153] ,
  \[1807] ,
  \[334] ,
  \[21947] ,
  \[335] ,
  \[6714] ,
  \[1471] ,
  \[7574] ,
  \[11698] ,
  \[336] ,
  \[21949] ,
  \[2669] ,
  \[337] ,
  \[22411] ,
  \[91] ,
  \[3861] ,
  \[338] ,
  \[92] ,
  \[21943] ,
  \[93] ,
  \[12891] ,
  \[94] ,
  \[21945] ,
  \[7579] ,
  \[95] ,
  \[10836] ,
  \[9238] ,
  \[6383] ,
  \[5524] ,
  \[96] ,
  \[13353] ,
  \[1478] ,
  \[10110] ,
  \[7913] ,
  \[22417] ,
  \[97] ,
  \[10840] ,
  \[8773] ,
  \[98] ,
  \[21951] ,
  \[12500] ,
  \[12898] ,
  \[13360] ,
  \[22413] ,
  \[8047] ,
  \[343] ,
  \[6722] ,
  \[22415] ,
  \[4334] ,
  \[12163] ,
  \[12893] ,
  \[344] ,
  \[21957] ,
  \[2677] ,
  \[11305] ,
  \[345] ,
  \[10848] ,
  \[12895] ,
  \[21959] ,
  \[22089] ,
  \[3142] ,
  \[21953] ,
  \[12172] ,
  \[5199] ,
  \[13702] ,
  \[12509] ,
  \[6391] ,
  \[21955] ,
  \[10846] ,
  \[8781] ,
  \[12503] ,
  \[1820] ,
  \[22427] ,
  \[21961] ,
  \[12510] ,
  \[22091] ,
  \[22429] ,
  \[13370] ,
  \[13708] ,
  \[5538] ,
  \[4342] ,
  \[8057] ,
  \[12179] ,
  \[1825] ,
  \[7591] ,
  \[6732] ,
  \[11316] ,
  \[9251] ,
  \[21967] ,
  \[2687] ,
  \[10857] ,
  \[21969] ,
  \[6006] ,
  \[9983] ,
  \[22431] ,
  \[10129] ,
  \[3152] ,
  \[21963] ,
  \[22093] ,
  \[10854] ,
  \[12181] ,
  \[3883] ,
  \[12519] ,
  \[10123] ,
  \[21965] ,
  \[7599] ,
  \[22095] ,
  \[5543] ,
  \[8791] ,
  \[12513] ,
  \[7203] ,
  \[1830] ,
  \[7933] ,
  \[21971] ,
  \[12520] ,
  \[8065] ,
  \[12187] ,
  \[13718] ,
  \[4351] ,
  \[361] ,
  \[6740] ,
  \[1105] ,
  \[12189] ,
  \[362] ,
  \[2695] ,
  \[363] ,
  \[364] ,
  \[21977] ,
  \[9991] ,
  \[11325] ,
  \[365] ,
  \[6015] ,
  \[10137] ,
  \[366] ,
  \[3160] ,
  \[21979] ,
  \[367] ,
  \[13388] ,
  \[8405] ,
  \[11332] ,
  \[368] ,
  \[5550] ,
  \[2303] ,
  \[21973] ,
  \[12529] ,
  \[6749] ,
  \[10863] ,
  \[21975] ,
  \[703] ,
  \[12523] ,
  \[10865] ,
  \[9269] ,
  \[2307] ,
  \[13383] ,
  \[13386] ,
  \[21981] ,
  \[1842] ,
  \[8075] ,
  \[12197] ,
  \[13728] ,
  \[10141] ,
  \[10871] ,
  \[3502] ,
  \[373] ,
  \[1847] ,
  \[374] ,
  \[3506] ,
  \[11335] ,
  \[375] ,
  \[12195] ,
  \[3170] ,
  \[10877] ,
  \[8415] ,
  \[10149] ,
  \[11341] ,
  \[12539] ,
  \[6759] ,
  \[10146] ,
  \[4705] ,
  \[12536] ,
  \[8083] ,
  \[13396] ,
  \[12535] ,
  \[1851] ,
  \[716] ,
  \[3178] ,
  \[1122] ,
  \[7955] ,
  \[13008] ,
  \[5900] ,
  \[7227] ,
  \[13737] ,
  \[12542] ,
  \[6033] ,
  \[10158] ,
  \[2320] ,
  \[8423] ,
  \[13736] ,
  \[21999] ,
  \[4378] ,
  \[3519] ,
  \[14208] ,
  \[11351] ,
  \[10154] ,
  \[10884] ,
  \[13012] ,
  \[5572] ,
  \[2325] ,
  \[723] ,
  \[12543] ,
  \[4716] ,
  \[8093] ,
  \[11358] ,
  \[3188] ,
  \[21609] ,
  \[12550] ,
  \[10892] ,
  \[391] ,
  \[1135] ,
  \[392] ,
  \[6771] ,
  \[393] ,
  \[5913] ,
  \[394] ,
  \[395] ,
  \[2330] ,
  \[8433] ,
  \[13746] ,
  \[1869] ,
  \[396] ,
  \[21611] ,
  \[3528] ,
  \[397] ,
  \[12557] ,
  \[398] ,
  \[10501] ,
  \[730] ,
  \[11361] ,
  \[2335] ,
  \[3196] ,
  \[14213] ,
  \[11368] ,
  \[4727] ,
  \[9633] ,
  \[1142] ,
  \[12560] ,
  \[7975] ,
  \[13028] ,
  \[10509] ,
  \[14220] ,
  \[21613] ,
  \[12561] ,
  \[21615] ,
  \[5923] ,
  \[8441] ,
  \[6053] ,
  \[11366] ,
  \[3536] ,
  \[1149] ,
  \[13756] ,
  \[13025] ,
  \[12900] ,
  \[13030] ,
  \[12567] ,
  \[2343] ,
  \[4002] ,
  \[7250] ,
  \[11703] ,
  \[5594] ,
  \[21627] ,
  \[12566] ,
  \[11705] ,
  \[4007] ,
  \[21629] ,
  \[4738] ,
  \[10181] ,
  \[14230] ,
  \[13037] ,
  \[21623] ,
  \[9645] ,
  \[11711] ,
  \[10514] ,
  \[11374] ,
  \[21625] ,
  \[7259] ,
  \[10516] ,
  \[8451] ,
  \[11376] ,
  \[1887] ,
  \[12903] ,
  \[3546] ,
  \[13763] ,
  \[6794] ,
  \[10520] ,
  \[11380] ,
  \[12905] ,
  \[21631] ,
  \[10522] ,
  \[6401] ,
  \[12911] ,
  \[4013] ,
  \[8458] ,
  \[13771] ,
  \[10186] ,
  \[11713] ,
  \[21637] ,
  \[2357] ,
  \[7993] ,
  \[10528] ,
  \[12575] ,
  \[14236] ,
  \[9653] ,
  \[12917] ,
  \[21633] ,
  \[4749] ,
  \[6070] ,
  \[12582] ,
  \[11389] ,
  \[11721] ,
  \[6409] ,
  \[21635] ,
  \[3554] ,
  \[7269] ,
  \[11383] ,
  \[14241] ,
  \[12913] ,
  \[6074] ,
  \[22107] ,
  \[10530] ,
  \[13046] ,
  \[5216] ,
  \[13775] ,
  \[22109] ,
  \[10199] ,
  \[11391] ,
  \[22103] ,
  \[13782] ,
  \[10193] ,
  \[762] ,
  \[8800] ,
  \[7609] ,
  \[22105] ,
  \[12583] ,
  \[10195] ,
  \[4025] ,
  \[21647] ,
  \[12586] ,
  \[10537] ,
  \[21649] ,
  \[2369] ,
  \[9663] ,
  \[22111] ,
  \[4029] ,
  \[10539] ,
  \[7277] ,
  \[12592] ,
  \[11399] ,
  \[5221] ,
  \[11731] ,
  \[5951] ,
  \[6419] ,
  \[3564] ,
  \[2705] ,
  \[8808] ,
  \[11393] ,
  \[14251] ,
  \[12923] ,
  \[22117] ,
  \[1511] ,
  \[5226] ,
  \[21651] ,
  \[22119] ,
  \[13060] ,
  \[4760] ,
  \[6087] ,
  \[13790] ,
  \[8476] ,
  \[1514] ,
  \[7617] ,
  \[22113] ,
  \[3903] ,
  \[22115] ,
  \[12593] ,
  \[4035] ,
  \[4765] ,
  \[11005] ,
  \[12596] ,
  \[6424] ,
  \[775] ,
  \[11740] ,
  \[10547] ,
  \[14256] ,
  \[9673] ,
  \[1182] ,
  \[12208] ,
  \[22121] ,
  \[13798] ,
  \[3572] ,
  \[7287] ,
  \[2713] ,
  \[12209] ,
  \[6429] ,
  \[12939] ,
  \[14262] ,
  \[8818] ,
  \[12203] ,
  \[12933] ,
  \[10545] ,
  \[13063] ,
  \[22127] ,
  \[11018] ,
  \[6095] ,
  \[13065] ,
  \[22129] ,
  \[4770] ,
  \[2382] ,
  \[7627] ,
  \[22123] ,
  \[782] ,
  \[13409] ,
  \[11013] ,
  \[1526] ,
  \[22125] ,
  \[11746] ,
  \[9681] ,
  \[10558] ,
  \[14263] ,
  \[4047] ,
  \[14266] ,
  \[21669] ,
  \[22131] ,
  \[12948] ,
  \[9684] ,
  \[12217] ,
  \[7296] ,
  \[5240] ,
  \[10559] ,
  \[5970] ,
  \[3582] ,
  \[2723] ,
  \[8826] ,
  \[789] ,
  \[13412] ,
  \[1195] ,
  \[10556] ,
  \[5245] ,
  \[13076] ,
  \[2728] ,
  \[21671] ,
  \[8494] ,
  \[7635] ,
  \[3921] ,
  \[13417] ,
  \[14277] ,
  \[6441] ,
  \[11753] ,
  \[4784] ,
  \[8101] ,
  \[1537] ,
  \[4055] ,
  \[794] ,
  \[11025] ,
  \[11755] ,
  \[10568] ,
  \[10900] ,
  \[14273] ,
  \[14276] ,
  \[3590] ,
  \[13415] ,
  \[12228] ,
  \[6446] ,
  \[12958] ,
  \[11762] ,
  \[13087] ,
  \[21673] ,
  \[4789] ,
  \[2733] ,
  \[8836] ,
  \[11761] ,
  \[2004] ,
  \[5252] ,
  \[10563] ,
  \[21675] ,
  \[403] ,
  \[404] ,
  \[10565] ,
  \[9699] ,
  \[405] ,
  \[10570] ,
  \[7645] ,
  \[22149] ,
  \[3599] ,
  \[10909] ,
  \[5988] ,
  \[6451] ,
  \[12961] ,
  \[9308] ,
  \[8111] ,
  \[4065] ,
  \[3206] ,
  \[14284] ,
  \[21687] ,
  \[13423] ,
  \[11035] ,
  \[1548] ,
  \[11765] ,
  \[10578] ,
  \[10910] ,
  \[14283] ,
  \[4796] ,
  \[21689] ,
  \[13425] ,
  \[8844] ,
  \[22151] ,
  \[21683] ,
  \[11771] ,
  \[12969] ,
  \[14292] ,
  \[2015] ,
  \[21685] ,
  \[13431] ,
  \[12234] ,
  \[2745] ,
  \[10576] ,
  \[8119] ,
  \[12963] ,
  \[414] ,
  \[7653] ,
  \[415] ,
  \[5266] ,
  \[416] ,
  \[21691] ,
  \[3940] ,
  \[12970] ,
  \[417] ,
  \[10919] ,
  \[14298] ,
  \[22153] ,
  \[14297] ,
  \[11044] ,
  \[3214] ,
  \[10913] ,
  \[22155] ,
  \[4074] ,
  \[11773] ,
  \[13434] ,
  \[6463] ,
  \[9319] ,
  \[21697] ,
  \[11775] ,
  \[2750] ,
  \[1559] ,
  \[3948] ,
  \[8854] ,
  \[13440] ,
  \[12247] ,
  \[10921] ,
  \[21693] ,
  \[11051] ,
  \[5271] ,
  \[11781] ,
  \[6800] ,
  \[10584] ,
  \[13442] ,
  \[12979] ,
  \[21695] ,
  \[2755] ,
  \[10586] ,
  \[8129] ,
  \[12243] ,
  \[12973] ,
  \[7663] ,
  \[22167] ,
  \[10927] ,
  \[22169] ,
  \[11787] ,
  \[13448] ,
  \[5278] ,
  \[10929] ,
  \[22163] ,
  \[4082] ,
  \[3223] ,
  \[0] ,
  \[6471] ,
  \[12981] ,
  \[5612] ,
  \[11053] ,
  \[22165] ,
  \[9328] ,
  \[8862] ,
  \[10597] ,
  \[2031] ,
  \[3958] ,
  \[22171] ,
  \[12257] ,
  \[11061] ,
  \[4422] ,
  \[8137] ,
  \[12989] ,
  \[13451] ,
  \[7671] ,
  \[12983] ,
  \[2767] ,
  \[1570] ,
  \[22177] ,
  \[436] ,
  \[22179] ,
  \[437] ,
  \[4091] ,
  \[438] ,
  \[22173] ,
  \[439] ,
  \[9336] ,
  \[6481] ,
  \[10206] ,
  \[22175] ,
  \[13454] ,
  \[8871] ,
  \[11796] ,
  \[10935] ,
  \[3966] ,
  \[11070] ,
  \[11407] ,
  \[22181] ,
  \[13460] ,
  \[12267] ,
  \[10211] ,
  \[5290] ,
  \[440] ,
  \[4431] ,
  \[441] ,
  \[8147] ,
  \[6489] ,
  \[442] ,
  \[13461] ,
  \[2775] ,
  \[7681] ,
  \[443] ,
  \[6822] ,
  \[11405] ,
  \[22187] ,
  \[10948] ,
  \[1581] ,
  \[12995] ,
  \[11077] ,
  \[22189] ,
  \[3241] ,
  \[12607] ,
  \[448] ,
  \[5630] ,
  \[22183] ,
  \[449] ,
  \[9346] ,
  \[12604] ,
  \[7689] ,
  \[22185] ,
  \[13464] ,
  \[3975] ,
  \[8881] ,
  \[12603] ,
  \[10215] ,
  \[8152] ,
  \[11080] ,
  \[22191] ,
  \[10952] ,
  \[13470] ,
  \[11082] ,
  \[450] ,
  \[2053] ,
  \[13807] ,
  \[451] ,
  \[5639] ,
  \[8157] ,
  \[6499] ,
  \[452] ,
  \[2785] ,
  \[11413] ,
  \[1926] ,
  \[453] ,
  \[12273] ,
  \[454] ,
  \[11415] ,
  \[455] ,
  \[11088] ,
  \[6105] ,
  \[456] ,
  \[457] ,
  \[9354] ,
  \[12617] ,
  \[11422] ,
  \[458] ,
  \[10959] ,
  \[12282] ,
  \[6838] ,
  \[13479] ,
  \[13811] ,
  \[12614] ,
  \[7699] ,
  \[3985] ,
  \[1597] ,
  \[12613] ,
  \[13473] ,
  \[7304] ,
  \[11090] ,
  \[8893] ,
  \[1202] ,
  \[12287] ,
  \[5649] ,
  \[12289] ,
  \[2794] ,
  \[11424] ,
  \[13481] ,
  \[463] ,
  \[9360] ,
  \[8169] ,
  \[6113] ,
  \[464] ,
  \[10238] ,
  \[1938] ,
  \[465] ,
  \[1209] ,
  \[11430] ,
  \[12628] ,
  \[4458] ,
  \[3261] ,
  \[13820] ,
  \[11432] ,
  \[10969] ,
  \[13487] ,
  \[11099] ,
  \[2404] ,
  \[3994] ,
  \[11096] ,
  \[10235] ,
  \[7314] ,
  \[2071] ,
  \[8174] ,
  \[10242] ,
  \[5657] ,
  \[12297] ,
  \[6851] ,
  \[8179] ,
  \[6123] ,
  \[474] ,
  \[8512] ,
  \[475] ,
  \[9372] ,
  \[12295] ,
  \[13826] ,
  \[1949] ,
  \[476] ,
  \[4467] ,
  \[12638] ,
  \[477] ,
  \[13100] ,
  \[3609] ,
  \[10979] ,
  \[13497] ,
  \[10976] ,
  \[7322] ,
  \[9379] ,
  \[5667] ,
  \[13838] ,
  \[6131] ,
  \[11443] ,
  \[14301] ,
  \[13103] ,
  \[10987] ,
  \[3618] ,
  \[13835] ,
  \[13110] ,
  \[14308] ,
  \[11451] ,
  \[3283] ,
  \[13112] ,
  \[12649] ,
  \[5672] ,
  \[13841] ,
  \[823] ,
  \[8191] ,
  \[2426] ,
  \[9389] ,
  \[21707] ,
  \[1960] ,
  \[5676] ,
  \[21709] ,
  \[7335] ,
  \[13847] ,
  \[6141] ,
  \[13849] ,
  \[14311] ,
  \[8199] ,
  \[4485] ,
  \[2097] ,
  \[3626] ,
  \[11455] ,
  \[6874] ,
  \[8533] ,
  \[10267] ,
  \[21711] ,
  \[4822] ,
  \[6149] ,
  \[12659] ,
  \[12654] ,
  \[103] ,
  \[10996] ,
  \[104] ,
  \[105] ,
  \[1241] ,
  \[1971] ,
  \[836] ,
  \[14316] ,
  \[13858] ,
  \[5689] ,
  \[9006] ,
  \[13129] ,
  \[11463] ,
  \[14321] ,
  \[10605] ,
  \[9739] ,
  \[13126] ,
  \[3638] ,
  \[13855] ,
  \[11472] ,
  \[4101] ,
  \[6887] ,
  \[14328] ,
  \[13132] ,
  \[2444] ,
  \[6159] ,
  \[11804] ,
  \[12664] ,
  \[843] ,
  \[114] ,
  \[5694] ,
  \[115] ,
  \[9742] ,
  \[116] ,
  \[21729] ,
  \[12670] ,
  \[117] ,
  \[1982] ,
  \[9014] ,
  \[13868] ,
  \[4109] ,
  \[5698] ,
  \[4839] ,
  \[3642] ,
  \[1254] ,
  \[5301] ,
  \[10614] ,
  \[7358] ,
  \[11473] ,
  \[14331] ,
  \[13864] ,
  \[11476] ,
  \[10288] ,
  \[13136] ,
  \[21731] ,
  \[3648] ,
  \[10622] ,
  \[8555] ,
  \[6167] ,
  \[13870] ,
  \[11482] ,
  \[850] ,
  \[121] ,
  \[14337] ,
  \[13142] ,
  \[122] ,
  \[12674] ,
  \[123] ,
  \[11813] ,
  \[14339] ,
  \[12673] ,
  \[124] ,
  \[10285] ,
  \[125] ,
  \[1261] ,
  \[11488] ,
  \[126] ,
  \[11820] ,
  \[127] ,
  \[10292] ,
  \[13878] ,
  \[128] ,
  \[6507] ,
  \[1993] ,
  \[4119] ,
  \[11822] ,
  \[21733] ,
  \[12682] ,
  \[12681] ,
  \[9027] ,
  \[21735] ,
  \[10626] ,
  \[13144] ,
  \[11486] ,
  \[1268] ,
  \[10630] ,
  \[22209] ,
  \[5317] ,
  \[10632] ,
  \[13150] ,
  \[3659] ,
  \[2462] ,
  \[6177] ,
  \[13880] ,
  \[10299] ,
  \[7707] ,
  \[11829] ,
  \[13152] ,
  \[7371] ,
  \[133] ,
  \[10296] ,
  \[134] ,
  \[21747] ,
  \[135] ,
  \[10638] ,
  \[12685] ,
  \[4127] ,
  \[21749] ,
  \[22211] ,
  \[1273] ,
  \[2802] ,
  \[13888] ,
  \[6517] ,
  \[21743] ,
  \[13887] ,
  \[12692] ,
  \[12691] ,
  \[11494] ,
  \[21745] ,
  \[8909] ,
  \[11496] ,
  \[10635] ,
  \[6185] ,
  \[11838] ,
  \[13155] ,
  \[21751] ,
  \[2471] ,
  \[8574] ,
  \[11107] ,
  \[4861] ,
  \[7717] ,
  \[22213] ,
  \[1615] ,
  \[13161] ,
  \[13891] ,
  \[22215] ,
  \[21757] ,
  \[11105] ,
  \[10648] ,
  \[12695] ,
  \[6525] ,
  \[4137] ,
  \[21759] ,
  \[2812] ,
  \[13898] ,
  \[21753] ,
  \[10644] ,
  \[1285] ,
  \[12309] ,
  \[21755] ,
  \[7389] ,
  \[13899] ,
  \[10646] ,
  \[13163] ,
  \[12306] ,
  \[22227] ,
  \[12305] ,
  \[6195] ,
  \[11848] ,
  \[13165] ,
  \[21761] ,
  \[7725] ,
  \[22229] ,
  \[3679] ,
  \[11119] ,
  \[151] ,
  \[22223] ,
  \[5339] ,
  \[152] ,
  \[882] ,
  \[13171] ,
  \[11113] ,
  \[153] ,
  \[22225] ,
  \[9050] ,
  \[11116] ,
  \[154] ,
  \[21767] ,
  \[155] ,
  \[4146] ,
  \[2820] ,
  \[156] ,
  \[6535] ,
  \[21769] ,
  \[2489] ,
  \[13505] ,
  \[157] ,
  \[22231] ,
  \[4878] ,
  \[158] ,
  \[21763] ,
  \[10654] ,
  \[13512] ,
  \[12319] ,
  \[21765] ,
  \[12316] ,
  \[22237] ,
  \[10660] ,
  \[12315] ,
  \[13175] ,
  \[21771] ,
  \[2829] ,
  \[7735] ,
  \[22239] ,
  \[11857] ,
  \[11129] ,
  \[22233] ,
  \[13181] ,
  \[163] ,
  \[22235] ,
  \[4154] ,
  \[11126] ,
  \[8931] ,
  \[164] ,
  \[6543] ,
  \[11125] ,
  \[165] ,
  \[11855] ,
  \[895] ,
  \[22241] ,
  \[13520] ,
  \[4889] ,
  \[12329] ,
  \[13189] ,
  \[8209] ,
  \[9401] ,
  \[13183] ,
  \[7013] ,
  \[7743] ,
  \[22247] ,
  \[3697] ,
  \[11138] ,
  \[11868] ,
  \[2839] ,
  \[22249] ,
  \[10672] ,
  \[22243] ,
  \[3303] ,
  \[13192] ,
  \[4163] ,
  \[13529] ,
  \[22245] ,
  \[6553] ,
  \[11135] ,
  \[2110] ,
  \[21789] ,
  \[13525] ,
  \[22251] ,
  \[13198] ,
  \[5361] ,
  \[8217] ,
  \[4503] ,
  \[13531] ,
  \[7753] ,
  \[7024] ,
  \[2848] ,
  \[9413] ,
  \[21791] ,
  \[13538] ,
  \[10681] ,
  \[1654] ,
  \[181] ,
  \[11879] ,
  \[12341] ,
  \[11144] ,
  \[182] ,
  \[6561] ,
  \[4173] ,
  \[183] ,
  \[11146] ,
  \[184] ,
  \[8952] ,
  \[185] ,
  \[186] ,
  \[187] ,
  \[11152] ,
  \[188] ,
  \[10689] ,
  \[21793] ,
  \[14007] ,
  \[8227] ,
  \[4513] ,
  \[21795] ,
  \[7761] ,
  \[2856] ,
  \[14004] ,
  \[2127] ,
  \[14003] ,
  \[11158] ,
  \[11888] ,
  \[6905] ,
  \[22269] ,
  \[3321] ,
  \[13547] ,
  \[4182] ,
  \[5711] ,
  \[6571] ,
  \[8960] ,
  \[193] ,
  \[194] ,
  \[13543] ,
  \[195] ,
  \[13545] ,
  \[22271] ,
  \[9094] ,
  \[8235] ,
  \[10699] ,
  \[14017] ,
  \[5719] ,
  \[4522] ,
  \[12359] ,
  \[6579] ,
  \[10693] ,
  \[5383] ,
  \[12353] ,
  \[14014] ,
  \[14013] ,
  \[1671] ,
  \[11898] ,
  \[4190] ,
  \[22273] ,
  \[13559] ,
  \[8970] ,
  \[22275] ,
  \[11166] ,
  \[13553] ,
  \[11895] ,
  \[4530] ,
  \[3339] ,
  \[8245] ,
  \[4199] ,
  \[14028] ,
  \[6920] ,
  \[5729] ,
  \[12369] ,
  \[2874] ,
  \[6589] ,
  \[8978] ,
  \[7781] ,
  \[7052] ,
  \[11506] ,
  \[14024] ,
  \[12366] ,
  \[22287] ,
  \[12365] ,
  \[10317] ,
  \[2149] ,
  \[22289] ,
  \[14025] ,
  \[10319] ,
  \[4539] ,
  \[22283] ,
  \[6928] ,
  \[13902] ,
  \[12709] ,
  \[22285] ,
  \[11175] ,
  \[1688] ,
  \[8253] ,
  \[2880] ,
  \[11518] ,
  \[22291] ,
  \[5737] ,
  \[13570] ,
  \[6597] ,
  \[14038] ,
  \[12379] ,
  \[13909] ,
  \[8988] ,
  \[6203] ,
  \[14034] ,
  \[7063] ,
  \[12376] ,
  \[22297] ,
  \[12375] ,
  \[14035] ,
  \[1693] ,
  \[11522] ,
  \[4549] ,
  \[22293] ,
  \[6938] ,
  \[12719] ,
  \[10323] ,
  \[9457] ,
  \[13579] ,
  \[11183] ,
  \[10326] ,
  \[22295] ,
  \[1698] ,
  \[5015] ,
  \[3357] ,
  \[8263] ,
  \[11190] ,
  \[1302] ,
  \[7405] ,
  \[5747] ,
  \[12387] ,
  \[11192] ,
  \[10331] ,
  \[8996] ,
  \[14047] ,
  \[7072] ,
  \[6213] ,
  \[8602] ,
  \[12386] ,
  \[11198] ,
  \[12390] ,
  \[13915] ,
  \[567] ,
  \[6946] ,
  \[4558] ,
  \[9464] ,
  \[13587] ,
  \[11199] ,
  \[902] ,
  \[13921] ,
  \[8271] ,
  \[10335] ,
  \[5755] ,
  \[12725] ,
  \[2171] ,
  \[2509] ,
  \[12730] ,
  \[12397] ,
  \[10341] ,
  \[11539] ,
  \[14057] ,
  \[909] ,
  \[12001] ,
  \[7080] ,
  \[13592] ,
  \[1315] ,
  \[6221] ;
assign
  \[8612]  = ~\[10774]  & (~v15 & v14),
  \[12396]  = ~\[5405]  | (v2 | (~v1 | v0)),
  \[11535]  = ~v12 | (~v11 | v9),
  \[10348]  = ~v7 | (~v5 | v4),
  \[14053]  = ~\[2097]  | (~v15 | (~v13 | v12)),
  \[4566]  = ~v2 & (v1 & ~v0),
  \[14056]  = v4 | (v3 | (~v2 | ~v0)),
  \[6956]  = ~\[11627]  & (~v15 & (v14 & ~v13)),
  \[13200]  = ~v3 | (~v1 | v0),
  \[4900]  = ~\[12649]  & (~v15 & (v14 & ~v13)),
  \[12737]  = v8 | (~v7 | ~v4),
  \[13597]  = ~v11 | ~v8,
  \[10344]  = ~v7 | (~v5 | v4),
  \[9477]  = ~v12 & (v7 & (v5 & ~v4)),
  \[3375]  = ~v12 & (v11 & ~v9),
  \[8281]  = ~\[10959]  & (v7 & (~v5 & ~v3)),
  \[4905]  = ~v6 & (~v5 & ~v8),
  \[5765]  = ~v6 & (~v5 & (~\[12217]  & ~v3)),
  \[12005]  = ~v7 | v5,
  \[1322]  = ~\[98]  & (~\[97]  & (~\[96]  & ~\[95] )),
  \[5037]  = ~v6 & (~v5 & ~v8),
  \[12740]  = v11 | (~v10 | ~v9),
  \[10352]  = ~v7 | (~v5 | v4),
  \[12012]  = ~v3 | (~v1 | v0),
  \[7427]  = v11 & (~v9 & ~v7),
  \[13937]  = v11 | (~v10 | ~v9),
  \[7090]  = ~\[11552]  & (~v15 & (v14 & ~v13)),
  \[6231]  = ~\[11986]  & (~v2 & (v1 & ~v0)),
  \[8620]  = ~v3 & (v2 & ~v1),
  \[8289]  = v12 & (~v10 & ~v9),
  \[3715]  = ~v10 & (~v9 & ~v12),
  \[584]  = ~\[14256]  & (~\[14213]  & ~\[14337] ),
  \[4575]  = ~v12 & (v11 & v8),
  \[11545]  = ~v12 | (~v11 | v9),
  \[6964]  = v3 & (v1 & ~v0),
  \[13206]  = ~v15 | (~v13 | ~\[3787] ),
  \[1329]  = ~\[94]  & (~\[93]  & (~\[92]  & ~\[91] )),
  \[14065]  = ~\[2071]  | (~v15 | (~v13 | v12)),
  \[9484]  = v5 & ~v4,
  \[4910]  = ~v3 & (v2 & ~v1),
  \[11552]  = ~v11 | ~v8,
  \[7098]  = ~v2 & (v1 & ~v0),
  \[6239]  = ~v13 & (v11 & ~v9),
  \[12749]  = v8 | (~v7 | ~v4),
  \[14072]  = ~v10 | ~v9,
  \[14071]  = ~\[2053]  | (v3 | (~v2 | v1)),
  \[5773]  = ~v12 & (v11 & ~v9),
  \[3385]  = ~\[13388]  & (v7 & ~v5),
  \[2526]  = ~v14 & (v13 & ~v12),
  \[8629]  = v12 & (~v10 & ~v9),
  \[21807]  = ~\[7707]  | (~\[7717]  | (v14 | ~v13)),
  \[12745]  = ~\[22109]  | (~\[22107]  | (~\[22105]  | ~\[22103] )),
  \[21471]  = ~\[10057]  | (v10 | ~v9),
  \[926]  = ~\[299]  & (~\[298]  & (~\[300]  & ~\[12494] )),
  \[21809]  = ~\[7689]  | (~\[7699]  | (v14 | ~v13)),
  \[12020]  = ~v2 | v1,
  \[13948]  = v11 | (~v10 | ~v9),
  \[2193]  = ~v6 & (~v5 & ~v8),
  \[21803]  = ~\[7743]  | (~\[7753]  | (v14 | ~v13)),
  \[12752]  = v11 | (~v10 | ~v9),
  \[13219]  = ~v3 | (~v1 | v0),
  \[21805]  = ~\[7725]  | (~\[7735]  | (v14 | ~v13)),
  \[8299]  = ~\[10952]  & (~v3 & (v2 & ~v1)),
  \[3725]  = ~v6 & (~v5 & (~\[13235]  & ~v3)),
  \[21477]  = ~v15 | (v13 | (v2 | v1)),
  \[4585]  = ~v6 & (~v5 & ~\[12806] ),
  \[13216]  = ~v15 | ~v13,
  \[21479]  = ~\[10028]  | (v11 | (~v10 | ~v8)),
  \[21811]  = ~\[7671]  | (~\[7681]  | (v14 | ~v13)),
  \[12028]  = ~v0 | ~v2,
  \[2531]  = ~v10 & (v8 & ~v7),
  \[597]  = ~\[464]  & (~\[463]  & (~\[465]  & ~\[14132] )),
  \[10702]  = ~v2 | v1,
  \[14075]  = ~v15 | (~v13 | v12),
  \[21473]  = ~\[10049]  | (v11 | ~v10),
  \[11561]  = ~v11 | ~v8,
  \[4922]  = ~\[12638]  & (~v15 & (v14 & ~v13)),
  \[6249]  = ~v6 & (~v5 & ~\[11976] ),
  \[14082]  = ~v10 | ~v9,
  \[21475]  = v14 | (v13 | (v2 | v1)),
  \[3394]  = ~\[13409]  & (~v12 & (v11 & ~v9)),
  \[14081]  = ~\[2031]  | (v3 | (~v2 | ~v0)),
  \[5783]  = ~v6 & (~v5 & (~\[12209]  & ~v3)),
  \[933]  = ~\[293]  & (~\[292]  & (~\[291]  & ~\[290] )),
  \[8639]  = ~\[10787]  & (~v2 & (v1 & ~v0)),
  \[204]  = ~\[11581]  & (~\[11579]  & ~\[11587] ),
  \[21817]  = ~\[7617]  | (~\[7627]  | (v14 | ~v13)),
  \[5055]  = ~v11 & (v10 & (v9 & ~v8)),
  \[205]  = ~\[11593]  & (~\[11591]  & (~v15 & v14)),
  \[11568]  = ~v6 | (~v5 | v4),
  \[206]  = ~\[11602]  & (~\[11600]  & (~v15 & v14)),
  \[3000]  = ~\[13597]  & (~v14 & (v13 & ~v12)),
  \[21481]  = ~v11 | (~v9 | ~\[10021] ),
  \[21819]  = ~\[7599]  | (~\[7609]  | (v14 | ~v13)),
  \[4927]  = ~v8 & (v7 & ~v5),
  \[12760]  = ~v11 | ~v8,
  \[207]  = ~\[11610]  & (~\[11608]  & (~v15 & v14)),
  \[13958]  = v11 | (~v10 | ~v9),
  \[13227]  = ~v2 | v1,
  \[21813]  = ~\[7653]  | (~\[7663]  | (v14 | ~v13)),
  \[1344]  = ~\[87]  & (~\[86]  & (~\[85]  & ~\[84] )),
  \[3733]  = ~v10 & (~v9 & ~v12),
  \[9107]  = ~v6 & v4,
  \[4593]  = ~v12 & (v11 & v8),
  \[21815]  = ~\[7635]  | (~\[7645]  | (v14 | ~v13)),
  \[6982]  = ~v2 & (v1 & ~v0),
  \[21487]  = v14 | (~v12 | (v2 | v1)),
  \[10378]  = ~v2 | (~v1 | v0),
  \[3008]  = v3 & (v1 & ~v0),
  \[21489]  = ~\[9991]  | (v10 | ~v9),
  \[21821]  = ~\[7574]  | (~\[7579]  | ~\[7591] ),
  \[14085]  = ~v15 | (~v13 | v12),
  \[12037]  = ~\[21975]  | (~\[21973]  | (~\[21971]  | ~\[21969] )),
  \[6257]  = ~v13 & (v11 & ~v9),
  \[10711]  = ~v0 | ~v2,
  \[21483]  = ~v15 | (~v12 | (v2 | v1)),
  \[940]  = ~\[289]  & (~\[288]  & (~\[287]  & ~\[286] )),
  \[4931]  = v1 & ~v0,
  \[2543]  = ~\[13811]  & (~v3 & (v2 & ~v1)),
  \[11571]  = ~v11 | (~v8 | v7),
  \[211]  = ~\[11649]  & (~\[11647]  & (~v15 & v14)),
  \[5791]  = ~v12 & (v11 & ~v9),
  \[8647]  = v12 & (~v10 & v8),
  \[12769]  = ~v11 | ~v8,
  \[212]  = ~\[11657]  & (~\[11655]  & (~v15 & v14)),
  \[11904]  = ~v0 | ~v2,
  \[21485]  = ~\[10007]  | (v15 | (~v14 | ~v13)),
  \[213]  = ~\[11666]  & (~\[11664]  & (~v15 & v14)),
  \[10376]  = ~\[21615]  | (~\[21613]  | (~\[21611]  | ~\[21609] )),
  \[214]  = ~\[11674]  & (~\[11672]  & (~v15 & v14)),
  \[21827]  = ~\[7519]  | (~\[7529]  | (v14 | ~v13)),
  \[9841]  = ~v8 & (v3 & ~v1),
  \[215]  = ~\[11688]  & ~\[11683] ,
  \[216]  = ~\[11689]  & (~v3 & (~\[11692]  & ~\[11698] )),
  \[21491]  = ~\[9983]  | (v11 | ~v10),
  \[21829]  = ~\[7501]  | (~\[7511]  | (v14 | ~v13)),
  \[7455]  = v1 & ~v0,
  \[217]  = ~\[11705]  & (~\[11703]  & (~v15 & v14)),
  \[9844]  = ~v14 & v12,
  \[13968]  = ~\[2215]  | (~v3 | (~v1 | v0)),
  \[218]  = ~\[11713]  & (~\[11711]  & (~v15 & v14)),
  \[4209]  = ~v6 & (~v5 & ~\[12995] ),
  \[21823]  = ~\[7552]  | (~\[7557]  | ~\[7569] ),
  \[11579]  = ~v3 | (~v1 | v0),
  \[12041]  = ~v6 | (~v5 | v4),
  \[3743]  = ~v6 & (~v5 & (~\[13227]  & ~v3)),
  \[21825]  = ~\[7537]  | (~\[7547]  | (v14 | ~v13)),
  \[13969]  = ~v10 | ~v9,
  \[11576]  = ~\[21877]  | (~\[21875]  | (~\[21873]  | ~\[21871] )),
  \[21497]  = ~\[9958]  | (~v8 | (v2 | ~v0)),
  \[13963]  = ~\[22365]  | (~\[22363]  | (~\[22361]  | ~\[22359] )),
  \[5405]  = ~v8 & (v7 & ~v5),
  \[14093]  = v8 | (~v7 | ~v4),
  \[10387]  = ~v2 | (~v1 | v0),
  \[3018]  = ~\[13587]  & (~v14 & (v13 & ~v12)),
  \[6995]  = ~v6 & ~v5,
  \[14096]  = v11 | (~v10 | ~v9),
  \[21499]  = ~v11 | (~v9 | ~\[9955] ),
  \[13235]  = ~v0 | ~v2,
  \[21831]  = ~\[7483]  | (~\[7493]  | (v14 | ~v13)),
  \[2551]  = ~v12 & (~v10 & v8),
  \[6267]  = ~v6 & (~v5 & (~\[11967]  & ~v2)),
  \[21493]  = v14 | (v13 | (v2 | ~v0)),
  \[11581]  = ~v6 | (~v5 | v4),
  \[8657]  = ~\[10777]  & (v7 & (~v5 & ~v3)),
  \[13972]  = ~v15 | (~v13 | v12),
  \[12779]  = ~v11 | (~v8 | v7),
  \[10383]  = v3 | (~v2 | (~v1 | v0)),
  \[11914]  = ~v4 | ~v7,
  \[21495]  = ~v15 | (v13 | (v2 | ~v0)),
  \[223]  = ~\[11762]  & (~v2 & (~\[11765]  & ~\[11771] )),
  \[4944]  = ~\[12628]  & (~v15 & (v14 & ~v13)),
  \[224]  = ~\[11775]  & (~\[11773]  & ~\[11781] ),
  \[954]  = ~\[282]  & (~\[281]  & (~\[280]  & ~\[279] )),
  \[12776]  = ~v6 | (~v5 | v4),
  \[225]  = ~v6 & (~v5 & (~\[11755]  & ~\[11761] )),
  \[10728]  = ~\[21697]  | (~\[21695]  | (~\[21693]  | ~\[21691] )),
  \[1361]  = ~\[10449]  & (~\[10416]  & ~\[10514] ),
  \[4217]  = ~v12 & (~v10 & v8),
  \[12050]  = v6 | ~v4,
  \[11587]  = ~\[7024]  | (~v11 | (~v8 | v7)),
  \[13248]  = ~v6 | (~v5 | v4),
  \[3751]  = ~v10 & (~v9 & ~v12),
  \[13978]  = ~\[2259]  | (~v3 | (~v1 | v0)),
  \[6607]  = ~\[11796]  & (~v2 & (v1 & ~v0)),
  \[4949]  = ~v8 & (v7 & ~v5),
  \[11921]  = ~\[21949]  | (~\[21947]  | ~\[21951] ),
  \[10724]  = ~v12 | (v10 | ~v8),
  \[6272]  = ~v15 & (v14 & ~v13),
  \[13979]  = ~v10 | ~v9,
  \[13244]  = ~\[22215]  | (~\[22213]  | (~\[22211]  | ~\[22209] )),
  \[3026]  = ~v2 & (v1 & ~v0),
  \[7803]  = ~v9 & (~v7 & ~v10),
  \[22307]  = ~\[2856]  | (~\[2848]  | (~v7 | v5)),
  \[13245]  = ~v2 | v1,
  \[2561]  = ~\[13826]  & (~v6 & (v4 & ~v3)),
  \[6276]  = ~v9 & ~v7,
  \[22309]  = ~\[2829]  | (~\[2839]  | (v14 | ~v13)),
  \[11591]  = ~\[7013]  | (v2 | (~v1 | v0)),
  \v16.0  = \[0] ,
  \[13982]  = ~v15 | (~v13 | v12),
  \[12789]  = ~v6 | (~v5 | v4),
  \[11924]  = ~\[1083]  | (~\[1090]  | (~\[1076]  | ~\[1063] )),
  \[12784]  = ~\[22117]  | (~\[22115]  | (~\[22113]  | ~\[22111] )),
  \[9130]  = ~v3 & (v2 & ~v1),
  \[4954]  = ~v2 & (v1 & ~v0),
  \[12056]  = ~v0 | ~v2,
  \[9861]  = ~v12 & (~v7 & (v6 & v4)),
  \[10738]  = ~v2 | v1,
  \[7474]  = ~v2 & (v1 & ~v0),
  \[10007]  = ~v2 & (~v1 & ~v12),
  \[6615]  = ~v13 & (~v10 & v8),
  \[11930]  = ~v4 | ~v7,
  \[21849]  = ~\[7322]  | (~\[7314]  | (~v7 | v5)),
  \[2569]  = ~v12 & (~v10 & v8),
  \[22311]  = ~v4 | (~v7 | (~\[2820]  | ~\[2812] )),
  \[3761]  = ~\[13219]  & (v7 & ~v5),
  \[11202]  = ~v6 | (~v5 | v4),
  \[2902]  = ~v14 & (v13 & ~v12),
  \[13988]  = ~\[2237]  | (v2 | (~v1 | v0)),
  \[1374]  = ~\[74]  & (~\[73]  & (~\[75]  & ~\[10376] )),
  \[12792]  = ~v11 | (~v8 | v7),
  \[10733]  = ~\[8731]  | (v3 | (~v2 | ~v0)),
  \[13989]  = ~v10 | ~v9,
  \[11593]  = v13 | (~v11 | ~v8),
  \[13254]  = ~\[3659]  | (~v15 | (~v13 | v12)),
  \[3036]  = ~\[13579]  & (~v14 & (v13 & ~v12)),
  \[10735]  = ~v12 | (v10 | ~v8),
  \[9869]  = ~v7 & (v6 & v4),
  \[1710]  = ~\[14241]  & (~v14 & (v13 & ~v12)),
  \[22317]  = ~\[2750]  | (~\[2755]  | ~\[2767] ),
  \[13256]  = v3 | (~v2 | v1),
  \[11208]  = ~\[7803]  | (v14 | (~v13 | v12)),
  \[11938]  = ~v4 | ~v7,
  \[21851]  = ~\[7304]  | (~\[7296]  | (~v7 | v5)),
  \[12068]  = ~v0 | ~v2,
  \[8674]  = ~v3 & (v2 & ~v1),
  \[12400]  = v15 | (~v14 | ~v12),
  \[22319]  = ~\[2728]  | (~\[2733]  | ~\[2745] ),
  \[5427]  = ~v8 & (~v6 & v4),
  \[10741]  = ~v6 | (~v5 | v4),
  \[22313]  = ~v4 | (~v7 | (~\[2802]  | ~\[2794] )),
  \[971]  = ~\[12282]  & (~\[12243]  & ~\[12359] ),
  \[13262]  = ~v15 | (~v13 | ~\[3697] ),
  \[6289]  = ~\[11958]  & (v3 & (v1 & ~v0)),
  \[13992]  = ~v15 | (~v13 | v12),
  \[22315]  = ~\[2775]  | (~\[2785]  | (v14 | ~v13)),
  \[5094]  = ~v4 & (~v2 & (v1 & ~v0)),
  \[7483]  = ~v10 & (~v9 & ~v12),
  \[12796]  = ~v1 | v0,
  \[12065]  = ~\[21979]  | (~\[21977]  | ~\[21981] ),
  \[1381]  = ~\[68]  & (~\[67]  & (~\[66]  & ~\[65] )),
  \[11210]  = ~v3 | (~v1 | v0),
  \[6625]  = ~v6 & (~v5 & ~\[11787] ),
  \[4237]  = ~v10 & (v8 & ~v7),
  \[10747]  = ~\[8707]  | (v15 | (~v14 | ~v12)),
  \[9143]  = ~v6 & ~v5,
  \[3770]  = ~v10 & (~v9 & (~v12 & ~\[13216] )),
  \[2579]  = ~\[13820]  & (~v3 & (v2 & ~v1)),
  \[12408]  = ~\[5383]  | (~v3 | (~v1 | v0)),
  \[22321]  = ~\[2713]  | (~\[2723]  | (v14 | ~v13)),
  \[11212]  = ~v6 | (~v5 | v4),
  \[13998]  = ~\[634]  | (~\[641]  | (~\[627]  | ~\[672] )),
  \[10749]  = ~v0 | ~v2,
  \[21853]  = ~\[7277]  | (~\[7287]  | (v15 | ~v14)),
  \[12071]  = ~v6 | (~v5 | v4),
  \[12409]  = ~v10 | ~v9,
  \[3044]  = v3 & (v1 & ~v0),
  \[21855]  = ~\[7259]  | (~\[7269]  | (v15 | ~v14)),
  \[13264]  = v3 | (~v2 | ~v0),
  \[1388]  = ~\[64]  & (~\[63]  & (~\[62]  & ~\[61] )),
  \[6294]  = ~v15 & (v14 & ~v13),
  \[7823]  = ~v10 & (~v9 & ~v12),
  \[22327]  = ~\[2659]  | (~\[2669]  | (v14 | ~v13)),
  \[11218]  = ~\[7781]  | (v14 | (~v13 | v12)),
  \[2918]  = ~v3 & (v2 & ~v1),
  \[1721]  = ~v6 & (~v5 & (~v8 & ~\[14236] )),
  \[11948]  = ~v6 | (~v5 | v4),
  \[3778]  = ~v2 & (v1 & ~v0),
  \[22329]  = ~\[2641]  | (~\[2651]  | (v14 | ~v13)),
  \[10752]  = ~v6 | (~v5 | v4),
  \[13270]  = ~v15 | (~v13 | ~\[3679] ),
  \[12077]  = ~\[6053]  | (v15 | (~v14 | v13)),
  \[8685]  = ~v10 & (v8 & ~v7),
  \[10021]  = ~v2 & (~v1 & ~v8),
  \[4971]  = ~v8 & (~v6 & v4),
  \[12412]  = v15 | (~v14 | ~v12),
  \[6298]  = ~v9 & ~v7,
  \[22323]  = ~\[2695]  | (~\[2705]  | (v14 | ~v13)),
  \[12079]  = v3 | (~v2 | v1),
  \[22325]  = ~\[2677]  | (~\[2687]  | (v14 | ~v13)),
  \[6633]  = ~v13 & (~v10 & v8),
  \[21867]  = ~\[7143]  | (~\[7153]  | (v15 | ~v14)),
  \[2587]  = ~v12 & (~v10 & v8),
  \[7493]  = ~\[11335]  & (~v3 & (v2 & v0)),
  \[10028]  = ~v2 & ~v1,
  \[10758]  = ~\[8685]  | (v15 | (~v14 | ~v12)),
  \[985]  = ~\[269]  & (~\[268]  & (~\[270]  & ~\[12179] )),
  \[256]  = ~\[12068]  & (~v3 & (~\[12071]  & ~\[12077] )),
  \[21869]  = ~v4 | (~v7 | (~\[7134]  | ~\[7126] )),
  \[13605]  = ~v11 | ~v8,
  \[12418]  = ~\[5361]  | (v3 | (~v2 | v1)),
  \[257]  = ~\[12079]  & (~\[12085]  & (v7 & ~v5)),
  \[22331]  = ~\[2623]  | (~\[2633]  | (v14 | ~v13)),
  \[13610]  = ~v0 | ~v2,
  \[258]  = ~\[12088]  & (~\[12094]  & (v7 & ~v5)),
  \[21863]  = ~\[7180]  | (~v11 | (~\[7176]  | ~\[7193] )),
  \[259]  = ~\[12100]  & (~\[12098]  & (~v14 & v13)),
  \[12419]  = ~v10 | ~v9,
  \[3054]  = ~\[13570]  & (~v14 & (v13 & ~v12)),
  \[21865]  = ~\[7170]  | (~\[7162]  | (~v7 | v5)),
  \[7833]  = ~\[11183]  & (v3 & (v1 & ~v0)),
  \[22337]  = ~\[2569]  | (~\[2579]  | (v14 | ~v13)),
  \[3787]  = ~v10 & (~v9 & ~v12),
  \[11958]  = ~v6 | (~v5 | v4),
  \[21871]  = ~v4 | (~v7 | (~\[7116]  | ~\[7108] )),
  \[12088]  = v3 | (~v2 | ~v0),
  \[1732]  = ~\[14230]  & (~v14 & (v13 & ~v12)),
  \[22339]  = ~\[2551]  | (~\[2561]  | (v14 | ~v13)),
  \[10762]  = ~\[8674]  | (~v7 | v5),
  \[260]  = ~\[12110]  & (~\[12108]  & (~v15 & v14)),
  \[12422]  = v15 | (~v14 | ~v12),
  \[261]  = ~\[12118]  & (~\[12116]  & (~v15 & v14)),
  \[22333]  = ~\[2605]  | (~\[2615]  | (v14 | ~v13)),
  \[5449]  = ~v8 & (~v6 & v4),
  \[7108]  = ~\[11545]  & (~v15 & v14),
  \[11224]  = ~v3 | (~v1 | v0),
  \[262]  = ~\[12127]  & (~\[12125]  & (~v14 & v13)),
  \[992]  = ~\[263]  & (~\[262]  & (~\[261]  & ~\[260] )),
  \[263]  = ~\[12130]  & (~v2 & (~\[12133]  & ~\[12139] )),
  \[22335]  = ~\[2587]  | (~\[2597]  | (v14 | ~v13)),
  \[1737]  = ~v6 & (~v5 & ~v8),
  \[9161]  = ~v6 & ~v5,
  \[21877]  = ~\[7052]  | ~\[7063] ,
  \[2597]  = ~v6 & (~v5 & (~\[13798]  & ~v3)),
  \[12085]  = ~\[6033]  | (v15 | ~v14),
  \[2931]  = ~v6 & v4,
  \[22341]  = ~\[2526]  | (~\[2531]  | ~\[2543] ),
  \[268]  = ~\[12189]  & (~\[12195]  & (~v6 & v4)),
  \[4259]  = ~v10 & (v8 & ~v7),
  \[3062]  = ~v2 & (v1 & ~v0),
  \[21873]  = ~v4 | (~v7 | (~\[7098]  | ~\[7090] )),
  \[269]  = ~\[12197]  & (~\[12203]  & (v7 & ~v5)),
  \[10764]  = ~v12 | (v10 | ~v8),
  \[999]  = ~\[259]  & (~\[258]  & (~\[257]  & ~\[256] )),
  \[13622]  = ~v11 | ~v8,
  \[12429]  = ~\[5339]  | (v3 | (~v2 | ~v0)),
  \[21875]  = ~v4 | (~v7 | (~\[7080]  | ~\[7072] )),
  \[7841]  = ~v10 & (~v9 & ~v13),
  \[604]  = ~\[458]  & (~\[457]  & (~\[456]  & ~\[455] )),
  \[13283]  = ~v15 | (~v13 | v12),
  \[12098]  = ~v4 | (~v7 | ~\[6006] ),
  \[12430]  = ~v10 | ~v9,
  \[1742]  = ~v3 & (v2 & ~v1),
  \[11967]  = ~v1 | v0,
  \[7116]  = ~v3 & (v2 & v0),
  \[270]  = ~\[12181]  & (~\[12187]  & (v7 & ~v5)),
  \[3402]  = ~v2 & (v1 & ~v0),
  \[13627]  = ~\[22297]  | (~\[22295]  | (~\[22293]  | ~\[22291] )),
  \[13291]  = ~v15 | ~v13,
  \[4993]  = ~v8 & (~v6 & v4),
  \[8310]  = ~v9 & (~v7 & (~v10 & ~\[10948] )),
  \[12094]  = ~\[6015]  | (v15 | ~v14),
  \[11233]  = v6 | ~v4,
  \[6653]  = ~v10 & (v8 & ~v7),
  \[11966]  = ~\[21959]  | (~\[21957]  | (~\[21955]  | ~\[21953] )),
  \[21887]  = ~\[6964]  | (~\[6956]  | (v6 | ~v4)),
  \[10777]  = ~v0 | ~v2,
  \[21889]  = ~\[6946]  | (~\[6938]  | (~v7 | v5)),
  \[8314]  = v5 & ~v4,
  \[3071]  = ~v12 & (v11 & v8),
  \[10049]  = ~v2 & (~v1 & ~v9),
  \[11241]  = ~v3 | (~v1 | v0),
  \[279]  = ~\[12289]  & (~\[12287]  & (~v14 & v13)),
  \[611]  = ~\[454]  & (~\[453]  & (~\[452]  & ~\[451] )),
  \[10774]  = ~v12 | (v10 | ~v8),
  \[9176]  = ~\[10493]  & (~v15 & v14),
  \[13632]  = ~\[2931]  | (v3 | (~v2 | ~v0)),
  \[12439]  = ~\[5317]  | (v3 | (~v2 | v1)),
  \[4603]  = ~v6 & (~v5 & (~\[12796]  & ~v2)),
  \[2215]  = ~v8 & (v7 & ~v5),
  \[7851]  = ~\[11175]  & (~v3 & (v2 & v0)),
  \[13294]  = ~v0 | ~v2,
  \[12433]  = v15 | (~v14 | ~v12),
  \[2946]  = ~\[13622]  & (~v14 & (v13 & ~v12)),
  \[21891]  = ~\[6928]  | (~\[6920]  | (~v7 | v5)),
  \[12440]  = ~v10 | ~v9,
  \[22359]  = ~\[2335]  | (~v15 | (~\[2343]  | ~\[2357] )),
  \[3411]  = ~v12 & (v11 & ~v9),
  \[7126]  = ~\[11535]  & (~v15 & v14),
  \[280]  = ~\[12297]  & (~\[12295]  & (~v14 & v13)),
  \[1754]  = ~\[14220]  & (~v14 & (v13 & ~v12)),
  \[281]  = ~\[12306]  & (~v11 & (~\[12309]  & ~\[12305] )),
  \[282]  = ~\[12316]  & (~v11 & (~\[12319]  & ~\[12315] )),
  \[8320]  = ~v3 & (v2 & v0),
  \[7859]  = ~v10 & (~v9 & ~v13),
  \[13634]  = v12 | (~v11 | ~v8),
  \[11976]  = ~v3 | (~v1 | v0),
  \[11250]  = ~v7 | v5,
  \[10057]  = ~v2 & (~v1 & ~v8),
  \[1759]  = ~v8 & (v7 & ~v5),
  \[286]  = ~\[12366]  & (~v11 & (~\[12369]  & ~\[12365] )),
  \[10787]  = ~v4 | ~v7,
  \[21501]  = ~v15 | (~v12 | (v2 | ~v0)),
  \[287]  = ~\[12376]  & (~v11 & (~\[12379]  & ~\[12375] )),
  \[22361]  = ~\[2325]  | (~\[2330]  | ~\[2320] ),
  \[3081]  = ~v6 & (~v5 & ~\[13559] ),
  \[9184]  = v3 & (v1 & ~v0),
  \[288]  = ~\[12387]  & (~v11 & (~\[12390]  & ~\[12386] )),
  \[289]  = ~\[12397]  & (~v11 & (~\[12400]  & ~\[12396] )),
  \[5471]  = ~v6 & (~v5 & ~v8),
  \[5809]  = ~v12 & (v11 & ~v9),
  \[12449]  = v3 | (~v2 | ~v0),
  \[2954]  = ~v3 & (v2 & ~v1),
  \[13641]  = ~\[2918]  | (~v6 | (~v5 | v4)),
  \[4614]  = ~\[12792]  & (v15 & (v13 & ~v12)),
  \[12443]  = v15 | (~v14 | ~v12),
  \[1030]  = ~\[12065]  & (~\[12037]  & (~\[12001]  & ~\[11966] )),
  \[14103]  = v8 | (~v7 | ~v4),
  \[7134]  = ~v3 & (v2 & ~v1),
  \[14106]  = v11 | (~v10 | ~v9),
  \[11257]  = ~\[21809]  | (~\[21807]  | (~\[21805]  | ~\[21803] )),
  \[4280]  = ~\[12958]  & (~v12 & (~v10 & v8)),
  \[627]  = ~\[449]  & (~\[448]  & (~\[450]  & ~\[13963] )),
  \[3421]  = ~\[13396]  & (~v6 & v4),
  \[1033]  = ~\[13132]  & (~\[12851]  & (~\[12529]  & ~\[12208] )),
  \[13648]  = ~v0 | ~v2,
  \[1763]  = v1 & ~v0,
  \[290]  = ~\[12409]  & (~v11 & (~\[12412]  & ~\[12408] )),
  \[11259]  = ~v3 | (~v1 | v0),
  \[291]  = ~\[12419]  & (~v11 & (~\[12422]  & ~\[12418] )),
  \[22363]  = ~\[2307]  | (~v3 | (~\[2303]  | ~\[2298] )),
  \[292]  = ~\[12430]  & (~v11 & (~\[12433]  & ~\[12429] )),
  \[7869]  = ~\[11166]  & (~v3 & (v2 & ~v1)),
  \[293]  = ~\[12440]  & (~v11 & (~\[12443]  & ~\[12439] )),
  \[22365]  = ~\[2281]  | (~\[2286]  | ~\[2276] ),
  \[8331]  = ~v9 & (~v7 & ~v10),
  \[11986]  = v6 | ~v4,
  \[13646]  = ~\[2902]  | (~v11 | (~v8 | v7)),
  \[6675]  = ~v10 & (v8 & ~v7),
  \[10797]  = ~\[1322]  | (~\[1329]  | (~\[1315]  | ~\[1302] )),
  \[4288]  = v3 & (v1 & ~v0),
  \[9194]  = ~\[10509]  & (~v15 & v14),
  \[298]  = ~\[12510]  & (~v11 & (~\[12513]  & ~\[12509] )),
  \[2963]  = ~v12 & (v11 & v8),
  \[299]  = ~\[12520]  & (~v11 & (~\[12523]  & ~\[12519] )),
  \[3093]  = ~v6 & ~v5,
  \[14117]  = v11 | (~v10 | ~v9),
  \[13651]  = ~v6 | (~v5 | v4),
  \[12454]  = v11 | (~v10 | ~v9),
  \[634]  = ~\[443]  & (~\[442]  & (~\[441]  & ~\[440] )),
  \[10795]  = ~\[21709]  | (~\[21707]  | (~\[21711]  | ~\[1285] )),
  \[14114]  = v8 | (~v7 | ~v4),
  \[4625]  = ~\[12789]  & (v3 & (v1 & ~v0)),
  \[2237]  = ~v8 & (v7 & ~v5),
  \[7143]  = v12 & (v11 & ~v9),
  \[11600]  = ~\[6995]  | (~v3 | (~v1 | v0)),
  \[21519]  = ~v12 | (~v15 | ~\[9869] ),
  \[3430]  = ~\[13383]  & (~v12 & (v11 & ~v9)),
  \[11602]  = v13 | (~v11 | ~v8),
  \[5488]  = ~\[12329]  & (~v15 & (v14 & v12)),
  \[13657]  = ~\[2880]  | (~v11 | (~v8 | v7)),
  \[7877]  = ~v10 & (~v9 & ~v12),
  \[1776]  = ~\[14208]  & (~v14 & (v13 & ~v12)),
  \[11993]  = ~v3 | (~v1 | v0),
  \[11266]  = ~v2 | v1,
  \[11608]  = ~\[6982]  | (v6 | ~v4),
  \[21521]  = ~\[9861]  | (v15 | (~v14 | ~v13)),
  \[3438]  = ~v2 & (v1 & ~v0),
  \[4298]  = ~\[12948]  & (v15 & (v13 & ~v12)),
  \[5827]  = ~v12 & (v11 & ~v9),
  \[10079]  = ~\[21477]  | (~\[21475]  | (~\[21473]  | ~\[21471] )),
  \[2973]  = ~v6 & (~v5 & (~\[13610]  & ~v3)),
  \[641]  = ~\[439]  & (~\[438]  & (~\[437]  & ~\[436] )),
  \[14127]  = v11 | (~v10 | ~v9),
  \[13661]  = ~\[2874]  | (~v7 | v5),
  \[5493]  = ~v6 & (~v5 & ~v8),
  \[14124]  = v8 | (~v7 | ~v4),
  \[7153]  = ~\[11522]  & (v7 & (~v5 & ~v3)),
  \[12466]  = v11 | (~v10 | (~v9 | v8)),
  \[4636]  = ~\[12779]  & (v15 & (v13 & ~v12)),
  \[1781]  = ~v8 & (v7 & ~v5),
  \[11610]  = v13 | (~v11 | ~v8),
  \[22389]  = ~\[2004]  | ~\[2015] ,
  \[5100]  = ~v15 & (v14 & ~v13),
  \[5498]  = ~v2 & (v1 & ~v0),
  \[21523]  = ~\[9844]  | (v7 | (~v6 | ~v4)),
  \[7887]  = ~\[11158]  & (~v2 & (v1 & ~v0)),
  \[14132]  = ~\[22395]  | (~\[22393]  | (~\[22391]  | ~\[22389] )),
  \[21525]  = ~\[9841]  | (v10 | ~v9),
  \[8350]  = ~v10 & ~v9,
  \[1786]  = ~v2 & (v1 & ~v0),
  \[10416]  = ~\[21629]  | (~\[21627]  | (~\[21625]  | ~\[21623] )),
  \[13663]  = v12 | (~v11 | ~v8),
  \[11275]  = ~v0 | ~v2,
  \[12806]  = ~v3 | (~v1 | v0),
  \[3447]  = ~v12 & (v11 & ~v9),
  \[6695]  = ~v13 & (~v10 & v8),
  \[22391]  = ~\[1982]  | ~\[1993] ,
  \[2982]  = ~\[13605]  & (~v14 & (v13 & ~v12)),
  \[14138]  = ~v10 | ~v9,
  \[11619]  = ~v11 | ~v8,
  \[14137]  = ~\[1869]  | (v2 | (~v1 | v0)),
  \[13672]  = ~v11 | ~v8,
  \[12479]  = v11 | (~v10 | (~v9 | v8)),
  \[7162]  = ~\[11518]  & (~v15 & v14),
  \[16]  = ~\[10129]  & (~v12 & (~v2 & v0)),
  \[17]  = ~v14 & (v12 & (~v2 & v0)),
  \[18]  = ~\[10137]  & (~v10 & (v9 & ~v8)),
  \[4647]  = ~\[12776]  & (~v2 & (v1 & ~v0)),
  \[2259]  = ~v8 & (~v6 & v4),
  \[22001]  = ~\[5881]  | (~\[5891]  | (v14 | ~v13)),
  \[7895]  = ~v10 & (~v9 & ~v13),
  \[19]  = ~\[10141]  & (~v11 & (v10 & ~v9)),
  \[1063]  = ~\[11921]  & (~\[11895]  & (~\[11855]  & ~\[11820] )),
  \[12817]  = ~v11 | ~v8,
  \[22393]  = ~\[1960]  | ~\[1971] ,
  \[7501]  = ~v10 & (~v9 & ~v12),
  \[10426]  = ~v11 | (~v8 | ~v12),
  \[22395]  = ~\[1938]  | ~\[1949] ,
  \[14141]  = v14 | (~v13 | v12),
  \[11285]  = v6 | ~v4,
  \[1798]  = ~\[14198]  & (~v14 & (v13 & ~v12)),
  \[5845]  = ~v12 & (v11 & ~v9),
  \[3457]  = ~v6 & (~v5 & ~\[13370] ),
  \[2990]  = ~v3 & (v2 & ~v1),
  \[20]  = ~v14 & (~v13 & (~\[10146]  & ~v7)),
  \[11627]  = ~v11 | ~v8,
  \[21]  = ~\[10149]  & (v15 & (~v13 & ~v7)),
  \[13680]  = ~v11 | ~v8,
  \[11292]  = ~\[21817]  | (~\[21815]  | (~\[21813]  | ~\[21811] )),
  \[22]  = ~\[10154]  & (~v11 & (v10 & v8)),
  \[14148]  = ~\[1926]  | (v7 | (~v6 | ~v5)),
  \[1404]  = ~\[57]  & (~\[56]  & (~\[55]  & ~\[54] )),
  \[22003]  = ~\[5863]  | (~\[5873]  | (v14 | ~v13)),
  \[12822]  = ~\[22125]  | (~\[22123]  | (~\[22121]  | ~\[22119] )),
  \[23]  = ~\[10158]  & (v11 & (v9 & ~v8)),
  \[7170]  = ~v3 & (v2 & ~v1),
  \[12489]  = v11 | (~v10 | ~v9),
  \[6311]  = ~\[11948]  & (~v2 & (v1 & ~v0)),
  \[8368]  = ~v10 & ~v9,
  \[22005]  = ~\[5845]  | (~\[5855]  | (v14 | ~v13)),
  \[10095]  = ~\[21485]  | (~\[21483]  | (~\[21481]  | ~\[21479] )),
  \[4656]  = ~\[12769]  & (v15 & (v13 & ~v12)),
  \[28]  = ~\[10186]  & (~v9 & (v3 & ~v1)),
  \[21549]  = ~v15 | (v13 | (~v3 | ~v0)),
  \[29]  = ~v14 & (~v13 & (v3 & ~v1)),
  \[7176]  = ~v15 & (v14 & v12),
  \[8707]  = ~v10 & (v8 & ~v7),
  \[11294]  = ~v0 | ~v2,
  \[6319]  = ~v13 & (v11 & ~v9),
  \[14152]  = ~v13 | v12,
  \[1076]  = ~\[224]  & (~\[223]  & (~\[225]  & ~\[11753] )),
  \[2605]  = ~v12 & (~v10 & v8),
  \[7511]  = ~\[11351]  & (~v3 & (v2 & ~v1)),
  \[12824]  = ~v3 | (~v1 | v0),
  \[14151]  = v11 | (~v10 | (~v9 | v8)),
  \[3465]  = ~v12 & (v11 & ~v9),
  \[10435]  = ~v11 | (~v8 | ~v12),
  \[9569]  = ~v6 & (v5 & ~v4),
  \[22017]  = ~\[5737]  | (~\[5747]  | (v14 | ~v13)),
  \[5855]  = ~\[12172]  & (~v2 & (v1 & ~v0)),
  \[13686]  = ~v4 | ~v7,
  \[30]  = v15 & (~v13 & (v3 & ~v1)),
  \[21551]  = ~v3 | (~v0 | (~v8 | ~\[9742] )),
  \[12100]  = v12 | (~v11 | v9),
  \[22019]  = ~\[5719]  | (~\[5729]  | (v14 | ~v13)),
  \[31]  = ~\[10195]  & (~v11 & v10),
  \[10441]  = ~v6 | (~v5 | v4),
  \[32]  = ~\[10199]  & (~v8 & (v3 & ~v1)),
  \[14158]  = ~v5 | ~v6,
  \[22013]  = ~\[5773]  | (~\[5783]  | (v14 | ~v13)),
  \[12832]  = ~v3 | (~v1 | v0),
  \[33]  = v15 & (v12 & (v3 & ~v1)),
  \[14157]  = v4 | (~v3 | (~v1 | v0)),
  \[7180]  = ~v9 & ~v7,
  \[12499]  = ~\[5160]  | (v8 | (~v7 | ~v4)),
  \[34]  = ~\[10206]  & (~v12 & (v3 & ~v1)),
  \[672]  = ~\[13835]  & (~\[13807]  & (~\[13771]  & ~\[13736] )),
  \[12494]  = ~\[22065]  | (~\[22063]  | (~\[22061]  | ~\[22059] )),
  \[7519]  = ~v10 & (~v9 & ~v12),
  \[22015]  = ~\[5755]  | (~\[5765]  | (v14 | ~v13)),
  \[35]  = ~v14 & (v12 & (v3 & ~v1)),
  \[4664]  = v3 & (v1 & ~v0),
  \[2276]  = ~\[13958]  & (v15 & (v13 & ~v12)),
  \[3805]  = ~v10 & (~v9 & ~v12),
  \[36]  = ~\[10211]  & (~v10 & (v9 & ~v8)),
  \[11635]  = ~v11 | ~v8,
  \[37]  = ~\[10215]  & (~v11 & (v10 & ~v9)),
  \[38]  = ~v14 & (~v13 & (v3 & v0)),
  \[12108]  = ~v4 | (~v7 | ~\[5988] ),
  \[22021]  = ~\[5698]  | (~v11 | (~\[5694]  | ~\[5711] )),
  \[1083]  = ~\[218]  & (~\[217]  & (~\[216]  & ~\[215] )),
  \[10449]  = ~\[21637]  | (~\[21635]  | (~\[21633]  | ~\[21631] )),
  \[21553]  = ~v11 | (~v9 | ~\[9739] ),
  \[11641]  = ~\[21889]  | (~\[21887]  | (~\[21891]  | ~\[1105] )),
  \[10444]  = ~v11 | (~v8 | v7),
  \[6329]  = ~\[11938]  & (v3 & (v1 & ~v0)),
  \[21555]  = ~v12 | (~v15 | (~v3 | ~v0)),
  \[2615]  = ~v6 & (~v5 & (~\[13790]  & ~v3)),
  \[5863]  = ~v12 & (v11 & ~v9),
  \[3475]  = ~v6 & (~v5 & (~\[13360]  & ~v2)),
  \[13694]  = ~\[22309]  | (~\[22307]  | (~\[22311]  | ~\[686] )),
  \[9579]  = ~v6 & (v5 & ~v4),
  \[22027]  = ~\[5639]  | (~\[5649]  | (v14 | ~v13)),
  \[13696]  = ~\[723]  | (~\[730]  | (~\[716]  | ~\[703] )),
  \[1421]  = ~\[10285]  & (~\[10267]  & ~\[10317] ),
  \[2281]  = ~v8 & (~v6 & v4),
  \[12110]  = v13 | (~v11 | v9),
  \[11647]  = ~\[6905]  | (v3 | (~v2 | v1)),
  \[10452]  = ~v3 | (~v1 | v0),
  \[13308]  = ~v15 | ~v13,
  \[5138]  = ~v3 & (v2 & v0),
  \[22023]  = ~\[5676]  | (~v11 | (~\[5672]  | ~\[5689] )),
  \[11649]  = v13 | (~v11 | ~v8),
  \[43]  = ~\[10242]  & (~v15 & (v14 & v13)),
  \[8387]  = v12 & (~v10 & ~v9),
  \[44]  = ~v14 & (v12 & (v3 & v0)),
  \[7529]  = ~\[11341]  & (v7 & (~v5 & ~v3)),
  \[22025]  = ~\[5657]  | (~\[5667]  | (v14 | ~v13)),
  \[11643]  = ~\[1142]  | (~\[1149]  | (~\[1135]  | ~\[1122] )),
  \[45]  = ~\[10238]  & (~v10 & (v9 & ~v8)),
  \[4674]  = ~\[12760]  & (v15 & (v13 & ~v12)),
  \[2286]  = ~v2 & (v1 & ~v0),
  \[21567]  = ~\[9681]  | (~v15 | v13),
  \[1090]  = ~\[214]  & (~\[213]  & (~\[212]  & ~\[211] )),
  \[7193]  = ~\[11506]  & (~v3 & (v2 & v0)),
  \[10457]  = ~v11 | (~v8 | v7),
  \[686]  = ~\[417]  & (~\[416]  & (~\[415]  & ~\[414] )),
  \[14166]  = ~\[1887]  | (v14 | (~v13 | v12)),
  \[21569]  = ~\[9673]  | (v11 | (~v10 | ~v8)),
  \[3480]  = v15 & (v13 & ~v12),
  \[12118]  = v13 | (~v11 | v9),
  \[12848]  = ~\[22129]  | (~\[22127]  | ~\[22131] ),
  \[6337]  = ~v13 & (v11 & ~v9),
  \[10459]  = v15 | (~v14 | ~v12),
  \[21563]  = ~\[9699]  | (v11 | (~v10 | v9)),
  \[2623]  = ~v12 & (~v10 & v8),
  \[10454]  = ~v6 | (~v5 | v4),
  \[21565]  = ~\[9684]  | (v7 | (~v6 | v5)),
  \[3484]  = ~v9 & ~v7,
  \[13311]  = ~\[22229]  | (~\[22227]  | (~\[22225]  | ~\[22223] )),
  \[5873]  = ~v6 & (~v5 & ~\[12163] ),
  \[12843]  = ~v11 | ~v8,
  \[9589]  = ~v6 & (v5 & ~v4),
  \[12116]  = ~v4 | (~v7 | ~\[5970] ),
  \[22037]  = ~\[5543]  | (~\[5550]  | ~\[5538] ),
  \[21571]  = ~\[9663]  | (~v11 | (~v9 | v8)),
  \[21909]  = ~\[6749]  | (~\[6759]  | (v15 | ~v14)),
  \[22039]  = ~\[5517]  | (~\[5524]  | ~\[5512] ),
  \[11657]  = v13 | (~v11 | ~v8),
  \[13318]  = ~v15 | ~v13,
  \[1434]  = ~\[44]  & (~\[43]  & (~\[45]  & ~\[10235] )),
  \[7537]  = ~v10 & (~v9 & ~v12),
  \[14177]  = v11 | (~v10 | ~v9),
  \[4682]  = ~v2 & (v1 & ~v0),
  \[8397]  = ~v6 & (~v5 & (~\[10900]  & ~v3)),
  \[3823]  = ~v10 & (~v9 & ~v12),
  \[12851]  = ~\[902]  | (~\[909]  | (~\[895]  | ~\[882] )),
  \[54]  = ~\[10288]  & (~v10 & (v9 & ~v8)),
  \[55]  = ~\[10292]  & (~v11 & (v10 & ~v9)),
  \[8731]  = ~v6 & v4,
  \[56]  = ~v14 & (~v13 & (~\[10296]  & ~v6)),
  \[21577]  = ~\[9633]  | (v14 | ~v12),
  \[11655]  = ~\[6887]  | (v3 | (~v2 | ~v0)),
  \[57]  = ~\[10299]  & (v15 & (~v13 & ~v6)),
  \[2298]  = ~\[13948]  & (v15 & (v13 & ~v12)),
  \[21911]  = ~v4 | (~v7 | (~\[6740]  | ~\[6732] )),
  \[22041]  = ~\[5493]  | (~\[5498]  | ~\[5488] ),
  \[12127]  = v12 | (~v11 | v9),
  \[6347]  = ~\[11930]  & (~v2 & (v1 & ~v0)),
  \[300]  = ~\[12500]  & (~v11 & (~\[12503]  & ~\[12499] )),
  \[21573]  = ~v12 | (~v15 | ~\[9653] ),
  \[2633]  = ~\[13782]  & (v7 & ~v5),
  \[301]  = ~\[12536]  & (~v11 & (~\[12539]  & ~\[12535] )),
  \[10464]  = ~\[9269]  | (v2 | (~v1 | v0)),
  \[5881]  = ~v12 & (v11 & ~v9),
  \[12859]  = ~v15 | (~v13 | ~\[4485] ),
  \[302]  = ~\[12543]  & (~v8 & (~\[12542]  & ~\[12550] )),
  \[21575]  = ~\[9645]  | (v15 | (~v14 | ~v13)),
  \[303]  = ~\[12561]  & (~v15 & (~\[12560]  & ~\[12557] )),
  \[10466]  = ~v11 | (~v8 | ~v12),
  \[12853]  = v3 | (~v2 | v1),
  \[304]  = ~\[12567]  & (~v7 & (~\[12566]  & ~\[12575] )),
  \[305]  = ~\[12583]  & (~v11 & (~\[12586]  & ~\[12582] )),
  \[9202]  = ~v2 & (v1 & ~v0),
  \[3497]  = ~\[13353]  & (v3 & (v1 & ~v0)),
  \[12125]  = ~v4 | (~v7 | (~\[5951]  | ~v3)),
  \[1441]  = ~\[38]  & (~\[37]  & (~\[36]  & ~\[35] )),
  \[306]  = ~\[12593]  & (~v11 & (~\[12596]  & ~\[12592] )),
  \[12130]  = ~v1 | v0,
  \[307]  = ~\[12604]  & (~v11 & (~\[12607]  & ~\[12603] )),
  \[61]  = ~\[10323]  & (~v15 & (v14 & v13)),
  \[308]  = ~\[12614]  & (~v11 & (~\[12617]  & ~\[12613] )),
  \[62]  = ~\[10326]  & (~v14 & (v12 & ~v6)),
  \[10809]  = ~v3 | (~v1 | v0),
  \[21913]  = ~v4 | (~v7 | (~\[6722]  | ~\[6714] )),
  \[7547]  = ~\[11325]  & (~v3 & (v2 & ~v1)),
  \[63]  = ~\[10331]  & (~v10 & (v9 & ~v8)),
  \[14187]  = v11 | (~v10 | ~v9),
  \[12861]  = v3 | (~v2 | ~v0),
  \[11664]  = ~\[6874]  | (v6 | ~v4),
  \[64]  = ~\[10335]  & (~v11 & (v10 & ~v9)),
  \[3104]  = ~v14 & (v13 & ~v12),
  \[10803]  = ~v4 | (~v7 | ~\[8602] ),
  \[21915]  = ~\[6695]  | (~\[6705]  | (v15 | ~v14)),
  \[65]  = ~v14 & (~v13 & ~\[10341] ),
  \[4694]  = ~\[12752]  & (~v15 & (v14 & ~v13)),
  \[8011]  = ~v10 & (~v9 & ~v13),
  \[11666]  = v13 | (~v11 | ~v8),
  \[66]  = ~\[10344]  & (v15 & ~v13),
  \[10805]  = ~v12 | (v10 | ~v8),
  \[21587]  = ~\[9589]  | (v11 | (~v10 | ~v8)),
  \[1448]  = ~\[34]  & (~\[33]  & (~\[32]  & ~\[31] )),
  \[67]  = ~\[10348]  & (~v11 & (v10 & v8)),
  \[13326]  = ~v15 | ~v13,
  \[6355]  = ~v13 & (~v10 & v8),
  \[68]  = ~\[10352]  & (v11 & (v9 & ~v8)),
  \[21589]  = ~\[9579]  | (~v11 | (~v9 | v8)),
  \[2641]  = ~v12 & (~v10 & v8),
  \[5160]  = ~v3 & (v2 & ~v1),
  \[12867]  = ~v15 | (~v13 | ~\[4467] ),
  \[11672]  = ~\[6851]  | (v3 | (~v2 | ~v0)),
  \[8746]  = ~\[10724]  & (~v15 & v14),
  \[5891]  = ~v6 & (~v5 & (~\[12153]  & ~v2)),
  \[12139]  = ~\[5923]  | (v14 | (~v13 | v12)),
  \[10473]  = ~\[9251]  | (~v3 | (~v1 | v0)),
  \[313]  = ~\[12682]  & (~v11 & (~\[12685]  & ~\[12681] )),
  \[12133]  = ~v6 | (~v5 | v4),
  \[7552]  = ~v14 & (v13 & ~v12),
  \[314]  = ~\[12692]  & (~v11 & (~\[12695]  & ~\[12691] )),
  \[10475]  = ~v11 | (~v8 | ~v12),
  \[21927]  = ~\[6579]  | (~\[6589]  | (v15 | ~v14)),
  \[315]  = ~\[12674]  & (~v15 & (~\[12673]  & ~\[12670] )),
  \[4306]  = ~v3 & (v2 & v0),
  \[9212]  = ~\[10501]  & (~v15 & v14),
  \[10817]  = ~v1 | v0,
  \[5896]  = ~v14 & (v13 & ~v12),
  \[21591]  = ~v12 | (~v15 | ~\[9569] ),
  \[21929]  = ~\[6561]  | (~\[6571]  | (v15 | ~v14)),
  \[22059]  = ~\[5290]  | ~\[5301] ,
  \[3841]  = ~v10 & (~v9 & ~v12),
  \[10481]  = ~\[9238]  | (v6 | ~v4),
  \[14198]  = v11 | (~v10 | ~v9),
  \[21923]  = ~\[6615]  | (~\[6625]  | (v15 | ~v14)),
  \[7557]  = ~v9 & (~v7 & ~v10),
  \[12872]  = ~\[4458]  | (v6 | ~v4),
  \[73]  = ~\[10383]  & (~v11 & (v10 & ~v9)),
  \[11674]  = v13 | (~v11 | ~v8),
  \[74]  = ~v13 & (~v3 & (~v14 & ~\[10387] )),
  \[21925]  = ~\[6597]  | (~\[6607]  | (v15 | ~v14)),
  \[75]  = ~\[10378]  & (v15 & (~v13 & ~v3)),
  \[10815]  = ~\[8574]  | (v15 | (~v14 | ~v12)),
  \[10820]  = ~v6 | (~v5 | v4),
  \[6365]  = ~\[11898]  & (~v3 & (v2 & v0)),
  \[13335]  = ~v15 | ~v13,
  \[21931]  = ~\[6543]  | (~\[6553]  | (v15 | ~v14)),
  \[2651]  = ~\[13775]  & (~v2 & (v1 & ~v0)),
  \[8754]  = ~v3 & (v2 & ~v1),
  \[22061]  = ~\[5271]  | (~\[5278]  | ~\[5266] ),
  \[12878]  = v3 | (~v2 | ~v0),
  \[13340]  = ~v6 | (~v5 | v4),
  \[10483]  = ~v11 | (~v8 | ~v12),
  \[12874]  = v12 | (~v11 | ~v8),
  \[9220]  = v3 & (v1 & ~v0),
  \[8029]  = ~v10 & (~v9 & ~v13),
  \[21937]  = ~\[6489]  | (~\[6499]  | (v15 | ~v14)),
  \[12146]  = ~v6 | (~v5 | v4),
  \[4316]  = ~\[12939]  & (v15 & (v13 & ~v12)),
  \[10828]  = ~v3 | (~v1 | v0),
  \[11688]  = ~\[6822]  | (~v11 | (~v8 | v7)),
  \[6705]  = ~\[11746]  & (v3 & (v1 & ~v0)),
  \[21939]  = ~\[6471]  | (~\[6481]  | (v15 | ~v14)),
  \[2659]  = ~v12 & (~v10 & v8),
  \[13348]  = ~\[22237]  | (~\[22235]  | (~\[22233]  | ~\[22231] )),
  \[21933]  = ~\[6525]  | (~\[6535]  | (v15 | ~v14)),
  \[9955]  = ~v8 & (~v2 & v0),
  \[1464]  = ~\[29]  & (~\[28]  & (~\[30]  & ~\[10181] )),
  \[22063]  = ~\[5245]  | (~\[5252]  | ~\[5240] ),
  \[11689]  = ~v0 | ~v2,
  \[5512]  = ~\[12353]  & (~v15 & (v14 & v12)),
  \[84]  = ~\[10459]  & (~\[10457]  & (~\[10454]  & ~\[10452] )),
  \[21935]  = ~\[6507]  | (~\[6517]  | (v15 | ~v14)),
  \[7569]  = ~\[11316]  & (~v3 & (v2 & v0)),
  \[22065]  = ~\[5221]  | (~\[5226]  | ~\[5216] ),
  \[11683]  = ~\[6838]  | (~v6 | (~v5 | v4)),
  \[85]  = ~\[10466]  & (~\[10464]  & (~v15 & v14)),
  \[10826]  = ~\[8555]  | (v15 | (~v14 | ~v12)),
  \[9958]  = ~v11 & v10,
  \[6373]  = ~v13 & (~v10 & v8),
  \[86]  = ~\[10475]  & (~\[10473]  & (~v15 & v14)),
  \[3126]  = ~v14 & (v13 & ~v12),
  \[22407]  = ~\[1807]  | (~v3 | (~\[1803]  | ~\[1798] )),
  \[87]  = ~\[10483]  & (~\[10481]  & (~v15 & v14)),
  \[10830]  = ~v6 | (~v5 | v4),
  \[8763]  = v12 & (~v10 & v8),
  \[21941]  = ~\[6446]  | (~\[6451]  | ~\[6463] ),
  \[22409]  = ~\[1781]  | (~\[1786]  | ~\[1776] ),
  \[5517]  = ~v7 & (v6 & v5),
  \[1803]  = ~v8 & (~v6 & v4),
  \[11692]  = ~v6 | (~v5 | v4),
  \[331]  = ~v6 & (~v5 & (~\[12853]  & ~\[12859] )),
  \[22403]  = ~\[1851]  | (~v3 | (~\[1847]  | ~\[1842] )),
  \[5182]  = ~v2 & (v1 & ~v0),
  \[332]  = ~v6 & (~v5 & (~\[12861]  & ~\[12867] )),
  \[10493]  = ~v11 | (~v8 | ~v12),
  \[12884]  = ~v15 | (~v13 | ~\[4431] ),
  \[333]  = ~\[12874]  & (~\[12872]  & (v15 & v13)),
  \[22405]  = ~\[1825]  | (~\[1830]  | ~\[1820] ),
  \[4324]  = ~v3 & (v2 & ~v1),
  \[12153]  = ~v1 | v0,
  \[1807]  = v1 & ~v0,
  \[334]  = ~\[12878]  & (~\[12884]  & (~v6 & v4)),
  \[21947]  = ~\[6391]  | (~\[6401]  | (v15 | ~v14)),
  \[335]  = ~\[12895]  & (~\[12893]  & ~\[12891] ),
  \[6714]  = ~\[11740]  & (~v15 & (v14 & ~v13)),
  \[1471]  = ~\[23]  & (~\[22]  & (~\[21]  & ~\[20] )),
  \[7574]  = ~v14 & (v13 & ~v12),
  \[11698]  = ~\[6800]  | (~v11 | (~v8 | v7)),
  \[336]  = ~\[12905]  & (~\[12903]  & (~\[12900]  & ~\[12898] )),
  \[21949]  = ~\[6373]  | (~\[6383]  | (v15 | ~v14)),
  \[2669]  = ~\[13763]  & (~v6 & v4),
  \[337]  = ~\[12913]  & (~\[12911]  & (v15 & v13)),
  \[22411]  = ~\[1763]  | (~v3 | (~\[1759]  | ~\[1754] )),
  \[91]  = ~\[10522]  & (~\[10520]  & (~v15 & v14)),
  \[3861]  = ~v9 & (~v7 & ~v10),
  \[338]  = ~\[12917]  & (~\[12923]  & (v7 & ~v5)),
  \[92]  = ~\[10530]  & (~\[10528]  & (~v15 & v14)),
  \[21943]  = ~\[6424]  | (~\[6429]  | ~\[6441] ),
  \[93]  = ~\[10539]  & (~\[10537]  & (~v15 & v14)),
  \[12891]  = ~\[4422]  | (~v6 | (~v5 | v4)),
  \[94]  = ~\[10547]  & (~\[10545]  & (~v15 & v14)),
  \[21945]  = ~\[6409]  | (~\[6419]  | (v15 | ~v14)),
  \[7579]  = ~v9 & (~v7 & ~v10),
  \[95]  = ~\[10559]  & (~v15 & (~\[10558]  & ~\[10556] )),
  \[10836]  = ~\[8533]  | (v15 | (~v14 | ~v12)),
  \[9238]  = ~v2 & (v1 & ~v0),
  \[6383]  = ~\[11914]  & (~v3 & (v2 & ~v1)),
  \[5524]  = ~v4 & (v3 & (v1 & ~v0)),
  \[96]  = ~\[10570]  & (~\[10568]  & (~\[10565]  & ~\[10563] )),
  \[13353]  = ~v6 | (~v5 | v4),
  \[1478]  = ~\[19]  & (~\[18]  & (~\[17]  & ~\[16] )),
  \[10110]  = ~\[21493]  | (~\[21491]  | (~\[21489]  | ~\[21487] )),
  \[7913]  = ~v10 & (~v9 & ~v13),
  \[22417]  = ~\[1693]  | (~\[1698]  | ~\[1688] ),
  \[97]  = ~\[10578]  & (~\[10576]  & (~v15 & v14)),
  \[10840]  = v2 | (~v1 | v0),
  \[8773]  = ~v6 & (~v5 & (~\[10711]  & ~v3)),
  \[98]  = ~\[10586]  & (~\[10584]  & (~v15 & v14)),
  \[21951]  = ~\[6355]  | (~\[6365]  | (v15 | ~v14)),
  \[12500]  = ~v10 | ~v9,
  \[12898]  = v3 | (~v2 | ~v0),
  \[13360]  = ~v1 | v0,
  \[22413]  = ~\[1737]  | (~\[1742]  | ~\[1732] ),
  \[8047]  = ~v10 & (~v9 & ~v13),
  \[343]  = ~\[12970]  & (~v2 & (~\[12973]  & ~\[12979] )),
  \[6722]  = ~v3 & (v2 & v0),
  \[22415]  = ~\[1710]  | ~\[1721] ,
  \[4334]  = ~\[12933]  & (~v12 & (~v10 & v8)),
  \[12163]  = ~v3 | (~v1 | v0),
  \[12893]  = ~v11 | (~v8 | v7),
  \[344]  = ~\[12983]  & (~\[12981]  & ~\[12989] ),
  \[21957]  = ~\[6298]  | (~v11 | (~\[6294]  | ~\[6311] )),
  \[2677]  = ~v12 & (~v10 & v8),
  \[11305]  = ~v6 | (~v5 | v4),
  \[345]  = ~v6 & (~v5 & (~\[12963]  & ~\[12969] )),
  \[10848]  = ~v3 | (~v1 | v0),
  \[12895]  = ~v15 | (~v13 | v12),
  \[21959]  = ~\[6276]  | (~v11 | (~\[6272]  | ~\[6289] )),
  \[22089]  = ~\[4949]  | (~\[4954]  | ~\[4944] ),
  \[3142]  = ~v2 & (v1 & ~v0),
  \[21953]  = ~\[6337]  | (~\[6347]  | (v15 | ~v14)),
  \[12172]  = v6 | ~v4,
  \[5199]  = ~v8 & (v7 & ~v5),
  \[13702]  = ~v11 | ~v8,
  \[12509]  = ~\[5199]  | (v3 | (~v2 | ~v0)),
  \[6391]  = ~v13 & (~v10 & v8),
  \[21955]  = ~\[6319]  | (~\[6329]  | (v15 | ~v14)),
  \[10846]  = ~\[8512]  | (v15 | (~v14 | ~v12)),
  \[8781]  = v12 & (~v10 & v8),
  \[12503]  = v15 | (~v14 | ~v12),
  \[1820]  = ~\[14187]  & (~v14 & (v13 & ~v12)),
  \[22427]  = ~\[1570]  | ~\[1581] ,
  \[21961]  = ~\[6257]  | (~\[6267]  | (v15 | ~v14)),
  \[12510]  = ~v10 | ~v9,
  \[22091]  = ~\[4931]  | (~v3 | (~\[4927]  | ~\[4922] )),
  \[22429]  = ~\[1548]  | ~\[1559] ,
  \[13370]  = ~v3 | (~v1 | v0),
  \[13708]  = ~v4 | ~v7,
  \[5538]  = ~\[12341]  & (~v15 & (v14 & v12)),
  \[4342]  = ~v2 & (v1 & ~v0),
  \[8057]  = ~\[11053]  & (v7 & ~v5),
  \[12179]  = ~\[22005]  | (~\[22003]  | (~\[22001]  | ~\[21999] )),
  \[1825]  = ~v8 & (~v6 & v4),
  \[7591]  = ~\[11305]  & (~v3 & (v2 & ~v1)),
  \[6732]  = ~\[11731]  & (~v15 & (v14 & ~v13)),
  \[11316]  = ~v6 | (~v5 | v4),
  \[9251]  = ~v6 & ~v5,
  \[21967]  = ~\[6203]  | (~\[6213]  | (v15 | ~v14)),
  \[2687]  = ~\[13756]  & (~v2 & (v1 & ~v0)),
  \[10857]  = v2 | (~v1 | v0),
  \[21969]  = ~\[6185]  | (~\[6195]  | (v15 | ~v14)),
  \[6006]  = ~v2 & (v1 & ~v0),
  \[9983]  = ~v9 & (~v2 & v0),
  \[22431]  = ~\[1526]  | ~\[1537] ,
  \[10129]  = v15 | (~v14 | ~v13),
  \[3152]  = ~\[13520]  & (~v14 & (v13 & ~v12)),
  \[21963]  = ~\[6239]  | (~\[6249]  | (v15 | ~v14)),
  \[22093]  = ~\[4905]  | (~\[4910]  | ~\[4900] ),
  \[10854]  = ~\[8494]  | (v15 | (~v14 | ~v12)),
  \[12181]  = ~v3 | (~v1 | v0),
  \[3883]  = ~v9 & (~v7 & ~v10),
  \[12519]  = ~\[5182]  | (v8 | (~v7 | ~v4)),
  \[10123]  = ~\[21501]  | (~\[21499]  | (~\[21497]  | ~\[21495] )),
  \[21965]  = ~\[6221]  | (~\[6231]  | (v15 | ~v14)),
  \[7599]  = ~v10 & (~v9 & ~v12),
  \[22095]  = ~\[4878]  | ~\[4889] ,
  \[5543]  = ~v7 & (v6 & v5),
  \[8791]  = ~v6 & (~v5 & (~\[10702]  & ~v3)),
  \[12513]  = v15 | (~v14 | ~v12),
  \[7203]  = v11 & (~v9 & ~v7),
  \[1830]  = ~v2 & (v1 & ~v0),
  \[7933]  = ~v9 & (~v7 & ~v10),
  \[21971]  = ~\[6167]  | (~\[6177]  | (v15 | ~v14)),
  \[12520]  = ~v10 | ~v9,
  \[8065]  = ~v10 & (~v9 & ~v13),
  \[12187]  = ~\[5791]  | (v14 | ~v13),
  \[13718]  = ~v6 | (~v5 | v4),
  \[4351]  = ~v12 & (v11 & v8),
  \[361]  = ~\[13136]  & (~\[13142]  & (v7 & v4)),
  \[6740]  = ~v3 & (v2 & ~v1),
  \[1105]  = ~\[207]  & (~\[206]  & (~\[205]  & ~\[204] )),
  \[12189]  = ~v3 | (~v1 | v0),
  \[362]  = ~\[13144]  & (~\[13150]  & (v7 & v4)),
  \[2695]  = ~v12 & (~v10 & v8),
  \[363]  = ~\[13152]  & (~v2 & (~\[13155]  & ~\[13161] )),
  \[364]  = ~\[13165]  & (~\[13163]  & ~\[13171] ),
  \[21977]  = ~\[6113]  | (~\[6123]  | (v15 | ~v14)),
  \[9991]  = ~v8 & (~v2 & v0),
  \[11325]  = ~v7 | v5,
  \[365]  = ~v6 & (~v5 & (~\[13175]  & ~\[13181] )),
  \[6015]  = ~v13 & (v11 & ~v9),
  \[10137]  = v7 | (~v6 | ~v4),
  \[366]  = ~v6 & (~v5 & (~\[13183]  & ~\[13189] )),
  \[3160]  = v3 & (v1 & ~v0),
  \[21979]  = ~\[6095]  | (~\[6105]  | (v15 | ~v14)),
  \[367]  = ~\[13192]  & (~\[13198]  & (~v6 & v4)),
  \[13388]  = ~v3 | (~v1 | v0),
  \[8405]  = v12 & (~v10 & ~v9),
  \[11332]  = ~\[21825]  | (~\[21823]  | (~\[21821]  | ~\[21819] )),
  \[368]  = ~\[13200]  & (~\[13206]  & (~v6 & v4)),
  \[5550]  = ~v4 & (~v2 & (v1 & ~v0)),
  \[2303]  = ~v6 & (~v5 & ~v8),
  \[21973]  = ~\[6149]  | (~\[6159]  | (v15 | ~v14)),
  \[12529]  = ~\[933]  | (~\[940]  | (~\[926]  | ~\[971] )),
  \[6749]  = ~v13 & (~v10 & v8),
  \[10863]  = ~\[8476]  | (v15 | (~v14 | ~v12)),
  \[21975]  = ~\[6131]  | (~\[6141]  | (v15 | ~v14)),
  \[703]  = ~\[13627]  & (~\[13592]  & ~\[13694] ),
  \[12523]  = v15 | (~v14 | v13),
  \[10865]  = ~v3 | (~v1 | v0),
  \[9269]  = ~v6 & ~v5,
  \[2307]  = v1 & ~v0,
  \[13383]  = ~v15 | ~v13,
  \[13386]  = ~\[22245]  | (~\[22243]  | (~\[22241]  | ~\[22239] )),
  \[21981]  = ~\[6074]  | (~v11 | (~\[6070]  | ~\[6087] )),
  \[1842]  = ~\[14177]  & (~v14 & (v13 & ~v12)),
  \[8075]  = ~\[11070]  & (~v2 & (v1 & ~v0)),
  \[12197]  = v2 | (~v1 | v0),
  \[13728]  = ~v6 | (~v5 | v4),
  \[10141]  = v7 | (~v6 | ~v4),
  \[10871]  = ~\[8458]  | (v15 | (~v14 | ~v12)),
  \[3502]  = v15 & (v13 & ~v12),
  \[373]  = ~\[13256]  & (~\[13262]  & (~v6 & v4)),
  \[1847]  = ~v6 & (~v5 & ~v8),
  \[374]  = ~\[13264]  & (~\[13270]  & (~v6 & v4)),
  \[3506]  = ~v9 & ~v7,
  \[11335]  = ~v4 | ~v7,
  \[375]  = ~\[13245]  & (~v3 & (~\[13248]  & ~\[13254] )),
  \[12195]  = ~\[5827]  | (v14 | ~v13),
  \[3170]  = ~\[13512]  & (~v14 & (v13 & ~v12)),
  \[10877]  = ~v7 | v5,
  \[8415]  = ~v6 & (~v5 & (~\[10892]  & ~v3)),
  \[10149]  = ~v6 | ~v4,
  \[11341]  = ~v0 | ~v2,
  \[12539]  = v15 | (~v14 | ~v12),
  \[6759]  = ~\[11721]  & (~v2 & (v1 & ~v0)),
  \[10146]  = ~v6 | ~v4,
  \[4705]  = ~\[12749]  & (~v3 & (v2 & v0)),
  \[12536]  = ~v10 | ~v9,
  \[8083]  = ~v10 & (~v9 & ~v13),
  \[13396]  = ~v3 | (~v1 | v0),
  \[12535]  = ~\[5138]  | (v8 | (~v7 | ~v4)),
  \[1851]  = v1 & ~v0,
  \[716]  = ~\[404]  & (~\[403]  & (~\[405]  & ~\[13525] )),
  \[3178]  = ~v2 & (v1 & ~v0),
  \[1122]  = ~\[11576]  & (~\[11539]  & ~\[11641] ),
  \[7955]  = ~v9 & (~v7 & ~v10),
  \[13008]  = ~v15 | ~v13,
  \[5900]  = ~v9 & ~v7,
  \[7227]  = ~v6 & v4,
  \[13737]  = ~v1 | v0,
  \[12542]  = ~v3 | (~v1 | v0),
  \[6033]  = ~v13 & (v11 & ~v9),
  \[10158]  = v7 | (~v6 | ~v4),
  \[2320]  = ~\[13937]  & (v15 & (v13 & ~v12)),
  \[8423]  = v12 & (~v10 & ~v9),
  \[13736]  = ~\[22319]  | (~\[22317]  | (~\[22315]  | ~\[22313] )),
  \[21999]  = ~\[5900]  | (~v11 | (~\[5896]  | ~\[5913] )),
  \[4378]  = ~v3 & (v2 & ~v1),
  \[3519]  = ~\[13340]  & (~v2 & (v1 & ~v0)),
  \[14208]  = v11 | (~v10 | ~v9),
  \[11351]  = ~v4 | ~v7,
  \[10154]  = v7 | (~v6 | ~v4),
  \[10884]  = ~v3 | (~v1 | v0),
  \[13012]  = ~v3 | (~v1 | v0),
  \[5572]  = v3 & (v1 & ~v0),
  \[2325]  = ~v6 & (~v5 & ~v8),
  \[723]  = ~\[398]  & (~\[397]  & (~\[396]  & ~\[395] )),
  \[12543]  = ~v4 | ~v7,
  \[4716]  = ~\[12740]  & (~v15 & (v14 & ~v13)),
  \[8093]  = ~\[11061]  & (~v6 & v4),
  \[11358]  = ~\[21829]  | (~\[21827]  | ~\[21831] ),
  \[3188]  = ~\[13505]  & (~v12 & (v11 & ~v9)),
  \[21609]  = ~v12 | (~v15 | (~\[9484]  | ~v7)),
  \[12550]  = ~\[5100]  | (v11 | (~v10 | ~v9)),
  \[10892]  = ~v2 | v1,
  \[391]  = ~v6 & (~v5 & (~\[13417]  & ~\[13423] )),
  \[1135]  = ~\[194]  & (~\[193]  & (~\[195]  & ~\[11472] )),
  \[392]  = ~v6 & (~v5 & (~\[13425]  & ~\[13431] )),
  \[6771]  = v7 & ~v5,
  \[393]  = ~\[13434]  & (~\[13440]  & (~v6 & v4)),
  \[5913]  = ~\[12146]  & (v3 & (v1 & ~v0)),
  \[394]  = ~\[13442]  & (~\[13448]  & (~v6 & v4)),
  \[395]  = ~\[13451]  & (~v3 & (~\[13454]  & ~\[13460] )),
  \[2330]  = ~v2 & (v1 & ~v0),
  \[8433]  = ~\[10884]  & (v7 & ~v5),
  \[13746]  = ~v3 | (~v1 | v0),
  \[1869]  = ~v6 & (~v5 & ~v8),
  \[396]  = ~\[13461]  & (~v3 & (~\[13464]  & ~\[13470] )),
  \[21611]  = ~\[9477]  | (v15 | (~v14 | ~v13)),
  \[3528]  = ~\[13335]  & (~v12 & (v11 & ~v9)),
  \[397]  = ~\[13473]  & (~\[13479]  & (v7 & ~v5)),
  \[12557]  = ~\[5094]  | (v7 | (~v6 | ~v5)),
  \[398]  = ~\[13481]  & (~\[13487]  & (v7 & ~v5)),
  \[10501]  = ~v11 | (~v8 | ~v12),
  \[730]  = ~\[394]  & (~\[393]  & (~\[392]  & ~\[391] )),
  \[11361]  = ~\[1202]  | (~\[1209]  | (~\[1195]  | ~\[1182] )),
  \[2335]  = v13 & ~v12,
  \[3196]  = ~v3 & (v2 & v0),
  \[14213]  = ~\[22409]  | (~\[22407]  | (~\[22405]  | ~\[22403] )),
  \[11368]  = ~v12 | (~v11 | v9),
  \[4727]  = ~\[12737]  & (~v3 & (v2 & ~v1)),
  \[9633]  = ~v7 & (v6 & ~v5),
  \[1142]  = ~\[188]  & (~\[187]  & (~\[186]  & ~\[185] )),
  \[12560]  = v11 | (~v10 | (~v9 | v8)),
  \[7975]  = ~v10 & (~v9 & ~v13),
  \[13028]  = ~\[22169]  | (~\[22167]  | (~\[22165]  | ~\[22163] )),
  \[10509]  = ~v11 | (~v8 | ~v12),
  \[14220]  = v11 | (~v10 | ~v9),
  \[21613]  = ~\[9464]  | (v14 | (~v12 | ~v7)),
  \[12561]  = ~v14 | v13,
  \[21615]  = ~\[9457]  | (v10 | (~v9 | v8)),
  \[5923]  = v11 & (~v9 & ~v7),
  \[8441]  = v12 & (~v10 & ~v9),
  \[6053]  = v11 & (~v9 & ~v7),
  \[11366]  = ~v4 | (~v7 | ~\[7474] ),
  \[3536]  = v3 & (v1 & ~v0),
  \[1149]  = ~\[184]  & (~\[183]  & (~\[182]  & ~\[181] )),
  \[13756]  = v6 | ~v4,
  \[13025]  = ~v15 | ~v13,
  \[12900]  = ~v6 | (~v5 | v4),
  \[13030]  = ~v3 | (~v1 | v0),
  \[12567]  = ~v5 | ~v6,
  \[2343]  = ~v11 & (v10 & (v9 & ~v8)),
  \[4002]  = ~v3 & (v2 & ~v1),
  \[7250]  = ~v3 & (v2 & ~v1),
  \[11703]  = ~\[6794]  | (~v7 | v5),
  \[5594]  = ~v2 & (v1 & ~v0),
  \[21627]  = ~\[9389]  | (~v15 | (~v12 | v3)),
  \[12566]  = v4 | (~v3 | (~v1 | v0)),
  \[11705]  = v13 | (~v11 | ~v8),
  \[4007]  = v13 & ~v12,
  \[21629]  = ~\[9372]  | ~\[9379] ,
  \[4738]  = ~\[12730]  & (~v15 & (v14 & ~v13)),
  \[10181]  = ~\[21525]  | (~\[21523]  | (~\[21521]  | ~\[21519] )),
  \[14230]  = v11 | (~v10 | ~v9),
  \[13037]  = ~v2 | v1,
  \[21623]  = ~\[9413]  | (v11 | (~v10 | ~v8)),
  \[9645]  = ~v12 & (~v7 & (v6 & ~v5)),
  \[11711]  = ~\[6771]  | (v3 | (~v2 | ~v0)),
  \[10514]  = ~\[21649]  | (~\[21647]  | (~\[21651]  | ~\[1344] )),
  \[11374]  = ~v4 | (~v7 | (~\[7455]  | ~v3)),
  \[21625]  = ~\[9401]  | (~v11 | (~v9 | v8)),
  \[7259]  = v12 & (v11 & ~v9),
  \[10516]  = ~\[1381]  | (~\[1388]  | (~\[1374]  | ~\[1361] )),
  \[8451]  = ~\[10877]  & (~v2 & (v1 & ~v0)),
  \[11376]  = ~v12 | (~v11 | v9),
  \[1887]  = ~v11 & (v10 & (v9 & ~v8)),
  \[12903]  = ~v11 | (~v8 | v7),
  \[3546]  = ~\[13326]  & (~v12 & (v11 & ~v9)),
  \[13763]  = ~v3 | (~v1 | v0),
  \[6794]  = ~v3 & (v2 & ~v1),
  \[10520]  = ~\[9161]  | (v3 | (~v2 | v1)),
  \[11380]  = ~v1 | v0,
  \[12905]  = ~v15 | (~v13 | v12),
  \[21631]  = ~\[9360]  | (~v2 | (~v1 | v0)),
  \[10522]  = ~v11 | (~v8 | ~v12),
  \[6401]  = ~\[11904]  & (v7 & (~v5 & ~v3)),
  \[12911]  = ~\[4378]  | (~v7 | v5),
  \[4013]  = ~v10 & (v8 & ~v7),
  \[8458]  = ~v10 & ~v9,
  \[13771]  = ~\[22327]  | (~\[22325]  | (~\[22323]  | ~\[22321] )),
  \[10186]  = v11 | ~v10,
  \[11713]  = v13 | (~v11 | ~v8),
  \[21637]  = ~\[9308]  | ~\[9319] ,
  \[2357]  = ~\[13921]  & (~v7 & (v6 & v5)),
  \[7993]  = ~v10 & (~v9 & ~v13),
  \[10528]  = ~\[9143]  | (v3 | (~v2 | ~v0)),
  \[12575]  = ~\[5055]  | (v15 | (~v14 | v13)),
  \[14236]  = v3 | (~v2 | ~v0),
  \[9653]  = ~v7 & (v6 & ~v5),
  \[12917]  = v3 | (~v2 | ~v0),
  \[21633]  = ~v4 | (~v7 | (~\[9354]  | ~\[9346] )),
  \[4749]  = ~\[12725]  & (~v8 & (v7 & ~v5)),
  \[6070]  = ~v15 & (v14 & ~v13),
  \[12582]  = ~\[5037]  | (v2 | (~v1 | v0)),
  \[11389]  = ~\[7427]  | (v15 | (~v14 | ~v12)),
  \[11721]  = ~v4 | ~v7,
  \[6409]  = ~v13 & (~v10 & v8),
  \[21635]  = ~v4 | (~v7 | (~\[9336]  | ~\[9328] )),
  \[3554]  = ~v2 & (v1 & ~v0),
  \[7269]  = ~v6 & (~v5 & (~\[11463]  & ~v3)),
  \[11383]  = ~v6 | (~v5 | v4),
  \[14241]  = v11 | (~v10 | ~v9),
  \[12913]  = v12 | (~v11 | ~v8),
  \[6074]  = ~v9 & ~v7,
  \[22107]  = ~\[4738]  | ~\[4749] ,
  \[10530]  = ~v11 | (~v8 | ~v12),
  \[13046]  = ~v0 | ~v2,
  \[5216]  = ~\[12489]  & (~v15 & (v14 & v12)),
  \[13775]  = ~v7 | v5,
  \[22109]  = ~\[4716]  | ~\[4727] ,
  \[10199]  = ~v11 | ~v9,
  \[11391]  = ~v3 | (~v1 | v0),
  \[22103]  = ~\[4789]  | (~\[4796]  | ~\[4784] ),
  \[13782]  = ~v3 | (~v1 | v0),
  \[10193]  = ~\[1471]  | (~\[1478]  | (~\[1464]  | ~\[1511] )),
  \[762]  = ~\[13412]  & (~\[13386]  & (~\[13348]  & ~\[13311] )),
  \[8800]  = ~\[10699]  & (~v15 & v14),
  \[7609]  = ~\[11294]  & (~v6 & (v4 & ~v3)),
  \[22105]  = ~\[4765]  | (~\[4770]  | ~\[4760] ),
  \[12583]  = ~v10 | ~v9,
  \[10195]  = ~v8 | (~v3 | v1),
  \[4025]  = ~\[13087]  & (~v3 & (v2 & v0)),
  \[21647]  = ~\[9220]  | (~\[9212]  | (v6 | ~v4)),
  \[12586]  = v15 | (~v14 | v13),
  \[10537]  = ~\[9130]  | (v6 | ~v4),
  \[21649]  = ~\[9202]  | (~\[9194]  | (~v7 | v5)),
  \[2369]  = ~v11 & (v10 & (v9 & ~v8)),
  \[9663]  = ~v7 & (v6 & ~v5),
  \[22111]  = ~\[4694]  | ~\[4705] ,
  \[4029]  = v13 & ~v12,
  \[10539]  = ~v11 | (~v8 | ~v12),
  \[7277]  = v12 & (v11 & ~v9),
  \[12592]  = ~\[5015]  | (~v3 | (~v1 | v0)),
  \[11399]  = ~\[7405]  | (v15 | (~v14 | ~v12)),
  \[5221]  = ~v8 & (v7 & ~v5),
  \[11731]  = ~v11 | ~v8,
  \[5951]  = v1 & ~v0,
  \[6419]  = ~\[11888]  & (~v3 & (v2 & ~v1)),
  \[3564]  = ~v10 & (~v9 & (~v12 & ~\[13318] )),
  \[2705]  = ~v6 & (~v5 & ~\[13746] ),
  \[8808]  = v3 & (v1 & ~v0),
  \[11393]  = ~v6 | (~v5 | v4),
  \[14251]  = v11 | (~v10 | ~v9),
  \[12923]  = ~v15 | (~v13 | ~\[4351] ),
  \[22117]  = ~\[4636]  | ~\[4647] ,
  \[1511]  = ~\[10123]  & (~\[10110]  & (~\[10095]  & ~\[10079] )),
  \[5226]  = ~v3 & (v2 & ~v1),
  \[21651]  = ~\[9184]  | (~\[9176]  | (~v7 | v5)),
  \[22119]  = ~\[4614]  | ~\[4625] ,
  \[13060]  = ~v15 | ~v13,
  \[4760]  = ~\[12719]  & (~v15 & (v14 & ~v13)),
  \[6087]  = ~\[12041]  & (~v3 & (v2 & ~v1)),
  \[13790]  = ~v2 | v1,
  \[8476]  = ~v10 & ~v9,
  \[1514]  = ~\[10797]  & (~\[10516]  & (~\[10319]  & ~\[10193] )),
  \[7617]  = ~v10 & (~v9 & ~v12),
  \[22113]  = ~v4 | (~v7 | (~\[4682]  | ~\[4674] )),
  \[3903]  = ~v10 & (~v9 & ~v12),
  \[22115]  = ~v4 | (~v7 | (~\[4664]  | ~\[4656] )),
  \[12593]  = ~v10 | ~v9,
  \[4035]  = ~v10 & (v8 & ~v7),
  \[4765]  = ~v8 & (v7 & ~v5),
  \[11005]  = ~v6 | (~v5 | v4),
  \[12596]  = v15 | (~v14 | v13),
  \[6424]  = ~v15 & (v14 & ~v13),
  \[775]  = ~\[374]  & (~\[373]  & (~\[375]  & ~\[13244] )),
  \[11740]  = ~v11 | ~v8,
  \[10547]  = ~v11 | (~v8 | ~v12),
  \[14256]  = ~\[22417]  | (~\[22415]  | (~\[22413]  | ~\[22411] )),
  \[9673]  = ~v7 & (v6 & ~v5),
  \[1182]  = ~\[11358]  & (~\[11332]  & (~\[11292]  & ~\[11257] )),
  \[12208]  = ~\[992]  | (~\[999]  | (~\[985]  | ~\[1030] )),
  \[22121]  = ~v15 | (~v13 | (~\[4593]  | ~\[4603] )),
  \[13798]  = ~v0 | ~v2,
  \[3572]  = ~v3 & (v2 & v0),
  \[7287]  = ~v6 & (~v5 & (~\[11455]  & ~v3)),
  \[2713]  = ~v12 & (~v10 & v8),
  \[12209]  = ~v2 | v1,
  \[6429]  = ~v10 & (v8 & ~v7),
  \[12939]  = ~v11 | ~v8,
  \[14262]  = ~\[1671]  | (v3 | (~v2 | ~v0)),
  \[8818]  = ~\[10689]  & (~v15 & v14),
  \[12203]  = ~\[5809]  | (v14 | ~v13),
  \[12933]  = ~v15 | ~v13,
  \[10545]  = ~\[9107]  | (v3 | (~v2 | ~v0)),
  \[13063]  = ~\[22177]  | (~\[22175]  | (~\[22173]  | ~\[22171] )),
  \[22127]  = ~v15 | (~v13 | (~\[4539]  | ~\[4549] )),
  \[11018]  = ~v6 | (~v5 | v4),
  \[6095]  = ~v13 & (v11 & ~v9),
  \[13065]  = ~v0 | ~v2,
  \[22129]  = ~\[4530]  | (~\[4522]  | (~v7 | v5)),
  \[4770]  = ~v3 & (v2 & ~v1),
  \[2382]  = ~v4 & (~v2 & (v1 & ~v0)),
  \[7627]  = ~\[11285]  & (~v3 & (v2 & ~v1)),
  \[22123]  = ~v15 | (~v13 | (~\[4575]  | ~\[4585] )),
  \[782]  = ~\[368]  & (~\[367]  & (~\[366]  & ~\[365] )),
  \[13409]  = ~v15 | ~v13,
  \[11013]  = ~\[21757]  | (~\[21755]  | (~\[21753]  | ~\[21751] )),
  \[1526]  = ~\[14311]  & (~v14 & (v13 & ~v12)),
  \[22125]  = ~\[4566]  | (~\[4558]  | (v6 | ~v4)),
  \[11746]  = ~v4 | ~v7,
  \[9681]  = ~v7 & (v6 & ~v5),
  \[10558]  = ~v11 | (~v8 | v7),
  \[14263]  = ~v10 | ~v9,
  \[4047]  = ~\[13076]  & (~v3 & (v2 & ~v1)),
  \[14266]  = v14 | (~v13 | v12),
  \[21669]  = ~v4 | (~v7 | (~\[9014]  | ~\[9006] )),
  \[22131]  = ~v15 | (~v13 | (~\[4503]  | ~\[4513] )),
  \[12948]  = ~v11 | ~v8,
  \[9684]  = ~v14 & ~v13,
  \[12217]  = ~v0 | ~v2,
  \[7296]  = ~\[11451]  & (~v15 & v14),
  \[5240]  = ~\[12479]  & (~v15 & (v14 & v12)),
  \[10559]  = ~v12 | ~v14,
  \[5970]  = ~v3 & (v2 & v0),
  \[3582]  = ~v10 & (~v9 & (~v12 & ~\[13308] )),
  \[2723]  = ~v6 & (~v5 & (~\[13737]  & ~v2)),
  \[8826]  = ~v2 & (v1 & ~v0),
  \[789]  = ~\[364]  & (~\[363]  & (~\[362]  & ~\[361] )),
  \[13412]  = ~\[22249]  | (~\[22247]  | ~\[22251] ),
  \[1195]  = ~\[164]  & (~\[163]  & (~\[165]  & ~\[11190] )),
  \[10556]  = ~\[9094]  | (~v6 | (~v5 | v4)),
  \[5245]  = ~v7 & (v6 & v5),
  \[13076]  = ~v6 | (~v5 | v4),
  \[2728]  = ~v14 & (v13 & ~v12),
  \[21671]  = ~v4 | (~v7 | (~\[8996]  | ~\[8988] )),
  \[8494]  = ~v10 & ~v9,
  \[7635]  = ~v10 & (~v9 & ~v12),
  \[3921]  = ~v12 & (~v10 & v8),
  \[13417]  = v3 | (~v2 | v1),
  \[14277]  = ~v13 | v12,
  \[6441]  = ~\[11879]  & (~v3 & (v2 & v0)),
  \[11753]  = ~\[21915]  | (~\[21913]  | (~\[21911]  | ~\[21909] )),
  \[4784]  = ~\[12709]  & (~v15 & (v14 & ~v13)),
  \[8101]  = ~v10 & (~v9 & ~v13),
  \[1537]  = ~\[14308]  & (~v3 & (v2 & v0)),
  \[4055]  = ~v12 & (~v10 & v8),
  \[794]  = ~\[14339]  & (~\[13998]  & (~\[13696]  & ~\[13415] )),
  \[11025]  = ~v1 | v0,
  \[11755]  = v2 | (~v1 | v0),
  \[10568]  = ~v11 | (~v8 | v7),
  \[10900]  = ~v0 | ~v2,
  \[14273]  = ~\[1654]  | (v7 | (~v6 | ~v5)),
  \[14276]  = v11 | (~v10 | (~v9 | v8)),
  \[3590]  = ~v3 & (v2 & ~v1),
  \[13415]  = ~\[782]  | (~\[789]  | (~\[775]  | ~\[762] )),
  \[12228]  = v6 | ~v4,
  \[6446]  = ~v15 & (v14 & ~v13),
  \[12958]  = ~v15 | ~v13,
  \[11762]  = ~v1 | v0,
  \[13087]  = ~v6 | (~v5 | v4),
  \[21673]  = ~v4 | (~v7 | (~\[8978]  | ~\[8970] )),
  \[4789]  = ~v7 & (v6 & v5),
  \[2733]  = ~v10 & (v8 & ~v7),
  \[8836]  = ~\[10681]  & (~v15 & v14),
  \[11761]  = ~\[6633]  | (v15 | ~v14),
  \[2004]  = ~\[14096]  & (~v14 & (v13 & ~v12)),
  \[5252]  = ~v4 & (~v3 & (v2 & v0)),
  \[10563]  = v3 | (~v2 | ~v0),
  \[21675]  = ~v4 | (~v7 | (~\[8960]  | ~\[8952] )),
  \[403]  = ~\[13543]  & ~\[13538] ,
  \[404]  = ~\[13547]  & (~\[13545]  & ~\[13553] ),
  \[10565]  = ~v6 | (~v5 | v4),
  \[9699]  = ~v7 & (v6 & ~v5),
  \[405]  = ~\[13531]  & (~\[13529]  & (~v14 & v13)),
  \[10570]  = v15 | (~v14 | ~v12),
  \[7645]  = ~v6 & (~v5 & (~\[11275]  & ~v3)),
  \[22149]  = ~v4 | (~v7 | (~\[4342]  | ~\[4334] )),
  \[3599]  = ~v10 & (~v9 & ~v12),
  \[10909]  = ~\[21735]  | (~\[21733]  | (~\[21731]  | ~\[21729] )),
  \[5988]  = ~v3 & (v2 & ~v1),
  \[6451]  = ~v10 & (v8 & ~v7),
  \[12961]  = ~\[22155]  | (~\[22153]  | (~\[22151]  | ~\[22149] )),
  \[9308]  = ~\[10444]  & (~v15 & (v14 & v12)),
  \[8111]  = ~\[11044]  & (~v2 & (v1 & ~v0)),
  \[4065]  = ~\[13065]  & (~v6 & (v4 & ~v3)),
  \[3206]  = ~\[13497]  & (~v12 & (v11 & ~v9)),
  \[14284]  = ~v5 | ~v6,
  \[21687]  = ~\[8844]  | (~\[8836]  | (v6 | ~v4)),
  \[13423]  = ~v15 | (~v13 | ~\[3357] ),
  \[11035]  = ~v3 | (~v1 | v0),
  \[1548]  = ~\[14331]  & (~v14 & (v13 & ~v12)),
  \[11765]  = ~v6 | (~v5 | v4),
  \[10578]  = ~v11 | (~v8 | ~v12),
  \[10910]  = ~v2 | v1,
  \[14283]  = v4 | (v3 | (~v2 | ~v0)),
  \[4796]  = ~v4 & (~v3 & (v2 & v0)),
  \[21689]  = ~\[8826]  | (~\[8818]  | (~v7 | v5)),
  \[13425]  = v3 | (~v2 | ~v0),
  \[8844]  = v3 & (v1 & ~v0),
  \[22151]  = ~v4 | (~v7 | (~\[4324]  | ~\[4316] )),
  \[21683]  = ~\[8871]  | (~\[8881]  | (v15 | ~v14)),
  \[11771]  = ~\[6675]  | (v15 | (~v14 | v13)),
  \[12969]  = ~v15 | (~v13 | ~\[4217] ),
  \[14292]  = ~\[1615]  | (v14 | (~v13 | v12)),
  \[2015]  = ~\[14093]  & (~v2 & (v1 & ~v0)),
  \[21685]  = ~\[8862]  | (~\[8854]  | (v6 | ~v4)),
  \[13431]  = ~v15 | (~v13 | ~\[3339] ),
  \[12234]  = ~v0 | ~v2,
  \[2745]  = ~\[13728]  & (v3 & (v1 & ~v0)),
  \[10576]  = ~\[9050]  | (~v7 | v5),
  \[8119]  = ~v10 & (~v9 & ~v13),
  \[12963]  = v2 | (~v1 | v0),
  \[414]  = ~\[13634]  & (~\[13632]  & (~v14 & v13)),
  \[7653]  = ~v10 & (~v9 & ~v12),
  \[415]  = ~\[13646]  & ~\[13641] ,
  \[5266]  = ~\[12466]  & (~v15 & (v14 & v12)),
  \[416]  = ~\[13648]  & (~v3 & (~\[13651]  & ~\[13657] )),
  \[21691]  = ~\[8808]  | (~\[8800]  | (~v7 | v5)),
  \[3940]  = ~\[13110]  & (~v12 & (~v10 & v8)),
  \[12970]  = ~v1 | v0,
  \[417]  = ~\[13663]  & (~\[13661]  & (~v14 & v13)),
  \[10919]  = ~\[8331]  | (v15 | (~v14 | ~v12)),
  \[14298]  = ~v10 | ~v9,
  \[22153]  = ~v4 | (~v7 | (~\[4306]  | ~\[4298] )),
  \[14297]  = ~\[1597]  | (v3 | (~v2 | v1)),
  \[11044]  = v6 | ~v4,
  \[3214]  = ~v3 & (v2 & ~v1),
  \[10913]  = ~v6 | (~v5 | v4),
  \[22155]  = ~v4 | (~v7 | (~\[4288]  | ~\[4280] )),
  \[4074]  = ~\[13060]  & (~v12 & (~v10 & v8)),
  \[11773]  = ~v3 | (~v1 | v0),
  \[13434]  = v3 | (~v2 | v1),
  \[6463]  = ~\[11868]  & (~v3 & (v2 & ~v1)),
  \[9319]  = ~\[10441]  & (~v2 & (v1 & ~v0)),
  \[21697]  = ~\[8754]  | (~\[8746]  | (v6 | ~v4)),
  \[11775]  = ~v6 | (~v5 | v4),
  \[2750]  = ~v14 & (v13 & ~v12),
  \[1559]  = ~\[14328]  & (~v3 & (v2 & ~v1)),
  \[3948]  = ~v3 & (v2 & ~v1),
  \[8854]  = ~\[10672]  & (~v15 & v14),
  \[13440]  = ~v15 | (~v13 | ~\[3321] ),
  \[12247]  = ~v6 | (~v5 | v4),
  \[10921]  = v3 | (~v2 | v1),
  \[21693]  = ~\[8781]  | (~\[8791]  | (v15 | ~v14)),
  \[11051]  = ~\[21765]  | (~\[21763]  | (~\[21761]  | ~\[21759] )),
  \[5271]  = ~v7 & (v6 & v5),
  \[11781]  = ~\[6653]  | (v15 | (~v14 | v13)),
  \[6800]  = ~v15 & (v14 & ~v13),
  \[10584]  = ~\[9027]  | (v3 | (~v2 | ~v0)),
  \[13442]  = v3 | (~v2 | ~v0),
  \[12979]  = ~\[4259]  | (~v15 | (~v13 | v12)),
  \[21695]  = ~\[8763]  | (~\[8773]  | (v15 | ~v14)),
  \[2755]  = ~v10 & (v8 & ~v7),
  \[10586]  = ~v11 | (~v8 | ~v12),
  \[8129]  = ~v6 & (~v5 & ~\[11035] ),
  \[12243]  = ~\[22019]  | (~\[22017]  | (~\[22015]  | ~\[22013] )),
  \[12973]  = ~v6 | (~v5 | v4),
  \[7663]  = ~v6 & (~v5 & (~\[11266]  & ~v3)),
  \[22167]  = ~v15 | (~v13 | (~\[4163]  | ~\[4173] )),
  \[10927]  = ~\[8368]  | (v15 | (~v14 | ~v12)),
  \[22169]  = ~\[4154]  | (~\[4146]  | (~v7 | v5)),
  \[11787]  = ~v3 | (~v1 | v0),
  \[13448]  = ~v15 | (~v13 | ~\[3303] ),
  \[5278]  = ~v4 & (~v3 & (v2 & ~v1)),
  \[10929]  = v3 | (~v2 | ~v0),
  \[22163]  = ~v15 | (~v13 | (~\[4199]  | ~\[4209] )),
  \[4082]  = ~v3 & (v2 & ~v1),
  \[3223]  = ~v12 & (v11 & ~v9),
  \[0]  = ~\[794]  | (~\[1033]  | (~\[1273]  | ~\[1514] )),
  \[6471]  = ~v13 & (~v10 & v8),
  \[12981]  = ~v3 | (~v1 | v0),
  \[5612]  = ~v3 & (v2 & v0),
  \[11053]  = ~v3 | (~v1 | v0),
  \[22165]  = ~\[4190]  | (~\[4182]  | (v6 | ~v4)),
  \[9328]  = ~\[10435]  & (~v15 & v14),
  \[8862]  = ~v2 & (v1 & ~v0),
  \[10597]  = ~v12 | (v10 | ~v8),
  \[2031]  = ~v8 & (v7 & ~v5),
  \[3958]  = ~v10 & (~v9 & (~v12 & ~\[13126] )),
  \[22171]  = ~v15 | (~v13 | (~\[4127]  | ~\[4137] )),
  \[12257]  = ~v6 | (~v5 | v4),
  \[11061]  = ~v3 | (~v1 | v0),
  \[4422]  = ~v3 & (v2 & ~v1),
  \[8137]  = ~v10 & (~v9 & ~v13),
  \[12989]  = ~\[4237]  | (~v15 | (~v13 | v12)),
  \[13451]  = ~v2 | v1,
  \[7671]  = ~v10 & (~v9 & ~v12),
  \[12983]  = ~v6 | (~v5 | v4),
  \[2767]  = ~\[13718]  & (~v2 & (v1 & ~v0)),
  \[1570]  = ~\[14321]  & (~v14 & (v13 & ~v12)),
  \[22177]  = ~\[4082]  | (~\[4074]  | (v6 | ~v4)),
  \[436]  = ~\[13838]  & (~v3 & (~\[13841]  & ~\[13847] )),
  \[22179]  = ~v15 | (~v13 | (~\[4055]  | ~\[4065] )),
  \[437]  = ~\[13849]  & (~\[13855]  & (v7 & ~v5)),
  \[4091]  = ~v12 & (~v10 & v8),
  \[438]  = ~\[13858]  & (~\[13864]  & (v7 & ~v5)),
  \[22173]  = ~v15 | (~v13 | (~\[4109]  | ~\[4119] )),
  \[439]  = ~\[13870]  & (~\[13868]  & (~v14 & v13)),
  \[9336]  = v3 & (v1 & ~v0),
  \[6481]  = ~\[11857]  & (~v6 & (v4 & ~v3)),
  \[10206]  = v15 | (~v14 | ~v13),
  \[22175]  = ~v15 | (~v13 | (~\[4091]  | ~\[4101] )),
  \[13454]  = ~v6 | (~v5 | v4),
  \[8871]  = v12 & (~v10 & v8),
  \[11796]  = v6 | ~v4,
  \[10935]  = ~\[8350]  | (v15 | (~v14 | ~v12)),
  \[3966]  = ~v2 & (v1 & ~v0),
  \[11070]  = ~v7 | v5,
  \[11407]  = ~v12 | (~v11 | v9),
  \[22181]  = ~\[4029]  | (~v15 | (~\[4035]  | ~\[4047] )),
  \[13460]  = ~\[3283]  | (~v15 | (~v13 | v12)),
  \[12267]  = ~v7 | v5,
  \[10211]  = ~v3 | ~v0,
  \[5290]  = ~\[12454]  & (~v15 & (v14 & v12)),
  \[440]  = ~\[13880]  & (~\[13878]  & (~v14 & v13)),
  \[4431]  = ~v12 & (v11 & v8),
  \[441]  = ~\[13888]  & (~v11 & (~\[13891]  & ~\[13887] )),
  \[8147]  = ~v6 & (~v5 & (~\[11025]  & ~v2)),
  \[6489]  = ~v13 & (~v10 & v8),
  \[442]  = ~\[13899]  & (~v11 & (~\[13902]  & ~\[13898] )),
  \[13461]  = ~v0 | ~v2,
  \[2775]  = ~v12 & (~v10 & v8),
  \[7681]  = ~\[11259]  & (v7 & ~v5),
  \[443]  = ~\[13915]  & ~\[13909] ,
  \[6822]  = ~v15 & (v14 & ~v13),
  \[11405]  = ~\[7389]  | (v2 | (~v1 | v0)),
  \[22187]  = ~v15 | (~v13 | (~\[3975]  | ~\[3985] )),
  \[10948]  = v15 | (~v14 | ~v12),
  \[1581]  = ~\[14316]  & (~v8 & (v7 & ~v5)),
  \[12995]  = ~v3 | (~v1 | v0),
  \[11077]  = ~\[21769]  | (~\[21767]  | ~\[21771] ),
  \[22189]  = ~v4 | (~v7 | (~\[3966]  | ~\[3958] )),
  \[3241]  = ~v12 & (v11 & ~v9),
  \[12607]  = v15 | (~v14 | v13),
  \[448]  = ~\[13979]  & (~v11 & (~\[13982]  & ~\[13978] )),
  \[5630]  = ~v3 & (v2 & ~v1),
  \[22183]  = ~\[4007]  | (~v15 | (~\[4013]  | ~\[4025] )),
  \[449]  = ~\[13989]  & (~v11 & (~\[13992]  & ~\[13988] )),
  \[9346]  = ~\[10426]  & (~v15 & v14),
  \[12604]  = ~v10 | ~v9,
  \[7689]  = ~v10 & (~v9 & ~v12),
  \[22185]  = ~\[4002]  | (~\[3994]  | (~v7 | v5)),
  \[13464]  = ~v6 | (~v5 | v4),
  \[3975]  = ~v12 & (~v10 & v8),
  \[8881]  = ~v6 & (~v5 & ~\[10660] ),
  \[12603]  = ~\[4993]  | (v2 | (~v1 | v0)),
  \[10215]  = ~v3 | ~v0,
  \[8152]  = ~v15 & (v14 & ~v13),
  \[11080]  = ~\[1261]  | (~\[1268]  | (~\[1254]  | ~\[1241] )),
  \[22191]  = ~v4 | (~v7 | (~\[3948]  | ~\[3940] )),
  \[10952]  = ~v7 | v5,
  \[13470]  = ~\[3261]  | (~v15 | (~v13 | v12)),
  \[11082]  = v3 | (~v2 | v1),
  \[450]  = ~\[13969]  & (~v11 & (~\[13972]  & ~\[13968] )),
  \[2053]  = ~v8 & (v7 & ~v5),
  \[13807]  = ~\[22335]  | (~\[22333]  | (~\[22331]  | ~\[22329] )),
  \[451]  = ~\[14004]  & (~v11 & (~\[14007]  & ~\[14003] )),
  \[5639]  = ~v12 & (v11 & ~v9),
  \[8157]  = ~v9 & (~v7 & ~v10),
  \[6499]  = ~\[11848]  & (~v3 & (v2 & ~v1)),
  \[452]  = ~\[14014]  & (~v11 & (~\[14017]  & ~\[14013] )),
  \[2785]  = ~\[13708]  & (v3 & (v1 & ~v0)),
  \[11413]  = ~\[7371]  | (~v3 | (~v1 | v0)),
  \[1926]  = ~v4 & (~v2 & (v1 & ~v0)),
  \[453]  = ~\[14025]  & (~v11 & (~\[14028]  & ~\[14024] )),
  \[12273]  = ~v0 | ~v2,
  \[454]  = ~\[14035]  & (~v11 & (~\[14038]  & ~\[14034] )),
  \[11415]  = ~v12 | (~v11 | v9),
  \[455]  = ~\[14053]  & ~\[14047] ,
  \[11088]  = ~\[8029]  | (v15 | ~v14),
  \[6105]  = ~\[12056]  & (~v6 & (v4 & ~v3)),
  \[456]  = ~\[14057]  & (~v7 & (~\[14056]  & ~\[14065] )),
  \[457]  = ~\[14072]  & (~v11 & (~\[14075]  & ~\[14071] )),
  \[9354]  = ~v2 & (v1 & ~v0),
  \[12617]  = v15 | (~v14 | v13),
  \[11422]  = ~\[7358]  | (v6 | ~v4),
  \[458]  = ~\[14082]  & (~v11 & (~\[14085]  & ~\[14081] )),
  \[10959]  = ~v0 | ~v2,
  \[12282]  = ~\[22027]  | (~\[22025]  | (~\[22023]  | ~\[22021] )),
  \[6838]  = ~v3 & (v2 & ~v1),
  \[13479]  = ~v15 | (~v13 | ~\[3241] ),
  \[13811]  = ~v6 | (~v5 | v4),
  \[12614]  = ~v10 | ~v9,
  \[7699]  = ~\[11250]  & (~v2 & (v1 & ~v0)),
  \[3985]  = ~\[13112]  & (v7 & (~v5 & ~v3)),
  \[1597]  = ~v8 & (v7 & ~v5),
  \[12613]  = ~\[4971]  | (~v3 | (~v1 | v0)),
  \[13473]  = v3 | (~v2 | v1),
  \[7304]  = v3 & (v1 & ~v0),
  \[11090]  = v3 | (~v2 | ~v0),
  \[8893]  = ~v6 & ~v5,
  \[1202]  = ~\[158]  & (~\[157]  & (~\[156]  & ~\[155] )),
  \[12287]  = ~v4 | (~v7 | ~\[5630] ),
  \[5649]  = ~\[12273]  & (v7 & (~v5 & ~v3)),
  \[12289]  = v12 | (~v11 | v9),
  \[2794]  = ~\[13702]  & (~v14 & (v13 & ~v12)),
  \[11424]  = ~v12 | (~v11 | v9),
  \[13481]  = v3 | (~v2 | ~v0),
  \[463]  = ~\[14152]  & (~v14 & (~\[14151]  & ~\[14148] )),
  \[9360]  = ~v14 & (v12 & ~v3),
  \[8169]  = ~\[11018]  & (v3 & (v1 & ~v0)),
  \[6113]  = ~v13 & (v11 & ~v9),
  \[464]  = ~\[14158]  & (~v7 & (~\[14157]  & ~\[14166] )),
  \[10238]  = v7 | (~v6 | v5),
  \[1938]  = ~\[14127]  & (~v14 & (v13 & ~v12)),
  \[465]  = ~\[14138]  & (~v11 & (~\[14141]  & ~\[14137] )),
  \[1209]  = ~\[154]  & (~\[153]  & (~\[152]  & ~\[151] )),
  \[11430]  = ~\[7335]  | (~v3 | (~v1 | v0)),
  \[12628]  = v11 | (~v10 | ~v9),
  \[4458]  = ~v3 & (v2 & ~v1),
  \[3261]  = v11 & (~v9 & ~v7),
  \[13820]  = v6 | ~v4,
  \[11432]  = ~v12 | (~v11 | v9),
  \[10969]  = ~v4 | ~v7,
  \[13487]  = ~v15 | (~v13 | ~\[3223] ),
  \[11099]  = v3 | (~v2 | v1),
  \[2404]  = v3 & (v1 & ~v0),
  \[3994]  = ~\[13100]  & (~v12 & (~v10 & v8)),
  \[11096]  = ~\[8011]  | (v15 | ~v14),
  \[10235]  = ~\[21555]  | (~\[21553]  | (~\[21551]  | ~\[21549] )),
  \[7314]  = ~\[11443]  & (~v15 & v14),
  \[2071]  = ~v11 & (v10 & (v9 & ~v8)),
  \[8174]  = ~v15 & (v14 & ~v13),
  \[10242]  = v12 | (~v3 | ~v0),
  \[5657]  = ~v12 & (v11 & ~v9),
  \[12297]  = v12 | (~v11 | v9),
  \[6851]  = ~v6 & v4,
  \[8179]  = ~v9 & (~v7 & ~v10),
  \[6123]  = ~\[12050]  & (~v3 & (v2 & ~v1)),
  \[474]  = ~\[14263]  & (~v11 & (~\[14266]  & ~\[14262] )),
  \[8512]  = ~v10 & ~v9,
  \[475]  = ~\[14277]  & (~v14 & (~\[14276]  & ~\[14273] )),
  \[9372]  = ~v15 & (v14 & (v13 & ~v12)),
  \[12295]  = ~v4 | (~v7 | ~\[5612] ),
  \[13826]  = ~v0 | ~v2,
  \[1949]  = ~\[14124]  & (v3 & (v1 & ~v0)),
  \[476]  = ~\[14284]  & (~v7 & (~\[14283]  & ~\[14292] )),
  \[4467]  = ~v12 & (v11 & v8),
  \[12638]  = v11 | (~v10 | ~v9),
  \[477]  = ~\[14298]  & (~v11 & (~\[14301]  & ~\[14297] )),
  \[13100]  = ~v15 | ~v13,
  \[3609]  = ~\[13294]  & (v7 & (~v5 & ~v3)),
  \[10979]  = ~v4 | ~v7,
  \[13497]  = ~v15 | ~v13,
  \[10976]  = ~\[21749]  | (~\[21747]  | (~\[21745]  | ~\[21743] )),
  \[7322]  = ~v2 & (v1 & ~v0),
  \[9379]  = ~v3 & (v2 & (v1 & ~v0)),
  \[5667]  = ~\[12267]  & (~v3 & (v2 & ~v1)),
  \[13838]  = ~v0 | ~v2,
  \[6131]  = ~v13 & (v11 & ~v9),
  \[11443]  = ~v12 | (~v11 | v9),
  \[14301]  = v14 | (~v13 | v12),
  \[13103]  = ~\[22185]  | (~\[22183]  | (~\[22181]  | ~\[22179] )),
  \[10987]  = ~v4 | ~v7,
  \[3618]  = ~v10 & (~v9 & (~v12 & ~\[13291] )),
  \[13835]  = ~\[22339]  | (~\[22337]  | ~\[22341] ),
  \[13110]  = ~v15 | ~v13,
  \[14308]  = v8 | (~v7 | ~v4),
  \[11451]  = ~v12 | (~v11 | v9),
  \[3283]  = v11 & (~v9 & ~v7),
  \[13112]  = ~v0 | ~v2,
  \[12649]  = v11 | (~v10 | ~v9),
  \[5672]  = ~v14 & (v13 & ~v12),
  \[13841]  = ~v6 | (~v5 | v4),
  \[823]  = ~\[13129]  & (~\[13103]  & (~\[13063]  & ~\[13028] )),
  \[8191]  = ~\[11005]  & (~v2 & (v1 & ~v0)),
  \[2426]  = ~v2 & (v1 & ~v0),
  \[9389]  = v2 & (v1 & ~v0),
  \[21707]  = ~\[8647]  | (~\[8657]  | (v15 | ~v14)),
  \[1960]  = ~\[14117]  & (v15 & (v13 & ~v12)),
  \[5676]  = ~v9 & ~v7,
  \[21709]  = ~\[8629]  | (~\[8639]  | (v15 | ~v14)),
  \[7335]  = ~v6 & v4,
  \[13847]  = ~\[2509]  | (v14 | (~v13 | v12)),
  \[6141]  = ~v6 & (~v5 & (~\[12028]  & ~v3)),
  \[13849]  = v3 | (~v2 | v1),
  \[14311]  = v11 | (~v10 | ~v9),
  \[8199]  = ~v10 & (~v9 & ~v13),
  \[4485]  = ~v12 & (v11 & v8),
  \[2097]  = ~v11 & (v10 & (v9 & ~v8)),
  \[3626]  = ~v3 & (v2 & ~v1),
  \[11455]  = ~v2 | v1,
  \[6874]  = ~v3 & (v2 & ~v1),
  \[8533]  = ~v9 & (~v7 & ~v10),
  \[10267]  = ~\[21569]  | (~\[21567]  | (~\[21565]  | ~\[21563] )),
  \[21711]  = ~v4 | (~v7 | (~\[8620]  | ~\[8612] )),
  \[4822]  = ~v4 & (~v3 & (v2 & ~v1)),
  \[6149]  = ~v13 & (v11 & ~v9),
  \[12659]  = v11 | (~v10 | ~v9),
  \[12654]  = v3 | (~v2 | ~v0),
  \[103]  = ~\[10635]  & (~v2 & (~\[10638]  & ~\[10644] )),
  \[10996]  = ~v4 | ~v7,
  \[104]  = ~\[10648]  & (~\[10646]  & ~\[10654] ),
  \[105]  = ~\[10632]  & (~\[10630]  & (~v15 & v14)),
  \[1241]  = ~\[11077]  & (~\[11051]  & (~\[11013]  & ~\[10976] )),
  \[1971]  = ~\[14114]  & (~v3 & (v2 & v0)),
  \[836]  = ~\[344]  & (~\[343]  & (~\[345]  & ~\[12961] )),
  \[14316]  = v3 | (~v2 | ~v0),
  \[13858]  = v3 | (~v2 | ~v0),
  \[5689]  = ~\[12257]  & (~v3 & (v2 & v0)),
  \[9006]  = ~\[10597]  & (~v15 & v14),
  \[13129]  = ~\[22189]  | (~\[22187]  | ~\[22191] ),
  \[11463]  = ~v0 | ~v2,
  \[14321]  = v11 | (~v10 | ~v9),
  \[10605]  = ~v11 | (~v8 | ~v12),
  \[9739]  = ~v8 & (v3 & v0),
  \[13126]  = ~v15 | ~v13,
  \[3638]  = ~v9 & (~v7 & (~v10 & ~\[13283] )),
  \[13855]  = ~\[2489]  | (v14 | ~v13),
  \[11472]  = ~\[21855]  | (~\[21853]  | (~\[21851]  | ~\[21849] )),
  \[4101]  = ~v6 & (~v5 & (~\[13046]  & ~v3)),
  \[6887]  = ~v6 & ~v5,
  \[14328]  = v8 | (~v7 | ~v4),
  \[13132]  = ~\[843]  | (~\[850]  | (~\[836]  | ~\[823] )),
  \[2444]  = ~v3 & (v2 & v0),
  \[6159]  = ~v6 & (~v5 & (~\[12020]  & ~v3)),
  \[11804]  = ~v3 | (~v1 | v0),
  \[12664]  = ~\[22095]  | (~\[22093]  | (~\[22091]  | ~\[22089] )),
  \[843]  = ~\[338]  & (~\[337]  & (~\[336]  & ~\[335] )),
  \[114]  = ~\[10735]  & (~\[10733]  & (~v15 & v14)),
  \[5694]  = ~v14 & (v13 & ~v12),
  \[115]  = ~\[10738]  & (~v3 & (~\[10741]  & ~\[10747] )),
  \[9742]  = ~v11 & v10,
  \[116]  = ~\[10749]  & (~v3 & (~\[10752]  & ~\[10758] )),
  \[21729]  = ~\[8441]  | (~\[8451]  | (v15 | ~v14)),
  \[12670]  = ~\[4822]  | (v7 | (~v6 | ~v5)),
  \[117]  = ~\[10764]  & (~\[10762]  & (~v15 & v14)),
  \[1982]  = ~\[14106]  & (v15 & (v13 & ~v12)),
  \[9014]  = ~v2 & (v1 & ~v0),
  \[13868]  = ~v4 | (~v7 | ~\[2462] ),
  \[4109]  = ~v12 & (~v10 & v8),
  \[5698]  = ~v9 & ~v7,
  \[4839]  = ~v8 & (~v6 & v4),
  \[3642]  = v5 & ~v4,
  \[1254]  = ~\[134]  & (~\[133]  & (~\[135]  & ~\[10909] )),
  \[5301]  = ~\[12449]  & (~v8 & (~v6 & v4)),
  \[10614]  = ~v11 | (~v8 | ~v12),
  \[7358]  = ~v2 & (v1 & ~v0),
  \[11473]  = ~v2 | v1,
  \[14331]  = v11 | (~v10 | ~v9),
  \[13864]  = ~\[2471]  | (v14 | ~v13),
  \[11476]  = ~v6 | (~v5 | v4),
  \[10288]  = v6 | (~v5 | v4),
  \[13136]  = v3 | (~v2 | ~v0),
  \[21731]  = ~\[8423]  | (~\[8433]  | (v15 | ~v14)),
  \[3648]  = ~v3 & (v2 & v0),
  \[10622]  = ~v12 | (v10 | ~v8),
  \[8555]  = ~v9 & (~v7 & ~v10),
  \[6167]  = ~v13 & (v11 & ~v9),
  \[13870]  = v12 | (v10 | ~v8),
  \[11482]  = ~\[7203]  | (v15 | (~v14 | ~v12)),
  \[850]  = ~\[334]  & (~\[333]  & (~\[332]  & ~\[331] )),
  \[121]  = ~\[10805]  & (~\[10803]  & (~v15 & v14)),
  \[14337]  = ~\[22429]  | (~\[22427]  | (~\[22431]  | ~\[567] )),
  \[13142]  = ~v15 | (~v13 | ~\[3921] ),
  \[122]  = ~\[10809]  & (~\[10815]  & (v7 & v4)),
  \[12674]  = ~v14 | v13,
  \[123]  = ~\[10817]  & (~v2 & (~\[10820]  & ~\[10826] )),
  \[11813]  = ~v7 | v5,
  \[14339]  = ~\[604]  | (~\[611]  | (~\[597]  | ~\[584] )),
  \[12673]  = v11 | (~v10 | (~v9 | v8)),
  \[124]  = ~\[10830]  & (~\[10828]  & ~\[10836] ),
  \[10285]  = ~\[21577]  | (~\[21575]  | (~\[21573]  | ~\[21571] )),
  \[125]  = ~v6 & (~v5 & (~\[10840]  & ~\[10846] )),
  \[1261]  = ~\[128]  & (~\[127]  & (~\[126]  & ~\[125] )),
  \[11488]  = ~v12 | (~v11 | v9),
  \[126]  = ~v6 & (~v5 & (~\[10848]  & ~\[10854] )),
  \[11820]  = ~\[21929]  | (~\[21927]  | (~\[21925]  | ~\[21923] )),
  \[127]  = ~\[10857]  & (~\[10863]  & (~v6 & v4)),
  \[10292]  = v6 | (~v5 | v4),
  \[13878]  = ~v4 | (~v7 | ~\[2444] ),
  \[128]  = ~\[10865]  & (~\[10871]  & (~v6 & v4)),
  \[6507]  = ~v13 & (~v10 & v8),
  \[1993]  = ~\[14103]  & (~v3 & (v2 & ~v1)),
  \[4119]  = ~v6 & (~v5 & (~\[13037]  & ~v3)),
  \[11822]  = ~v3 | (~v1 | v0),
  \[21733]  = ~\[8405]  | (~\[8415]  | (v15 | ~v14)),
  \[12682]  = ~v10 | ~v9,
  \[12681]  = ~\[4861]  | (v3 | (~v2 | v1)),
  \[9027]  = v7 & ~v5,
  \[21735]  = ~\[8387]  | (~\[8397]  | (v15 | ~v14)),
  \[10626]  = ~\[21675]  | (~\[21673]  | (~\[21671]  | ~\[21669] )),
  \[13144]  = ~v3 | (~v1 | v0),
  \[11486]  = ~\[7250]  | (v6 | ~v4),
  \[1268]  = ~\[124]  & (~\[123]  & (~\[122]  & ~\[121] )),
  \[10630]  = ~\[8893]  | (v2 | (~v1 | v0)),
  \[22209]  = ~\[3778]  | (~\[3770]  | (~v7 | v5)),
  \[5317]  = ~v8 & (~v6 & v4),
  \[10632]  = ~v12 | (v10 | ~v8),
  \[13150]  = ~v15 | (~v13 | ~\[3903] ),
  \[3659]  = ~v9 & (~v7 & ~v10),
  \[2462]  = ~v3 & (v2 & ~v1),
  \[6177]  = ~\[12012]  & (v7 & ~v5),
  \[13880]  = v12 | (v10 | ~v8),
  \[10299]  = ~v5 | v4,
  \[7707]  = ~v10 & (~v9 & ~v12),
  \[11829]  = ~v2 | v1,
  \[13152]  = ~v1 | v0,
  \[7371]  = ~v6 & ~v5,
  \[133]  = ~\[10921]  & (~\[10927]  & (~v6 & v4)),
  \[10296]  = ~v5 | v4,
  \[134]  = ~\[10929]  & (~\[10935]  & (~v6 & v4)),
  \[21747]  = ~\[8271]  | (~\[8281]  | (v15 | ~v14)),
  \[135]  = ~\[10910]  & (~v3 & (~\[10913]  & ~\[10919] )),
  \[10638]  = ~v6 | (~v5 | v4),
  \[12685]  = v15 | (~v14 | v13),
  \[4127]  = ~v12 & (~v10 & v8),
  \[21749]  = ~\[8253]  | (~\[8263]  | (v15 | ~v14)),
  \[22211]  = ~v15 | (~v13 | (~\[3751]  | ~\[3761] )),
  \[1273]  = ~\[11924]  & (~\[11643]  & (~\[11361]  & ~\[11080] )),
  \[2802]  = ~v3 & (v2 & v0),
  \[13888]  = ~v10 | ~v9,
  \[6517]  = ~v6 & (~v5 & (~\[11838]  & ~v3)),
  \[21743]  = ~\[8314]  | (~v6 | (~\[8320]  | ~\[8310] )),
  \[13887]  = ~\[2426]  | (v8 | (~v7 | ~v4)),
  \[12692]  = ~v10 | ~v9,
  \[12691]  = ~\[4839]  | (v3 | (~v2 | ~v0)),
  \[11494]  = ~\[7227]  | (v3 | (~v2 | ~v0)),
  \[21745]  = ~\[8289]  | (~\[8299]  | (v15 | ~v14)),
  \[8909]  = ~v10 & (v8 & ~v7),
  \[11496]  = ~v12 | (~v11 | v9),
  \[10635]  = ~v1 | v0,
  \[6185]  = ~v13 & (v11 & ~v9),
  \[11838]  = ~v0 | ~v2,
  \[13155]  = ~v6 | (~v5 | v4),
  \[21751]  = ~\[8235]  | (~\[8245]  | (v15 | ~v14)),
  \[2471]  = ~v12 & (~v10 & v8),
  \[8574]  = ~v10 & ~v9,
  \[11107]  = v3 | (~v2 | ~v0),
  \[4861]  = ~v8 & (~v6 & v4),
  \[7717]  = ~\[11241]  & (~v6 & v4),
  \[22213]  = ~v15 | (~v13 | (~\[3733]  | ~\[3743] )),
  \[1615]  = ~v11 & (v10 & (v9 & ~v8)),
  \[13161]  = ~\[3883]  | (~v15 | (~v13 | v12)),
  \[13891]  = ~v15 | (~v13 | v12),
  \[22215]  = ~v15 | (~v13 | (~\[3715]  | ~\[3725] )),
  \[21757]  = ~\[8174]  | (~\[8179]  | ~\[8191] ),
  \[11105]  = ~\[7993]  | (v15 | ~v14),
  \[10648]  = ~v6 | (~v5 | v4),
  \[12695]  = v15 | (~v14 | v13),
  \[6525]  = ~v13 & (~v10 & v8),
  \[4137]  = ~\[13030]  & (v7 & ~v5),
  \[21759]  = ~\[8152]  | (~\[8157]  | ~\[8169] ),
  \[2812]  = ~\[13672]  & (~v14 & (v13 & ~v12)),
  \[13898]  = ~\[2404]  | (v8 | (~v7 | ~v4)),
  \[21753]  = ~\[8217]  | (~\[8227]  | (v15 | ~v14)),
  \[10644]  = ~\[8931]  | (v15 | (~v14 | ~v12)),
  \[1285]  = ~\[117]  & (~\[116]  & (~\[115]  & ~\[114] )),
  \[12309]  = v15 | (~v14 | ~v12),
  \[21755]  = ~\[8199]  | (~\[8209]  | (v15 | ~v14)),
  \[7389]  = ~v6 & ~v5,
  \[13899]  = ~v10 | ~v9,
  \[10646]  = ~v3 | (~v1 | v0),
  \[13163]  = ~v3 | (~v1 | v0),
  \[12306]  = ~v10 | ~v9,
  \[22227]  = ~v15 | (~v13 | (~\[3599]  | ~\[3609] )),
  \[12305]  = ~\[5594]  | (v8 | (~v7 | ~v4)),
  \[6195]  = ~\[12005]  & (~v2 & (v1 & ~v0)),
  \[11848]  = v6 | ~v4,
  \[13165]  = ~v6 | (~v5 | v4),
  \[21761]  = ~\[8137]  | (~\[8147]  | (v15 | ~v14)),
  \[7725]  = ~v10 & (~v9 & ~v12),
  \[22229]  = ~v4 | (~v7 | (~\[3590]  | ~\[3582] )),
  \[3679]  = ~v10 & (~v9 & ~v12),
  \[11119]  = ~v6 | (~v5 | v4),
  \[151]  = ~v6 & (~v5 & (~\[11082]  & ~\[11088] )),
  \[22223]  = ~\[3642]  | (~v6 | (~\[3648]  | ~\[3638] )),
  \[5339]  = ~v6 & (~v5 & ~v8),
  \[152]  = ~v6 & (~v5 & (~\[11090]  & ~\[11096] )),
  \[882]  = ~\[12848]  & (~\[12822]  & (~\[12784]  & ~\[12745] )),
  \[13171]  = ~\[3861]  | (~v15 | (~v13 | v12)),
  \[11113]  = ~\[7975]  | (v15 | ~v14),
  \[153]  = ~\[11099]  & (~\[11105]  & (~v6 & v4)),
  \[22225]  = ~\[3626]  | (~\[3618]  | (~v7 | v5)),
  \[9050]  = ~v3 & (v2 & ~v1),
  \[11116]  = ~v2 | v1,
  \[154]  = ~\[11107]  & (~\[11113]  & (~v6 & v4)),
  \[21767]  = ~\[8083]  | (~\[8093]  | (v15 | ~v14)),
  \[155]  = ~\[11116]  & (~v3 & (~\[11119]  & ~\[11125] )),
  \[4146]  = ~\[13025]  & (~v12 & (~v10 & v8)),
  \[2820]  = ~v3 & (v2 & ~v1),
  \[156]  = ~\[11126]  & (~v3 & (~\[11129]  & ~\[11135] )),
  \[6535]  = ~v6 & (~v5 & (~\[11829]  & ~v3)),
  \[21769]  = ~\[8065]  | (~\[8075]  | (v15 | ~v14)),
  \[2489]  = ~v12 & (~v10 & v8),
  \[13505]  = ~v15 | ~v13,
  \[157]  = ~\[11138]  & (~\[11144]  & (v7 & ~v5)),
  \[22231]  = ~v4 | (~v7 | (~\[3572]  | ~\[3564] )),
  \[4878]  = ~\[12659]  & (~v15 & (v14 & ~v13)),
  \[158]  = ~\[11146]  & (~\[11152]  & (v7 & ~v5)),
  \[21763]  = ~\[8119]  | (~\[8129]  | (v15 | ~v14)),
  \[10654]  = ~\[8909]  | (v15 | (~v14 | ~v12)),
  \[13512]  = ~v11 | ~v8,
  \[12319]  = v15 | (~v14 | ~v12),
  \[21765]  = ~\[8101]  | (~\[8111]  | (v15 | ~v14)),
  \[12316]  = ~v10 | ~v9,
  \[22237]  = ~\[3506]  | (~v11 | (~\[3502]  | ~\[3519] )),
  \[10660]  = ~v3 | (~v1 | v0),
  \[12315]  = ~\[5572]  | (v8 | (~v7 | ~v4)),
  \[13175]  = v2 | (~v1 | v0),
  \[21771]  = ~\[8047]  | (~\[8057]  | (v15 | ~v14)),
  \[2829]  = ~v12 & (~v10 & v8),
  \[7735]  = ~\[11233]  & (~v2 & (v1 & ~v0)),
  \[22239]  = ~\[3484]  | (~v11 | (~\[3480]  | ~\[3497] )),
  \[11857]  = ~v0 | ~v2,
  \[11129]  = ~v6 | (~v5 | v4),
  \[22233]  = ~v4 | (~v7 | (~\[3554]  | ~\[3546] )),
  \[13181]  = ~v15 | (~v13 | ~\[3841] ),
  \[163]  = ~\[11199]  & (~v2 & (~\[11202]  & ~\[11208] )),
  \[22235]  = ~v4 | (~v7 | (~\[3536]  | ~\[3528] )),
  \[4154]  = ~v2 & (v1 & ~v0),
  \[11126]  = ~v0 | ~v2,
  \[8931]  = ~v10 & (v8 & ~v7),
  \[164]  = ~\[11212]  & (~\[11210]  & ~\[11218] ),
  \[6543]  = ~v13 & (~v10 & v8),
  \[11125]  = ~\[7955]  | (v15 | (~v14 | v13)),
  \[165]  = ~v6 & (~v5 & (~\[11192]  & ~\[11198] )),
  \[11855]  = ~\[21937]  | (~\[21935]  | (~\[21933]  | ~\[21931] )),
  \[895]  = ~\[314]  & (~\[313]  & (~\[315]  & ~\[12664] )),
  \[22241]  = ~v15 | (~v13 | (~\[3465]  | ~\[3475] )),
  \[13520]  = ~v11 | ~v8,
  \[4889]  = ~v6 & (~v5 & (~v8 & ~\[12654] )),
  \[12329]  = v11 | (~v10 | ~v9),
  \[13189]  = ~v15 | (~v13 | ~\[3823] ),
  \[8209]  = ~\[10996]  & (v3 & (v1 & ~v0)),
  \[9401]  = ~v3 & (v2 & (v1 & ~v0)),
  \[13183]  = ~v3 | (~v1 | v0),
  \[7013]  = ~v6 & ~v5,
  \[7743]  = ~v10 & (~v9 & ~v12),
  \[22247]  = ~v15 | (~v13 | (~\[3411]  | ~\[3421] )),
  \[3697]  = ~v10 & (~v9 & ~v12),
  \[11138]  = v3 | (~v2 | v1),
  \[11868]  = ~v6 | (~v5 | v4),
  \[2839]  = ~\[13686]  & (~v2 & (v1 & ~v0)),
  \[22249]  = ~\[3402]  | (~\[3394]  | (~v7 | v5)),
  \[10672]  = ~v12 | (v10 | ~v8),
  \[22243]  = ~v15 | (~v13 | (~\[3447]  | ~\[3457] )),
  \[3303]  = ~v12 & (v11 & ~v9),
  \[13192]  = v2 | (~v1 | v0),
  \[4163]  = ~v12 & (~v10 & v8),
  \[13529]  = ~\[3093]  | (v2 | (~v1 | v0)),
  \[22245]  = ~\[3438]  | (~\[3430]  | (v6 | ~v4)),
  \[6553]  = ~\[11822]  & (v7 & ~v5),
  \[11135]  = ~\[7933]  | (v15 | (~v14 | v13)),
  \[2110]  = ~v4 & (~v3 & (v2 & ~v1)),
  \[21789]  = ~\[7877]  | (~\[7887]  | (v14 | ~v13)),
  \[13525]  = ~\[22275]  | (~\[22273]  | (~\[22271]  | ~\[22269] )),
  \[22251]  = ~v15 | (~v13 | (~\[3375]  | ~\[3385] )),
  \[13198]  = ~v15 | (~v13 | ~\[3805] ),
  \[5361]  = ~v6 & (~v5 & ~v8),
  \[8217]  = v12 & (~v10 & ~v9),
  \[4503]  = ~v12 & (v11 & v8),
  \[13531]  = v12 | (~v11 | ~v8),
  \[7753]  = ~v6 & (~v5 & ~\[11224] ),
  \[7024]  = ~v15 & (v14 & ~v13),
  \[2848]  = ~\[13680]  & (~v14 & (v13 & ~v12)),
  \[9413]  = ~v3 & (v2 & (v1 & ~v0)),
  \[21791]  = ~\[7859]  | (~\[7869]  | (v15 | ~v14)),
  \[13538]  = ~\[3142]  | (~v6 | (~v5 | v4)),
  \[10681]  = ~v12 | (v10 | ~v8),
  \[1654]  = ~v4 & (~v3 & (v2 & ~v1)),
  \[181]  = ~\[11368]  & (~\[11366]  & (~v15 & v14)),
  \[11879]  = ~v6 | (~v5 | v4),
  \[12341]  = v11 | (~v10 | (~v9 | v8)),
  \[11144]  = ~\[7913]  | (v15 | ~v14),
  \[182]  = ~\[11376]  & (~\[11374]  & (~v15 & v14)),
  \[6561]  = ~v13 & (~v10 & v8),
  \[4173]  = ~\[13012]  & (~v6 & v4),
  \[183]  = ~\[11380]  & (~v2 & (~\[11383]  & ~\[11389] )),
  \[11146]  = v3 | (~v2 | ~v0),
  \[184]  = ~\[11393]  & (~\[11391]  & ~\[11399] ),
  \[8952]  = ~\[10622]  & (~v15 & v14),
  \[185]  = ~\[11407]  & (~\[11405]  & (~v15 & v14)),
  \[186]  = ~\[11415]  & (~\[11413]  & (~v15 & v14)),
  \[187]  = ~\[11424]  & (~\[11422]  & (~v15 & v14)),
  \[11152]  = ~\[7895]  | (v15 | ~v14),
  \[188]  = ~\[11432]  & (~\[11430]  & (~v15 & v14)),
  \[10689]  = ~v12 | (v10 | ~v8),
  \[21793]  = ~\[7841]  | (~\[7851]  | (v15 | ~v14)),
  \[14007]  = ~v15 | (~v13 | v12),
  \[8227]  = ~\[10987]  & (~v3 & (v2 & v0)),
  \[4513]  = ~\[12824]  & (v7 & ~v5),
  \[21795]  = ~\[7823]  | (~\[7833]  | (v14 | ~v13)),
  \[7761]  = ~v10 & (~v9 & ~v12),
  \[2856]  = ~v3 & (v2 & v0),
  \[14004]  = ~v10 | ~v9,
  \[2127]  = ~v8 & (~v6 & v4),
  \[14003]  = ~\[2193]  | (v3 | (~v2 | v1)),
  \[11158]  = ~v4 | ~v7,
  \[11888]  = ~v7 | v5,
  \[6905]  = ~v6 & ~v5,
  \[22269]  = ~v4 | (~v7 | (~\[3214]  | ~\[3206] )),
  \[3321]  = ~v12 & (v11 & ~v9),
  \[13547]  = ~v6 | (~v5 | v4),
  \[4182]  = ~\[13008]  & (~v12 & (~v10 & v8)),
  \[5711]  = ~\[12247]  & (~v3 & (v2 & ~v1)),
  \[6571]  = ~\[11813]  & (~v2 & (v1 & ~v0)),
  \[8960]  = v3 & (v1 & ~v0),
  \[193]  = ~\[11488]  & (~\[11486]  & (~v15 & v14)),
  \[194]  = ~\[11496]  & (~\[11494]  & (~v15 & v14)),
  \[13543]  = ~\[3126]  | (~v11 | (~v8 | v7)),
  \[195]  = ~\[11473]  & (~v3 & (~\[11476]  & ~\[11482] )),
  \[13545]  = ~v3 | (~v1 | v0),
  \[22271]  = ~v4 | (~v7 | (~\[3196]  | ~\[3188] )),
  \[9094]  = ~v3 & (v2 & ~v1),
  \[8235]  = v12 & (~v10 & ~v9),
  \[10699]  = ~v12 | (v10 | ~v8),
  \[14017]  = ~v15 | (~v13 | v12),
  \[5719]  = ~v12 & (v11 & ~v9),
  \[4522]  = ~\[12843]  & (v15 & (v13 & ~v12)),
  \[12359]  = ~\[22039]  | (~\[22037]  | (~\[22041]  | ~\[954] )),
  \[6579]  = ~v13 & (~v10 & v8),
  \[10693]  = ~\[21689]  | (~\[21687]  | (~\[21685]  | ~\[21683] )),
  \[5383]  = ~v8 & (v7 & ~v5),
  \[12353]  = v11 | (~v10 | (~v9 | v8)),
  \[14014]  = ~v10 | ~v9,
  \[14013]  = ~\[2171]  | (v3 | (~v2 | ~v0)),
  \[1671]  = ~v8 & (~v6 & v4),
  \[11898]  = ~v4 | ~v7,
  \[4190]  = ~v2 & (v1 & ~v0),
  \[22273]  = ~v4 | (~v7 | (~\[3178]  | ~\[3170] )),
  \[13559]  = ~v3 | (~v1 | v0),
  \[8970]  = ~\[10614]  & (~v15 & v14),
  \[22275]  = ~v4 | (~v7 | (~\[3160]  | ~\[3152] )),
  \[11166]  = ~v4 | ~v7,
  \[13553]  = ~\[3104]  | (~v11 | (~v8 | v7)),
  \[11895]  = ~\[21945]  | (~\[21943]  | (~\[21941]  | ~\[21939] )),
  \[4530]  = ~v2 & (v1 & ~v0),
  \[3339]  = ~v12 & (v11 & ~v9),
  \[8245]  = ~\[10979]  & (~v3 & (v2 & ~v1)),
  \[4199]  = ~v12 & (~v10 & v8),
  \[14028]  = ~v15 | (~v13 | v12),
  \[6920]  = ~\[11619]  & (~v15 & (v14 & ~v13)),
  \[5729]  = ~\[12234]  & (~v6 & (v4 & ~v3)),
  \[12369]  = v15 | (~v14 | ~v12),
  \[2874]  = ~v3 & (v2 & ~v1),
  \[6589]  = ~\[11804]  & (~v6 & v4),
  \[8978]  = ~v3 & (v2 & v0),
  \[7781]  = ~v9 & (~v7 & ~v10),
  \[7052]  = ~\[11571]  & (~v15 & (v14 & ~v13)),
  \[11506]  = ~v6 | (~v5 | v4),
  \[14024]  = ~\[2149]  | (v3 | (~v2 | v1)),
  \[12366]  = ~v10 | ~v9,
  \[22287]  = ~\[3044]  | (~\[3036]  | (v6 | ~v4)),
  \[12365]  = ~\[5471]  | (~v3 | (~v1 | v0)),
  \[10317]  = ~\[21589]  | (~\[21587]  | (~\[21591]  | ~\[1404] )),
  \[2149]  = ~v8 & (~v6 & v4),
  \[22289]  = ~\[3026]  | (~\[3018]  | (~v7 | v5)),
  \[14025]  = ~v10 | ~v9,
  \[10319]  = ~\[1441]  | (~\[1448]  | (~\[1434]  | ~\[1421] )),
  \[4539]  = ~v12 & (v11 & v8),
  \[22283]  = ~\[3071]  | (~\[3081]  | (v14 | ~v13)),
  \[6928]  = v3 & (v1 & ~v0),
  \[13902]  = ~v15 | (~v13 | v12),
  \[12709]  = v11 | (~v10 | (~v9 | v8)),
  \[22285]  = ~\[3062]  | (~\[3054]  | (v6 | ~v4)),
  \[11175]  = ~v4 | ~v7,
  \[1688]  = ~\[14251]  & (~v14 & (v13 & ~v12)),
  \[8253]  = ~v10 & (~v9 & ~v13),
  \[2880]  = ~v14 & (v13 & ~v12),
  \[11518]  = ~v12 | (~v11 | v9),
  \[22291]  = ~\[3008]  | (~\[3000]  | (~v7 | v5)),
  \[5737]  = ~v12 & (v11 & ~v9),
  \[13570]  = ~v11 | ~v8,
  \[6597]  = ~v13 & (~v10 & v8),
  \[14038]  = ~v15 | (~v13 | v12),
  \[12379]  = v15 | (~v14 | ~v12),
  \[13909]  = ~\[2382]  | (v7 | (~v6 | ~v5)),
  \[8988]  = ~\[10605]  & (~v15 & v14),
  \[6203]  = ~v13 & (v11 & ~v9),
  \[14034]  = ~\[2127]  | (v3 | (~v2 | ~v0)),
  \[7063]  = ~\[11568]  & (~v2 & (v1 & ~v0)),
  \[12376]  = ~v10 | ~v9,
  \[22297]  = ~\[2954]  | (~\[2946]  | (v6 | ~v4)),
  \[12375]  = ~\[5449]  | (v2 | (~v1 | v0)),
  \[14035]  = ~v10 | ~v9,
  \[1693]  = ~v8 & (~v6 & v4),
  \[11522]  = ~v0 | ~v2,
  \[4549]  = ~\[12832]  & (~v6 & v4),
  \[22293]  = ~\[2990]  | (~\[2982]  | (v6 | v5)),
  \[6938]  = ~\[11635]  & (~v15 & (v14 & ~v13)),
  \[12719]  = v11 | (~v10 | ~v9),
  \[10323]  = v12 | (v6 | (~v5 | v4)),
  \[9457]  = ~v3 & (v2 & (v1 & ~v0)),
  \[13579]  = ~v11 | ~v8,
  \[11183]  = ~v4 | ~v7,
  \[10326]  = ~v5 | v4,
  \[22295]  = ~\[2963]  | (~\[2973]  | (v14 | ~v13)),
  \[1698]  = ~v3 & (v2 & ~v1),
  \[5015]  = ~v6 & (~v5 & ~v8),
  \[3357]  = ~v12 & (v11 & ~v9),
  \[8263]  = ~\[10969]  & (~v2 & (v1 & ~v0)),
  \[11190]  = ~\[21795]  | (~\[21793]  | (~\[21791]  | ~\[21789] )),
  \[1302]  = ~\[10728]  & (~\[10693]  & ~\[10795] ),
  \[7405]  = v11 & (~v9 & ~v7),
  \[5747]  = ~\[12228]  & (~v3 & (v2 & ~v1)),
  \[12387]  = ~v10 | ~v9,
  \[11192]  = v2 | (~v1 | v0),
  \[10331]  = ~v7 | (~v5 | v4),
  \[8996]  = ~v3 & (v2 & ~v1),
  \[14047]  = ~\[2110]  | (v7 | (~v6 | ~v5)),
  \[7072]  = ~\[11561]  & (~v15 & (v14 & ~v13)),
  \[6213]  = ~\[11993]  & (~v6 & v4),
  \[8602]  = ~v3 & (v2 & v0),
  \[12386]  = ~\[5427]  | (~v3 | (~v1 | v0)),
  \[11198]  = ~\[7761]  | (v14 | ~v13),
  \[12390]  = v15 | (~v14 | ~v12),
  \[13915]  = ~\[2369]  | (~v15 | (~v13 | v12)),
  \[567]  = ~\[477]  & (~\[476]  & (~\[475]  & ~\[474] )),
  \[6946]  = ~v2 & (v1 & ~v0),
  \[4558]  = ~\[12817]  & (v15 & (v13 & ~v12)),
  \[9464]  = v5 & ~v4,
  \[13587]  = ~v11 | ~v8,
  \[11199]  = ~v1 | v0,
  \[902]  = ~\[308]  & (~\[307]  & (~\[306]  & ~\[305] )),
  \[13921]  = v4 | (~v3 | (~v1 | v0)),
  \[8271]  = v12 & (~v10 & ~v9),
  \[10335]  = ~v7 | (~v5 | v4),
  \[5755]  = ~v12 & (v11 & ~v9),
  \[12725]  = v3 | (~v2 | ~v0),
  \[2171]  = ~v6 & (~v5 & ~v8),
  \[2509]  = ~v10 & (v8 & ~v7),
  \[12730]  = v11 | (~v10 | ~v9),
  \[12397]  = ~v10 | ~v9,
  \[10341]  = ~v7 | (~v5 | v4),
  \[11539]  = ~\[21869]  | (~\[21867]  | (~\[21865]  | ~\[21863] )),
  \[14057]  = ~v5 | ~v6,
  \[909]  = ~\[304]  & (~\[303]  & (~\[302]  & ~\[301] )),
  \[12001]  = ~\[21967]  | (~\[21965]  | (~\[21963]  | ~\[21961] )),
  \[7080]  = v3 & (v1 & ~v0),
  \[13592]  = ~\[22289]  | (~\[22287]  | (~\[22285]  | ~\[22283] )),
  \[1315]  = ~\[104]  & (~\[103]  & (~\[105]  & ~\[10626] )),
  \[6221]  = ~v13 & (v11 & ~v9);
endmodule

