//NOTE: no-implementation module stub

module lmi_watchb (
    input wire DATAUPI,
    input wire DATADOWNI,
    input wire C_IADDR_A,
    input wire C_IREAD_I_N,
    input wire IX_VAL,
    input wire IX_MISS_S_R,
    input wire C_DADDR_E,
    input wire C_DREAD_E,
    input wire C_DWRITE_E,
    input wire C_DBYEN_E,
    input wire CP0_XCPN_M,
    input wire DC_VAL,
    input wire DC_MISS_W_R,
    input wire X_HALT_R,
    input wire DATAUPI_buf,
    input wire DATADOWNI_buf,
    input wire C_IADDR_A_buf,
    input wire C_IREAD_I_N_buf,
    input wire IX_VAL_buf,
    input wire IX_MISS_S_R_buf,
    input wire C_DADDR_E_buf,
    input wire C_DREAD_E_buf,
    input wire C_DWRITE_E_buf,
    input wire C_DBYEN_E_buf,
    input wire CP0_XCPN_M_buf,
    input wire DC_VAL_buf,
    input wire DC_MISS_W_R_buf,
    input wire X_HALT_R_buf
);

endmodule
