//NOTE: no-implementation module stub

module mux32 (
    output wire OUT,
    input wire THRU,
    input wire IN,
    input wire EN1,
    input wire DIS1,
    input wire DIS2
);

endmodule
