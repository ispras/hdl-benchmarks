//NOTE: no-implementation module stub

module REG9L (
    input wire DSPCLK,
    input wire CLKovfenb,
    input wire MRovfwe,
    input wire [8:0] MACin,
    output reg [8:0] MRovf
);

endmodule
