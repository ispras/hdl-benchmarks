`timescale 1 ps / 1 ps

module cascade (midas_macys,kappa_rufus_outwire);
  input midas_macys;
  output kappa_rufus_outwire;
endmodule
