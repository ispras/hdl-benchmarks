//NOTE: no-implementation module stub

module MEMC (
    input `ifdef FD_EVB PERICLK, `else DSPCLK, `endif
    input GRST,
    input STBY,
    input [15:0] DMDin,
    input PPclr_h,
    input GO_Ex,
    input GO_Cx,
    input redoM_h,
    input redoSTI_h,
    input redoLD_h,
    input IDLE_ST,
    input [3:0] DMOVL_dsp,
    input [7:4] PMOVL_dsp,
    input Pread_R,
    input Pwrite_R,
    input Dread_R,
    input Dwrite_R,
    input IOcmd_R,
    input IOread_R,
    input IOwrite_R,
    input Dummy_R,
    input Dummy_E,
    input [13:5] DMA_R,
    input [13:12] PMA_R,
    input [13:0] DMA,
    input [13:5] DMAin,
    input [13:12] PMAin,
    input SREQ,
    input STEAL,
    input DMSreqx_wr,
    input PMSreqx_wr,
    input DMSreqx_rd,
    input PMSreqx_rd,
    input BOOT,
    input [3:0] PMOVL,
    input [3:0] DMOVL,
    input DSreqx,
    input DRDcyc,
    input T_selECM,
    input BM_cyc,
    input ECYC,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input PM_bdry_sel,
    input SP0_EN,
    input selAUTO0,
    input selFSDIV0,
    input selSCLKDIV0,
    input selSCTL0,
    input selMWORD0,
    input AUTO0_we,
    input FSDIV0_we,
    input SCLKDIV0_we,
    input SCTL0_we,
    input MWORD0_we,
    input SP1_EN,
    input selAUTO1,
    input selFSDIV1,
    input selSCLKDIV1,
    input selSCTL1,
    input selMWORD1,
    input AUTO1_we,
    input FSDIV1_we,
    input SCLKDIV1_we,
    input SCTL1_we,
    input MWORD1_we,
    input selPFTYPE,
    input selPDATA,
    input selPIMASK,
    input selPINT,
    input PFTYPE_we,
    input PDATA_we,
    input PIMASK_we,
    input PINT_we,
    input selTPERIOD,
    input selTCOUNT,
    input selTSCALE,
    input TPERIOD_we,
    input TCOUNT_we,
    input TSCALE_we,
    input Pread_Ei,
    input Pwrite_Ei,
    input Dread_Ei,
    input Dwrite_Ei,
    input IOcmd_Ei,
    input IOread_Ei,
    input IOwrite_Ei,
    input WSCR_we,
    input WSCR_ext_we,
    input selWSCR,
    input selWSCR_ext,
    input EXTC_Eg,
    input [3:0] ECMWAIT,
    input [1:0] ECMAWAIT,
    input selCKR,
    input CKR_we,
    input [2:0] DWWAIT,
    input [2:0] DRWAIT,
    input selDCTL,
    input selDOVL,
    input DCTL_we,
    input DOVL_we,
    input selSYSR,
    input ldSREG_E,
    input MMR_web,
    input TB_EN,
    input DwriteI_Eg,
    input PwriteI_Eg,
    input STI_Cg,
    input LDaST_Eg,
    input BIASRND,
    input accPM_Eg,
    input accDM_Eg,
    input PMo_cs0,
    input PMo_cs1,
    input PMo_cs2,
    input PMo_cs3,
    input PMo_cs4,
    input PMo_cs5,
    input PMo_cs6,
    input PMo_cs7,
    input PMo_web,
    input PMo_oe0_K,
    input PMo_oe1_K,
    input PMo_oe2_K,
    input PMo_oe3_K,
    input PMo_oe4_K,
    input PMo_oe5_K,
    input PMo_oe6_K,
    input PMo_oe7_K,
    input DM_cs,
    input DMo_cs0,
    input DMo_cs1,
    input DMo_cs2,
    input DMo_cs3,
    input DMo_cs4,
    input DMo_cs5,
    input DMo_cs6,
    input DMo_cs7,
    input DMo_web,
    input DM_oe_K,
    input DMo_oe0_K,
    input DMo_oe1_K,
    input DMo_oe2_K,
    input DMo_oe3_K,
    input DMo_oe4_K,
    input DMo_oe5_K,
    input DMo_oe6_K,
    input DMo_oe7_K,
    input selBIAD,
    input selBEAD,
    input selBCTL,
    input selBCNT,
    input selBOVL,
    input BCNT_we,
    input BCTL_we,
    input BOVL_we,
    input BIAD_we,
    input BEAD_we,
    input selIVER
);

endmodule
