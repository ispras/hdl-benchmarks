//NOTE: no-implementation module stub

module IDMA (
    input T_IRDn,
    input T_IWRn,
    input T_ISn,
    input T_IAL,
    input T_BMODE,
    input T_MMAP,
    input T_selECM,
    input PM_bdry_sel,
    input STBY,
    input Awake_h,
    input P_RSTn,
    input GRST,
    `ifdef FD_EVB
    input PERICLK,
    `else
    input DSPCLK,
    `endif
    input GO_Fx,
    input GO_Ex,
    input IDLE_ST_h,
    input ICE_ST_h,
    input ICE_ST,
    input [15:0] DMDin,
    input [7:0] PMOVL_dsp,
    input [3:0] DMOVL_dsp,
    input [13:12] CMAin,
    input redoIF_h,
    input [2:0] DWWAIT,
    input [2:0] DRWAIT,
    input DCTL_we,
    input DOVL_we,
    input MMR_web,
    input STEAL,
    input DSack,
    input DSreqx,
    input [23:0] IDR,
    input accCM_R,
    input accCM_E,
    input wrCM_R,
    input BDMA_end,
    input BDMA_boot,
    input BCMRD_cyc,
    input [11:0] BOVL,
    input [23:0] BRdataBUF,
    input BCM_cyc,
    input BSreqx,
    input BM_cyc,
    input ECYC,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input IACKn,
    input BOOT,
    input [14:0] DCTL,
    input [11:0] DOVL,
    input [3:0] PMOVL,
    input [3:0] DMOVL,
    input idmaDMD_oe,
    input idmaPMD_oe,
    input [15:0] idmaPMD_do,
    input DSreq,
    input DWRcyc,
    input PWRcyc,
    input DRDcyc,
    input PRDcyc,
    input CM_cs,
    input CM_web,
    input CM_oe_K,
    input CMo_cs0,
    input CMo_cs1,
    input CMo_cs2,
    input CMo_cs3,
    input CMo_cs4,
    input CMo_cs5,
    input CMo_cs6,
    input CMo_cs7,
    input CMo_oe0_K,
    input CMo_oe1_K,
    input CMo_oe2_K,
    input CMo_oe3_K,
    input CMo_oe4_K,
    input CMo_oe5_K,
    input CMo_oe6_K,
    input CMo_oe7_K,
    input [15:0] T_IAD,
    input [15:0] IAD_do,
    input IAD_oe,
    input [15:0] PMDin,
    input [23:0] CM_rd,
    input [23:0] CM_wd,
    input GO_STEAL
);

endmodule
