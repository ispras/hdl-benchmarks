




`ifdef LINE_SIZE 
`define LBUS_LINE_SIZE `LINE_SIZE 
`define LBUS_LINE_ADDR_HI `LINE_ADDR_HI 
`define LBUS_LINE_CTR_FIRST `LINE_CTR_FIRST 
`else 
`define LBUS_LINE_SIZE 4 
`define LBUS_LINE_ADDR_HI 3 
`define LBUS_LINE_CTR_FIRST 2'b00 
`endif 



`define LBM_XTION_FIELD 47:44 
`define LBM_DATAPOS_FIELD 43:36 
`define LBM_LENGTH_FIELD 43:36 
`define LBM_BYTEEN_FIELD 39:36 
`define LBM_IRDYDEL_FIELD 35:32 
`define LBM_ADDR_FIELD 31:0 
`define LBM_DATA_FIELD 31:0 



`define LBT_TRDYPOS_FIELD 43:36 
`define LBT_TRDYDEL_FIELD 35:32 
`define LBT_SELDEL_FIELD 33:32 
`define LBT_BASEADDR_FIELD 31:0 



`define LBM_NOOP 4'b0000 
`define LBM_READDATA 4'b0001 
`define LBM_WRITEDATA 4'b0010 
`define LBM_READSINGLE 4'b0011 
`define LBM_WRITESINGLE 4'b0100 
`define LBM_READLINEL 4'b0101 
`define LBM_READLINEI 4'b0110 
`define LBM_WRITELINE 4'b0111 
`define LBM_READBURSTF 4'b1000 
`define LBM_READBURSTU 4'b1001 
`define LBM_WRITEBURSTF 4'b1010 
`define LBM_WRITEBURSTU 4'b1011 
`define LBM_IDLE 4'b1100 
`define LBM_FINISH 4'b1111 



`define LBT_SETBASEADDR 4'b0000 
`define LBT_SETSELDELAY 4'b0001 
`define LBT_SETTRDYDELAY 4'b0010 
`define LBT_EXCLUDEADDR 4'b0011 


