module bitwise_and_1_4_1(a, b, c);
  input a;
  input [3:0] b;
  output c;
  assign c = a & b;
endmodule
