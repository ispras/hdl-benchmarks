//NOTE: no-implementation module stub

module DAG (
    input DSPCLK,
    input T_RST,
    input GO_Ex,
    input GO_Cx,
    input EX_en,
    input STBY,
    input [7:0] MTIreg_E,
    input [7:0] MTLreg_E,
    input [7:0] MTMreg_E,
    input [7:0] MFIreg_E,
    input [7:0] MFLreg_E,
    input [7:0] MFMreg_E,
    input MFDAG1_E,
    input Post1_E,
    input imAddr_R,
    input DAG1D_R,
    input DAG2D_R,
    input DAG1_EN,
    input Double_R,
    input idBR_R,
    input Post2_E,
    input MFDAG2_E,
    input DAG2_EN,
    input DAG2P_R,
    input DMAen_R,
    input [3:0] IRE,
    input [17:0] IR,
    input MSTAT,
    input redoSTI_h,
    input redoEX_h,
    input PwriteI_Eg,
    input DwriteI_Eg,
    input accPM_E,
    input redoM_h,
    input STEAL,
    input T0Sreqx,
    input T1Sreqx,
    input R0Sreqx,
    input R1Sreqx,
    input SREQ,
    input T0sack,
    input T1sack,
    input R0sack,
    input R1sack,
    input [2:0] R0IREG,
    input [2:0] R1IREG,
    input [2:0] T0IREG,
    input [2:0] T1IREG,
    input [1:0] R0MREG,
    input [1:0] R1MREG,
    input [1:0] T0MREG,
    input [1:0] T1MREG,
    input DSreqx,
    input BOOT,
    input [14:0] DCTL,
    input [15:0] DMDid,
    input BSreqx,
    input BPM_cyc,
    input BDM_cyc,
    input [13:0] BIAD,
    input BM_cyc,
    input ECYC,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input T0wrap,
    input T1wrap,
    input R0wrap,
    input R1wrap,
    input [13:0] DMA_R,
    input [13:0] DMA,
    input [13:0] PMA_R,
    input [13:0] PMA,
    input [13:0] DMAin,
    input [13:0] PMAin,
    output [15:0] dagDMD_do
);

endmodule
