//NOTE: no-implementation module stub

module BDMA (
    input BSreqx,
    input BSack,
    input T_MMAP,
    input T_BMODE,
    input [7:0] T_ED,
    input P_RSTn,
    input GRST,
    input PM_bdry_sel,
    input ENS12,
    input ECS12,
    input ENS13,
    input ECS13,
    input ENS14,
    input ECS14,
    input ENS0,
    `ifdef FD_EVB
    input PERICLK,
    `else
    input DSPCLK,
    `endif
    input [23:0] CM_rd,
    input [15:0] PMDin,
    input [15:0] DMDin,
    input BOOT,
    input GO_STEAL,
    input BCNT_we,
    input BCTL_we,
    input BOVL_we,
    input BIAD_we,
    input BEAD_we,
    input selBCNT,
    input selBCTL,
    input selBOVL,
    input selBIAD,
    input selBEAD,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input BDMWR_cyc,
    input BPMWR_cyc,
    input BDMRD_cyc,
    input BPMRD_cyc,
    input BSreq,
    input BDMAmode,
    input [7:0] BMpage,
    input [13:0] BEAD,
    input [7:0] BWdataBUF,
    input BDIR,
    input BWRn,
    input BWend,
    input BDMA_end,
    input BDMA_boot,
    input BCM_cyc,
    input BCMRD_cyc,
    input [23:0] BRdataBUF,
    input [11:0] BOVL,
    input BM_cyc,
    input T_BDMA,
    input BPM_cyc,
    input BDM_cyc,
    input [13:0] BIAD,
    input BRST,
    input [15:0] BDMAmmio,
    input bdmaDMD_oe,
    input bdmaPMD_oe
);

endmodule
