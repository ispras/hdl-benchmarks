//NOTE: no-implementation module stub

module REG8L (
    input wire DSPCLK,
    input wire CLKSErenb,
    input wire SErwe,
    input wire [7:0] SEin,
    output reg [7:0] SEr
);

endmodule
