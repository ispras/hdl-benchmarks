// IWLS benchmark module "rot" printed on Wed May 29 17:28:07 2002
module rot(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8);
input
  z0,
  z1,
  z2,
  z3,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  a1,
  a2,
  a3,
  a4,
  b0,
  b1,
  b2,
  b3,
  b4,
  c0,
  c1,
  c2,
  c3,
  c4,
  d0,
  d1,
  d2,
  d3,
  d4,
  e0,
  e1,
  e2,
  e3,
  e4,
  f0,
  f1,
  f2,
  f3,
  g0,
  g1,
  g2,
  g3,
  h0,
  h1,
  h2,
  h3,
  i0,
  i1,
  i2,
  i3,
  j0,
  j1,
  j2,
  j3,
  k0,
  k1,
  k2,
  k3,
  l0,
  l1,
  l2,
  l3,
  m0,
  m1,
  m2,
  m3,
  n0,
  n1,
  n2,
  n3,
  o0,
  o1,
  o2,
  o3,
  p0,
  p1,
  p2,
  p3,
  q0,
  q1,
  q2,
  q3,
  r0,
  r1,
  r2,
  r3,
  s0,
  s1,
  s2,
  s3,
  t0,
  t1,
  t2,
  t3,
  u0,
  u1,
  u2,
  u3,
  v0,
  v1,
  v2,
  v3,
  w0,
  w1,
  w2,
  w3,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3;
output
  z4,
  z5,
  z6,
  z7,
  a5,
  a6,
  a7,
  a8,
  b5,
  b6,
  b7,
  b8,
  c5,
  c6,
  c7,
  c8,
  d5,
  d6,
  d7,
  d8,
  e5,
  e6,
  e7,
  e8,
  f4,
  f5,
  f6,
  f7,
  f8,
  g4,
  g5,
  g6,
  g7,
  g8,
  h4,
  h5,
  h6,
  h7,
  h8,
  i4,
  i5,
  i6,
  i7,
  j4,
  j5,
  j6,
  j7,
  k4,
  k5,
  k6,
  k7,
  l4,
  l5,
  l6,
  l7,
  m4,
  m5,
  m6,
  m7,
  n4,
  n5,
  n6,
  n7,
  o4,
  o5,
  o6,
  o7,
  p4,
  p5,
  p6,
  p7,
  q4,
  q5,
  q6,
  q7,
  r4,
  r5,
  r6,
  r7,
  s4,
  s5,
  s6,
  s7,
  t4,
  t5,
  t6,
  t7,
  u4,
  u5,
  u6,
  u7,
  v4,
  v5,
  v6,
  v7,
  w4,
  w5,
  w6,
  w7,
  x4,
  x5,
  x6,
  x7,
  y4,
  y5,
  y6,
  y7;
wire
  j13,
  j14,
  j15,
  j16,
  j17,
  r12,
  r13,
  r14,
  r15,
  r16,
  z12,
  z13,
  z14,
  z15,
  z16,
  c13,
  c14,
  c15,
  c16,
  c17,
  k13,
  k14,
  k15,
  k16,
  k17,
  \[6] ,
  s12,
  s13,
  s14,
  s15,
  s16,
  d13,
  d14,
  d15,
  d16,
  d17,
  l12,
  l13,
  l14,
  l15,
  l16,
  l17,
  t12,
  t13,
  t14,
  t15,
  t16,
  e13,
  e14,
  e15,
  e16,
  e17,
  m12,
  m13,
  m14,
  m15,
  m16,
  m17,
  u12,
  u13,
  u14,
  u15,
  u16,
  f13,
  f14,
  f15,
  f16,
  f17,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  v12,
  v13,
  v14,
  v15,
  v16,
  g13,
  g14,
  g15,
  g16,
  g17,
  o12,
  o13,
  o14,
  o15,
  o16,
  o17,
  w12,
  w13,
  w14,
  w15,
  w16,
  h13,
  h14,
  h15,
  h16,
  h17,
  p12,
  p13,
  p14,
  p15,
  p16,
  p17,
  x12,
  x13,
  x14,
  x15,
  x16,
  a13,
  a14,
  a15,
  a16,
  a17,
  \[50] ,
  i13,
  i14,
  i15,
  i16,
  i17,
  q12,
  q13,
  q14,
  q15,
  q16,
  q17,
  y12,
  y13,
  y14,
  y15,
  y16,
  b13,
  b14,
  b15,
  b16,
  b17;
assign
  z4 = c13,
  z5 = a14,
  z6 = x14,
  z7 = q15,
  j13 = (l2 & (~d1 & ~c1)) | (~q17 & l2),
  j14 = (~g16 & (~q2 & r0)) | ((~g16 & (~p2 & r0)) | ((~g16 & (~l2 & r0)) | o16)),
  j15 = h16 & ~s16,
  j16 = r16 & a2,
  j17 = w16 & v16,
  r12 = v16 & w1,
  r13 = (l16 & j16) | ((l16 & j0) | ((~k16 & j16) | ((~k16 & j0) | ((j16 & i16) | (i16 & j0))))),
  r14 = (~g16 & (~e16 & (~g17 & c3))) | ((~e16 & (~g17 & (c3 & b3))) | (e16 & a3)),
  r15 = c4 | j17,
  r16 = t3 | (o3 | n3),
  z12 = (~y15 & (b & ~x15)) | ((y15 & (~b & ~x15)) | (x15 & d2)),
  z13 = (l3 & (t0 & g0)) | a17,
  z14 = (~y3 & (o1 & (~h17 & (~i17 & m1)))) | ((~y3 & (o1 & (~s1 & (~i17 & m1)))) | ((~y3 & (o1 & (~i17 & q2))) | ((~y3 & (o1 & (~i17 & p2))) | ((~y3 & (o1 & (~i17 & ~l2))) | ((~y3 & (o1 & (~i17 & ~q))) | ((~h17 & (~i17 & (m1 & i1))) | ((~s1 & (~i17 & (m1 & i1))) | ((~i17 & (q2 & i1)) | ((~i17 & (p2 & i1)) | ((~i17 & (~l2 & i1)) | (~i17 & (i1 & ~q)))))))))))),
  z15 = (~e17 & (m3 & (~i3 & h3))) | (~e17 & e3),
  z16 = (~z0 & (~y0 & (x0 & ~w0))) | ((~z0 & (y0 & (~x0 & ~w0))) | (z0 & w0)),
  c13 = b4 & v0,
  c14 = (q2 & m2) | ((m2 & m1) | (m2 & r0)),
  c15 = (~k1 & k17) | (~k17 & q3),
  c16 = (~c17 & (d16 & (~g16 & m3))) | ((e16 & (d16 & (~g16 & m3))) | ((~c17 & (i3 & h3)) | ((e16 & (i3 & h3)) | ((~c17 & d17) | (e16 & d17))))),
  c17 = ~a3 & ~z2,
  k13 = (~q17 & l2) | (l2 & ~d1),
  k14 = ~k2 & ~m0,
  k15 = (~h16 & ~r16) | s16,
  k16 = ~a17 & (m0 & (l0 & k0)),
  k17 = (q2 & (p2 & (~m2 & q))) | ((o17 & ~q2) | (o17 & ~p2)),
  \[6]  = ~o3,
  s12 = (l2 & (~h2 & (~g2 & (q16 & (~t2 & ~a))))) | ((l2 & (~h2 & (~g2 & (q16 & (t1 & ~a))))) | ((l2 & (~h2 & (~g2 & (m16 & (~t2 & ~a))))) | ((l2 & (~h2 & (~g2 & (m16 & (t1 & ~a))))) | ((l2 & (~g2 & (~f2 & (q16 & (~t2 & ~a))))) | ((l2 & (~g2 & (~f2 & (q16 & (t1 & ~a))))) | ((l2 & (~g2 & (~f2 & (m16 & (~t2 & ~a))))) | ((l2 & (~g2 & (~f2 & (m16 & (t1 & ~a))))) | ((~l2 & (z1 & (q16 & (~t2 & ~a)))) | ((~l2 & (z1 & (q16 & (t1 & ~a)))) | ((~l2 & (z1 & (m16 & (~t2 & ~a)))) | ((~l2 & (z1 & (m16 & (t1 & ~a)))) | ((~h2 & (~f2 & (q16 & (~t2 & ~a)))) | ((~h2 & (~f2 & (q16 & (t1 & ~a)))) | ((~h2 & (~f2 & (m16 & (~t2 & ~a)))) | ((~h2 & (~f2 & (m16 & (t1 & ~a)))) | ((~h2 & (z1 & (q16 & (~t2 & ~a)))) | ((~h2 & (z1 & (q16 & (t1 & ~a)))) | ((~h2 & (z1 & (m16 & (~t2 & ~a)))) | ((~h2 & (z1 & (m16 & (t1 & ~a)))) | ((~g2 & (z1 & (q16 & (~t2 & ~a)))) | ((~g2 & (z1 & (q16 & (t1 & ~a)))) | ((~g2 & (z1 & (m16 & (~t2 & ~a)))) | ((~g2 & (z1 & (m16 & (t1 & ~a)))) | ((~f2 & (z1 & (q16 & (~t2 & ~a)))) | ((~f2 & (z1 & (q16 & (t1 & ~a)))) | ((~f2 & (z1 & (m16 & (~t2 & ~a)))) | (~f2 & (z1 & (m16 & (t1 & ~a)))))))))))))))))))))))))))))),
  s13 = p16 & (~i16 & ~o16),
  s14 = (~o0 & (~e16 & d3)) | (g17 & c3),
  s15 = ~w16 & (v16 & (x2 & ~w2)),
  s16 = (u15 & n1) | ((~b2 & n1) | ((~s1 & n1) | (r1 & n1))),
  d13 = (~d1 & c1) | (d1 & ~c1),
  d14 = m2 & (~y1 & (x1 & w1)),
  d15 = (~l1 & (k1 & k17)) | ((l1 & (~k1 & k17)) | (~k17 & r3)),
  d16 = (~i3 & h3) | (i3 & ~h3),
  d17 = c17 & (~e16 & (t0 & ~h0)),
  l12 = (~y & (\x  & j1)) | ((y & e0) | (~\x  & e0)),
  l13 = (~q17 & l2) | (l2 & ~c1),
  l14 = (~i3 & (m2 & ~k2)) | ((h3 & (m2 & ~k2)) | ((p2 & ~k2) | (~k2 & ~m0))),
  l15 = (l3 & (a4 & (~u16 & (y3 & (~h16 & (~u15 & (~s16 & t16))))))) | ((l3 & (a4 & (~u16 & (y3 & (~h16 & (~u15 & (~s16 & p16))))))) | ((s & (a4 & (~u16 & (y3 & (~h16 & (~u15 & (~s16 & t16))))))) | ((s & (a4 & (~u16 & (y3 & (~h16 & (~u15 & (~s16 & p16))))))) | ((l3 & (a4 & (~u16 & (~v2 & (~h16 & (~u15 & t16)))))) | ((l3 & (a4 & (~u16 & (~v2 & (~h16 & (~u15 & p16)))))) | ((s & (a4 & (~u16 & (~v2 & (~h16 & (~u15 & t16)))))) | ((s & (a4 & (~u16 & (~v2 & (~h16 & (~u15 & p16)))))) | ((a4 & (y3 & (~u2 & (~h16 & (~u15 & (~s16 & t16)))))) | ((a4 & (y3 & (~u2 & (~h16 & (~u15 & (~s16 & p16)))))) | ((a4 & (~f16 & (y3 & (h16 & (~u15 & ~s16))))) | ((a4 & (g16 & (y3 & (h16 & (~u15 & ~s16))))) | ((a4 & (y3 & (~y2 & (h16 & (~u15 & ~s16))))) | ((a4 & (~v2 & (~u2 & (~h16 & (~u15 & t16))))) | ((a4 & (~v2 & (~u2 & (~h16 & (~u15 & p16))))) | ((a4 & (~f16 & (~v2 & (h16 & ~u15)))) | ((a4 & (g16 & (~v2 & (h16 & ~u15)))) | ((a4 & (~y2 & (~v2 & (h16 & ~u15)))) | ((a4 & (~q16 & (h16 & ~u15))) | ((a4 & (~q16 & (~u15 & s16))) | ((a4 & (~q16 & (~u15 & t16))) | ((a4 & (~q16 & (~u15 & p16))) | (a4 & (~v2 & (~u15 & s16)))))))))))))))))))))))),
  l16 = n3 & (t0 & ~h0),
  l17 = (q2 & (p2 & (~m2 & p))) | n17,
  t12 = (~h2 & (~f2 & (~t1 & (~a & t2)))) | (t2 & a1),
  t13 = (j16 & ~o3) | m17,
  t14 = (x16 & (l2 & ~k2)) | m17,
  t15 = (~v16 & w2) | ~a4,
  t16 = e4 & i1,
  e13 = (~e1 & (d1 & c1)) | ((e1 & ~d1) | (e1 & ~c1)),
  e14 = (~q2 & p2) | (q2 & ~p2),
  e15 = t16 & y3,
  e16 = (l2 & (o0 & (c17 & (~g16 & (~c3 & b3))))) | ((l2 & (o0 & (c17 & (~c3 & (b3 & ~a3))))) | ((l2 & (o0 & (c17 & (~c3 & (b3 & z2))))) | ((l2 & (o0 & (c17 & (~g16 & d3)))) | ((l2 & (o0 & (c17 & (d3 & ~a3)))) | ((l2 & (o0 & (c17 & (d3 & z2)))) | ((c17 & (~g16 & (~d3 & (~c3 & ~b3)))) | ((c17 & (~d3 & (~c3 & (~b3 & ~a3)))) | (c17 & (~d3 & (~c3 & (~b3 & z2))))))))))),
  e17 = ~u15 & (b2 & v1),
  m12 = (~y1 & p0) | (y1 & k1),
  m13 = e1 & (d1 & (c1 & n)),
  m14 = (y16 & h3) | (d17 | o16),
  m15 = (d4 & ~s1) | ((j17 & ~s1) | (u15 & ~s1)),
  m16 = (~z3 & (h16 & (f16 & (~g16 & (~u15 & y2))))) | ((~l3 & (~s & (~z3 & (~u15 & u2)))) | ((~z3 & (~u15 & (s16 & v2))) | ((~z3 & (~u15 & (u16 & u2))) | ((~z3 & (~u15 & (~y3 & v2))) | ((~w16 & (v16 & w2)) | (~x2 & w2)))))),
  m17 = ~p17 & (~z16 & j2),
  u12 = (~q & (~p & (~o & (~g2 & (~s1 & (~r1 & (~q1 & (h2 & ~f17)))))))) | ((~q & (~p & (~o & (~g2 & (~s1 & (~r1 & (~q1 & (h2 & a)))))))) | ((~q & (~p & (~o & (g2 & (~h1 & (~g1 & (~f1 & (h2 & ~f17)))))))) | ((~q & (~p & (~o & (g2 & (~h1 & (~g1 & (~f1 & (h2 & a)))))))) | ((g2 & (~s1 & (~r1 & (~q1 & (~h1 & (~g1 & (~f1 & (~h2 & a)))))))) | ((~g2 & (~s1 & (~r1 & (~q1 & (~h2 & a))))) | ((~g2 & (~s1 & (~r1 & (~q1 & (o0 & ~f17))))) | ((~g2 & (~s1 & (~r1 & (~q1 & (o0 & a))))) | ((g2 & (~h1 & (~g1 & (~f1 & (o0 & ~f17))))) | ((g2 & (~h1 & (~g1 & (~f1 & (o0 & a))))) | ((~s1 & (~r1 & (~q1 & (~h2 & (~l2 & a))))) | ((~q & (~p & (~o & (h2 & ~l2)))) | (o0 & ~l2)))))))))))),
  u13 = (~c17 & k0) | ((h0 & k0) | ((~j16 & k0) | l2)),
  u14 = ~p17 & (t0 & g0),
  u15 = (~w16 & w2) | ((~v16 & x2) | (~x2 & w2)),
  u16 = (u15 & s0) | ((~b2 & s0) | (s1 & s0)),
  f13 = (l2 & (~e1 & (~d1 & ~c1))) | (~q17 & l2),
  f14 = (q2 & m2) | ((p2 & m2) | (m2 & r0)),
  f15 = ~u15 & ~m1,
  f16 = a16 | z15,
  f17 = (~h2 & (~g2 & f2)) | (h2 & (~g2 & ~f2)),
  n12 = u15 | v2,
  n13 = (s1 & (~r1 & ~f)) | ((s1 & (~r1 & ~e)) | ((s1 & (~r1 & ~d)) | ((b1 & ~f) | ((b1 & ~e) | (b1 & ~d))))),
  n14 = (~y16 & (~i3 & h3)) | ((y16 & i3) | d17),
  n15 = (d4 & (s1 & ~r1)) | ((j17 & (s1 & ~r1)) | (u15 & (s1 & ~r1))),
  n16 = (h17 & ~p12) | (f0 & a),
  n17 = (~q2 & (m2 & (~y1 & (x1 & r0)))) | (~p2 & (m2 & (~y1 & (x1 & r0)))),
  v12 = (h17 & (p12 & ~a)) | (f0 & ~a),
  v13 = (~q16 & (u2 & l0)) | ((f17 & l2) | ((~j16 & l0) | ((~s0 & l0) | z1))),
  v14 = ~z0 & ~y0,
  v15 = ~x0 & ~w0,
  v16 = y1 & (x1 & m2),
  g13 = (l2 & (~e1 & ~d1)) | (~q17 & l2),
  g14 = (~p0 & l17) | (~l17 & v3),
  g15 = o17 | i1,
  g16 = h17 & r1,
  g17 = (c3 & o0) | (b3 & o0),
  o12 = (~s0 & (u2 & (h0 & ~g0))) | ((s0 & (u2 & (u & ~t))) | u15),
  o13 = (~l2 & (h2 & (g2 & ~f2))) | a,
  o14 = (~e16 & (~d16 & z2)) | ((~e16 & (~c16 & z2)) | ((~s0 & (c16 & ~h0)) | ((s0 & (c16 & ~u)) | (~d16 & (c16 & z2))))),
  o15 = (~p3 & r) | ((k3 & r) | (s2 & u0)),
  o16 = ~l3 & (t0 & (h0 & ~g0)),
  o17 = m2 & (y1 & ~x1),
  w12 = (~s0 & (~o12 & (i0 & x15))) | ((s0 & (~o12 & (v & x15))) | ((~b16 & (n2 & ~x15)) | ((b16 & (~n2 & ~x15)) | ((f16 & (y2 & x15)) | ((~n12 & (o12 & x15)) | (n12 & (~o12 & x15))))))),
  w13 = (~i3 & (l2 & (~q & (p & (~o & ~o16))))) | ((h3 & (l2 & (~q & (p & (~o & ~o16))))) | ((p2 & (l2 & (~q & (p & ~o16)))) | ((m2 & (~y1 & (x1 & (~w1 & ~o16)))) | (~o16 & m0)))),
  w14 = ~x0 & ~w0,
  w15 = (~w2 & u15) | (~w2 & ~x2),
  w16 = (~s0 & (u2 & (~h0 & (x2 & (~w2 & (~d0 & ~m)))))) | ((~s0 & (u2 & (~h0 & (x2 & (~w2 & (d0 & ~k)))))) | ((s0 & (u2 & (~u & (x2 & (~w2 & (~d0 & ~m)))))) | ((s0 & (u2 & (~u & (x2 & (~w2 & (d0 & ~k)))))) | ((~s0 & (u2 & (~h0 & (u3 & ~h)))) | ((s0 & (u2 & (~u & (u3 & ~h)))) | ((u3 & ~i) | ((~d0 & ~l) | ((d0 & ~j) | ~g)))))))),
  h13 = (l2 & (~e1 & ~c1)) | (~q17 & l2),
  h14 = (~q0 & (p0 & l17)) | ((q0 & (~p0 & l17)) | (~l17 & w3)),
  h15 = (x15 & u2) | ((~l3 & s) | h16),
  h16 = f16 & (~g16 & (~e17 & g3)),
  h17 = (h2 & (f17 & (o2 & (l2 & (~s1 & (r1 & ~p1)))))) | ((h2 & (f17 & (o2 & (l2 & (s1 & (~r1 & ~p1)))))) | ((f2 & (f17 & (o2 & (l2 & (~s1 & (r1 & ~p1)))))) | ((f2 & (f17 & (o2 & (l2 & (s1 & (~r1 & ~p1)))))) | ((h2 & (o2 & (z1 & (~s1 & (r1 & ~p1))))) | ((h2 & (o2 & (z1 & (s1 & (~r1 & ~p1))))) | ((f2 & (o2 & (z1 & (~s1 & (r1 & ~p1))))) | (f2 & (o2 & (z1 & (s1 & (~r1 & ~p1))))))))))),
  p12 = (~s0 & (u2 & h0)) | ((s0 & (u2 & u)) | (u15 & c2)),
  p13 = (f2 & (~l2 & h2)) | (~l2 & (h2 & ~g2)),
  p14 = (~e16 & (~s0 & (~g16 & (a3 & h0)))) | ((~e16 & (~s0 & (a3 & (z2 & h0)))) | ((~e16 & (s0 & (~g16 & (a3 & u)))) | ((~e16 & (s0 & (a3 & (z2 & u)))) | ((~s0 & (~g16 & (c16 & (a3 & h0)))) | ((~s0 & (c16 & (a3 & (z2 & h0)))) | ((s0 & (~g16 & (c16 & (a3 & u)))) | ((s0 & (c16 & (a3 & (z2 & u)))) | ((~e16 & (~g16 & (~c16 & a3))) | ((~e16 & (~c16 & (a3 & z2))) | ((~s0 & (c16 & (i0 & ~h0))) | ((s0 & (c16 & (v & ~u))) | (d16 & c16)))))))))))),
  p15 = p3 & j3,
  p16 = (~l16 & (k16 & j16)) | (k16 & j0),
  p17 = (u1 & (~z0 & (~y0 & (~x0 & ~w0)))) | ((u1 & (~z0 & (y0 & (~x0 & w0)))) | ((u1 & (z0 & (~y0 & (x0 & ~w0)))) | (u1 & (z0 & (y0 & (x0 & w0)))))),
  x12 = (b16 & (~o2 & (~n2 & ~x15))) | ((a16 & (z15 & (y2 & x15))) | ((~b16 & (o2 & ~x15)) | ((o2 & (n2 & ~x15)) | ((~n12 & (o12 & x15)) | (n12 & (~o12 & x15)))))),
  x13 = p16 & n3,
  x14 = ~z0 & ~y0,
  x15 = ~q16 & m16,
  x16 = ~q & (~p & o),
  a5 = m2,
  a6 = b14,
  a7 = y0,
  a8 = r15,
  b5 = d13,
  b6 = c14,
  b7 = z0,
  b8 = s15,
  c5 = e13,
  c6 = d14,
  c7 = y14,
  c8 = t15,
  d5 = f13,
  d6 = \[50] ,
  d7 = z14,
  d8 = u15,
  e5 = g13,
  e6 = e14,
  e7 = a15,
  e8 = v15,
  f4 = l12,
  f5 = h13,
  f6 = f14,
  f7 = b15,
  f8 = w0,
  g4 = m12,
  g5 = i13,
  g6 = g14,
  g7 = c15,
  a13 = (y15 & (~c & (b & ~x15))) | ((~y15 & (c & ~x15)) | ((c & (~b & ~x15)) | (x15 & e2))),
  g8 = x0,
  a14 = l16 | (u15 | (k2 | i2)),
  a15 = (l3 & (z3 & (y3 & t16))) | (s & (z3 & (y3 & t16))),
  a16 = (~e17 & (m3 & (i3 & ~h3))) | (~e17 & f3),
  a17 = (p17 & j2) | (z16 & j2),
  h4 = n12,
  h5 = j13,
  h6 = h14,
  h7 = d15,
  h8 = w15,
  i4 = o12,
  i5 = k13,
  i6 = i14,
  i7 = e15,
  \[50]  = ~p2,
  j4 = p12,
  j5 = l13,
  j6 = j14,
  j7 = f15,
  i13 = (~q17 & l2) | (l2 & ~e1),
  i14 = p16 & l3,
  i15 = ~h16 & (~s16 & r16),
  i16 = (c17 & (t0 & (j16 & (~l3 & ~h0)))) | ((q16 & (t0 & (j16 & ~l3))) | ((~u2 & (t0 & (j16 & ~l3))) | ((~s0 & (z3 & ~h0)) | ((~s0 & (u15 & ~h0)) | ((s0 & (z3 & ~u)) | ((s0 & (u15 & ~u)) | ((b17 & j16) | ((d16 & ~y16) | ((a17 & ~z16) | ((a17 & ~x16) | (a17 & ~l2))))))))))),
  i17 = q2 & (p2 & (l2 & q)),
  k4 = s3,
  k5 = l2,
  k6 = k14,
  k7 = g15,
  l4 = \[6] ,
  l5 = m13,
  l6 = l14,
  l7 = h15,
  m4 = t3,
  m5 = n13,
  m6 = m14,
  m7 = i15,
  q12 = (o17 & (e1 & (d1 & c1))) | ((v16 & ~w1) | ((o17 & ~n) | n17)),
  q13 = (g2 & l2) | ((g2 & ~h2) | ((f2 & l2) | ((f2 & ~h2) | (~l2 & ~h2)))),
  q14 = (~e16 & (~g17 & b3)) | (e16 & z2),
  q15 = (~d0 & k) | (d0 & m),
  q16 = ~n16 & r2,
  q17 = q & (~p & n),
  n4 = q12,
  n5 = o13,
  n6 = n14,
  n7 = j15,
  o4 = r12,
  o5 = p13,
  o6 = o14,
  o7 = k15,
  p4 = s12,
  p5 = q13,
  p6 = p14,
  p7 = l15,
  y12 = (o2 & (~n16 & m16)) | ((o2 & (~n16 & r2)) | ((n2 & (~n16 & m16)) | ((n2 & (~n16 & r2)) | ((~n16 & (m16 & ~y15)) | (~n16 & (~y15 & r2)))))),
  y13 = (~x16 & k2) | ((~l2 & k2) | b17),
  y14 = (~y3 & (o1 & (~h17 & ~i17))) | ((~y3 & (o1 & (~s1 & ~i17))) | ((~h17 & (~i17 & m1)) | (~s1 & (~i17 & m1)))),
  y15 = (f & (e & (d & a))) | ((~n & a) | ((~s1 & a) | (r1 & a))),
  y16 = (c17 & (~e16 & (~g16 & m3))) | (c17 & (~e16 & (i3 & h3))),
  q4 = t12,
  q5 = r13,
  q6 = q14,
  q7 = m15,
  r4 = u12,
  r5 = s13,
  r6 = r14,
  r7 = n15,
  s4 = v12,
  s5 = t13,
  s6 = s14,
  s7 = w,
  t4 = w12,
  t5 = u13,
  t6 = t14,
  t7 = z,
  u4 = x12,
  u5 = v13,
  u6 = u14,
  u7 = a0,
  v4 = y12,
  v5 = w13,
  v6 = v14,
  v7 = b0,
  w4 = z12,
  w5 = x13,
  w6 = y0,
  w7 = c0,
  b13 = (~x3 & v0) | a,
  b14 = (y & (~\x  & e0)) | ((~y & n0) | (\x  & n0)),
  b15 = (q2 & m2) | ((p2 & m2) | (m2 & m1)),
  b16 = (o2 & y15) | (n2 & y15),
  b17 = p17 & (~l2 & (t0 & g0)),
  x4 = a13,
  x5 = y13,
  x6 = w14,
  x7 = o15,
  y4 = b13,
  y5 = z13,
  y6 = w0,
  y7 = p15;
endmodule

