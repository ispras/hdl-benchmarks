// IWLS benchmark module "dalu" printed on Wed May 29 16:32:29 2002
module dalu(inA15, inA14, inA13, inA12, inA11, inA10, inA9, inA8, inA7, inA6, inA5, inA4, inA3, inA2, inA1, inA0, inB15, inB14, inB13, inB12, inB11, inB10, inB9, inB8, inB7, inB6, inB5, inB4, inB3, inB2, inB1, inB0, inC15, inC14, inC13, inC12, inC11, inC10, inC9, inC8, inC7, inC6, inC5, inC4, inC3, inC2, inC1, inC0, inD15, inD14, inD13, inD12, inD11, inD10, inD9, inD8, inD7, inD6, inD5, inD4, inD3, inD2, inD1, inD0, opsel3, opsel2, opsel1, opsel0, musel4, musel3, musel2, musel1, sh2, sh1, sh0, O15, O14, O13, O12, O11, O10, O9, O8, O7, O6, O5, O4, O3, O2, O1, O0);
input
  inA0,
  inA1,
  inA2,
  inA3,
  inA4,
  inA5,
  inA6,
  inA7,
  inA8,
  inA9,
  inB0,
  inB1,
  inB2,
  inB3,
  inB4,
  inB5,
  inB6,
  inB7,
  inB8,
  inB9,
  inC0,
  inC1,
  inC2,
  inC3,
  inC4,
  inC5,
  inC6,
  inC7,
  inC8,
  inC9,
  inD0,
  inD1,
  inD2,
  inD3,
  inD4,
  inD5,
  inD6,
  inD7,
  inD8,
  inD9,
  inA10,
  inA11,
  inA12,
  inA13,
  inA14,
  inA15,
  inB10,
  inB11,
  inB12,
  inB13,
  inB14,
  inB15,
  inC10,
  inC11,
  inC12,
  inC13,
  inC14,
  inC15,
  inD10,
  inD11,
  inD12,
  inD13,
  inD14,
  inD15,
  musel1,
  musel2,
  musel3,
  musel4,
  sh0,
  sh1,
  sh2,
  opsel0,
  opsel1,
  opsel2,
  opsel3;
output
  O10,
  O11,
  O12,
  O13,
  O14,
  O15,
  O0,
  O1,
  O2,
  O3,
  O4,
  O5,
  O6,
  O7,
  O8,
  O9;
wire
  \[60] ,
  \[61] ,
  \[5928] ,
  \[8586] ,
  \[5542] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[8491] ,
  \[66] ,
  \[67] ,
  \[5835] ,
  \[69] ,
  \[8418] ,
  \[9529] ,
  \[6082] ,
  \[5645] ,
  \[9337] ,
  \[0] ,
  \[5933] ,
  \[5740] ,
  \[1] ,
  \[6008] ,
  \[9433] ,
  \[2] ,
  \[3] ,
  \[1478] ,
  \[4] ,
  \[5] ,
  \[71] ,
  \[6105] ,
  \[6] ,
  \[72] ,
  \[5840] ,
  \[7] ,
  \[73] ,
  \[1382] ,
  \[5554] ,
  \[8] ,
  \[74] ,
  \[5748] ,
  \[1400] ,
  \[5555] ,
  \[9] ,
  \[75] ,
  \[76] ,
  \[1115] ,
  \[8905] ,
  \[5844] ,
  \[77] ,
  \[8520] ,
  \[78] ,
  \[5653] ,
  \[5849] ,
  \[1502] ,
  \[6094] ,
  \[1580] ,
  \[6114] ,
  \[8335] ,
  \[82] ,
  \[5563] ,
  \[83] ,
  \[9449] ,
  \[84] ,
  \[5758] ,
  \[85] ,
  \[9545] ,
  \[5854] ,
  \[9353] ,
  \[88] ,
  \[8917] ,
  \[5663] ,
  \[89] ,
  \[5950] ,
  \[5859] ,
  \[9932] ,
  \[10] ,
  e10,
  e14,
  \[11] ,
  \[12] ,
  \[12790] ,
  \[13] ,
  \[1592] ,
  \[5957] ,
  \[14] ,
  \[8440] ,
  \[15] ,
  \[5573] ,
  \[17] ,
  \[19] ,
  \[467] ,
  \[96] ,
  \[5671] ,
  \[97] ,
  \[1616] ,
  \[5865] ,
  \[8540] ,
  \[98] ,
  \[1424] ,
  \[8929] ,
  \[102] ,
  \[1520] ,
  \[103] ,
  \[104] ,
  \[20] ,
  \[5771] ,
  \[9369] ,
  \[105] ,
  \[6038] ,
  \[21] ,
  \[106] ,
  \[6039] ,
  \[950] ,
  \[107] ,
  \[9465] ,
  \[23] ,
  \[1332] ,
  \[5967] ,
  \[5581] ,
  \[24] ,
  \[25] ,
  \[9561] ,
  \[5870] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[5681] ,
  \[5875] ,
  \[8263] ,
  \[8360] ,
  \[5609] ,
  \[30] ,
  \[5704] ,
  \[5781] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[5591] ,
  \[34] ,
  \[1630] ,
  \[35] ,
  \[8941] ,
  \[36] ,
  \[1538] ,
  \[484] ,
  \[5881] ,
  \[37] ,
  \[38] ,
  \[5789] ,
  \[8464] ,
  \[39] ,
  \[1442] ,
  \[5807] ,
  \[1349] ,
  \[6052] ,
  \[9577] ,
  \[5599] ,
  \[9401] ,
  \[5886] ,
  \[9385] ,
  \[5617] ,
  \[5904] ,
  \[5694] ,
  \[8562] ,
  \[5712] ,
  \[9674] ,
  \[9481] ,
  \[40] ,
  \[41] ,
  \[9677] ,
  \[42] ,
  \[5909] ,
  \[8181] ,
  \[43] ,
  \[44] ,
  \[5988] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[9776] ,
  \[782] ,
  \[48] ,
  \[5799] ,
  \[5893] ,
  \[49] ,
  \[5817] ,
  \[9779] ,
  e2,
  e6,
  e9,
  \[6063] ,
  \[5627] ,
  \[5898] ,
  \[8286] ,
  \[5722] ,
  \[5993] ,
  \[50] ,
  \[5917] ,
  \[5994] ,
  \[9417] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[1556] ,
  \[9513] ,
  \[5998] ,
  pgx3,
  \[9497] ,
  \[55] ,
  \[1364] ,
  \[56] ,
  \[8388] ,
  \[57] ,
  \[1460] ,
  \[5825] ,
  \[58] ,
  \[59] ,
  \[9883] ,
  \[5635] ,
  \[5922] ,
  \[5730] ,
  \[8313] ;
assign
  \[60]  = \[57]  & ~sh1,
  \[61]  = 0,
  \[5928]  = (\[45]  & \[9561] ) | (~\[9561]  & ~\[5849] ),
  \[8586]  = (\[38]  & inB1) | (\[21]  & inD1),
  \[5542]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA15))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC15))) | ((~\[42]  & (~musel2 & (~inB15 & ~inA15))) | ((~\[42]  & (musel2 & (~inC15 & ~inB15))) | ((~\[40]  & (~musel2 & (~inD15 & ~inA15))) | ((~\[40]  & (musel2 & (~inD15 & ~inC15))) | ((~musel2 & (~inD15 & (~inB15 & ~inA15))) | ((musel2 & (~inD15 & (~inC15 & ~inB15))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB15)) | ((~\[40]  & (\[30]  & ~inD15)) | ((\[30]  & (~inD15 & ~inB15)) | musel4))))))))))),
  \[62]  = 0,
  \[63]  = 0,
  \[64]  = ~\[5933]  | \[5849] ,
  \[65]  = ~pgx3 | ~\[5865] ,
  \[8491]  = (\[38]  & inB5) | (\[21]  & inD5),
  \[66]  = \[5998] ,
  \[67]  = ~\[12790]  | ~\[5886] ,
  \[5835]  = (\[43]  & inC0) | \[1364] ,
  \[69]  = \[5663]  | ~\[5653] ,
  \[8418]  = (\[38]  & inB8) | (\[21]  & inD8),
  \[9529]  = (\[34]  & inA3) | (\[27]  & inC3),
  \[6082]  = \[5781]  | ~\[5771] ,
  \[5645]  = (\[43]  & inC10) | \[1556] ,
  \[9337]  = (\[34]  & inA15) | (\[27]  & inC15),
  \[0]  = (\[31]  & (~\[8905]  & \[5854] )) | ((\[29]  & \[5555] ) | \[83] ),
  \[5933]  = (\[45]  & \[9577] ) | (~\[9577]  & ~\[5849] ),
  \[5740]  = (\[43]  & inC5) | \[1460] ,
  \[1]  = (\[85]  & \[8263] ) | ((\[83]  & \[5950] ) | ((\[31]  & \[8905] ) | (\[29]  & ~e14))),
  \[6008]  = \[5645]  | ~\[5635] ,
  \[9433]  = (\[34]  & inA9) | (\[27]  & inC9),
  \[2]  = (~\[107]  & (~\[85]  & \[83] )) | ((\[96]  & (~\[65]  & \[31] )) | ((\[96]  & (\[31]  & \[5859] )) | ((\[107]  & \[8263] ) | ((\[85]  & \[8286] ) | (\[29]  & \[5967] ))))),
  \[3]  = (~\[106]  & (~\[105]  & (~\[104]  & (\[20]  & \[8181] )))) | ((\[65]  & (\[31]  & pgx3)) | ((\[65]  & (\[31]  & \[5865] )) | ((\[106]  & \[8286] ) | ((\[105]  & \[8313] ) | ((\[104]  & \[8263] ) | ((\[36]  & \[24] ) | (\[24]  & \[5609] ))))))),
  \[1478]  = (\[35]  & (~\[9481]  & inC6)) | ((\[39]  & \[9481] ) | (\[37]  & inA6)),
  \[4]  = (\[88]  & (\[31]  & \[5893] )) | ((\[55]  & (\[17]  & \[8263] )) | ((\[54]  & (\[17]  & \[8286] )) | ((\[53]  & (\[17]  & \[8313] )) | ((\[50]  & (\[17]  & \[8181] )) | ((\[17]  & (\[8335]  & ~\[5950] )) | (\[29]  & \[5993] )))))),
  \[5]  = (\[60]  & (\[17]  & \[8263] )) | ((\[58]  & (\[17]  & \[8181] )) | ((\[55]  & (\[17]  & \[8286] )) | ((\[54]  & (\[17]  & \[8313] )) | ((\[53]  & (\[17]  & \[8335] )) | ((\[17]  & (\[8360]  & ~\[5950] )) | ((\[84]  & \[17] ) | ((\[31]  & \[8917] ) | (\[29]  & ~e10)))))))),
  \[71]  = 0,
  \[6105]  = \[5817]  | ~\[5807] ,
  \[6]  = (\[66]  & (\[31]  & \[5904] )) | ((\[60]  & (\[17]  & \[8286] )) | ((\[58]  & (\[17]  & \[8263] )) | ((\[55]  & (\[17]  & \[8313] )) | ((\[54]  & (\[17]  & \[8335] )) | ((\[107]  & \[8360] ) | ((\[85]  & \[8388] ) | ((\[84]  & \[17] ) | (\[29]  & ~e9)))))))),
  \[72]  = 0,
  \[5840]  = 0,
  \[7]  = (\[60]  & (\[20]  & \[8313] )) | ((\[58]  & (\[20]  & \[8286] )) | ((\[55]  & (\[20]  & \[8335] )) | ((\[31]  & (\[5998]  & \[5909] )) | ((\[106]  & \[8388] ) | ((\[105]  & \[8418] ) | ((\[104]  & \[8360] ) | ((\[84]  & \[20] ) | (~\[77]  & \[24] )))))))),
  \[73]  = ~opsel2 | opsel3,
  \[1382]  = (\[35]  & (~\[9561]  & inC1)) | ((\[39]  & \[9561] ) | (\[37]  & inA1)),
  \[5554]  = (\[43]  & inC15) | \[1630] ,
  \[8]  = (~\[89]  & (\[31]  & ~\[5870] )) | ((\[89]  & (\[31]  & \[5870] )) | ((\[60]  & (\[17]  & \[8335] )) | ((\[58]  & (\[17]  & \[8313] )) | ((\[55]  & (\[17]  & \[8360] )) | ((\[54]  & (\[17]  & \[8388] )) | ((\[53]  & (\[17]  & \[8418] )) | ((\[17]  & (\[8440]  & ~\[5950] )) | ((\[84]  & \[17] ) | (\[29]  & \[6038] ))))))))),
  \[74]  = 0,
  \[5748]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA4))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC4))) | ((~\[42]  & (~musel2 & (~inB4 & ~inA4))) | ((~\[42]  & (musel2 & (~inC4 & ~inB4))) | ((~\[40]  & (~musel2 & (~inD4 & ~inA4))) | ((~\[40]  & (musel2 & (~inD4 & ~inC4))) | ((~musel2 & (~inD4 & (~inB4 & ~inA4))) | ((musel2 & (~inD4 & (~inC4 & ~inB4))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB4)) | ((~\[40]  & (\[30]  & ~inD4)) | ((\[30]  & (~inD4 & ~inB4)) | musel4))))))))))),
  \[1400]  = (\[35]  & (~\[9545]  & inC2)) | ((\[39]  & \[9545] ) | (\[37]  & inA2)),
  \[5555]  = \[5554]  | ~\[5542] ,
  \[9]  = (\[60]  & (\[17]  & \[8360] )) | ((\[59]  & (\[17]  & \[8263] )) | ((\[58]  & (\[17]  & \[8335] )) | ((\[55]  & (\[17]  & \[8388] )) | ((\[54]  & (\[17]  & \[8418] )) | ((\[107]  & \[8440] ) | ((\[85]  & \[8464] ) | ((\[31]  & \[8929] ) | (\[29]  & ~e6)))))))),
  \[75]  = 0,
  \[76]  = ~\[9677] ,
  \[1115]  = 0,
  \[8905]  = (~\[96]  & ~\[5854] ) | (\[96]  & \[5854] ),
  \[5844]  = 0,
  \[77]  = ~\[9883] ,
  \[8520]  = (\[38]  & inB4) | (\[21]  & inD4),
  \[78]  = ~\[9779] ,
  \[5653]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA9))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC9))) | ((~\[42]  & (~musel2 & (~inB9 & ~inA9))) | ((~\[42]  & (musel2 & (~inC9 & ~inB9))) | ((~\[40]  & (~musel2 & (~inD9 & ~inA9))) | ((~\[40]  & (musel2 & (~inD9 & ~inC9))) | ((~musel2 & (~inD9 & (~inB9 & ~inA9))) | ((musel2 & (~inD9 & (~inC9 & ~inB9))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB9)) | ((~\[40]  & (\[30]  & ~inD9)) | ((\[30]  & (~inD9 & ~inB9)) | musel4))))))))))),
  \[5849]  = \[19]  | ~\[9337] ,
  \[1502]  = (\[35]  & (~\[9465]  & inC7)) | ((\[39]  & \[9465] ) | (\[37]  & inA7)),
  \[6094]  = \[5799]  | ~\[5789] ,
  \[1580]  = (\[35]  & (~\[9401]  & inC11)) | ((\[39]  & \[9401] ) | (\[37]  & inA11)),
  \[6114]  = opsel0 | opsel1,
  \[8335]  = (\[38]  & inB11) | (\[21]  & inD11),
  \[82]  = \[64]  | ~\[5928] ,
  \[5563]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA14))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC14))) | ((~\[42]  & (~musel2 & (~inB14 & ~inA14))) | ((~\[42]  & (musel2 & (~inC14 & ~inB14))) | ((~\[40]  & (~musel2 & (~inD14 & ~inA14))) | ((~\[40]  & (musel2 & (~inD14 & ~inC14))) | ((~musel2 & (~inD14 & (~inB14 & ~inA14))) | ((musel2 & (~inD14 & (~inC14 & ~inB14))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB14)) | ((~\[40]  & (\[30]  & ~inD14)) | ((\[30]  & (~inD14 & ~inB14)) | musel4))))))))))),
  \[83]  = \[17]  & \[8181] ,
  \[9449]  = (\[34]  & inA8) | (\[27]  & inC8),
  \[84]  = \[59]  & \[8181] ,
  \[5758]  = (\[43]  & inC4) | \[1442] ,
  \[85]  = \[17]  & ~\[5950] ,
  \[9545]  = (\[34]  & inA2) | (\[27]  & inC2),
  \[5854]  = (\[45]  & \[9353] ) | (~\[5849]  & ~\[9353] ),
  \[9353]  = (\[34]  & inA14) | (\[27]  & inC14),
  \[88]  = \[8917]  | ~\[5898] ,
  \[8917]  = \[97]  & \[5898] ,
  \[5663]  = (\[43]  & inC9) | \[1538] ,
  \[89]  = \[8929]  | ~\[5875] ,
  \[5950]  = (sh0 & ~sh1) | (\[57]  | \[52] ),
  \[5859]  = (\[45]  & \[9369] ) | (~\[9369]  & ~\[5849] ),
  \[9932]  = 0,
  \[10]  = (~\[67]  & (\[31]  & ~\[5881] )) | ((\[67]  & (\[31]  & \[5881] )) | ((\[60]  & (\[17]  & \[8388] )) | ((\[59]  & (\[17]  & \[8286] )) | ((\[58]  & (\[17]  & \[8360] )) | ((\[55]  & (\[17]  & \[8418] )) | ((\[54]  & (\[17]  & \[8440] )) | ((\[107]  & \[8464] ) | ((\[85]  & \[8491] ) | (\[29]  & \[6063] ))))))))),
  e10 = ~\[6008] ,
  e14 = \[33] ,
  \[11]  = (\[60]  & (\[20]  & \[8418] )) | ((\[59]  & (\[20]  & \[8313] )) | ((\[58]  & (\[20]  & \[8388] )) | ((\[55]  & (\[20]  & \[8440] )) | ((\[31]  & (~\[12790]  & \[5886] )) | ((\[31]  & (\[12790]  & ~\[5886] )) | ((\[106]  & \[8491] ) | ((\[105]  & \[8520] ) | ((\[104]  & \[8464] ) | (~\[78]  & \[24] ))))))))),
  \[12]  = (\[31]  & (~\[8941]  & (~\[12790]  & \[5922] ))) | ((\[60]  & (\[17]  & \[8440] )) | ((\[59]  & (\[17]  & \[8335] )) | ((\[58]  & (\[17]  & \[8418] )) | ((\[55]  & (\[17]  & \[8464] )) | ((\[54]  & (\[17]  & \[8491] )) | ((\[53]  & (\[17]  & \[8520] )) | ((\[31]  & (~\[12790]  & \[5917] )) | ((\[17]  & (\[8540]  & ~\[5950] )) | (\[29]  & \[6082] ))))))))),
  \[12790]  = ~\[82]  & (\[5922]  & \[5917] ),
  \[13]  = (\[60]  & (\[17]  & \[8464] )) | ((\[59]  & (\[17]  & \[8360] )) | ((\[58]  & (\[17]  & \[8440] )) | ((\[55]  & (\[17]  & \[8491] )) | ((\[54]  & (\[17]  & \[8520] )) | ((\[107]  & \[8540] ) | ((\[85]  & \[8562] ) | ((\[31]  & \[8941] ) | (\[29]  & ~e2)))))))),
  \[1592]  = (\[35]  & (~\[9369]  & inC13)) | ((\[39]  & \[9369] ) | (\[37]  & inA13)),
  \[5957]  = ~sh0 | ~sh2,
  \[14]  = (~\[64]  & (\[31]  & ~\[5928] )) | ((\[64]  & (\[31]  & \[5928] )) | ((\[60]  & (\[17]  & \[8491] )) | ((\[59]  & (\[17]  & \[8388] )) | ((\[58]  & (\[17]  & \[8464] )) | ((\[55]  & (\[17]  & \[8520] )) | ((\[54]  & (\[17]  & \[8540] )) | ((\[107]  & \[8562] ) | ((\[85]  & \[8586] ) | (\[29]  & \[6105] ))))))))),
  \[8440]  = (\[38]  & inB7) | (\[21]  & inD7),
  \[15]  = (\[85]  & (\[38]  & inB0)) | ((\[85]  & (\[21]  & inD0)) | ((\[64]  & (\[31]  & \[5933] )) | ((\[64]  & (\[31]  & ~\[5849] )) | ((\[60]  & (\[17]  & \[8520] )) | ((\[59]  & (\[17]  & \[8418] )) | ((\[58]  & (\[17]  & \[8491] )) | ((\[55]  & (\[17]  & \[8540] )) | ((\[54]  & (\[17]  & \[8562] )) | ((\[107]  & \[8586] ) | (~\[76]  & \[29] )))))))))),
  \[5573]  = (\[43]  & inC14) | \[1616] ,
  \[17]  = (~\[6114]  & \[1349] ) | \[102] ,
  \[19]  = musel3 | ~musel4,
  \[467]  = \[17] ,
  \[96]  = \[65]  | ~\[5859] ,
  \[5671]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA8))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC8))) | ((~\[42]  & (~musel2 & (~inB8 & ~inA8))) | ((~\[42]  & (musel2 & (~inC8 & ~inB8))) | ((~\[40]  & (~musel2 & (~inD8 & ~inA8))) | ((~\[40]  & (musel2 & (~inD8 & ~inC8))) | ((~musel2 & (~inD8 & (~inB8 & ~inA8))) | ((musel2 & (~inD8 & (~inC8 & ~inB8))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB8)) | ((~\[40]  & (\[30]  & ~inD8)) | ((\[30]  & (~inD8 & ~inB8)) | musel4))))))))))),
  \[97]  = \[66] ,
  \[1616]  = (\[35]  & (~\[9353]  & inC14)) | ((\[39]  & \[9353] ) | (\[37]  & inA14)),
  \[5865]  = (\[45]  & \[9385] ) | (~\[9385]  & ~\[5849] ),
  \[8540]  = (\[38]  & inB3) | (\[21]  & inD3),
  \[98]  = \[67]  | ~\[5881] ,
  \[1424]  = (\[35]  & (~\[9529]  & inC3)) | ((\[39]  & \[9529] ) | (\[37]  & inA3)),
  \[8929]  = (~\[98]  & ~\[5875] ) | (\[98]  & \[5875] ),
  \[102]  = ~\[73]  & \[6114] ,
  \[1520]  = (\[35]  & (~\[9449]  & inC8)) | ((\[39]  & \[9449] ) | (\[37]  & inA8)),
  \[103]  = ~opsel2 & opsel3,
  \[104]  = \[54]  & \[20] ,
  \[20]  = \[102]  | \[467] ,
  \[5771]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA3))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC3))) | ((~\[42]  & (~musel2 & (~inB3 & ~inA3))) | ((~\[42]  & (musel2 & (~inC3 & ~inB3))) | ((~\[40]  & (~musel2 & (~inD3 & ~inA3))) | ((~\[40]  & (musel2 & (~inD3 & ~inC3))) | ((~musel2 & (~inD3 & (~inB3 & ~inA3))) | ((musel2 & (~inD3 & (~inC3 & ~inB3))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB3)) | ((~\[40]  & (\[30]  & ~inD3)) | ((\[30]  & (~inD3 & ~inB3)) | musel4))))))))))),
  \[9369]  = (\[34]  & inA13) | (\[27]  & inC13),
  \[105]  = \[20]  & ~\[5950] ,
  \[6038]  = \[5704]  | ~\[5694] ,
  \[21]  = (\[35]  & musel1) | ~\[25] ,
  \[106]  = \[53]  & \[20] ,
  \[6039]  = 0,
  \[950]  = 0,
  \[107]  = \[53]  & \[17] ,
  \[9465]  = (\[34]  & inA7) | (\[27]  & inC7),
  \[23]  = musel1 | musel2,
  \[1332]  = (\[35]  & (~\[9385]  & inC12)) | ((\[39]  & \[9385] ) | (\[37]  & inA12)),
  \[5967]  = ~\[5581]  | \[5591] ,
  \[5581]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA13))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC13))) | ((~\[42]  & (~musel2 & (~inB13 & ~inA13))) | ((~\[42]  & (musel2 & (~inC13 & ~inB13))) | ((~\[40]  & (~musel2 & (~inD13 & ~inA13))) | ((~\[40]  & (musel2 & (~inD13 & ~inC13))) | ((~musel2 & (~inD13 & (~inB13 & ~inA13))) | ((musel2 & (~inD13 & (~inC13 & ~inB13))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB13)) | ((~\[40]  & (\[30]  & ~inD13)) | ((\[30]  & (~inD13 & ~inB13)) | musel4))))))))))),
  \[24]  = \[29] ,
  \[25]  = \[23]  | \[19] ,
  \[9561]  = (\[34]  & inA1) | (\[27]  & inC1),
  \[5870]  = (\[45]  & \[9465] ) | (~\[9465]  & ~\[5849] ),
  \[26]  = musel3 & ~musel4,
  O10 = \[5] ,
  O11 = \[4] ,
  O12 = \[3] ,
  \[27]  = ~musel1 & musel2,
  O13 = \[2] ,
  O14 = \[1] ,
  O15 = \[0] ,
  \[28]  = ~\[5563]  | \[5573] ,
  \[29]  = (\[103]  & (\[6114]  & ~opsel0)) | (\[6114]  & \[1349] ),
  \[5681]  = (\[43]  & inC8) | \[1520] ,
  \[5875]  = (\[45]  & \[9481] ) | (~\[9481]  & ~\[5849] ),
  \[8263]  = (\[38]  & inB14) | (\[21]  & inD14),
  \[8360]  = (\[38]  & inB10) | (\[21]  & inD10),
  \[5609]  = (\[43]  & inC12) | \[1332] ,
  \[30]  = ~musel1 | musel3,
  \[5704]  = (\[43]  & inC7) | \[1502] ,
  \[5781]  = (\[43]  & inC3) | \[1424] ,
  \[31]  = (\[6114]  & (~opsel2 & ~opsel3)) | (~\[73]  & ~\[6114] ),
  \[32]  = 0,
  \[33]  = ~\[28] ,
  \[5591]  = (\[43]  & inC13) | \[1592] ,
  \[34]  = musel1 & ~musel2,
  \[1630]  = (\[35]  & (~\[9337]  & inC15)) | ((\[39]  & \[9337] ) | (\[37]  & inA15)),
  O0 = \[15] ,
  \[35]  = \[26]  & musel2,
  O1 = \[14] ,
  O2 = \[13] ,
  O3 = \[12] ,
  O4 = \[11] ,
  O5 = \[10] ,
  O6 = \[9] ,
  O7 = \[8] ,
  O8 = \[7] ,
  O9 = \[6] ,
  \[8941]  = (~\[82]  & ~\[5922] ) | (\[82]  & \[5922] ),
  \[36]  = ~\[5599] ,
  \[1538]  = (\[35]  & (~\[9433]  & inC9)) | ((\[39]  & \[9433] ) | (\[37]  & inA9)),
  \[484]  = 0,
  \[5881]  = (\[45]  & \[9497] ) | (~\[9497]  & ~\[5849] ),
  \[37]  = \[27]  & \[26] ,
  \[38]  = (\[34]  & \[26] ) | \[37] ,
  \[5789]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA2))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC2))) | ((~\[42]  & (~musel2 & (~inB2 & ~inA2))) | ((~\[42]  & (musel2 & (~inC2 & ~inB2))) | ((~\[40]  & (~musel2 & (~inD2 & ~inA2))) | ((~\[40]  & (musel2 & (~inD2 & ~inC2))) | ((~musel2 & (~inD2 & (~inB2 & ~inA2))) | ((musel2 & (~inD2 & (~inC2 & ~inB2))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB2)) | ((~\[40]  & (\[30]  & ~inD2)) | ((\[30]  & (~inD2 & ~inB2)) | musel4))))))))))),
  \[8464]  = (\[38]  & inB6) | (\[21]  & inD6),
  \[39]  = \[26]  & musel1,
  \[1442]  = (\[35]  & (~\[9513]  & inC4)) | ((\[39]  & \[9513] ) | (\[37]  & inA4)),
  \[5807]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA1))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC1))) | ((~\[42]  & (~musel2 & (~inB1 & ~inA1))) | ((~\[42]  & (musel2 & (~inC1 & ~inB1))) | ((~\[40]  & (~musel2 & (~inD1 & ~inA1))) | ((~\[40]  & (musel2 & (~inD1 & ~inC1))) | ((~musel2 & (~inD1 & (~inB1 & ~inA1))) | ((musel2 & (~inD1 & (~inC1 & ~inB1))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB1)) | ((~\[40]  & (\[30]  & ~inD1)) | ((\[30]  & (~inD1 & ~inB1)) | musel4))))))))))),
  \[1349]  = \[103]  & ~opsel1,
  \[6052]  = \[5722]  | ~\[5712] ,
  \[9577]  = (\[34]  & inA0) | (\[27]  & inC0),
  \[5599]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA12))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC12))) | ((~\[42]  & (~musel2 & (~inB12 & ~inA12))) | ((~\[42]  & (musel2 & (~inC12 & ~inB12))) | ((~\[40]  & (~musel2 & (~inD12 & ~inA12))) | ((~\[40]  & (musel2 & (~inD12 & ~inC12))) | ((~musel2 & (~inD12 & (~inB12 & ~inA12))) | ((musel2 & (~inD12 & (~inC12 & ~inB12))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB12)) | ((~\[40]  & (\[30]  & ~inD12)) | ((\[30]  & (~inD12 & ~inB12)) | musel4))))))))))),
  \[9401]  = (\[34]  & inA11) | (\[27]  & inC11),
  \[5886]  = (\[45]  & \[9513] ) | (~\[9513]  & ~\[5849] ),
  \[9385]  = (\[34]  & inA12) | (\[27]  & inC12),
  \[5617]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA11))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC11))) | ((~\[42]  & (~musel2 & (~inB11 & ~inA11))) | ((~\[42]  & (musel2 & (~inC11 & ~inB11))) | ((~\[40]  & (~musel2 & (~inD11 & ~inA11))) | ((~\[40]  & (musel2 & (~inD11 & ~inC11))) | ((~musel2 & (~inD11 & (~inB11 & ~inA11))) | ((musel2 & (~inD11 & (~inC11 & ~inB11))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB11)) | ((~\[40]  & (\[30]  & ~inD11)) | ((\[30]  & (~inD11 & ~inB11)) | musel4))))))))))),
  \[5904]  = (\[45]  & \[9433] ) | (~\[9433]  & ~\[5849] ),
  \[5694]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA7))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC7))) | ((~\[42]  & (~musel2 & (~inB7 & ~inA7))) | ((~\[42]  & (musel2 & (~inC7 & ~inB7))) | ((~\[40]  & (~musel2 & (~inD7 & ~inA7))) | ((~\[40]  & (musel2 & (~inD7 & ~inC7))) | ((~musel2 & (~inD7 & (~inB7 & ~inA7))) | ((musel2 & (~inD7 & (~inC7 & ~inB7))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB7)) | ((~\[40]  & (\[30]  & ~inD7)) | ((\[30]  & (~inD7 & ~inB7)) | musel4))))))))))),
  \[8562]  = (\[38]  & inB2) | (\[21]  & inD2),
  \[5712]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA6))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC6))) | ((~\[42]  & (~musel2 & (~inB6 & ~inA6))) | ((~\[42]  & (musel2 & (~inC6 & ~inB6))) | ((~\[40]  & (~musel2 & (~inD6 & ~inA6))) | ((~\[40]  & (musel2 & (~inD6 & ~inC6))) | ((~musel2 & (~inD6 & (~inB6 & ~inA6))) | ((musel2 & (~inD6 & (~inC6 & ~inB6))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB6)) | ((~\[40]  & (\[30]  & ~inD6)) | ((\[30]  & (~inD6 & ~inB6)) | musel4))))))))))),
  \[9674]  = 0,
  \[9481]  = (\[34]  & inA6) | (\[27]  & inC6),
  \[40]  = \[27]  & ~musel3,
  \[41]  = 0,
  \[9677]  = \[5835]  | ~\[5825] ,
  \[42]  = ~\[23]  & musel3,
  \[5909]  = (\[45]  & \[9449] ) | (~\[9449]  & ~\[5849] ),
  \[8181]  = (\[38]  & inB15) | (\[21]  & inD15),
  \[43]  = ~\[25] ,
  \[44]  = 0,
  \[5988]  = ~sh0 | ~sh1,
  \[45]  = ~\[19]  & \[5849] ,
  \[46]  = 0,
  \[47]  = 0,
  \[9776]  = 0,
  \[782]  = 0,
  \[48]  = 0,
  \[5799]  = (\[43]  & inC2) | \[1400] ,
  \[5893]  = (\[45]  & \[9401] ) | (~\[9401]  & ~\[5849] ),
  \[49]  = 0,
  \[5817]  = (\[43]  & inC1) | \[1382] ,
  \[9779]  = \[5758]  | ~\[5748] ,
  e2 = ~\[6094] ,
  e6 = ~\[6052] ,
  e9 = ~\[69] ,
  \[6063]  = \[5740]  | ~\[5730] ,
  \[5627]  = (\[43]  & inC11) | \[1580] ,
  \[5898]  = (\[45]  & \[9417] ) | (~\[9417]  & ~\[5849] ),
  \[8286]  = (\[38]  & inB13) | (\[21]  & inD13),
  \[5722]  = (\[43]  & inC6) | \[1478] ,
  \[5993]  = \[5627]  | ~\[5617] ,
  \[50]  = \[5988]  & sh2,
  \[5917]  = (\[45]  & \[9529] ) | (~\[9529]  & ~\[5849] ),
  \[5994]  = 0,
  \[9417]  = (\[34]  & inA10) | (\[27]  & inC10),
  \[52]  = sh1 & ~sh2,
  \[53]  = \[5950]  & (~sh1 & ~sh2),
  \[54]  = \[52]  & ~sh0,
  \[1556]  = (\[35]  & (~\[9417]  & inC10)) | ((\[39]  & \[9417] ) | (\[37]  & inA10)),
  \[9513]  = (\[34]  & inA4) | (\[27]  & inC4),
  \[5998]  = ~\[12790]  | (~\[5909]  | (~\[5904]  | (~\[5898]  | ~\[5893] ))),
  pgx3 = ~\[5998]  & (\[5886]  & (\[5881]  & (\[5875]  & \[5870] ))),
  \[9497]  = (\[34]  & inA5) | (\[27]  & inC5),
  \[55]  = ~\[5988]  & \[5950] ,
  \[1364]  = (\[35]  & (~\[9577]  & inC0)) | ((\[39]  & \[9577] ) | (\[37]  & inA0)),
  \[56]  = 0,
  \[8388]  = (\[38]  & inB9) | (\[21]  & inD9),
  \[57]  = ~sh0 & sh2,
  \[1460]  = (\[35]  & (~\[9497]  & inC5)) | ((\[39]  & \[9497] ) | (\[37]  & inA5)),
  \[5825]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA0))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC0))) | ((~\[42]  & (~musel2 & (~inB0 & ~inA0))) | ((~\[42]  & (musel2 & (~inC0 & ~inB0))) | ((~\[40]  & (~musel2 & (~inD0 & ~inA0))) | ((~\[40]  & (musel2 & (~inD0 & ~inC0))) | ((~musel2 & (~inD0 & (~inB0 & ~inA0))) | ((musel2 & (~inD0 & (~inC0 & ~inB0))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB0)) | ((~\[40]  & (\[30]  & ~inD0)) | ((\[30]  & (~inD0 & ~inB0)) | musel4))))))))))),
  \[58]  = ~\[5957]  & \[5950] ,
  \[59]  = \[50]  & sh1,
  \[9883]  = \[5681]  | ~\[5671] ,
  \[5635]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA10))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC10))) | ((~\[42]  & (~musel2 & (~inB10 & ~inA10))) | ((~\[42]  & (musel2 & (~inC10 & ~inB10))) | ((~\[40]  & (~musel2 & (~inD10 & ~inA10))) | ((~\[40]  & (musel2 & (~inD10 & ~inC10))) | ((~musel2 & (~inD10 & (~inB10 & ~inA10))) | ((musel2 & (~inD10 & (~inC10 & ~inB10))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB10)) | ((~\[40]  & (\[30]  & ~inD10)) | ((\[30]  & (~inD10 & ~inB10)) | musel4))))))))))),
  \[5922]  = (\[45]  & \[9545] ) | (~\[9545]  & ~\[5849] ),
  \[5730]  = (~\[42]  & (~\[40]  & (~musel2 & ~inA5))) | ((~\[42]  & (~\[40]  & (musel2 & ~inC5))) | ((~\[42]  & (~musel2 & (~inB5 & ~inA5))) | ((~\[42]  & (musel2 & (~inC5 & ~inB5))) | ((~\[40]  & (~musel2 & (~inD5 & ~inA5))) | ((~\[40]  & (musel2 & (~inD5 & ~inC5))) | ((~musel2 & (~inD5 & (~inB5 & ~inA5))) | ((musel2 & (~inD5 & (~inC5 & ~inB5))) | ((~\[42]  & (~\[40]  & \[30] )) | ((~\[42]  & (\[30]  & ~inB5)) | ((~\[40]  & (\[30]  & ~inD5)) | ((\[30]  & (~inD5 & ~inB5)) | musel4))))))))))),
  \[8313]  = (\[38]  & inB12) | (\[21]  & inD12);
endmodule

