module reduce_and_1(a, b);
  input a;
  output b;
  assign b = &a;
endmodule
