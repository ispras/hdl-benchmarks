//NOTE: no-implementation module stub

module XSCIOM5 (
    inout wire IO,
    input wire I,
    input wire E,
    output wire O,
    input wire FEB
);
endmodule

module XC (
    output wire O,
    input wire I
);
endmodule

module XCU8 (
    output wire O,
    input wire I
);
endmodule

module XCD8 (
    output wire O,
    input wire I
);
endmodule

module INV1 (
    output wire O,
    input wire I
);
endmodule

module AN2P (
    output wire O,
    input wire I1,
    input wire I2
);
endmodule

module BUF4 (
    output wire O,
    input wire I
);
endmodule

module YC04T (
    output wire O,
    input wire I,
    input wire E
);
endmodule

module YC04A (
    output wire O,
    input wire I,
    input wire E
);
endmodule

module OR2P (
    output wire O,
    input wire I1,
    input wire I2
);
endmodule

module AO12P (
    output wire O,
    input wire A1,
    input wire B1,
    input wire B2
);
endmodule

module ZCC04A (
    inout wire IO,
    output wire O,
    input wire I,
    input wire E
);
endmodule

module INV2 (
    output wire O,
    input wire I
);
endmodule
