// IWLS benchmark module "vda" printed on Wed May 29 17:30:36 2002
module vda(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q;
output
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  a1,
  b0,
  b1,
  c0,
  c1,
  d0,
  d1,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0;
wire
  \[59] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[130] ,
  \[19] ,
  \[131] ,
  \[132] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[0] ,
  \[136] ,
  \[1] ,
  \[137] ,
  \[64] ,
  \[20] ,
  \[65] ,
  \[21] ,
  \[3] ,
  \[66] ,
  \[22] ,
  \[4] ,
  \[67] ,
  \[23] ,
  \[68] ,
  \[24] ,
  \[6] ,
  \[25] ,
  \[7] ,
  \[26] ,
  \[8] ,
  \[27] ,
  \[9] ,
  \[28] ,
  \[140] ,
  \[29] ,
  \[143] ,
  \[70] ,
  \[100] ,
  \[71] ,
  \[101] ,
  \[72] ,
  \[102] ,
  \[73] ,
  \[74] ,
  \[30] ,
  \[75] ,
  \[31] ,
  \[105] ,
  \[76] ,
  \[32] ,
  \[106] ,
  \[77] ,
  \[33] ,
  \[107] ,
  \[78] ,
  \[34] ,
  a6,
  \[108] ,
  \[79] ,
  \[35] ,
  \[109] ,
  \[36] ,
  \[37] ,
  d5,
  \[38] ,
  e5,
  \[39] ,
  g5,
  g6,
  h4,
  h6,
  h7,
  \[80] ,
  \[110] ,
  \[81] ,
  j5,
  j6,
  \[111] ,
  j7,
  \[82] ,
  k5,
  k6,
  \[112] ,
  \[83] ,
  l5,
  l6,
  \[113] ,
  \[84] ,
  \[40] ,
  m4,
  m6,
  \[85] ,
  \[41] ,
  n4,
  n5,
  n6,
  \[115] ,
  \[86] ,
  \[42] ,
  o4,
  o5,
  o6,
  \[87] ,
  \[43] ,
  p4,
  p5,
  \[88] ,
  \[44] ,
  q5,
  \[118] ,
  \[89] ,
  \[45] ,
  r4,
  r6,
  \[119] ,
  \[46] ,
  s5,
  s6,
  \[47] ,
  t5,
  t6,
  \[48] ,
  u5,
  u6,
  \[49] ,
  v4,
  w4,
  w5,
  w6,
  x5,
  \[90] ,
  y5,
  \[91] ,
  z4,
  z5,
  \[121] ,
  \[122] ,
  \[123] ,
  \[50] ,
  \[124] ,
  \[95] ,
  \[51] ,
  \[125] ,
  \[96] ,
  \[52] ,
  \[126] ,
  \[53] ,
  \[127] ,
  \[54] ,
  \[10] ,
  \[128] ,
  \[55] ,
  \[11] ,
  \[129] ,
  \[56] ,
  \[12] ,
  \[13] ,
  \[14] ;
assign
  \[59]  = \[52]  | \[50] ,
  \[15]  = \[131]  | (\[130]  | (\[128]  | (\[127]  | (\[124]  | (\[118]  | (\[113]  | (\[105]  | (\[83]  | (\[70]  | (\[50]  | (r4 | (g5 | (o5 | (m4 | (n6 | \[35] ))))))))))))))),
  \[16]  = (e5 & (~i & ~c)) | ((\[8]  & p) | (\[131]  | (\[127]  | (\[119]  | (\[115]  | (\[101]  | (\[100]  | (\[90]  | (\[82]  | (\[68]  | (\[54]  | (z4 | (h7 | (j5 | (p5 | (s5 | (w5 | (h6 | (l6 | (m6 | (\[38]  | (\[37]  | \[11] )))))))))))))))))))))),
  \[17]  = (\[46]  & (\[44]  & (~m & ~c))) | (\[131]  | (\[129]  | (\[126]  | (\[119]  | (\[96]  | (\[85]  | (\[77]  | (\[64]  | (\[55]  | (\[48]  | (y5 | (v4 | (u6 | (d5 | (w5 | (j6 | t6)))))))))))))))),
  \[18]  = \[128]  | d5,
  \[130]  = (\[87]  & (\[41]  & ~g)) | ((\[53]  & (\[43]  & g)) | (e5 | l5)),
  \[19]  = \[102]  | (\[62]  | (\[38]  | (\[37]  | (\[36]  | \[18] )))),
  \[131]  = (\[51]  & (\[41]  & m)) | (p4 | w4),
  \[132]  = \[45]  & a,
  r = \[0] ,
  s = \[1] ,
  t = \[6] ,
  \[60]  = (\[143]  & (~i & d)) | ((\[109]  & (k & g)) | ((\[109]  & (i & g)) | (\[109]  & (g & c)))),
  u = \[3] ,
  v = \[4] ,
  w = \[6] ,
  \x  = \[6] ,
  y = \[7] ,
  z = \[8] ,
  \[61]  = ~o & n,
  \[62]  = (\[87]  & (\[41]  & g)) | (\[49]  & (\[42]  & g)),
  \[0]  = \[84]  | (\[62]  | (n5 | \[6] )),
  \[136]  = \[46]  & \[42] ,
  \[1]  = \[107]  | (d5 | (j7 | \[35] )),
  \[137]  = \[44]  & \[39] ,
  \[64]  = s5 | z5,
  \[20]  = \[123]  | (\[101]  | (\[96]  | (\[89]  | (\[82]  | (\[79]  | (\[54]  | u5)))))),
  \[65]  = (\[132]  & (\[80]  & e)) | (\[111]  & (~g6 & e)),
  \[21]  = \[96]  | (\[83]  | (\[78]  | (\[54]  | (\[52]  | (z5 | (g6 | (h4 | \[37] ))))))),
  \[3]  = \[95]  | (\[76]  | (j5 | \[11] )),
  \[66]  = o & n,
  \[22]  = \[123]  | (\[102]  | (\[101]  | (\[89]  | (n4 | \[37] )))),
  \[4]  = j6 | \[7] ,
  \[67]  = \[40]  & ~i,
  \[23]  = \[122]  | (\[121]  | (\[101]  | (\[72]  | (\[50]  | (x5 | (j6 | (\[18]  | \[10] ))))))),
  \[68]  = n6 | t6,
  \[24]  = \[125]  | (\[102]  | (\[62]  | r6)),
  \[6]  = \[96]  | (\[86]  | (\[85]  | (\[83]  | (\[82]  | \[56] )))),
  \[25]  = \[124]  | (\[123]  | (\[91]  | (\[86]  | \[85] ))),
  \[7]  = \[60]  | (m4 | (n5 | (\[9]  | \[3] ))),
  \[26]  = \[112]  | (\[95]  | (\[84]  | (\[83]  | (\[78]  | (\[76]  | (\[52]  | (\[48]  | (m4 | (x5 | \[8] ))))))))),
  \[8]  = \[45]  & (\[41]  & ~l),
  \[27]  = \[85]  | \[24] ,
  \[9]  = \[112]  | \[62] ,
  \[28]  = \[122]  | (\[121]  | (\[90]  | (\[72]  | (\[50]  | (j5 | (t5 | (z5 | (j6 | \[10] )))))))),
  \[140]  = \[61]  & \[47] ,
  \[29]  = \[122]  | (\[102]  | (\[85]  | (r6 | l6))),
  \[143]  = \[74]  & \[42] ,
  \[70]  = \[55]  | \[54] ,
  \[100]  = w6 | r4,
  \[71]  = \[64]  | x5,
  \[101]  = \[36]  | \[34] ,
  \[72]  = (\[88]  & (\[81]  & (j & ~f))) | ((\[88]  & (\[81]  & (j & ~c))) | (\[88]  & (\[81]  & (j & b)))),
  \[102]  = \[86]  | \[78] ,
  \[73]  = \[44]  & \[42] ,
  \[74]  = \[43]  & ~o,
  \[30]  = \[124]  | (\[91]  | (\[70]  | (\[62]  | (\[56]  | s5)))),
  \[75]  = \[41]  & \[39] ,
  \[31]  = \[83]  | (\[59]  | k6),
  \[105]  = (\[137]  & \[53] ) | (p5 | n4),
  \[76]  = k5 | u6,
  \[32]  = \[125]  | (\[83]  | (\[59]  | r6)),
  \[106]  = (\[88]  & (\[49]  & (m & (~j & ~f)))) | ((\[88]  & (\[49]  & (m & (~j & ~c)))) | ((\[88]  & (\[49]  & (m & (~j & b)))) | (\[75]  & (\[67]  & (~k & (g & ~c)))))),
  \[77]  = m4 | j5,
  \[33]  = \[125]  | (\[121]  | (\[68]  | (\[59]  | (\[56]  | (\[55]  | (s5 | \[11] )))))),
  \[107]  = (~\[88]  & (\[67]  & (\[66]  & (~l5 & (~o6 & ~l))))) | ((\[132]  & (\[80]  & (~f & ~e))) | ((\[87]  & (\[66]  & ~l5)) | (\[108]  & \[66] ))),
  \[78]  = \[56]  | n5,
  \[34]  = \[73]  & \[47] ,
  a0 = \[9] ,
  a1 = \[35] ,
  a6 = \[143]  & i,
  \[108]  = \[51]  & \[45] ,
  \[79]  = \[71]  | \[59] ,
  \[35]  = \[73]  & \[51] ,
  b0 = \[10] ,
  b1 = \[36] ,
  \[109]  = \[75]  & \[40] ,
  \[36]  = l5 & j,
  c0 = \[11] ,
  c1 = \[37] ,
  \[37]  = (\[53]  & \[49] ) | s6,
  d0 = \[12] ,
  d1 = \[38] ,
  d5 = \[46]  & (\[45]  & \[44] ),
  \[38]  = \[140]  & \[53] ,
  e0 = \[13] ,
  e5 = \[49]  & (q & ~g),
  \[39]  = p & ~l,
  f0 = \[14] ,
  g0 = \[15] ,
  g5 = \[47]  & (\[42]  & n),
  g6 = \[111]  & (f & ~b),
  h0 = \[16] ,
  h4 = \[73]  & (\[46]  & c),
  h6 = \[108]  & \[44] ,
  h7 = \[75]  & (\[42]  & k),
  \[80]  = \[47]  & \[41] ,
  i0 = \[17] ,
  \[110]  = \[51]  & \[42] ,
  \[81]  = \[67]  & \[49] ,
  j0 = \[18] ,
  j5 = \[137]  & \[40] ,
  j6 = \[61]  & (\[46]  & \[45] ),
  \[111]  = \[73]  & \[39] ,
  j7 = \[73]  & (p & (~f & ~e)),
  \[82]  = n4 | h4,
  k0 = \[19] ,
  k5 = z4 & n,
  k6 = \[80]  & \[53] ,
  \[112]  = \[11]  | \[10] ,
  \[83]  = \[65]  | m6,
  l0 = \[20] ,
  l5 = \[87]  & (\[66]  & h),
  l6 = \[137]  & \[45] ,
  \[113]  = (\[80]  & ~a) | j7,
  \[84]  = \[68]  | j6,
  \[40]  = ~q & m,
  m0 = \[21] ,
  m4 = \[143]  & (~i & ~d),
  m6 = \[136]  & \[41] ,
  \[85]  = \[72]  | h6,
  \[41]  = o & ~n,
  n0 = \[22] ,
  n4 = \[108]  & \[41] ,
  n5 = \[110]  & (\[41]  & g),
  n6 = \[74]  & (\[45]  & ~f),
  \[115]  = (\[53]  & (\[46]  & \[41] )) | y5,
  \[86]  = \[79]  | \[70] ,
  \[42]  = q & ~m,
  o0 = \[23] ,
  o4 = \[110]  & (\[41]  & ~g),
  o5 = \[51]  & (\[40]  & ~n),
  o6 = \[81]  & (h & (f & (c & ~b))),
  \[87]  = \[46]  & \[40] ,
  \[43]  = \[39]  & n,
  p0 = \[24] ,
  p4 = \[110]  & \[61] ,
  p5 = \[80]  & \[40] ,
  \[88]  = h & e,
  \[44]  = ~o & ~n,
  q0 = \[25] ,
  q5 = \[53]  & (\[51]  & \[44] ),
  \[118]  = (\[74]  & \[40] ) | s6,
  \[89]  = \[38]  | \[35] ,
  \[45]  = ~q & ~m,
  r0 = \[26] ,
  r4 = \[49]  & (\[40]  & i),
  r6 = \[110]  & \[66] ,
  \[119]  = (\[132]  & (\[41]  & (l & (f & ~e)))) | (\[111]  & (f & (~e & b))),
  \[46]  = ~p & ~l,
  s0 = \[27] ,
  s5 = \[140]  & \[40] ,
  s6 = \[47]  & (\[45]  & \[44] ),
  \[47]  = ~p & l,
  t0 = \[28] ,
  t5 = \[80]  & \[42] ,
  t6 = \[74]  & (\[45]  & f),
  \[48]  = (\[74]  & (\[53]  & ~g)) | (\[109]  & ~g),
  u0 = \[29] ,
  u5 = \[61]  & (\[53]  & \[51] ),
  u6 = g5 & ~o,
  \[49]  = \[43]  & o,
  v0 = \[30] ,
  v4 = \[44]  & (\[40]  & l),
  w0 = \[31] ,
  w4 = \[53]  & (\[47]  & \[44] ),
  w5 = \[136]  & \[66] ,
  w6 = \[66]  & (\[45]  & ~p),
  x0 = \[32] ,
  x5 = \[75]  & \[53] ,
  \[90]  = \[60]  | k6,
  y0 = \[33] ,
  y5 = \[66]  & (\[45]  & ~l),
  \[91]  = \[77]  | \[76] ,
  z0 = \[34] ,
  z4 = \[53]  & (\[46]  & ~o),
  z5 = \[87]  & \[44] ,
  \[121]  = (\[8]  & ~p) | \[65] ,
  \[122]  = \[82]  | \[62] ,
  \[123]  = \[84]  | \[9] ,
  \[50]  = q5 | a6,
  \[124]  = \[90]  | \[8] ,
  \[95]  = k6 | r6,
  \[51]  = p & l,
  \[125]  = \[91]  | \[60] ,
  \[96]  = l6 | \[8] ,
  \[52]  = (w6 & y5) | p5,
  \[126]  = (\[87]  & \[61] ) | \[100] ,
  \[53]  = q & m,
  \[127]  = (\[108]  & \[61] ) | \[106] ,
  \[54]  = \[48]  | t5,
  \[10]  = \[75]  & (\[42]  & ~k),
  \[128]  = (\[66]  & (\[47]  & \[40] )) | \[107] ,
  \[55]  = u5 | g6,
  \[11]  = \[136]  & \[61] ,
  \[129]  = (\[140]  & \[45] ) | (\[105]  | o6),
  \[56]  = w5 | o4,
  \[12]  = (\[61]  & (\[40]  & p)) | (\[129]  | (\[128]  | (\[115]  | (\[113]  | (\[95]  | (\[89]  | (\[85]  | (s6 | (o5 | (v4 | (w4 | (h7 | (q5 | (s5 | (t5 | (o4 | (g6 | (n5 | \[34] )))))))))))))))))),
  \[13]  = \[130]  | (\[127]  | (\[126]  | (\[95]  | (\[89]  | (\[77]  | (\[71]  | (\[62]  | (\[48]  | (z4 | (g5 | (o5 | (v4 | (h7 | (o6 | (q5 | (o4 | n6)))))))))))))))),
  \[14]  = \[130]  | (\[129]  | (\[126]  | (\[119]  | (\[118]  | (\[115]  | (\[112]  | (\[106]  | (\[89]  | (\[84]  | (\[78]  | (\[60]  | (p4 | (k5 | (u5 | (x5 | a6)))))))))))))));
endmodule

