`timescale 1 ps / 1 ps

module carry_sum (sin, cin, sout, cout);
  input sin;
  input cin;
  output sout;
  output cout;
endmodule
