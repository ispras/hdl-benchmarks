// IWLS benchmark module "i8" printed on Wed May 29 17:26:52 2002
module i8(\V133(3) , \V133(1) , \V133(2) , \V133(0) , \V133(5) , \V133(10) , \V133(6) , \V133(7) , \V133(8) , \V47(31) , \V47(30) , \V47(29) , \V47(28) , \V47(27) , \V47(26) , \V47(25) , \V47(24) , \V47(23) , \V47(22) , \V47(21) , \V47(20) , \V47(19) , \V47(18) , \V47(17) , \V47(16) , \V47(15) , \V47(14) , \V47(13) , \V47(12) , \V47(11) , \V47(10) , \V47(9) , \V47(8) , \V47(7) , \V47(6) , \V47(5) , \V47(4) , \V47(3) , \V47(2) , \V47(1) , \V47(0) , \V84(11) , \V84(10) , \V84(9) , \V84(8) , \V84(7) , \V84(6) , \V84(5) , \V84(4) , \V84(3) , \V84(2) , \V84(1) , \V15(14) , \V15(13) , \V15(12) , \V15(11) , \V15(10) , \V15(9) , \V15(8) , \V15(7) , \V15(6) , \V15(5) , \V15(4) , \V15(3) , \V15(2) , \V15(1) , \V15(0) , \V84(31) , \V84(30) , \V84(29) , \V84(28) , \V84(27) , \V84(26) , \V84(25) , \V84(24) , \V84(23) , \V84(22) , \V84(21) , \V84(20) , \V84(19) , \V84(18) , \V84(17) , \V84(16) , \V84(15) , \V84(14) , \V84(13) , \V84(12) , \V84(0) , \V48(0) , \V49(0) , \V116(0) , \V50(0) , \V52(0) , \V51(0) , \V116(2) , \V133(9) , \V116(1) , \V116(8) , \V116(7) , \V116(6) , \V116(5) , \V116(4) , \V116(3) , \V116(9) , \V116(11) , \V116(10) , \V116(12) , \V116(15) , \V116(14) , \V116(13) , \V116(16) , \V116(31) , \V116(30) , \V116(29) , \V116(28) , \V116(27) , \V116(26) , \V116(25) , \V116(24) , \V116(23) , \V116(22) , \V116(21) , \V116(20) , \V116(19) , \V116(18) , \V116(17) , \V121(16) , \V119(0) , \V121(17) , \V122(0) , \V133(4) , \V118(0) , \V118(1) , \V134(0) , \V136(1) , \V136(0) , \V142(5) , \V142(4) , \V142(3) , \V142(2) , \V142(1) , \V142(0) , \V143(0) , \V145(1) , \V145(0) , \V146(0) , \V149(2) , \V149(1) , \V149(0) , \V150(0) , \V165(14) , \V165(13) , \V165(12) , \V165(11) , \V165(10) , \V165(9) , \V165(8) , \V165(7) , \V165(6) , \V165(5) , \V165(4) , \V165(3) , \V165(2) , \V165(1) , \V165(0) , \V197(31) , \V197(30) , \V197(29) , \V197(28) , \V197(27) , \V197(26) , \V197(25) , \V197(24) , \V197(23) , \V197(22) , \V197(21) , \V197(20) , \V197(19) , \V197(18) , \V197(17) , \V197(16) , \V197(15) , \V197(14) , \V197(13) , \V197(12) , \V197(11) , \V197(10) , \V197(9) , \V197(8) , \V197(7) , \V197(6) , \V197(5) , \V197(4) , \V197(3) , \V197(2) , \V197(1) , \V197(0) , \V212(14) , \V212(13) , \V212(12) , \V212(11) , \V212(10) , \V212(9) , \V212(8) , \V212(7) , \V212(6) , \V212(5) , \V212(4) , \V212(3) , \V212(2) , \V212(1) , \V212(0) , \V213(0) , \V214(0) );
input
  \V116(12) ,
  \V133(5) ,
  \V116(15) ,
  \V133(4) ,
  \V116(14) ,
  \V133(1) ,
  \V133(0) ,
  \V133(7) ,
  \V133(6) ,
  \V116(3) ,
  \V133(9) ,
  \V116(2) ,
  \V133(8) ,
  \V116(5) ,
  \V116(4) ,
  \V116(1) ,
  \V116(0) ,
  \V116(7) ,
  \V116(6) ,
  \V116(9) ,
  \V116(8) ,
  \V116(31) ,
  \V116(30) ,
  \V118(1) ,
  \V118(0) ,
  \V84(13) ,
  \V84(12) ,
  \V84(15) ,
  \V84(14) ,
  \V15(13) ,
  \V15(12) ,
  \V84(11) ,
  \V84(10) ,
  \V15(14) ,
  \V15(11) ,
  \V15(10) ,
  \V84(17) ,
  \V84(16) ,
  \V84(19) ,
  \V84(18) ,
  \V84(23) ,
  \V84(22) ,
  \V84(25) ,
  \V84(24) ,
  \V84(21) ,
  \V84(20) ,
  \V84(27) ,
  \V84(26) ,
  \V84(29) ,
  \V84(28) ,
  \V47(13) ,
  \V47(12) ,
  \V47(15) ,
  \V47(14) ,
  \V84(31) ,
  \V84(30) ,
  \V47(11) ,
  \V47(10) ,
  \V47(17) ,
  \V47(16) ,
  \V47(19) ,
  \V47(18) ,
  \V47(23) ,
  \V47(22) ,
  \V47(25) ,
  \V47(24) ,
  \V122(0) ,
  \V47(21) ,
  \V47(20) ,
  \V47(27) ,
  \V47(26) ,
  \V47(29) ,
  \V47(28) ,
  \V84(0) ,
  \V84(1) ,
  \V47(31) ,
  \V84(2) ,
  \V47(30) ,
  \V84(3) ,
  \V84(4) ,
  \V84(5) ,
  \V84(6) ,
  \V84(7) ,
  \V84(8) ,
  \V84(9) ,
  \V48(0) ,
  \V50(0) ,
  \V52(0) ,
  \V133(10) ,
  \V119(0) ,
  \V47(0) ,
  \V47(1) ,
  \V47(2) ,
  \V47(3) ,
  \V47(4) ,
  \V47(5) ,
  \V47(6) ,
  \V47(7) ,
  \V47(8) ,
  \V47(9) ,
  \V49(0) ,
  \V121(17) ,
  \V121(16) ,
  \V51(0) ,
  \V116(27) ,
  \V116(26) ,
  \V116(29) ,
  \V116(28) ,
  \V15(0) ,
  \V15(1) ,
  \V15(2) ,
  \V15(3) ,
  \V15(4) ,
  \V15(5) ,
  \V15(6) ,
  \V116(21) ,
  \V15(7) ,
  \V116(20) ,
  \V15(8) ,
  \V116(23) ,
  \V15(9) ,
  \V116(22) ,
  \V116(25) ,
  \V116(24) ,
  \V116(17) ,
  \V116(16) ,
  \V116(19) ,
  \V116(18) ,
  \V116(11) ,
  \V116(10) ,
  \V133(3) ,
  \V116(13) ,
  \V133(2) ;
output
  \V212(3) ,
  \V212(2) ,
  \V212(5) ,
  \V212(4) ,
  \V212(1) ,
  \V212(0) ,
  \V212(7) ,
  \V212(6) ,
  \V212(9) ,
  \V212(8) ,
  \V214(0) ,
  \V143(0) ,
  \V145(1) ,
  \V145(0) ,
  \V149(2) ,
  \V149(1) ,
  \V149(0) ,
  \V134(0) ,
  \V136(1) ,
  \V136(0) ,
  \V165(11) ,
  \V197(3) ,
  \V165(10) ,
  \V197(2) ,
  \V165(13) ,
  \V197(5) ,
  \V165(12) ,
  \V197(4) ,
  \V197(27) ,
  \V197(26) ,
  \V165(14) ,
  \V197(29) ,
  \V197(1) ,
  \V197(28) ,
  \V197(0) ,
  \V197(7) ,
  \V197(6) ,
  \V197(21) ,
  \V197(9) ,
  \V197(20) ,
  \V197(8) ,
  \V197(23) ,
  \V197(22) ,
  \V197(25) ,
  \V197(24) ,
  \V213(0) ,
  \V197(17) ,
  \V197(16) ,
  \V197(19) ,
  \V197(18) ,
  \V197(11) ,
  \V197(10) ,
  \V197(13) ,
  \V197(12) ,
  \V197(15) ,
  \V197(14) ,
  \V142(3) ,
  \V142(2) ,
  \V142(5) ,
  \V142(4) ,
  \V197(31) ,
  \V142(1) ,
  \V197(30) ,
  \V142(0) ,
  \V165(3) ,
  \V212(11) ,
  \V165(2) ,
  \V212(10) ,
  \V165(5) ,
  \V212(13) ,
  \V165(4) ,
  \V212(12) ,
  \V146(0) ,
  \V212(14) ,
  \V165(1) ,
  \V165(0) ,
  \V165(7) ,
  \V165(6) ,
  \V165(9) ,
  \V165(8) ,
  \V150(0) ;
wire
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  V215,
  V219,
  V222,
  V223,
  V224,
  V226,
  V228,
  V229,
  V230,
  V231,
  V236,
  V237,
  V238,
  V239,
  V240,
  V241,
  V242,
  V243,
  V244,
  V245,
  V246,
  V247,
  V248,
  V249,
  V250,
  V251,
  V252,
  V253,
  V254,
  V255,
  V256,
  V257,
  V258,
  V259,
  V260,
  V261,
  V262,
  V263,
  V264,
  V265,
  V266,
  V268,
  V270,
  V272,
  V274,
  V276,
  V278,
  V280,
  V282,
  V284,
  V286,
  V288,
  V290,
  V292,
  V294,
  V296,
  V298,
  V300,
  V302,
  V304,
  V306,
  V308,
  V310,
  V312,
  V314,
  V324,
  V325,
  V326,
  V327,
  V328,
  V329,
  V330,
  V331,
  V332,
  V333,
  V334,
  V335,
  V336,
  V337,
  V338,
  V339,
  V340,
  V341,
  V342,
  V343,
  V344,
  V345,
  V346,
  V347,
  V348,
  V349,
  V350,
  V351,
  V352,
  V353,
  V354,
  V356,
  V357,
  V358,
  V359,
  V360,
  V361,
  V362,
  V363,
  V364,
  V365,
  V366,
  V367,
  V368,
  V369,
  V370,
  V371,
  V372,
  V373,
  V374,
  V375,
  V376,
  V377,
  V378,
  V379,
  V380,
  V381,
  V382,
  V383,
  V384,
  V385,
  V386,
  V388,
  V389,
  V390,
  V391,
  V392,
  V393,
  V394,
  V395,
  V396,
  V397,
  V398,
  V399,
  V400,
  V401,
  V402,
  V403,
  V404,
  V405,
  V406,
  V407,
  V408,
  V409,
  V410,
  V411,
  V412,
  V413,
  V414,
  V415,
  V416,
  V417,
  V418,
  V419,
  V420,
  V422,
  V424,
  V426,
  V428,
  V430,
  V432,
  V434,
  V436,
  V438,
  V440,
  V442,
  V444,
  V446,
  V448,
  V450,
  V452,
  V454,
  V456,
  V458,
  V460,
  V462,
  V464,
  V466,
  V468,
  V470,
  V472,
  V474,
  V476,
  V478,
  V480,
  V482,
  V484,
  V487,
  V488,
  V489,
  V490,
  V491,
  V492,
  V493,
  V494,
  V495,
  V496,
  V497,
  V498,
  V499,
  \V235(3) ,
  \V235(2) ,
  V500,
  V501,
  V502,
  V503,
  V504,
  V505,
  V506,
  V507,
  V508,
  V509,
  V510,
  V511,
  V512,
  V513,
  V514,
  V515,
  V516,
  V517,
  V518,
  \V235(1) ,
  V520,
  V521,
  V522,
  V523,
  V524,
  V525,
  V526,
  V527,
  V528,
  V529,
  \V235(0) ,
  V530,
  V531,
  V532,
  V533,
  V534,
  V535,
  V536,
  V537,
  V538,
  V539,
  V540,
  V541,
  V542,
  V543,
  V544,
  V545,
  V546,
  V547,
  V548,
  V549,
  V550,
  V551,
  V553,
  V554,
  V555,
  V557,
  V558,
  V560,
  V561,
  V563,
  V564,
  V566,
  V568,
  V569,
  V570,
  V571,
  V573,
  V574,
  V575,
  V577,
  V578,
  V580,
  V581,
  V583,
  V584,
  V585,
  V587,
  V588,
  V589,
  V591,
  V592,
  V593,
  V594,
  V595,
  V596,
  V597,
  V598,
  V599,
  V601,
  V602,
  V603,
  V604,
  V605,
  V606,
  V607,
  V609,
  V610,
  V611,
  V612,
  V613,
  V614,
  V616,
  V617,
  V618,
  V619,
  V620,
  V621,
  V622,
  V623,
  V625,
  V626,
  V628,
  V630,
  V631,
  V632,
  V633,
  V635,
  V636,
  V637,
  V639,
  V640,
  V642,
  V643,
  V644,
  V645,
  V647,
  V648,
  V650,
  V651,
  V653,
  V654,
  V656,
  V658,
  V659,
  V661,
  V662,
  V663,
  V664,
  V665,
  V667,
  V668,
  V669,
  V670,
  V672,
  V673,
  V674,
  V675,
  V677,
  V678,
  V679,
  V680,
  V682,
  V683,
  V684,
  V686,
  V687,
  V688,
  V689,
  V691,
  V692,
  V693,
  V694,
  V695,
  V697,
  V698,
  V700,
  V701,
  V703,
  V704,
  V706,
  V707,
  V709,
  V711,
  V712,
  V714,
  V715,
  V716,
  V717,
  V718,
  V719,
  V720,
  V721,
  V722,
  V723,
  V724,
  V725,
  V726,
  V727,
  V728,
  V729,
  V730,
  V732,
  V733,
  V734,
  V735,
  V736,
  V737,
  V738,
  V739,
  V740,
  V741,
  V742,
  V743,
  V744,
  V745,
  V746,
  V747,
  V749,
  V750,
  V751,
  V752,
  V753,
  V754,
  V755,
  V756,
  V757,
  V758,
  V759,
  V760,
  V761,
  V762,
  V763,
  V764,
  V766,
  V767,
  V768,
  V769,
  V770,
  V771,
  V772,
  V773,
  V774,
  V775,
  V776,
  V777,
  V778,
  V779,
  V780,
  V781,
  V783,
  V784,
  V785,
  V786,
  V787,
  V788,
  V789,
  V790,
  V791,
  V792,
  V793,
  V794,
  V795,
  V796,
  V797,
  V799,
  V800,
  V801,
  V802,
  V803,
  V804,
  V805,
  V806,
  V807,
  V808,
  V809,
  V810,
  V811,
  V812,
  V813,
  V814,
  V816,
  V817,
  V818,
  V819,
  V820,
  V821,
  V822,
  V823,
  V824,
  V825,
  V826,
  V827,
  V828,
  V829,
  V830,
  V831,
  V832,
  V833,
  V834,
  V835,
  V836,
  V837,
  V838,
  V839,
  V840,
  V841,
  V842,
  V843,
  V844,
  V845,
  V846,
  V847,
  V848,
  V849,
  V850,
  V851,
  V852,
  V853,
  V854,
  V855,
  V856,
  V857,
  V858,
  V859,
  V860,
  V861,
  V862,
  V863,
  V865,
  V866,
  V867,
  V868,
  V869,
  V870,
  V871,
  V872,
  V873,
  V874,
  V875,
  V876,
  V877,
  V878,
  V879,
  V880,
  V881,
  V882,
  V883,
  V884,
  V885,
  V886,
  V887,
  V888,
  V889,
  V890,
  V891,
  V892,
  V893,
  V894,
  V895,
  V896,
  V897,
  V899,
  V900,
  V901,
  V902,
  V903,
  V904,
  V905,
  V906,
  V907,
  V908,
  V909,
  V910,
  V911,
  V912,
  V913,
  V914,
  V915,
  V916,
  V917,
  V918,
  V919,
  V920,
  V921,
  V922,
  V923,
  V924,
  V925,
  V926,
  V927,
  V928,
  V929,
  V930,
  V931,
  V933,
  V934,
  V935,
  V936,
  V937,
  V938,
  V939,
  V940,
  V941,
  V942,
  V943,
  V944,
  V945,
  V946,
  V947,
  V948,
  V949,
  V950,
  V951,
  V952,
  V953,
  V954,
  V955,
  V956,
  V957,
  V958,
  V959,
  V960,
  V961,
  V962,
  V963,
  V964,
  V965,
  V967,
  V968,
  V969,
  V970,
  V971,
  V972,
  V973,
  V974,
  V975,
  V976,
  V977,
  V978,
  V979,
  V980,
  V981,
  V982,
  V983,
  V984,
  V985,
  V986,
  V987,
  V988,
  V989,
  V990,
  V991,
  V992,
  V993,
  V994,
  V995,
  V996,
  V997,
  V998,
  V999,
  V1001,
  V1002,
  V1003,
  V1004,
  V1005,
  V1006,
  V1007,
  V1008,
  V1009,
  V1010,
  V1011,
  V1012,
  V1013,
  V1014,
  V1015,
  V1016,
  V1017,
  V1018,
  V1019,
  V1020,
  V1021,
  V1022,
  V1023,
  V1024,
  V1025,
  V1026,
  V1027,
  V1028,
  V1029,
  V1030,
  V1031,
  V1032,
  V1034,
  V1035,
  V1036,
  V1037,
  V1038,
  V1039,
  V1040,
  V1041,
  V1042,
  V1043,
  V1044,
  V1045,
  V1046,
  V1047,
  V1048,
  V1049,
  V1050,
  V1051,
  V1052,
  V1053,
  V1054,
  V1055,
  V1056,
  V1057,
  V1058,
  V1059,
  V1060,
  V1061,
  V1062,
  V1063,
  V1064,
  V1065,
  V1066,
  V1067,
  V1068,
  V1069,
  V1070,
  V1071,
  V1072,
  V1073,
  V1074,
  V1075,
  V1076,
  V1077,
  V1078,
  V1079,
  V1080,
  V1081,
  V1083,
  V1084,
  V1085,
  V1086,
  V1087,
  V1088,
  V1089,
  V1090,
  V1091,
  V1092,
  V1093,
  V1094,
  V1095,
  V1096,
  V1097,
  V1098,
  V1100,
  V1101,
  V1102,
  V1103,
  V1104,
  V1105,
  V1106,
  V1107,
  V1108,
  V1109,
  V1110,
  V1111,
  V1112,
  V1113,
  V1114,
  V1116,
  V1117,
  V1119,
  V1120,
  V1121,
  V1122,
  V1123,
  V1124,
  V1125,
  V1126,
  V1127,
  V1128,
  V1129,
  V1130,
  V1131,
  V1132,
  V1133,
  V1134,
  V1135,
  V1137,
  V1139,
  V1141,
  V1143,
  V1144,
  V1146,
  V1147,
  V1149,
  V1150,
  V1151,
  V1153,
  V1154,
  V1156,
  \V485(27) ,
  \V485(26) ,
  \V485(29) ,
  \V485(28) ,
  \V485(21) ,
  \V485(20) ,
  \V485(23) ,
  \V485(22) ,
  \V485(25) ,
  \V485(24) ,
  \V485(17) ,
  \V485(16) ,
  \V485(19) ,
  \V485(18) ,
  \V322(3) ,
  \V485(11) ,
  \V322(2) ,
  \V485(10) ,
  \V322(5) ,
  \V485(13) ,
  \V322(4) ,
  \V485(12) ,
  \V485(15) ,
  \V485(14) ,
  \V322(1) ,
  \V322(0) ,
  \V322(7) ,
  \V322(6) ,
  \V322(9) ,
  \V322(8) ,
  \V485(31) ,
  \V485(30) ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \V322(27) ,
  \[51] ,
  \V322(26) ,
  \[52] ,
  \V322(29) ,
  \[53] ,
  \V322(28) ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \V322(21) ,
  \V322(20) ,
  \V322(23) ,
  \V322(22) ,
  \V322(25) ,
  \V322(24) ,
  \[60] ,
  \V322(17) ,
  \[61] ,
  \V322(16) ,
  \[62] ,
  \V322(19) ,
  \[63] ,
  \V322(18) ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \V322(11) ,
  \V322(10) ,
  \V322(13) ,
  \V322(12) ,
  \V322(15) ,
  \V322(14) ,
  \[70] ,
  \[71] ,
  \V485(3) ,
  \[72] ,
  \V485(2) ,
  \[73] ,
  \V485(5) ,
  \[74] ,
  \V485(4) ,
  \[75] ,
  \[76] ,
  \[77] ,
  \V485(1) ,
  \[78] ,
  \V485(0) ,
  \[79] ,
  \V485(7) ,
  \V485(6) ,
  \V485(9) ,
  \[80] ,
  \V485(8) ,
  \V322(30) ;
assign
  \[0]  = V568 | (V566 | (V564 | (V561 | (V558 | V555)))),
  \[1]  = V588 | (V584 | (V591 | (V577 | (V574 | V570)))),
  \[2]  = V592 | (V589 | (V585 | (V581 | (V578 | (V575 | V571))))),
  \[3]  = V616 | (V609 | (V602 | V594)),
  \[4]  = V617 | (V610 | (V603 | V595)),
  \[5]  = V618 | (V611 | (V604 | V596)),
  \[6]  = V619 | (V612 | (V605 | V597)),
  \[7]  = V620 | (V613 | (V606 | V598)),
  \[8]  = V621 | (V614 | (V607 | V599)),
  \[9]  = V630 | (V628 | (V626 | V623)),
  V215 = \V133(2)  & (\V133(1)  & \V133(3) ),
  V219 = ~\V133(10)  & (~\V133(5)  & ~\V133(0) ),
  V222 = ~\V133(6)  & (~\V133(10)  & (~\V133(5)  & (~\V133(2)  & \V133(1) ))),
  V223 = \V133(7)  & (~\V133(10)  & ~\V133(0) ),
  V224 = \V133(8)  & (~\V133(10)  & \V133(1) ),
  V226 = ~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) )),
  V228 = ~\V133(6)  & (~\V133(10)  & (~\V133(5)  & (\V133(0)  & (\V133(2)  & ~\V133(1) )))),
  V229 = \V133(8)  & (~\V133(10)  & (\V133(2)  & ~\V133(1) )),
  V230 = ~\V133(6)  & (~\V133(10)  & (~\V133(5)  & (~\V133(2)  & ~\V133(1) ))),
  V231 = \V133(7)  & (~\V133(10)  & (~\V133(2)  & ~\V133(1) )),
  V236 = \V47(31)  & \V235(0) ,
  V237 = \V47(30)  & \V235(0) ,
  V238 = \V47(29)  & \V235(0) ,
  V239 = \V47(28)  & \V235(0) ,
  V240 = \V47(27)  & \V235(0) ,
  V241 = \V47(26)  & \V235(0) ,
  V242 = \V47(25)  & \V235(0) ,
  V243 = \V47(24)  & \V235(0) ,
  V244 = \V47(23)  & \V235(0) ,
  V245 = \V47(22)  & \V235(0) ,
  V246 = \V47(21)  & \V235(0) ,
  V247 = \V47(20)  & \V235(0) ,
  V248 = \V47(19)  & \V235(0) ,
  V249 = \V47(18)  & \V235(0) ,
  V250 = \V47(17)  & \V235(0) ,
  V251 = \V47(16)  & \V235(0) ,
  V252 = \V47(15)  & \V235(0) ,
  V253 = \V47(14)  & \V235(0) ,
  V254 = \V47(13)  & \V235(0) ,
  V255 = \V47(12)  & \V235(0) ,
  V256 = \V47(11)  & \V235(0) ,
  V257 = \V47(10)  & \V235(0) ,
  V258 = \V47(9)  & \V235(0) ,
  V259 = \V47(8)  & \V235(0) ,
  V260 = \V47(7)  & \V235(0) ,
  V261 = \V47(6)  & \V235(0) ,
  V262 = \V47(5)  & \V235(0) ,
  V263 = \V47(4)  & \V235(0) ,
  V264 = \V47(3)  & \V235(0) ,
  V265 = \V47(2)  & \V235(0) ,
  V266 = \V47(1)  & \V235(0) ,
  V268 = \V235(1)  & (~\V235(0)  & \V47(23) ),
  V270 = \V235(1)  & (~\V235(0)  & \V47(22) ),
  V272 = \V235(1)  & (~\V235(0)  & \V47(21) ),
  V274 = \V235(1)  & (~\V235(0)  & \V47(20) ),
  V276 = \V235(1)  & (~\V235(0)  & \V47(19) ),
  V278 = \V235(1)  & (~\V235(0)  & \V47(18) ),
  V280 = \V235(1)  & (~\V235(0)  & \V47(17) ),
  V282 = \V235(1)  & (~\V235(0)  & \V47(16) ),
  V284 = \V235(1)  & (~\V235(0)  & \V47(15) ),
  \V212(3)  = \[75] ,
  V286 = \V235(1)  & (~\V235(0)  & \V47(14) ),
  V288 = \V235(1)  & (~\V235(0)  & \V47(13) ),
  V290 = \V235(1)  & (~\V235(0)  & \V47(12) ),
  V292 = \V235(1)  & (~\V235(0)  & \V47(11) ),
  V294 = \V235(1)  & (~\V235(0)  & \V47(10) ),
  \V212(2)  = \[76] ,
  V296 = \V235(1)  & (~\V235(0)  & \V47(9) ),
  V298 = \V235(1)  & (~\V235(0)  & \V47(8) ),
  \V212(5)  = \[73] ,
  \V212(4)  = \[74] ,
  \V212(1)  = \[77] ,
  \V212(0)  = \[78] ,
  V300 = \V235(1)  & (~\V235(0)  & \V47(7) ),
  V302 = \V235(1)  & (~\V235(0)  & \V47(6) ),
  V304 = \V235(1)  & (~\V235(0)  & \V47(5) ),
  V306 = \V235(1)  & (~\V235(0)  & \V47(4) ),
  V308 = \V235(1)  & (~\V235(0)  & \V47(3) ),
  V310 = \V235(1)  & (~\V235(0)  & \V47(2) ),
  V312 = \V235(1)  & (~\V235(0)  & \V47(1) ),
  V314 = \V235(1)  & (~\V235(0)  & \V47(0) ),
  V324 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(20) )),
  V325 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(19) )),
  V326 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(18) )),
  V327 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(17) )),
  V328 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(16) )),
  V329 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(15) )),
  V330 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(14) )),
  V331 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(13) )),
  V332 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(12) )),
  V333 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(11) )),
  V334 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(10) )),
  V335 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(9) )),
  V336 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(8) )),
  V337 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(7) )),
  V338 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(6) )),
  V339 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(5) )),
  V340 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(4) )),
  V341 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(3) )),
  V342 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(2) )),
  V343 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(1) )),
  V344 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(11) )),
  V345 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(10) )),
  \V212(7)  = \[71] ,
  V346 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(9) )),
  V347 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(8) )),
  V348 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(7) )),
  V349 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(6) )),
  V350 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(5) )),
  V351 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(4) )),
  V352 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(3) )),
  V353 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(2) )),
  V354 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(1) )),
  \V212(6)  = \[72] ,
  V356 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(16) ))),
  V357 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(15) ))),
  V358 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(14) ))),
  V359 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(13) ))),
  V360 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(12) ))),
  V361 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(11) ))),
  V362 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(10) ))),
  V363 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(9) ))),
  V364 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(8) ))),
  V365 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(7) ))),
  \V212(9)  = \[69] ,
  V366 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(6) ))),
  V367 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(5) ))),
  V368 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(4) ))),
  V369 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(3) ))),
  V370 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(2) ))),
  V371 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(1) ))),
  V372 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(14) ))),
  V373 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(13) ))),
  V374 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(12) ))),
  V375 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(11) ))),
  \V212(8)  = \[70] ,
  V376 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(10) ))),
  V377 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(9) ))),
  V378 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(8) ))),
  V379 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(7) ))),
  V380 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(6) ))),
  V381 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(5) ))),
  V382 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(4) ))),
  V383 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(3) ))),
  V384 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(2) ))),
  V385 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(1) ))),
  V386 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V15(0) ))),
  V388 = ~\V235(3)  & (~\V235(2)  & (~\V235(1)  & ~\V235(0) )),
  V389 = \V84(31)  & \V235(0) ,
  V390 = \V84(30)  & \V235(0) ,
  V391 = \V84(29)  & \V235(0) ,
  V392 = \V84(28)  & \V235(0) ,
  V393 = \V84(27)  & \V235(0) ,
  V394 = \V84(26)  & \V235(0) ,
  V395 = \V84(25)  & \V235(0) ,
  V396 = \V84(24)  & \V235(0) ,
  V397 = \V84(23)  & \V235(0) ,
  V398 = \V84(22)  & \V235(0) ,
  V399 = \V84(21)  & \V235(0) ,
  \V214(0)  = \[80] ,
  V400 = \V84(20)  & \V235(0) ,
  V401 = \V84(19)  & \V235(0) ,
  V402 = \V84(18)  & \V235(0) ,
  V403 = \V84(17)  & \V235(0) ,
  V404 = \V84(16)  & \V235(0) ,
  V405 = \V84(15)  & \V235(0) ,
  V406 = \V84(14)  & \V235(0) ,
  V407 = \V84(13)  & \V235(0) ,
  V408 = \V84(12)  & \V235(0) ,
  V409 = \V84(11)  & \V235(0) ,
  V410 = \V84(10)  & \V235(0) ,
  V411 = \V84(9)  & \V235(0) ,
  V412 = \V84(8)  & \V235(0) ,
  V413 = \V84(7)  & \V235(0) ,
  V414 = \V84(6)  & \V235(0) ,
  V415 = \V84(5)  & \V235(0) ,
  V416 = \V84(4)  & \V235(0) ,
  V417 = \V84(3)  & \V235(0) ,
  V418 = \V84(2)  & \V235(0) ,
  V419 = \V84(1)  & \V235(0) ,
  V420 = \V84(0)  & \V235(0) ,
  V422 = \V235(1)  & (~\V235(0)  & \V84(23) ),
  V424 = \V235(1)  & (~\V235(0)  & \V84(22) ),
  V426 = \V235(1)  & (~\V235(0)  & \V84(21) ),
  V428 = \V235(1)  & (~\V235(0)  & \V84(20) ),
  V430 = \V235(1)  & (~\V235(0)  & \V84(19) ),
  V432 = \V235(1)  & (~\V235(0)  & \V84(18) ),
  V434 = \V235(1)  & (~\V235(0)  & \V84(17) ),
  V436 = \V235(1)  & (~\V235(0)  & \V84(16) ),
  V438 = \V235(1)  & (~\V235(0)  & \V84(15) ),
  V440 = \V235(1)  & (~\V235(0)  & \V84(14) ),
  V442 = \V235(1)  & (~\V235(0)  & \V84(13) ),
  V444 = \V235(1)  & (~\V235(0)  & \V84(12) ),
  V446 = \V235(1)  & (~\V235(0)  & \V84(11) ),
  V448 = \V235(1)  & (~\V235(0)  & \V84(10) ),
  V450 = \V235(1)  & (~\V235(0)  & \V84(9) ),
  V452 = \V235(1)  & (~\V235(0)  & \V84(8) ),
  V454 = \V235(1)  & (~\V235(0)  & \V84(7) ),
  V456 = \V235(1)  & (~\V235(0)  & \V84(6) ),
  V458 = \V235(1)  & (~\V235(0)  & \V84(5) ),
  V460 = \V235(1)  & (~\V235(0)  & \V84(4) ),
  V462 = \V235(1)  & (~\V235(0)  & \V84(3) ),
  V464 = \V235(1)  & (~\V235(0)  & \V84(2) ),
  V466 = \V235(1)  & (~\V235(0)  & \V84(1) ),
  V468 = \V235(1)  & (~\V235(0)  & \V84(0) ),
  V470 = \V235(1)  & (~\V235(0)  & \V47(31) ),
  V472 = \V235(1)  & (~\V235(0)  & \V47(30) ),
  V474 = \V235(1)  & (~\V235(0)  & \V47(29) ),
  V476 = \V235(1)  & (~\V235(0)  & \V47(28) ),
  V478 = \V235(1)  & (~\V235(0)  & \V47(27) ),
  V480 = \V235(1)  & (~\V235(0)  & \V47(26) ),
  V482 = \V235(1)  & (~\V235(0)  & \V47(25) ),
  V484 = \V235(1)  & (~\V235(0)  & \V47(24) ),
  V487 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(20) )),
  V488 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(19) )),
  V489 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(18) )),
  V490 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(17) )),
  V491 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(16) )),
  V492 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(15) )),
  V493 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(14) )),
  V494 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(13) )),
  V495 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(12) )),
  V496 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(11) )),
  V497 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(10) )),
  V498 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(9) )),
  V499 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(8) )),
  \V235(3)  = V230 | V231,
  \V235(2)  = V228 | (V226 | V229),
  V500 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(7) )),
  V501 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(6) )),
  V502 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(5) )),
  V503 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(4) )),
  V504 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(3) )),
  V505 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(2) )),
  V506 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(1) )),
  V507 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(0) )),
  V508 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(31) )),
  V509 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(30) )),
  V510 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(29) )),
  V511 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(28) )),
  V512 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(27) )),
  V513 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(26) )),
  V514 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(25) )),
  V515 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(24) )),
  V516 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(23) )),
  V517 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(22) )),
  V518 = \V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(21) )),
  \V235(1)  = V223 | (V219 | (V222 | V224)),
  V520 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(16) ))),
  V521 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(15) ))),
  V522 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(14) ))),
  V523 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(13) ))),
  V524 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(12) ))),
  V525 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(11) ))),
  V526 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(10) ))),
  V527 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(9) ))),
  V528 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(8) ))),
  V529 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(7) ))),
  \V235(0)  = V215 | \V133(10) ,
  V530 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(6) ))),
  V531 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(5) ))),
  V532 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(4) ))),
  V533 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(3) ))),
  V534 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(2) ))),
  V535 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(1) ))),
  V536 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V84(0) ))),
  V537 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(31) ))),
  V538 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(30) ))),
  V539 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(29) ))),
  V540 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(28) ))),
  V541 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(27) ))),
  V542 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(26) ))),
  V543 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(25) ))),
  V544 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(24) ))),
  V545 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(23) ))),
  V546 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(22) ))),
  V547 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(21) ))),
  V548 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(20) ))),
  V549 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(19) ))),
  V550 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(18) ))),
  V551 = \V235(3)  & (~\V235(2)  & (~\V235(1)  & (~\V235(0)  & \V47(17) ))),
  V553 = ~\V235(3)  & (~\V235(2)  & (~\V235(1)  & ~\V235(0) )),
  V554 = ~\V133(9)  & (\V133(7)  & (~\V133(10)  & ~\V133(1) )),
  V555 = \V48(0)  & V554,
  V557 = ~\V133(9)  & (\V133(7)  & (~\V133(10)  & ~\V133(2) )),
  V558 = V557 & (~V554 & \V48(0) ),
  V560 = ~\V133(9)  & (~\V133(7)  & ~\V133(10) ),
  V561 = V560 & (~V557 & (~V554 & \V49(0) )),
  V563 = \V133(9)  & ~\V133(10) ,
  V564 = V563 & (~V560 & (~V557 & (~V554 & \V116(0) ))),
  V566 = ~V563 & (~V560 & (~V557 & (~V554 & (\V84(0)  & \V133(10) )))),
  V568 = ~V563 & (~V560 & (~V557 & (~V554 & ~\V133(10) ))),
  V569 = ~\V133(4)  & (~\V133(9)  & (~\V133(8)  & (\V133(2)  & \V133(1) ))),
  V570 = \V322(1)  & V569,
  V571 = \V322(0)  & V569,
  V573 = ~\V133(9)  & (~\V133(8)  & \V133(7) ),
  V574 = V573 & (~V569 & \V322(1) ),
  V575 = V573 & (~V569 & \V322(0) ),
  V577 = ~V573 & (~V569 & (\V322(1)  & \V133(10) )),
  V578 = ~V573 & (~V569 & (\V322(0)  & \V133(10) )),
  V580 = ~\V133(9)  & (\V133(8)  & ~\V133(10) ),
  V581 = V580 & (~V573 & (~V569 & (\V50(0)  & ~\V133(10) ))),
  V583 = ~\V133(9)  & (~\V133(7)  & (~\V133(10)  & ~\V133(1) )),
  V584 = V583 & (~V580 & (~V573 & (~V569 & (\V52(0)  & ~\V133(10) )))),
  V585 = V583 & (~V580 & (~V573 & (~V569 & (\V51(0)  & ~\V133(10) )))),
  V587 = ~\V133(9)  & (~\V133(7)  & (~\V133(10)  & ~\V133(2) )),
  V588 = V587 & (~V583 & (~V580 & (~V573 & (~V569 & (\V52(0)  & ~\V133(10) ))))),
  V589 = V587 & (~V583 & (~V580 & (~V573 & (~V569 & (\V51(0)  & ~\V133(10) ))))),
  V591 = ~V587 & (~V583 & (~V580 & (~V573 & (~V569 & (\V133(9)  & (\V116(2)  & ~\V133(10) )))))),
  V592 = ~V587 & (~V583 & (~V580 & (~V573 & (~V569 & (\V116(1)  & (\V133(9)  & ~\V133(10) )))))),
  V593 = ~\V133(4)  & (~\V133(9)  & ~\V133(6) ),
  V594 = \V322(7)  & V593,
  V595 = \V322(6)  & V593,
  V596 = \V322(5)  & V593,
  V597 = \V322(4)  & V593,
  V598 = \V322(3)  & V593,
  V599 = \V322(2)  & V593,
  V601 = ~\V133(9)  & \V133(7) ,
  V602 = V601 & (~V593 & \V322(7) ),
  V603 = V601 & (~V593 & \V322(6) ),
  V604 = V601 & (~V593 & \V322(5) ),
  V605 = V601 & (~V593 & \V322(4) ),
  V606 = V601 & (~V593 & \V322(3) ),
  V607 = V601 & (~V593 & \V322(2) ),
  V609 = ~V601 & (~V593 & (\V322(7)  & \V133(10) )),
  V610 = ~V601 & (~V593 & (\V322(6)  & \V133(10) )),
  V611 = ~V601 & (~V593 & (\V322(5)  & \V133(10) )),
  V612 = ~V601 & (~V593 & (\V322(4)  & \V133(10) )),
  V613 = ~V601 & (~V593 & (\V322(3)  & \V133(10) )),
  V614 = ~V601 & (~V593 & (\V322(2)  & \V133(10) )),
  V616 = ~V601 & (~V593 & (\V116(8)  & (\V133(9)  & ~\V133(10) ))),
  V617 = ~V601 & (~V593 & (\V116(7)  & (\V133(9)  & ~\V133(10) ))),
  V618 = ~V601 & (~V593 & (\V116(6)  & (\V133(9)  & ~\V133(10) ))),
  V619 = ~V601 & (~V593 & (\V116(5)  & (\V133(9)  & ~\V133(10) ))),
  V620 = ~V601 & (~V593 & (\V116(4)  & (\V133(9)  & ~\V133(10) ))),
  V621 = ~V601 & (~V593 & (\V116(3)  & (\V133(9)  & ~\V133(10) ))),
  V622 = ~\V133(4)  & ~\V133(9) ,
  V623 = \V322(8)  & V622,
  V625 = ~\V133(9)  & \V133(7) ,
  V626 = V625 & (~V622 & \V322(8) ),
  V628 = ~V625 & (~V622 & (\V322(8)  & \V133(10) )),
  V630 = ~V625 & (~V622 & (\V116(9)  & (\V133(9)  & ~\V133(10) ))),
  V631 = ~\V133(4)  & (~\V133(9)  & ~\V133(6) ),
  V632 = \V322(10)  & V631,
  V633 = \V322(9)  & V631,
  V635 = ~\V133(9)  & \V133(7) ,
  V636 = V635 & (~V631 & \V322(10) ),
  V637 = V635 & (~V631 & \V322(9) ),
  V639 = ~V635 & (~V631 & (\V322(10)  & \V133(10) )),
  V640 = ~V635 & (~V631 & (\V322(9)  & \V133(10) )),
  V642 = ~V635 & (~V631 & (\V116(11)  & (\V133(9)  & ~\V133(10) ))),
  V643 = ~V635 & (~V631 & (\V116(10)  & (\V133(9)  & ~\V133(10) ))),
  V644 = ~\V133(4)  & (~\V133(9)  & ~\V133(1) ),
  V645 = \V322(11)  & V644,
  V647 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & ~\V133(2) )),
  V648 = V647 & (~V644 & \V322(11) ),
  V650 = ~\V133(4)  & (~\V133(9)  & \V133(3) ),
  V651 = V650 & (~V647 & (~V644 & \V322(11) )),
  V653 = ~\V133(9)  & \V133(7) ,
  V654 = V653 & (~V650 & (~V647 & (~V644 & \V322(11) ))),
  V656 = ~V653 & (~V650 & (~V647 & (~V644 & (\V322(11)  & \V133(10) )))),
  V658 = \V133(9)  & ~\V133(10) ,
  V659 = V658 & (~V653 & (~V650 & (~V647 & (~V644 & (\V116(12)  & ~\V133(10) ))))),
  V661 = ~V658 & (~V653 & (~V650 & (~V647 & (~V644 & (~\V133(4)  & (~\V133(9)  & (\V84(12)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V662 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & ~\V133(1) )),
  V663 = \V322(14)  & V662,
  V664 = \V322(13)  & V662,
  V665 = \V322(12)  & V662,
  V667 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & ~\V133(2) )),
  V668 = V667 & (~V662 & \V322(14) ),
  V669 = V667 & (~V662 & \V322(13) ),
  V670 = V667 & (~V662 & \V322(12) ),
  V672 = ~\V133(4)  & (~\V133(9)  & \V133(3) ),
  V673 = V672 & (~V667 & (~V662 & \V322(14) )),
  V674 = V672 & (~V667 & (~V662 & \V322(13) )),
  V675 = V672 & (~V667 & (~V662 & \V322(12) )),
  V677 = ~\V133(9)  & \V133(7) ,
  V678 = V677 & (~V672 & (~V667 & (~V662 & \V322(14) ))),
  V679 = V677 & (~V672 & (~V667 & (~V662 & \V322(13) ))),
  V680 = V677 & (~V672 & (~V667 & (~V662 & \V322(12) ))),
  V682 = ~V677 & (~V672 & (~V667 & (~V662 & (\V322(14)  & \V133(10) )))),
  V683 = ~V677 & (~V672 & (~V667 & (~V662 & (\V322(13)  & \V133(10) )))),
  V684 = ~V677 & (~V672 & (~V667 & (~V662 & (\V322(12)  & \V133(10) )))),
  V686 = \V133(9)  & ~\V133(10) ,
  V687 = V686 & (~V677 & (~V672 & (~V667 & (~V662 & (\V116(15)  & ~\V133(10) ))))),
  V688 = V686 & (~V677 & (~V672 & (~V667 & (~V662 & (\V116(14)  & ~\V133(10) ))))),
  V689 = V686 & (~V677 & (~V672 & (~V667 & (~V662 & (\V116(13)  & ~\V133(10) ))))),
  V691 = ~V686 & (~V677 & (~V672 & (~V667 & (~V662 & (~\V133(4)  & (~\V133(9)  & (\V84(15)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V692 = ~V686 & (~V677 & (~V672 & (~V667 & (~V662 & (~\V133(4)  & (~\V133(9)  & (\V84(14)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V693 = ~V686 & (~V677 & (~V672 & (~V667 & (~V662 & (~\V133(4)  & (~\V133(9)  & (\V84(13)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V694 = ~\V133(4)  & (~\V133(9)  & (~\V133(2)  & ~\V133(1) )),
  V695 = \V322(15)  & V694,
  V697 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & ~\V133(1) )),
  V698 = V697 & (~V694 & \V322(15) ),
  \V143(0)  = \[9] ,
  V700 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & ~\V133(2) )),
  V701 = V700 & (~V697 & (~V694 & \V322(15) )),
  V703 = ~\V133(4)  & (~\V133(9)  & \V133(3) ),
  V704 = V703 & (~V700 & (~V697 & (~V694 & \V322(15) ))),
  V706 = ~\V133(9)  & \V133(7) ,
  V707 = V706 & (~V703 & (~V700 & (~V697 & (~V694 & \V322(15) )))),
  V709 = ~V706 & (~V703 & (~V700 & (~V697 & (~V694 & (\V322(15)  & \V133(10) ))))),
  V711 = \V133(9)  & ~\V133(10) ,
  V712 = V711 & (~V706 & (~V703 & (~V700 & (~V697 & (~V694 & (\V116(16)  & ~\V133(10) )))))),
  V714 = ~V711 & (~V706 & (~V703 & (~V700 & (~V697 & (~V694 & (~\V133(4)  & (~\V133(9)  & (\V84(16)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) )))))))))))),
  V715 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & ~\V133(1) )),
  V716 = \V322(30)  & V715,
  V717 = \V322(29)  & V715,
  V718 = \V322(28)  & V715,
  V719 = \V322(27)  & V715,
  V720 = \V322(26)  & V715,
  V721 = \V322(25)  & V715,
  V722 = \V322(24)  & V715,
  V723 = \V322(23)  & V715,
  V724 = \V322(22)  & V715,
  V725 = \V322(21)  & V715,
  V726 = \V322(20)  & V715,
  V727 = \V322(19)  & V715,
  V728 = \V322(18)  & V715,
  V729 = \V322(17)  & V715,
  V730 = \V322(16)  & V715,
  V732 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & ~\V133(2) )),
  V733 = V732 & (~V715 & \V322(30) ),
  V734 = V732 & (~V715 & \V322(29) ),
  V735 = V732 & (~V715 & \V322(28) ),
  V736 = V732 & (~V715 & \V322(27) ),
  V737 = V732 & (~V715 & \V322(26) ),
  V738 = V732 & (~V715 & \V322(25) ),
  V739 = V732 & (~V715 & \V322(24) ),
  V740 = V732 & (~V715 & \V322(23) ),
  V741 = V732 & (~V715 & \V322(22) ),
  V742 = V732 & (~V715 & \V322(21) ),
  V743 = V732 & (~V715 & \V322(20) ),
  V744 = V732 & (~V715 & \V322(19) ),
  V745 = V732 & (~V715 & \V322(18) ),
  V746 = V732 & (~V715 & \V322(17) ),
  V747 = V732 & (~V715 & \V322(16) ),
  V749 = ~\V133(4)  & (~\V133(9)  & \V133(3) ),
  V750 = V749 & (~V732 & (~V715 & \V322(30) )),
  V751 = V749 & (~V732 & (~V715 & \V322(29) )),
  V752 = V749 & (~V732 & (~V715 & \V322(28) )),
  V753 = V749 & (~V732 & (~V715 & \V322(27) )),
  V754 = V749 & (~V732 & (~V715 & \V322(26) )),
  V755 = V749 & (~V732 & (~V715 & \V322(25) )),
  V756 = V749 & (~V732 & (~V715 & \V322(24) )),
  V757 = V749 & (~V732 & (~V715 & \V322(23) )),
  V758 = V749 & (~V732 & (~V715 & \V322(22) )),
  V759 = V749 & (~V732 & (~V715 & \V322(21) )),
  V760 = V749 & (~V732 & (~V715 & \V322(20) )),
  V761 = V749 & (~V732 & (~V715 & \V322(19) )),
  V762 = V749 & (~V732 & (~V715 & \V322(18) )),
  V763 = V749 & (~V732 & (~V715 & \V322(17) )),
  V764 = V749 & (~V732 & (~V715 & \V322(16) )),
  V766 = ~\V133(9)  & \V133(7) ,
  V767 = V766 & (~V749 & (~V732 & (~V715 & \V322(30) ))),
  V768 = V766 & (~V749 & (~V732 & (~V715 & \V322(29) ))),
  V769 = V766 & (~V749 & (~V732 & (~V715 & \V322(28) ))),
  V770 = V766 & (~V749 & (~V732 & (~V715 & \V322(27) ))),
  V771 = V766 & (~V749 & (~V732 & (~V715 & \V322(26) ))),
  V772 = V766 & (~V749 & (~V732 & (~V715 & \V322(25) ))),
  V773 = V766 & (~V749 & (~V732 & (~V715 & \V322(24) ))),
  V774 = V766 & (~V749 & (~V732 & (~V715 & \V322(23) ))),
  V775 = V766 & (~V749 & (~V732 & (~V715 & \V322(22) ))),
  V776 = V766 & (~V749 & (~V732 & (~V715 & \V322(21) ))),
  V777 = V766 & (~V749 & (~V732 & (~V715 & \V322(20) ))),
  V778 = V766 & (~V749 & (~V732 & (~V715 & \V322(19) ))),
  V779 = V766 & (~V749 & (~V732 & (~V715 & \V322(18) ))),
  V780 = V766 & (~V749 & (~V732 & (~V715 & \V322(17) ))),
  V781 = V766 & (~V749 & (~V732 & (~V715 & \V322(16) ))),
  V783 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(30)  & \V133(10) )))),
  V784 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(29)  & \V133(10) )))),
  V785 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(28)  & \V133(10) )))),
  V786 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(27)  & \V133(10) )))),
  V787 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(26)  & \V133(10) )))),
  V788 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(25)  & \V133(10) )))),
  V789 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(24)  & \V133(10) )))),
  V790 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(23)  & \V133(10) )))),
  V791 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(22)  & \V133(10) )))),
  V792 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(21)  & \V133(10) )))),
  V793 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(20)  & \V133(10) )))),
  V794 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(19)  & \V133(10) )))),
  V795 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(18)  & \V133(10) )))),
  V796 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(17)  & \V133(10) )))),
  V797 = ~V766 & (~V749 & (~V732 & (~V715 & (\V322(16)  & \V133(10) )))),
  V799 = \V133(9)  & ~\V133(10) ,
  \V145(1)  = \[10] ,
  \V145(0)  = \[11] ,
  V800 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(31)  & ~\V133(10) ))))),
  V801 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(30)  & ~\V133(10) ))))),
  V802 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(29)  & ~\V133(10) ))))),
  V803 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(28)  & ~\V133(10) ))))),
  V804 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(27)  & ~\V133(10) ))))),
  V805 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(26)  & ~\V133(10) ))))),
  V806 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(25)  & ~\V133(10) ))))),
  V807 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(24)  & ~\V133(10) ))))),
  V808 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(23)  & ~\V133(10) ))))),
  V809 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(22)  & ~\V133(10) ))))),
  V810 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(21)  & ~\V133(10) ))))),
  V811 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(20)  & ~\V133(10) ))))),
  V812 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(19)  & ~\V133(10) ))))),
  V813 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(18)  & ~\V133(10) ))))),
  V814 = V799 & (~V766 & (~V749 & (~V732 & (~V715 & (\V116(17)  & ~\V133(10) ))))),
  V816 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(31)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V817 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(30)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V818 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(29)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V819 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(28)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V820 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(27)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V821 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(26)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V822 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(25)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V823 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(24)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V824 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(23)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V825 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(22)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V826 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(21)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V827 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(20)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V828 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(19)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V829 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(18)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V830 = ~V799 & (~V766 & (~V749 & (~V732 & (~V715 & (~\V133(4)  & (~\V133(9)  & (\V84(17)  & (~\V133(7)  & (~\V133(10)  & (\V133(2)  & (\V133(1)  & ~\V133(3) ))))))))))),
  V831 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & (~\V133(5)  & ~\V133(1) ))),
  V832 = \V485(31)  & V831,
  V833 = \V485(30)  & V831,
  V834 = \V485(29)  & V831,
  V835 = \V485(28)  & V831,
  V836 = \V485(27)  & V831,
  V837 = \V485(26)  & V831,
  V838 = \V485(25)  & V831,
  V839 = \V485(24)  & V831,
  V840 = \V485(23)  & V831,
  V841 = \V485(22)  & V831,
  V842 = \V485(21)  & V831,
  V843 = \V485(20)  & V831,
  V844 = \V485(19)  & V831,
  V845 = \V485(18)  & V831,
  V846 = \V485(17)  & V831,
  V847 = \V485(16)  & V831,
  V848 = \V485(15)  & V831,
  V849 = \V485(14)  & V831,
  V850 = \V485(13)  & V831,
  V851 = \V485(12)  & V831,
  V852 = \V485(11)  & V831,
  V853 = \V485(10)  & V831,
  V854 = \V485(9)  & V831,
  V855 = \V485(8)  & V831,
  V856 = \V485(7)  & V831,
  V857 = \V485(6)  & V831,
  V858 = \V485(5)  & V831,
  V859 = \V485(4)  & V831,
  V860 = \V485(3)  & V831,
  V861 = \V485(2)  & V831,
  V862 = \V485(1)  & V831,
  V863 = \V485(0)  & V831,
  V865 = ~\V118(0)  & (~\V133(9)  & (\V133(5)  & (\V133(0)  & ~\V133(1) ))),
  V866 = V865 & (~V831 & \V485(31) ),
  V867 = V865 & (~V831 & \V485(30) ),
  V868 = V865 & (~V831 & \V485(29) ),
  V869 = V865 & (~V831 & \V485(28) ),
  V870 = V865 & (~V831 & \V485(27) ),
  V871 = V865 & (~V831 & \V485(26) ),
  V872 = V865 & (~V831 & \V485(25) ),
  V873 = V865 & (~V831 & \V485(24) ),
  V874 = V865 & (~V831 & \V485(23) ),
  V875 = V865 & (~V831 & \V485(22) ),
  V876 = V865 & (~V831 & \V485(21) ),
  V877 = V865 & (~V831 & \V485(20) ),
  V878 = V865 & (~V831 & \V485(19) ),
  V879 = V865 & (~V831 & \V485(18) ),
  V880 = V865 & (~V831 & \V485(17) ),
  V881 = V865 & (~V831 & \V485(16) ),
  V882 = V865 & (~V831 & \V485(15) ),
  V883 = V865 & (~V831 & \V485(14) ),
  V884 = V865 & (~V831 & \V485(13) ),
  V885 = V865 & (~V831 & \V485(12) ),
  V886 = V865 & (~V831 & \V485(11) ),
  V887 = V865 & (~V831 & \V485(10) ),
  V888 = V865 & (~V831 & \V485(9) ),
  V889 = V865 & (~V831 & \V485(8) ),
  V890 = V865 & (~V831 & \V485(7) ),
  V891 = V865 & (~V831 & \V485(6) ),
  V892 = V865 & (~V831 & \V485(5) ),
  V893 = V865 & (~V831 & \V485(4) ),
  V894 = V865 & (~V831 & \V485(3) ),
  V895 = V865 & (~V831 & \V485(2) ),
  V896 = V865 & (~V831 & \V485(1) ),
  V897 = V865 & (~V831 & \V485(0) ),
  V899 = ~\V133(9)  & (\V133(5)  & (~\V133(0)  & ~\V133(1) )),
  V900 = V899 & (~V865 & (~V831 & \V485(31) )),
  V901 = V899 & (~V865 & (~V831 & \V485(30) )),
  V902 = V899 & (~V865 & (~V831 & \V485(29) )),
  V903 = V899 & (~V865 & (~V831 & \V485(28) )),
  V904 = V899 & (~V865 & (~V831 & \V485(27) )),
  V905 = V899 & (~V865 & (~V831 & \V485(26) )),
  V906 = V899 & (~V865 & (~V831 & \V485(25) )),
  V907 = V899 & (~V865 & (~V831 & \V485(24) )),
  V908 = V899 & (~V865 & (~V831 & \V485(23) )),
  V909 = V899 & (~V865 & (~V831 & \V485(22) )),
  V910 = V899 & (~V865 & (~V831 & \V485(21) )),
  V911 = V899 & (~V865 & (~V831 & \V485(20) )),
  V912 = V899 & (~V865 & (~V831 & \V485(19) )),
  V913 = V899 & (~V865 & (~V831 & \V485(18) )),
  V914 = V899 & (~V865 & (~V831 & \V485(17) )),
  V915 = V899 & (~V865 & (~V831 & \V485(16) )),
  V916 = V899 & (~V865 & (~V831 & \V485(15) )),
  V917 = V899 & (~V865 & (~V831 & \V485(14) )),
  V918 = V899 & (~V865 & (~V831 & \V485(13) )),
  V919 = V899 & (~V865 & (~V831 & \V485(12) )),
  V920 = V899 & (~V865 & (~V831 & \V485(11) )),
  V921 = V899 & (~V865 & (~V831 & \V485(10) )),
  V922 = V899 & (~V865 & (~V831 & \V485(9) )),
  V923 = V899 & (~V865 & (~V831 & \V485(8) )),
  V924 = V899 & (~V865 & (~V831 & \V485(7) )),
  V925 = V899 & (~V865 & (~V831 & \V485(6) )),
  V926 = V899 & (~V865 & (~V831 & \V485(5) )),
  V927 = V899 & (~V865 & (~V831 & \V485(4) )),
  V928 = V899 & (~V865 & (~V831 & \V485(3) )),
  V929 = V899 & (~V865 & (~V831 & \V485(2) )),
  V930 = V899 & (~V865 & (~V831 & \V485(1) )),
  V931 = V899 & (~V865 & (~V831 & \V485(0) )),
  V933 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & (\V133(2)  & (\V133(1)  & \V133(3) )))),
  V934 = V933 & (~V899 & (~V865 & (~V831 & \V485(31) ))),
  V935 = V933 & (~V899 & (~V865 & (~V831 & \V485(30) ))),
  V936 = V933 & (~V899 & (~V865 & (~V831 & \V485(29) ))),
  V937 = V933 & (~V899 & (~V865 & (~V831 & \V485(28) ))),
  V938 = V933 & (~V899 & (~V865 & (~V831 & \V485(27) ))),
  V939 = V933 & (~V899 & (~V865 & (~V831 & \V485(26) ))),
  V940 = V933 & (~V899 & (~V865 & (~V831 & \V485(25) ))),
  V941 = V933 & (~V899 & (~V865 & (~V831 & \V485(24) ))),
  V942 = V933 & (~V899 & (~V865 & (~V831 & \V485(23) ))),
  V943 = V933 & (~V899 & (~V865 & (~V831 & \V485(22) ))),
  V944 = V933 & (~V899 & (~V865 & (~V831 & \V485(21) ))),
  V945 = V933 & (~V899 & (~V865 & (~V831 & \V485(20) ))),
  V946 = V933 & (~V899 & (~V865 & (~V831 & \V485(19) ))),
  V947 = V933 & (~V899 & (~V865 & (~V831 & \V485(18) ))),
  V948 = V933 & (~V899 & (~V865 & (~V831 & \V485(17) ))),
  V949 = V933 & (~V899 & (~V865 & (~V831 & \V485(16) ))),
  V950 = V933 & (~V899 & (~V865 & (~V831 & \V485(15) ))),
  V951 = V933 & (~V899 & (~V865 & (~V831 & \V485(14) ))),
  V952 = V933 & (~V899 & (~V865 & (~V831 & \V485(13) ))),
  V953 = V933 & (~V899 & (~V865 & (~V831 & \V485(12) ))),
  V954 = V933 & (~V899 & (~V865 & (~V831 & \V485(11) ))),
  V955 = V933 & (~V899 & (~V865 & (~V831 & \V485(10) ))),
  V956 = V933 & (~V899 & (~V865 & (~V831 & \V485(9) ))),
  V957 = V933 & (~V899 & (~V865 & (~V831 & \V485(8) ))),
  V958 = V933 & (~V899 & (~V865 & (~V831 & \V485(7) ))),
  V959 = V933 & (~V899 & (~V865 & (~V831 & \V485(6) ))),
  \V149(2)  = \[13] ,
  V960 = V933 & (~V899 & (~V865 & (~V831 & \V485(5) ))),
  V961 = V933 & (~V899 & (~V865 & (~V831 & \V485(4) ))),
  V962 = V933 & (~V899 & (~V865 & (~V831 & \V485(3) ))),
  V963 = V933 & (~V899 & (~V865 & (~V831 & \V485(2) ))),
  V964 = V933 & (~V899 & (~V865 & (~V831 & \V485(1) ))),
  V965 = V933 & (~V899 & (~V865 & (~V831 & \V485(0) ))),
  V967 = ~\V133(9)  & (\V133(7)  & ~\V133(1) ),
  V968 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(31) )))),
  V969 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(30) )))),
  V970 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(29) )))),
  V971 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(28) )))),
  V972 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(27) )))),
  V973 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(26) )))),
  V974 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(25) )))),
  V975 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(24) )))),
  V976 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(23) )))),
  V977 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(22) )))),
  V978 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(21) )))),
  V979 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(20) )))),
  V980 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(19) )))),
  V981 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(18) )))),
  V982 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(17) )))),
  V983 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(16) )))),
  V984 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(15) )))),
  V985 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(14) )))),
  V986 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(13) )))),
  V987 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(12) )))),
  V988 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(11) )))),
  V989 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(10) )))),
  V990 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(9) )))),
  V991 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(8) )))),
  V992 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(7) )))),
  V993 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(6) )))),
  V994 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(5) )))),
  V995 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(4) )))),
  V996 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(3) )))),
  V997 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(2) )))),
  V998 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(1) )))),
  V999 = V967 & (~V933 & (~V899 & (~V865 & (~V831 & \V485(0) )))),
  \V149(1)  = \[14] ,
  \V149(0)  = \[15] ,
  V1001 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(31)  & \V133(10) ))))),
  V1002 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(30)  & \V133(10) ))))),
  V1003 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(29)  & \V133(10) ))))),
  V1004 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(28)  & \V133(10) ))))),
  V1005 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(27)  & \V133(10) ))))),
  V1006 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(26)  & \V133(10) ))))),
  V1007 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(25)  & \V133(10) ))))),
  V1008 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(24)  & \V133(10) ))))),
  V1009 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(23)  & \V133(10) ))))),
  V1010 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(22)  & \V133(10) ))))),
  V1011 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(21)  & \V133(10) ))))),
  V1012 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(20)  & \V133(10) ))))),
  V1013 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(19)  & \V133(10) ))))),
  V1014 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(18)  & \V133(10) ))))),
  V1015 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(17)  & \V133(10) ))))),
  V1016 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(16)  & \V133(10) ))))),
  V1017 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(15)  & \V133(10) ))))),
  V1018 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(14)  & \V133(10) ))))),
  V1019 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(13)  & \V133(10) ))))),
  V1020 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(12)  & \V133(10) ))))),
  V1021 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(11)  & \V133(10) ))))),
  V1022 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(10)  & \V133(10) ))))),
  V1023 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(9)  & \V133(10) ))))),
  V1024 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(8)  & \V133(10) ))))),
  V1025 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(7)  & \V133(10) ))))),
  V1026 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(6)  & \V133(10) ))))),
  V1027 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(5)  & \V133(10) ))))),
  V1028 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(4)  & \V133(10) ))))),
  V1029 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(3)  & \V133(10) ))))),
  V1030 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(2)  & \V133(10) ))))),
  V1031 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(1)  & \V133(10) ))))),
  V1032 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V485(0)  & \V133(10) ))))),
  V1034 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(31)  & (\V133(9)  & ~\V133(10) )))))),
  V1035 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(30)  & (\V133(9)  & ~\V133(10) )))))),
  V1036 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(29)  & (\V133(9)  & ~\V133(10) )))))),
  V1037 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(28)  & (\V133(9)  & ~\V133(10) )))))),
  V1038 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(27)  & (\V133(9)  & ~\V133(10) )))))),
  V1039 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(26)  & (\V133(9)  & ~\V133(10) )))))),
  V1040 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(25)  & (\V133(9)  & ~\V133(10) )))))),
  V1041 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(24)  & (\V133(9)  & ~\V133(10) )))))),
  V1042 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(23)  & (\V133(9)  & ~\V133(10) )))))),
  V1043 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(22)  & (\V133(9)  & ~\V133(10) )))))),
  V1044 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(21)  & (\V133(9)  & ~\V133(10) )))))),
  V1045 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(20)  & (\V133(9)  & ~\V133(10) )))))),
  V1046 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(19)  & (\V133(9)  & ~\V133(10) )))))),
  V1047 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(18)  & (\V133(9)  & ~\V133(10) )))))),
  V1048 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(17)  & (\V133(9)  & ~\V133(10) )))))),
  V1049 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(16)  & (\V133(9)  & ~\V133(10) )))))),
  V1050 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(15)  & (\V133(9)  & ~\V133(10) )))))),
  V1051 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(14)  & (\V133(9)  & ~\V133(10) )))))),
  V1052 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(13)  & (\V133(9)  & ~\V133(10) )))))),
  V1053 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(12)  & (\V133(9)  & ~\V133(10) )))))),
  V1054 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(11)  & (\V133(9)  & ~\V133(10) )))))),
  V1055 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(10)  & (\V133(9)  & ~\V133(10) )))))),
  V1056 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(9)  & (\V133(9)  & ~\V133(10) )))))),
  V1057 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(8)  & (\V133(9)  & ~\V133(10) )))))),
  V1058 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(7)  & (\V133(9)  & ~\V133(10) )))))),
  V1059 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(6)  & (\V133(9)  & ~\V133(10) )))))),
  V1060 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(5)  & (\V133(9)  & ~\V133(10) )))))),
  V1061 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(4)  & (\V133(9)  & ~\V133(10) )))))),
  V1062 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(3)  & (\V133(9)  & ~\V133(10) )))))),
  V1063 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V133(9)  & (\V116(2)  & ~\V133(10) )))))),
  V1064 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V116(1)  & (\V133(9)  & ~\V133(10) )))))),
  V1065 = ~V967 & (~V933 & (~V899 & (~V865 & (~V831 & (\V133(9)  & (\V116(0)  & ~\V133(10) )))))),
  V1066 = ~\V133(4)  & (~\V133(9)  & (~\V133(6)  & (~\V133(5)  & (~\V133(2)  & ~\V133(1) )))),
  V1067 = \V84(31)  & V1066,
  V1068 = \V84(30)  & V1066,
  V1069 = \V84(29)  & V1066,
  V1070 = \V84(28)  & V1066,
  V1071 = \V84(27)  & V1066,
  V1072 = \V84(26)  & V1066,
  V1073 = \V84(25)  & V1066,
  V1074 = \V84(24)  & V1066,
  V1075 = \V84(23)  & V1066,
  V1076 = \V84(22)  & V1066,
  V1077 = \V84(21)  & V1066,
  V1078 = \V84(20)  & V1066,
  V1079 = \V84(19)  & V1066,
  V1080 = \V84(18)  & V1066,
  V1081 = \V84(17)  & V1066,
  V1083 = ~\V133(9)  & (\V133(7)  & (~\V133(2)  & ~\V133(1) )),
  V1084 = V1083 & (~V1066 & \V84(31) ),
  V1085 = V1083 & (~V1066 & \V84(30) ),
  V1086 = V1083 & (~V1066 & \V84(29) ),
  V1087 = V1083 & (~V1066 & \V84(28) ),
  V1088 = V1083 & (~V1066 & \V84(27) ),
  V1089 = V1083 & (~V1066 & \V84(26) ),
  V1090 = V1083 & (~V1066 & \V84(25) ),
  V1091 = V1083 & (~V1066 & \V84(24) ),
  V1092 = V1083 & (~V1066 & \V84(23) ),
  V1093 = V1083 & (~V1066 & \V84(22) ),
  V1094 = V1083 & (~V1066 & \V84(21) ),
  V1095 = V1083 & (~V1066 & \V84(20) ),
  V1096 = V1083 & (~V1066 & \V84(19) ),
  V1097 = V1083 & (~V1066 & \V84(18) ),
  V1098 = V1083 & (~V1066 & \V84(17) ),
  V1100 = ~V1083 & (~V1066 & (\V84(31)  & \V133(10) )),
  V1101 = ~V1083 & (~V1066 & (\V84(30)  & \V133(10) )),
  V1102 = ~V1083 & (~V1066 & (\V84(29)  & \V133(10) )),
  V1103 = ~V1083 & (~V1066 & (\V84(28)  & \V133(10) )),
  V1104 = ~V1083 & (~V1066 & (\V84(27)  & \V133(10) )),
  V1105 = ~V1083 & (~V1066 & (\V84(26)  & \V133(10) )),
  V1106 = ~V1083 & (~V1066 & (\V84(25)  & \V133(10) )),
  V1107 = ~V1083 & (~V1066 & (\V84(24)  & \V133(10) )),
  V1108 = ~V1083 & (~V1066 & (\V84(23)  & \V133(10) )),
  V1109 = ~V1083 & (~V1066 & (\V84(22)  & \V133(10) )),
  V1110 = ~V1083 & (~V1066 & (\V84(21)  & \V133(10) )),
  V1111 = ~V1083 & (~V1066 & (\V84(20)  & \V133(10) )),
  V1112 = ~V1083 & (~V1066 & (\V84(19)  & \V133(10) )),
  V1113 = ~V1083 & (~V1066 & (\V84(18)  & \V133(10) )),
  V1114 = ~V1083 & (~V1066 & (\V84(17)  & \V133(10) )),
  V1116 = ~\V118(1)  & (~\V118(0)  & (~\V133(9)  & (~\V133(7)  & (~\V133(10)  & (\V133(5)  & (~\V133(2)  & ~\V133(1) )))))),
  V1117 = V1116 & (~V1083 & (~V1066 & ~\V133(10) )),
  V1119 = ~V1116 & (~V1083 & (~V1066 & (\V116(14)  & (\V133(9)  & ~\V133(10) )))),
  V1120 = ~V1116 & (~V1083 & (~V1066 & (\V116(13)  & (\V133(9)  & ~\V133(10) )))),
  V1121 = ~V1116 & (~V1083 & (~V1066 & (\V116(12)  & (\V133(9)  & ~\V133(10) )))),
  V1122 = ~V1116 & (~V1083 & (~V1066 & (\V116(11)  & (\V133(9)  & ~\V133(10) )))),
  V1123 = ~V1116 & (~V1083 & (~V1066 & (\V116(10)  & (\V133(9)  & ~\V133(10) )))),
  V1124 = ~V1116 & (~V1083 & (~V1066 & (\V116(9)  & (\V133(9)  & ~\V133(10) )))),
  V1125 = ~V1116 & (~V1083 & (~V1066 & (\V116(8)  & (\V133(9)  & ~\V133(10) )))),
  V1126 = ~V1116 & (~V1083 & (~V1066 & (\V116(7)  & (\V133(9)  & ~\V133(10) )))),
  V1127 = ~V1116 & (~V1083 & (~V1066 & (\V116(6)  & (\V133(9)  & ~\V133(10) )))),
  V1128 = ~V1116 & (~V1083 & (~V1066 & (\V116(5)  & (\V133(9)  & ~\V133(10) )))),
  V1129 = ~V1116 & (~V1083 & (~V1066 & (\V116(4)  & (\V133(9)  & ~\V133(10) )))),
  V1130 = ~V1116 & (~V1083 & (~V1066 & (\V116(3)  & (\V133(9)  & ~\V133(10) )))),
  V1131 = ~V1116 & (~V1083 & (~V1066 & (\V133(9)  & (\V116(2)  & ~\V133(10) )))),
  V1132 = ~V1116 & (~V1083 & (~V1066 & (\V116(1)  & (\V133(9)  & ~\V133(10) )))),
  V1133 = ~V1116 & (~V1083 & (~V1066 & (\V133(9)  & (\V116(0)  & ~\V133(10) )))),
  V1134 = ~\V133(9)  & (~\V133(8)  & (\V133(7)  & ~\V133(10) )),
  V1135 = \V121(16)  & V1134,
  V1137 = \V133(9)  & ~\V133(10) ,
  V1139 = ~\V133(10)  & (\V133(2)  & \V133(1) ),
  V1141 = ~V1139 & (~V1137 & (~V1134 & (\V119(0)  & \V133(10) ))),
  V1143 = ~\V133(9)  & (\V133(8)  & ~\V133(10) ),
  V1144 = V1143 & (~V1139 & (~V1137 & (~V1134 & ~\V133(10) ))),
  V1146 = ~\V133(9)  & (~\V133(7)  & (~\V133(10)  & ~\V133(1) )),
  V1147 = V1146 & (~V1143 & (~V1139 & (~V1137 & (~V1134 & ~\V133(10) )))),
  V1149 = ~V1146 & (~V1143 & (~V1139 & (~V1137 & (~V1134 & ~\V133(10) )))),
  V1150 = ~\V133(9)  & (\V133(7)  & ~\V133(10) ),
  V1151 = \V121(17)  & V1150,
  V1153 = ~\V133(9)  & (~\V133(10)  & (\V133(2)  & \V133(1) )),
  V1154 = V1153 & ~V1150,
  V1156 = ~V1153 & (~V1150 & (\V122(0)  & \V133(10) )),
  \V485(27)  = V553 | (V524 | (V491 | (V430 | V393))),
  \V134(0)  = \[0] ,
  \V485(26)  = V553 | (V525 | (V492 | (V432 | V394))),
  \V485(29)  = V553 | (V522 | (V489 | (V426 | V391))),
  \V485(28)  = V553 | (V523 | (V490 | (V428 | V392))),
  \V485(21)  = V553 | (V530 | (V497 | (V442 | V399))),
  \V485(20)  = V553 | (V531 | (V498 | (V444 | V400))),
  \V485(23)  = V553 | (V528 | (V495 | (V438 | V397))),
  \V485(22)  = V553 | (V529 | (V496 | (V440 | V398))),
  \V485(25)  = V553 | (V526 | (V493 | (V434 | V395))),
  \V485(24)  = V553 | (V527 | (V494 | (V436 | V396))),
  \V136(1)  = \[1] ,
  \V485(17)  = V553 | (V534 | (V501 | (V450 | V403))),
  \V136(0)  = \[2] ,
  \V485(16)  = V553 | (V535 | (V502 | (V452 | V404))),
  \V485(19)  = V553 | (V532 | (V499 | (V446 | V401))),
  \V485(18)  = V553 | (V533 | (V500 | (V448 | V402))),
  \V322(3)  = V383 | (V351 | (V388 | V263)),
  \V485(11)  = V553 | (V540 | (V507 | (V462 | V409))),
  \V322(2)  = V384 | (V352 | (V388 | V264)),
  \V485(10)  = V553 | (V541 | (V508 | (V464 | V410))),
  \V322(5)  = V381 | (V349 | (V388 | V261)),
  \V485(13)  = V553 | (V538 | (V505 | (V458 | V407))),
  \V322(4)  = V382 | (V350 | (V388 | V262)),
  \V485(12)  = V553 | (V539 | (V506 | (V460 | V408))),
  \V485(15)  = V553 | (V536 | (V503 | (V454 | V405))),
  \V485(14)  = V553 | (V537 | (V504 | (V456 | V406))),
  \V322(1)  = V385 | (V353 | (V388 | V265)),
  \V322(0)  = V386 | (V354 | (V388 | V266)),
  \V322(7)  = V388 | (V379 | (V347 | (V314 | V259))),
  \V322(6)  = V380 | (V348 | (V388 | V260)),
  \V322(9)  = V388 | (V377 | (V345 | (V310 | V257))),
  \V322(8)  = V388 | (V378 | (V346 | (V312 | V258))),
  \V165(11)  = \[20] ,
  \V197(3)  = \[60] ,
  \V165(10)  = \[21] ,
  \V197(2)  = \[61] ,
  \V165(13)  = \[18] ,
  \V197(5)  = \[58] ,
  \V165(12)  = \[19] ,
  \V197(4)  = \[59] ,
  \V197(27)  = \[36] ,
  \V197(26)  = \[37] ,
  \V165(14)  = \[17] ,
  \V197(29)  = \[34] ,
  \V197(1)  = \[62] ,
  \V197(28)  = \[35] ,
  \V485(31)  = V553 | (V520 | (V487 | (V422 | V389))),
  \V197(0)  = \[63] ,
  \V485(30)  = V553 | (V521 | (V488 | (V424 | V390))),
  \V197(7)  = \[56] ,
  \V197(6)  = \[57] ,
  \V197(21)  = \[42] ,
  \V197(9)  = \[54] ,
  \V197(20)  = \[43] ,
  \V197(8)  = \[55] ,
  \V197(23)  = \[40] ,
  \V197(22)  = \[41] ,
  \V197(25)  = \[38] ,
  \V197(24)  = \[39] ,
  \V213(0)  = \[79] ,
  \V197(17)  = \[46] ,
  \V197(16)  = \[47] ,
  \V197(19)  = \[44] ,
  \V197(18)  = \[45] ,
  \[10]  = V642 | (V639 | (V636 | V632)),
  \[11]  = V643 | (V640 | (V637 | V633)),
  \[12]  = V661 | (V659 | (V656 | (V654 | (V651 | (V648 | V645))))),
  \[13]  = V691 | (V687 | (V682 | (V678 | (V673 | (V668 | V663))))),
  \[14]  = V692 | (V688 | (V683 | (V679 | (V674 | (V669 | V664))))),
  \[15]  = V693 | (V689 | (V684 | (V680 | (V675 | (V670 | V665))))),
  \[16]  = V714 | (V712 | (V709 | (V707 | (V704 | (V701 | (V698 | V695)))))),
  \V197(11)  = \[52] ,
  \[17]  = V816 | (V800 | (V783 | (V767 | (V750 | (V733 | V716))))),
  \V197(10)  = \[53] ,
  \[18]  = V817 | (V801 | (V784 | (V768 | (V751 | (V734 | V717))))),
  \V197(13)  = \[50] ,
  \[19]  = V818 | (V802 | (V785 | (V769 | (V752 | (V735 | V718))))),
  \V197(12)  = \[51] ,
  \V197(15)  = \[48] ,
  \V197(14)  = \[49] ,
  \[20]  = V819 | (V803 | (V786 | (V770 | (V753 | (V736 | V719))))),
  \[21]  = V820 | (V804 | (V787 | (V771 | (V754 | (V737 | V720))))),
  \[22]  = V821 | (V805 | (V788 | (V772 | (V755 | (V738 | V721))))),
  \[23]  = V822 | (V806 | (V789 | (V773 | (V756 | (V739 | V722))))),
  \[24]  = V823 | (V807 | (V790 | (V774 | (V757 | (V740 | V723))))),
  \[25]  = V824 | (V808 | (V791 | (V775 | (V758 | (V741 | V724))))),
  \[26]  = V825 | (V809 | (V792 | (V776 | (V759 | (V742 | V725))))),
  \[27]  = V826 | (V810 | (V793 | (V777 | (V760 | (V743 | V726))))),
  \[28]  = V827 | (V811 | (V794 | (V778 | (V761 | (V744 | V727))))),
  \[29]  = V828 | (V812 | (V795 | (V779 | (V762 | (V745 | V728))))),
  \[30]  = V829 | (V813 | (V796 | (V780 | (V763 | (V746 | V729))))),
  \V142(3)  = \[5] ,
  \[31]  = V830 | (V814 | (V797 | (V781 | (V764 | (V747 | V730))))),
  \V142(2)  = \[6] ,
  \[32]  = V1034 | (V1001 | (V968 | (V934 | (V900 | (V866 | V832))))),
  \V142(5)  = \[3] ,
  \[33]  = V1035 | (V1002 | (V969 | (V935 | (V901 | (V867 | V833))))),
  \V142(4)  = \[4] ,
  \[34]  = V1036 | (V1003 | (V970 | (V936 | (V902 | (V868 | V834))))),
  \[35]  = V1037 | (V1004 | (V971 | (V937 | (V903 | (V869 | V835))))),
  \[36]  = V1038 | (V1005 | (V972 | (V938 | (V904 | (V870 | V836))))),
  \V197(31)  = \[32] ,
  \V142(1)  = \[7] ,
  \[37]  = V1039 | (V1006 | (V973 | (V939 | (V905 | (V871 | V837))))),
  \V197(30)  = \[33] ,
  \V142(0)  = \[8] ,
  \[38]  = V1040 | (V1007 | (V974 | (V940 | (V906 | (V872 | V838))))),
  \[39]  = V1041 | (V1008 | (V975 | (V941 | (V907 | (V873 | V839))))),
  \[40]  = V1042 | (V1009 | (V976 | (V942 | (V908 | (V874 | V840))))),
  \[41]  = V1043 | (V1010 | (V977 | (V943 | (V909 | (V875 | V841))))),
  \[42]  = V1044 | (V1011 | (V978 | (V944 | (V910 | (V876 | V842))))),
  \[43]  = V1045 | (V1012 | (V979 | (V945 | (V911 | (V877 | V843))))),
  \[44]  = V1046 | (V1013 | (V980 | (V946 | (V912 | (V878 | V844))))),
  \[45]  = V1047 | (V1014 | (V981 | (V947 | (V913 | (V879 | V845))))),
  \[46]  = V1048 | (V1015 | (V982 | (V948 | (V914 | (V880 | V846))))),
  \[47]  = V1049 | (V1016 | (V983 | (V949 | (V915 | (V881 | V847))))),
  \[48]  = V1050 | (V1017 | (V984 | (V950 | (V916 | (V882 | V848))))),
  \[49]  = V1051 | (V1018 | (V985 | (V951 | (V917 | (V883 | V849))))),
  \[50]  = V1052 | (V1019 | (V986 | (V952 | (V918 | (V884 | V850))))),
  \V322(27)  = V388 | (V359 | (V327 | (V274 | V239))),
  \[51]  = V1053 | (V1020 | (V987 | (V953 | (V919 | (V885 | V851))))),
  \V322(26)  = V388 | (V360 | (V328 | (V276 | V240))),
  \[52]  = V1054 | (V1021 | (V988 | (V954 | (V920 | (V886 | V852))))),
  \V322(29)  = V388 | (V357 | (V325 | (V270 | V237))),
  \[53]  = V1055 | (V1022 | (V989 | (V955 | (V921 | (V887 | V853))))),
  \V322(28)  = V388 | (V358 | (V326 | (V272 | V238))),
  \[54]  = V1056 | (V1023 | (V990 | (V956 | (V922 | (V888 | V854))))),
  \V165(3)  = \[28] ,
  \V212(11)  = \[67] ,
  \[55]  = V1057 | (V1024 | (V991 | (V957 | (V923 | (V889 | V855))))),
  \V165(2)  = \[29] ,
  \V212(10)  = \[68] ,
  \[56]  = V1058 | (V1025 | (V992 | (V958 | (V924 | (V890 | V856))))),
  \V165(5)  = \[26] ,
  \V212(13)  = \[65] ,
  \[57]  = V1059 | (V1026 | (V993 | (V959 | (V925 | (V891 | V857))))),
  \V165(4)  = \[27] ,
  \V212(12)  = \[66] ,
  \[58]  = V1060 | (V1027 | (V994 | (V960 | (V926 | (V892 | V858))))),
  \V146(0)  = \[12] ,
  \[59]  = V1061 | (V1028 | (V995 | (V961 | (V927 | (V893 | V859))))),
  \V212(14)  = \[64] ,
  \V322(21)  = V388 | (V365 | (V333 | (V286 | V245))),
  \V165(1)  = \[30] ,
  \V322(20)  = V388 | (V366 | (V334 | (V288 | V246))),
  \V165(0)  = \[31] ,
  \V322(23)  = V388 | (V363 | (V331 | (V282 | V243))),
  \V322(22)  = V388 | (V364 | (V332 | (V284 | V244))),
  \V322(25)  = V388 | (V361 | (V329 | (V278 | V241))),
  \V322(24)  = V388 | (V362 | (V330 | (V280 | V242))),
  \[60]  = V1062 | (V1029 | (V996 | (V962 | (V928 | (V894 | V860))))),
  \V322(17)  = V388 | (V369 | (V337 | (V294 | V249))),
  \V165(7)  = \[24] ,
  \[61]  = V1063 | (V1030 | (V997 | (V963 | (V929 | (V895 | V861))))),
  \V322(16)  = V388 | (V370 | (V338 | (V296 | V250))),
  \V165(6)  = \[25] ,
  \[62]  = V1064 | (V1031 | (V998 | (V964 | (V930 | (V896 | V862))))),
  \V322(19)  = V388 | (V367 | (V335 | (V290 | V247))),
  \V165(9)  = \[22] ,
  \[63]  = V1065 | (V1032 | (V999 | (V965 | (V931 | (V897 | V863))))),
  \V322(18)  = V388 | (V368 | (V336 | (V292 | V248))),
  \V165(8)  = \[23] ,
  \[64]  = V1119 | (V1117 | (V1100 | (V1084 | V1067))),
  \[65]  = V1120 | (V1117 | (V1101 | (V1085 | V1068))),
  \[66]  = V1121 | (V1117 | (V1102 | (V1086 | V1069))),
  \[67]  = V1122 | (V1117 | (V1103 | (V1087 | V1070))),
  \[68]  = V1123 | (V1117 | (V1104 | (V1088 | V1071))),
  \[69]  = V1124 | (V1117 | (V1105 | (V1089 | V1072))),
  \V322(11)  = V388 | (V375 | (V343 | (V306 | V255))),
  \V322(10)  = V388 | (V376 | (V344 | (V308 | V256))),
  \V322(13)  = V388 | (V373 | (V341 | (V302 | V253))),
  \V322(12)  = V388 | (V374 | (V342 | (V304 | V254))),
  \V322(15)  = V388 | (V371 | (V339 | (V298 | V251))),
  \V322(14)  = V388 | (V372 | (V340 | (V300 | V252))),
  \[70]  = V1125 | (V1117 | (V1106 | (V1090 | V1073))),
  \[71]  = V1126 | (V1117 | (V1107 | (V1091 | V1074))),
  \V485(3)  = V553 | (V548 | (V515 | (V478 | V417))),
  \[72]  = V1127 | (V1117 | (V1108 | (V1092 | V1075))),
  \V485(2)  = V553 | (V549 | (V516 | (V480 | V418))),
  \[73]  = V1128 | (V1117 | (V1109 | (V1093 | V1076))),
  \V485(5)  = V553 | (V546 | (V513 | (V474 | V415))),
  \[74]  = V1129 | (V1117 | (V1110 | (V1094 | V1077))),
  \V485(4)  = V553 | (V547 | (V514 | (V476 | V416))),
  \[75]  = V1130 | (V1117 | (V1111 | (V1095 | V1078))),
  \[76]  = V1131 | (V1117 | (V1112 | (V1096 | V1079))),
  \[77]  = V1132 | (V1117 | (V1113 | (V1097 | V1080))),
  \V485(1)  = V553 | (V550 | (V517 | (V482 | V419))),
  \[78]  = V1133 | (V1117 | (V1114 | (V1098 | V1081))),
  \V485(0)  = V553 | (V551 | (V518 | (V484 | V420))),
  \[79]  = V1144 | (V1141 | (V1147 | (V1149 | V1135))),
  \V485(7)  = V553 | (V544 | (V511 | (V470 | V413))),
  \V485(6)  = V553 | (V545 | (V512 | (V472 | V414))),
  \V485(9)  = V553 | (V542 | (V509 | (V466 | V411))),
  \[80]  = V1156 | (V1154 | V1151),
  \V485(8)  = V553 | (V543 | (V510 | (V468 | V412))),
  \V322(30)  = V388 | (V356 | (V324 | (V268 | V236))),
  \V150(0)  = \[16] ;
endmodule

