//NOTE: no-implementation module stub

module RTBmem (
    input DSPCLK,
    input [4:0] BTB_wa,
    input RTB_web,
    input PWRDn,
    input [11:0] RTB_wd,
    input [4:0] BTB_ra,
    output [11:0] RTB_rd
);

endmodule
